magic
tech gf180mcuD
magscale 1 10
timestamp 1757859636
<< error_p >>
rect -48 1465 -37 1511
rect -48 553 -37 599
rect -48 433 -37 479
rect -48 -479 -37 -433
rect -48 -599 -37 -553
rect -48 -1511 -37 -1465
<< nwell >>
rect -300 -1642 300 1642
<< pmos >>
rect -50 632 50 1432
rect -50 -400 50 400
rect -50 -1432 50 -632
<< pdiff >>
rect -138 1419 -50 1432
rect -138 645 -125 1419
rect -79 645 -50 1419
rect -138 632 -50 645
rect 50 1419 138 1432
rect 50 645 79 1419
rect 125 645 138 1419
rect 50 632 138 645
rect -138 387 -50 400
rect -138 -387 -125 387
rect -79 -387 -50 387
rect -138 -400 -50 -387
rect 50 387 138 400
rect 50 -387 79 387
rect 125 -387 138 387
rect 50 -400 138 -387
rect -138 -645 -50 -632
rect -138 -1419 -125 -645
rect -79 -1419 -50 -645
rect -138 -1432 -50 -1419
rect 50 -645 138 -632
rect 50 -1419 79 -645
rect 125 -1419 138 -645
rect 50 -1432 138 -1419
<< pdiffc >>
rect -125 645 -79 1419
rect 79 645 125 1419
rect -125 -387 -79 387
rect 79 -387 125 387
rect -125 -1419 -79 -645
rect 79 -1419 125 -645
<< nsubdiff >>
rect -276 1546 276 1618
rect -276 1502 -204 1546
rect -276 -1502 -263 1502
rect -217 -1502 -204 1502
rect 204 1502 276 1546
rect -276 -1546 -204 -1502
rect 204 -1502 217 1502
rect 263 -1502 276 1502
rect 204 -1546 276 -1502
rect -276 -1618 276 -1546
<< nsubdiffcont >>
rect -263 -1502 -217 1502
rect 217 -1502 263 1502
<< polysilicon >>
rect -50 1511 50 1524
rect -50 1465 -37 1511
rect 37 1465 50 1511
rect -50 1432 50 1465
rect -50 599 50 632
rect -50 553 -37 599
rect 37 553 50 599
rect -50 540 50 553
rect -50 479 50 492
rect -50 433 -37 479
rect 37 433 50 479
rect -50 400 50 433
rect -50 -433 50 -400
rect -50 -479 -37 -433
rect 37 -479 50 -433
rect -50 -492 50 -479
rect -50 -553 50 -540
rect -50 -599 -37 -553
rect 37 -599 50 -553
rect -50 -632 50 -599
rect -50 -1465 50 -1432
rect -50 -1511 -37 -1465
rect 37 -1511 50 -1465
rect -50 -1524 50 -1511
<< polycontact >>
rect -37 1465 37 1511
rect -37 553 37 599
rect -37 433 37 479
rect -37 -479 37 -433
rect -37 -599 37 -553
rect -37 -1511 37 -1465
<< metal1 >>
rect -263 1559 263 1605
rect -263 1502 -217 1559
rect -48 1465 -37 1511
rect 37 1465 48 1511
rect 217 1502 263 1559
rect -125 1419 -79 1430
rect -125 634 -79 645
rect 79 1419 125 1430
rect 79 634 125 645
rect -48 553 -37 599
rect 37 553 48 599
rect -48 433 -37 479
rect 37 433 48 479
rect -125 387 -79 398
rect -125 -398 -79 -387
rect 79 387 125 398
rect 79 -398 125 -387
rect -48 -479 -37 -433
rect 37 -479 48 -433
rect -48 -599 -37 -553
rect 37 -599 48 -553
rect -125 -645 -79 -634
rect -125 -1430 -79 -1419
rect 79 -645 125 -634
rect 79 -1430 125 -1419
rect -263 -1559 -217 -1502
rect -48 -1511 -37 -1465
rect 37 -1511 48 -1465
rect 217 -1559 263 -1502
rect -263 -1605 263 -1559
<< properties >>
string FIXED_BBOX -240 -1582 240 1582
string gencell pfet_03v3
string library gf180mcu
string parameters w 4 l 0.5 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
