magic
tech gf180mcuD
magscale 1 10
timestamp 1756981609
<< nwell >>
rect -654 -310 654 310
<< pmos >>
rect -404 -100 -204 100
rect -100 -100 100 100
rect 204 -100 404 100
<< pdiff >>
rect -492 87 -404 100
rect -492 -87 -479 87
rect -433 -87 -404 87
rect -492 -100 -404 -87
rect -204 87 -100 100
rect -204 -87 -175 87
rect -129 -87 -100 87
rect -204 -100 -100 -87
rect 100 87 204 100
rect 100 -87 129 87
rect 175 -87 204 87
rect 100 -100 204 -87
rect 404 87 492 100
rect 404 -87 433 87
rect 479 -87 492 87
rect 404 -100 492 -87
<< pdiffc >>
rect -479 -87 -433 87
rect -175 -87 -129 87
rect 129 -87 175 87
rect 433 -87 479 87
<< nsubdiff >>
rect -630 214 630 286
rect -630 170 -558 214
rect -630 -170 -617 170
rect -571 -170 -558 170
rect 558 170 630 214
rect -630 -214 -558 -170
rect 558 -170 571 170
rect 617 -170 630 170
rect 558 -214 630 -170
rect -630 -286 630 -214
<< nsubdiffcont >>
rect -617 -170 -571 170
rect 571 -170 617 170
<< polysilicon >>
rect -404 179 -204 192
rect -404 133 -391 179
rect -217 133 -204 179
rect -404 100 -204 133
rect -100 179 100 192
rect -100 133 -87 179
rect 87 133 100 179
rect -100 100 100 133
rect 204 179 404 192
rect 204 133 217 179
rect 391 133 404 179
rect 204 100 404 133
rect -404 -133 -204 -100
rect -404 -179 -391 -133
rect -217 -179 -204 -133
rect -404 -192 -204 -179
rect -100 -133 100 -100
rect -100 -179 -87 -133
rect 87 -179 100 -133
rect -100 -192 100 -179
rect 204 -133 404 -100
rect 204 -179 217 -133
rect 391 -179 404 -133
rect 204 -192 404 -179
<< polycontact >>
rect -391 133 -217 179
rect -87 133 87 179
rect 217 133 391 179
rect -391 -179 -217 -133
rect -87 -179 87 -133
rect 217 -179 391 -133
<< metal1 >>
rect -617 227 617 273
rect -617 170 -571 227
rect -402 133 -391 179
rect -217 133 -206 179
rect -98 133 -87 179
rect 87 133 98 179
rect 206 133 217 179
rect 391 133 402 179
rect 571 170 617 227
rect -479 87 -433 98
rect -479 -98 -433 -87
rect -175 87 -129 98
rect -175 -98 -129 -87
rect 129 87 175 98
rect 129 -98 175 -87
rect 433 87 479 98
rect 433 -98 479 -87
rect -617 -227 -571 -170
rect -402 -179 -391 -133
rect -217 -179 -206 -133
rect -98 -179 -87 -133
rect 87 -179 98 -133
rect 206 -179 217 -133
rect 391 -179 402 -133
rect 571 -227 617 -170
rect -617 -273 617 -227
<< properties >>
string FIXED_BBOX -594 -250 594 250
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
