* NGSPICE file created from xschem_diffpairtest.ext - technology: gf180mcuD

.subckt nfet_03v3_3TMVZR a_n934_n336#
X0 a_n204_n150# a_n404_n242# a_n508_n150# a_n934_n336# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X1 a_n508_n150# a_n708_n242# a_n796_n150# a_n934_n336# nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X2 a_404_n150# a_204_n242# a_100_n150# a_n934_n336# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X3 a_100_n150# a_n100_n242# a_n204_n150# a_n934_n336# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X4 a_708_n150# a_508_n242# a_404_n150# a_n934_n336# nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
.ends

.subckt xschem_diffpairtest
XXM9 VSUBS nfet_03v3_3TMVZR
XXM20 VSUBS nfet_03v3_3TMVZR
XXM10 VSUBS nfet_03v3_3TMVZR
XXM21 VSUBS nfet_03v3_3TMVZR
.ends

