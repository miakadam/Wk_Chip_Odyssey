magic
tech gf180mcuD
magscale 1 10
timestamp 1756981609
<< error_p >>
rect -130 113 -119 159
rect 54 113 65 159
rect -130 -159 -119 -113
rect 54 -159 65 -113
<< nwell >>
rect -382 -290 382 290
<< pmos >>
rect -132 -80 -52 80
rect 52 -80 132 80
<< pdiff >>
rect -220 67 -132 80
rect -220 -67 -207 67
rect -161 -67 -132 67
rect -220 -80 -132 -67
rect -52 67 52 80
rect -52 -67 -23 67
rect 23 -67 52 67
rect -52 -80 52 -67
rect 132 67 220 80
rect 132 -67 161 67
rect 207 -67 220 67
rect 132 -80 220 -67
<< pdiffc >>
rect -207 -67 -161 67
rect -23 -67 23 67
rect 161 -67 207 67
<< nsubdiff >>
rect -358 194 358 266
rect -358 150 -286 194
rect -358 -150 -345 150
rect -299 -150 -286 150
rect 286 150 358 194
rect -358 -194 -286 -150
rect 286 -150 299 150
rect 345 -150 358 150
rect 286 -194 358 -150
rect -358 -266 358 -194
<< nsubdiffcont >>
rect -345 -150 -299 150
rect 299 -150 345 150
<< polysilicon >>
rect -132 159 -52 172
rect -132 113 -119 159
rect -65 113 -52 159
rect -132 80 -52 113
rect 52 159 132 172
rect 52 113 65 159
rect 119 113 132 159
rect 52 80 132 113
rect -132 -113 -52 -80
rect -132 -159 -119 -113
rect -65 -159 -52 -113
rect -132 -172 -52 -159
rect 52 -113 132 -80
rect 52 -159 65 -113
rect 119 -159 132 -113
rect 52 -172 132 -159
<< polycontact >>
rect -119 113 -65 159
rect 65 113 119 159
rect -119 -159 -65 -113
rect 65 -159 119 -113
<< metal1 >>
rect -345 207 345 253
rect -345 150 -299 207
rect -130 113 -119 159
rect -65 113 -54 159
rect 54 113 65 159
rect 119 113 130 159
rect 299 150 345 207
rect -207 67 -161 78
rect -207 -78 -161 -67
rect -23 67 23 78
rect -23 -78 23 -67
rect 161 67 207 78
rect 161 -78 207 -67
rect -345 -207 -299 -150
rect -130 -159 -119 -113
rect -65 -159 -54 -113
rect 54 -159 65 -113
rect 119 -159 130 -113
rect 299 -207 345 -150
rect -345 -253 345 -207
<< properties >>
string FIXED_BBOX -322 -230 322 230
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.8 l 0.4 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
