magic
tech gf180mcuD
magscale 1 10
timestamp 1758099978
<< metal1 >>
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 5430 5716 5512 5728
rect 14902 5716 14984 5728
rect 24374 5717 24456 5729
rect 33846 5717 33928 5729
rect 43318 5717 43400 5729
rect 52790 5717 52872 5729
rect 5430 5660 5444 5716
rect 5500 5660 5644 5716
rect 14902 5660 14916 5716
rect 14972 5660 15116 5716
rect 24374 5661 24388 5717
rect 24444 5661 24588 5717
rect 33846 5661 33860 5717
rect 33916 5661 34060 5717
rect 43318 5661 43332 5717
rect 43388 5661 43532 5717
rect 52790 5661 52804 5717
rect 52860 5661 53004 5717
rect 5430 5648 5512 5660
rect 14902 5648 14984 5660
rect 24374 5649 24456 5661
rect 33846 5649 33928 5661
rect 43318 5649 43400 5661
rect 52790 5649 52872 5661
rect 230 2890 234 4510
rect 47784 4311 48004 4321
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 47784 3501 48004 3511
rect 940 3346 1020 3356
rect 940 3290 952 3346
rect 1008 3290 1020 3346
rect 940 3280 1020 3290
rect 1156 2431 1166 2507
rect 1246 2431 1256 2507
rect 5478 2092 5556 2103
rect 14950 2092 15028 2103
rect 24422 2093 24500 2104
rect 33894 2093 33972 2104
rect 43366 2093 43444 2104
rect 52838 2093 52916 2104
rect 24422 2092 24844 2093
rect 5478 2091 5900 2092
rect 5478 2037 5490 2091
rect 5544 2037 5900 2091
rect 5478 2036 5900 2037
rect 14950 2091 15372 2092
rect 14950 2037 14962 2091
rect 15016 2037 15372 2091
rect 14950 2036 15372 2037
rect 24422 2038 24434 2092
rect 24488 2038 24844 2092
rect 24422 2037 24844 2038
rect 33894 2092 34316 2093
rect 33894 2038 33906 2092
rect 33960 2038 34316 2092
rect 33894 2037 34316 2038
rect 43366 2092 43788 2093
rect 43366 2038 43378 2092
rect 43432 2038 43788 2092
rect 43366 2037 43788 2038
rect 52838 2092 53260 2093
rect 52838 2038 52850 2092
rect 52904 2038 53260 2092
rect 52838 2037 53260 2038
rect 5478 2025 5556 2036
rect 14950 2025 15028 2036
rect 24422 2026 24500 2037
rect 33894 2026 33972 2037
rect 43366 2026 43444 2037
rect 52838 2026 52916 2037
rect 5529 1305 5615 1317
rect 15001 1305 15087 1317
rect 24473 1306 24559 1318
rect 33945 1306 34031 1318
rect 43417 1306 43503 1318
rect 52889 1306 52975 1318
rect 5529 1249 5541 1305
rect 5597 1249 5661 1305
rect 15001 1249 15013 1305
rect 15069 1249 15133 1305
rect 24473 1250 24485 1306
rect 24541 1250 24605 1306
rect 33945 1250 33957 1306
rect 34013 1250 34077 1306
rect 43417 1250 43429 1306
rect 43485 1250 43549 1306
rect 52889 1250 52901 1306
rect 52957 1250 53021 1306
rect 5529 1237 5615 1249
rect 15001 1237 15087 1249
rect 24473 1238 24559 1250
rect 33945 1238 34031 1250
rect 43417 1238 43503 1250
rect 52889 1238 52975 1250
rect 230 30 234 1150
rect 4814 230 4824 1030
rect 5124 230 5134 1030
rect 5324 30 9706 430
rect 14286 230 14296 1030
rect 14596 230 14606 1030
rect 14796 30 19178 430
rect 23758 231 23768 1031
rect 24068 231 24078 1031
rect 24268 31 28650 431
rect 33230 231 33240 1031
rect 33540 231 33550 1031
rect 33740 31 38122 431
rect 42702 231 42712 1031
rect 43012 231 43022 1031
rect 43212 31 47594 431
rect 52174 231 52184 1031
rect 52484 231 52494 1031
<< via1 >>
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 24588 8884 24644 8940
rect 34060 8884 34116 8940
rect 43532 8884 43588 8940
rect 53004 8884 53060 8940
rect 5444 5660 5500 5716
rect 14916 5660 14972 5716
rect 24388 5661 24444 5717
rect 33860 5661 33916 5717
rect 43332 5661 43388 5717
rect 52804 5661 52860 5717
rect 4824 3510 5124 4310
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 952 3290 1008 3346
rect 1166 2431 1246 2507
rect 5490 2037 5544 2091
rect 14962 2037 15016 2091
rect 24434 2038 24488 2092
rect 33906 2038 33960 2092
rect 43378 2038 43432 2092
rect 52850 2038 52904 2092
rect 5541 1249 5597 1305
rect 15013 1249 15069 1305
rect 24485 1250 24541 1306
rect 33957 1250 34013 1306
rect 43429 1250 43485 1306
rect 52901 1250 52957 1306
rect 4824 230 5124 1030
rect 14296 230 14596 1030
rect 23768 231 24068 1031
rect 33240 231 33540 1031
rect 42712 231 43012 1031
rect 52184 231 52484 1031
<< metal2 >>
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 56846 6619 56902 9891
rect 9056 6562 9542 6618
rect 18528 6562 19014 6618
rect 28000 6563 28486 6619
rect 37472 6563 37958 6619
rect 46944 6563 47430 6619
rect 56416 6563 56902 6619
rect 5430 5716 5512 5728
rect 5430 5660 5444 5716
rect 5500 5660 5512 5716
rect 5430 5648 5512 5660
rect 4814 4310 5134 4320
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 4814 3500 5134 3510
rect 940 3346 1020 3356
rect 940 3290 952 3346
rect 1008 3290 1020 3346
rect 9486 3290 9542 6562
rect 14902 5716 14984 5728
rect 14902 5660 14916 5716
rect 14972 5660 14984 5716
rect 14902 5648 14984 5660
rect 9896 4310 10116 4320
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 9896 3500 10116 3510
rect 14286 4310 14606 4320
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 14286 3500 14606 3510
rect 18958 3290 19014 6562
rect 24374 5717 24456 5729
rect 24374 5661 24388 5717
rect 24444 5661 24456 5717
rect 24374 5649 24456 5661
rect 19368 4311 19588 4321
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 19368 3501 19588 3511
rect 23758 4311 24078 4321
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 23758 3501 24078 3511
rect 28430 3291 28486 6563
rect 33846 5717 33928 5729
rect 33846 5661 33860 5717
rect 33916 5661 33928 5717
rect 33846 5649 33928 5661
rect 28840 4311 29060 4321
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 28840 3501 29060 3511
rect 33230 4311 33550 4321
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 33230 3501 33550 3511
rect 37902 3291 37958 6563
rect 43318 5717 43400 5729
rect 43318 5661 43332 5717
rect 43388 5661 43400 5717
rect 43318 5649 43400 5661
rect 38312 4311 38532 4321
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 38312 3501 38532 3511
rect 42702 4311 43022 4321
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 42702 3501 43022 3511
rect 47374 3291 47430 6563
rect 52790 5717 52872 5729
rect 52790 5661 52804 5717
rect 52860 5661 52872 5717
rect 52790 5649 52872 5661
rect 47784 4311 48004 4321
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 47784 3501 48004 3511
rect 52174 4311 52494 4321
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 52174 3501 52494 3511
rect 940 3280 1020 3290
rect 1156 2507 1256 2517
rect 1156 2431 1166 2507
rect 1246 2431 1256 2507
rect 1156 2421 1256 2431
rect 5478 2092 5556 2103
rect 14950 2092 15028 2103
rect 24422 2093 24500 2104
rect 33894 2093 33972 2104
rect 43366 2093 43444 2104
rect 52838 2093 52916 2104
rect 5368 2091 5556 2092
rect 5368 2037 5490 2091
rect 5544 2037 5556 2091
rect 5368 2036 5556 2037
rect 14840 2091 15028 2092
rect 14840 2037 14962 2091
rect 15016 2037 15028 2091
rect 24312 2092 24500 2093
rect 24312 2038 24434 2092
rect 24488 2038 24500 2092
rect 24312 2037 24500 2038
rect 33784 2092 33972 2093
rect 33784 2038 33906 2092
rect 33960 2038 33972 2092
rect 33784 2037 33972 2038
rect 43256 2092 43444 2093
rect 43256 2038 43378 2092
rect 43432 2038 43444 2092
rect 43256 2037 43444 2038
rect 52728 2092 52916 2093
rect 52728 2038 52850 2092
rect 52904 2038 52916 2092
rect 52728 2037 52916 2038
rect 14840 2036 15028 2037
rect 5478 2025 5556 2036
rect 14950 2025 15028 2036
rect 24422 2026 24500 2037
rect 33894 2026 33972 2037
rect 43366 2026 43444 2037
rect 52838 2026 52916 2037
rect -446 1792 122 1848
rect 9082 1793 9650 1849
rect 18554 1793 19122 1849
rect 28026 1794 28594 1850
rect 37498 1794 38066 1850
rect 46970 1794 47538 1850
rect -441 -51 -385 1792
rect 5529 1305 5615 1317
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 4814 1030 5134 1040
rect -441 -181 -385 -171
rect 10 -370 66 850
rect 4814 230 4824 1030
rect 5124 230 5134 1030
rect 4814 220 5134 230
rect 9087 -50 9143 1793
rect 15001 1305 15087 1317
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 14286 1030 14606 1040
rect 9087 -180 9143 -170
rect 9482 -370 9538 850
rect 14286 230 14296 1030
rect 14596 230 14606 1030
rect 14286 220 14606 230
rect 18559 -50 18615 1793
rect 24473 1306 24559 1318
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 23758 1031 24078 1041
rect 18559 -180 18615 -170
rect 18954 -370 19010 850
rect 23758 231 23768 1031
rect 24068 231 24078 1031
rect 23758 221 24078 231
rect 28031 -49 28087 1794
rect 33945 1306 34031 1318
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 33230 1031 33550 1041
rect 28031 -179 28087 -169
rect 28426 -369 28482 851
rect 33230 231 33240 1031
rect 33540 231 33550 1031
rect 33230 221 33550 231
rect 37503 -49 37559 1794
rect 43417 1306 43503 1318
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 42702 1031 43022 1041
rect 37503 -179 37559 -169
rect 37898 -369 37954 851
rect 42702 231 42712 1031
rect 43012 231 43022 1031
rect 42702 221 43022 231
rect 46975 -49 47031 1794
rect 52889 1306 52975 1318
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 52174 1031 52494 1041
rect 46975 -179 47031 -169
rect 47370 -369 47426 851
rect 52174 231 52184 1031
rect 52484 231 52494 1031
rect 52174 221 52494 231
<< via2 >>
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 24588 8884 24644 8940
rect 34060 8884 34116 8940
rect 43532 8884 43588 8940
rect 53004 8884 53060 8940
rect 5444 5660 5500 5716
rect 4824 3510 5124 4310
rect 952 3290 1008 3346
rect 14916 5660 14972 5716
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 24388 5661 24444 5717
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 33860 5661 33916 5717
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 43332 5661 43388 5717
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 52804 5661 52860 5717
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 1166 2431 1246 2507
rect 5541 1249 5597 1305
rect -441 -171 -385 -51
rect 4824 230 5124 1030
rect 15013 1249 15069 1305
rect 9087 -170 9143 -50
rect 14296 230 14596 1030
rect 24485 1250 24541 1306
rect 18559 -170 18615 -50
rect 23768 231 24068 1031
rect 33957 1250 34013 1306
rect 28031 -169 28087 -49
rect 33240 231 33540 1031
rect 43429 1250 43485 1306
rect 37503 -169 37559 -49
rect 42712 231 43012 1031
rect 52901 1250 52957 1306
rect 46975 -169 47031 -49
rect 52184 231 52484 1031
<< metal3 >>
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 5430 5716 5512 5728
rect 3058 5660 5444 5716
rect 5500 5709 5512 5716
rect 14902 5716 14984 5728
rect 14902 5709 14916 5716
rect 5500 5660 14916 5709
rect 14972 5709 14984 5716
rect 24374 5717 24456 5729
rect 24374 5709 24388 5717
rect 14972 5661 24388 5709
rect 24444 5709 24456 5717
rect 33846 5717 33928 5729
rect 33846 5709 33860 5717
rect 24444 5661 33860 5709
rect 33916 5709 33928 5717
rect 43318 5717 43400 5729
rect 43318 5709 43332 5717
rect 33916 5661 43332 5709
rect 43388 5709 43400 5717
rect 52790 5717 52872 5729
rect 52790 5709 52804 5717
rect 43388 5661 52804 5709
rect 52860 5661 52872 5717
rect 14972 5660 52872 5661
rect 3058 5655 52872 5660
rect 5430 5649 52872 5655
rect 5430 5648 52790 5649
rect 4814 4310 5134 4320
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 4814 3500 5134 3510
rect 9896 4310 10116 4320
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 9896 3500 10116 3510
rect 14286 4310 14606 4320
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 14286 3500 14606 3510
rect 19368 4311 19588 4321
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 19368 3501 19588 3511
rect 23758 4311 24078 4321
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 23758 3501 24078 3511
rect 28840 4311 29060 4321
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 28840 3501 29060 3511
rect 33230 4311 33550 4321
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 33230 3501 33550 3511
rect 38312 4311 38532 4321
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 38312 3501 38532 3511
rect 42702 4311 43022 4321
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 42702 3501 43022 3511
rect 47784 4311 48004 4321
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 47784 3501 48004 3511
rect 52174 4311 52494 4321
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 52174 3501 52494 3511
rect 940 3346 1020 3356
rect 940 3290 952 3346
rect 1008 3290 1020 3346
rect 940 2517 1020 3290
rect 940 2507 1256 2517
rect 940 2431 1166 2507
rect 1246 2431 1256 2507
rect 940 2421 1256 2431
rect 5529 1305 5615 1317
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 15001 1305 15087 1317
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 24473 1306 24559 1318
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 33945 1306 34031 1318
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 43417 1306 43503 1318
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 52889 1306 52975 1318
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 4814 1030 5134 1040
rect 4814 230 4824 1030
rect 5124 230 5134 1030
rect 4814 220 5134 230
rect 14286 1030 14606 1040
rect 14286 230 14296 1030
rect 14596 230 14606 1030
rect 14286 220 14606 230
rect 23758 1031 24078 1041
rect 23758 231 23768 1031
rect 24068 231 24078 1031
rect 23758 221 24078 231
rect 33230 1031 33550 1041
rect 33230 231 33240 1031
rect 33540 231 33550 1031
rect 33230 221 33550 231
rect 42702 1031 43022 1041
rect 42702 231 42712 1031
rect 43012 231 43022 1031
rect 42702 221 43022 231
rect 52174 1031 52494 1041
rect 52174 231 52184 1031
rect 52484 231 52494 1031
rect 52174 221 52494 231
rect 9077 -51 9087 -50
rect -689 -169 -441 -51
rect -451 -171 -441 -169
rect -385 -169 9087 -51
rect -385 -171 -375 -169
rect 9077 -170 9087 -169
rect 9143 -51 9153 -50
rect 18549 -51 18559 -50
rect 9143 -169 18559 -51
rect 9143 -170 9153 -169
rect 18549 -170 18559 -169
rect 18615 -51 18625 -50
rect 28021 -51 28031 -49
rect 18615 -169 28031 -51
rect 28087 -51 28097 -49
rect 37493 -51 37503 -49
rect 28087 -169 37503 -51
rect 37559 -51 37569 -49
rect 46965 -51 46975 -49
rect 37559 -169 46975 -51
rect 47031 -169 47041 -49
rect 18615 -170 18625 -169
<< via3 >>
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 24588 8884 24644 8940
rect 34060 8884 34116 8940
rect 43532 8884 43588 8940
rect 53004 8884 53060 8940
rect 4824 3510 5124 4310
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 5541 1249 5597 1305
rect 15013 1249 15069 1305
rect 24485 1250 24541 1306
rect 33957 1250 34013 1306
rect 43429 1250 43485 1306
rect 52901 1250 52957 1306
rect 4824 230 5124 1030
rect 14296 230 14596 1030
rect 23768 231 24068 1031
rect 33240 231 33540 1031
rect 42712 231 43012 1031
rect 52184 231 52484 1031
<< metal4 >>
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 4814 4310 5134 4320
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 4814 3500 5134 3510
rect 9896 4310 10116 4320
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 9896 3500 10116 3510
rect 14286 4310 14606 4320
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 14286 3500 14606 3510
rect 19368 4311 19588 4321
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 19368 3501 19588 3511
rect 23758 4311 24078 4321
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 23758 3501 24078 3511
rect 28840 4311 29060 4321
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 28840 3501 29060 3511
rect 33230 4311 33550 4321
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 33230 3501 33550 3511
rect 38312 4311 38532 4321
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 38312 3501 38532 3511
rect 42702 4311 43022 4321
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 42702 3501 43022 3511
rect 47784 4311 48004 4321
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 47784 3501 48004 3511
rect 52174 4311 52494 4321
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 52174 3501 52494 3511
rect 5529 1305 5615 1317
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 15001 1305 15087 1317
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 24473 1306 24559 1318
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 33945 1306 34031 1318
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 43417 1306 43503 1318
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 52889 1306 52975 1318
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 5782 1040 7078 1237
rect 15254 1040 16550 1237
rect 24726 1041 26022 1238
rect 34198 1041 35494 1238
rect 43670 1041 44966 1238
rect 53142 1041 54438 1238
rect 4814 1030 7078 1040
rect 4814 230 4824 1030
rect 5124 230 7078 1030
rect 4814 220 7078 230
rect 14286 1030 16550 1040
rect 14286 230 14296 1030
rect 14596 230 16550 1030
rect 14286 220 16550 230
rect 23758 1031 26022 1041
rect 23758 231 23768 1031
rect 24068 231 26022 1031
rect 23758 221 26022 231
rect 33230 1031 35494 1041
rect 33230 231 33240 1031
rect 33540 231 35494 1031
rect 33230 221 35494 231
rect 42702 1031 44966 1041
rect 42702 231 42712 1031
rect 43012 231 44966 1031
rect 42702 221 44966 231
rect 52174 1031 54438 1041
rect 52174 231 52184 1031
rect 52484 231 54438 1031
rect 52174 221 54438 231
<< via4 >>
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 24588 8884 24644 8940
rect 34060 8884 34116 8940
rect 43532 8884 43588 8940
rect 53004 8884 53060 8940
rect 4824 3510 5124 4310
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 5541 1249 5597 1305
rect 15013 1249 15069 1305
rect 24485 1250 24541 1306
rect 33957 1250 34013 1306
rect 43429 1250 43485 1306
rect 52901 1250 52957 1306
<< metal5 >>
rect 5630 8939 5782 9031
rect 5630 8883 5644 8939
rect 5700 8883 5782 8939
rect 5630 8871 5782 8883
rect 15102 8939 15254 9031
rect 15102 8883 15116 8939
rect 15172 8883 15254 8939
rect 15102 8871 15254 8883
rect 24574 8940 24726 9032
rect 24574 8884 24588 8940
rect 24644 8884 24726 8940
rect 24574 8872 24726 8884
rect 34046 8940 34198 9032
rect 34046 8884 34060 8940
rect 34116 8884 34198 8940
rect 34046 8872 34198 8884
rect 43518 8940 43670 9032
rect 43518 8884 43532 8940
rect 43588 8884 43670 8940
rect 43518 8872 43670 8884
rect 52990 8940 53142 9032
rect 52990 8884 53004 8940
rect 53060 8884 53142 8940
rect 52990 8872 53142 8884
rect 4814 4310 5782 4320
rect 4814 3510 4824 4310
rect 5124 3510 5782 4310
rect 4814 3500 5782 3510
rect 9082 4310 10116 4320
rect 9082 3510 9906 4310
rect 10106 3510 10116 4310
rect 9082 3500 10116 3510
rect 14286 4310 15254 4320
rect 14286 3510 14296 4310
rect 14596 3510 15254 4310
rect 14286 3500 15254 3510
rect 18554 4311 19588 4321
rect 18554 3511 19378 4311
rect 19578 3511 19588 4311
rect 18554 3501 19588 3511
rect 23758 4311 24726 4321
rect 23758 3511 23768 4311
rect 24068 3511 24726 4311
rect 23758 3501 24726 3511
rect 28026 4311 29060 4321
rect 28026 3511 28850 4311
rect 29050 3511 29060 4311
rect 28026 3501 29060 3511
rect 33230 4311 34198 4321
rect 33230 3511 33240 4311
rect 33540 3511 34198 4311
rect 33230 3501 34198 3511
rect 37498 4311 38532 4321
rect 37498 3511 38322 4311
rect 38522 3511 38532 4311
rect 37498 3501 38532 3511
rect 42702 4311 43670 4321
rect 42702 3511 42712 4311
rect 43012 3511 43670 4311
rect 42702 3501 43670 3511
rect 46970 4311 48004 4321
rect 46970 3511 47794 4311
rect 47994 3511 48004 4311
rect 46970 3501 48004 3511
rect 52174 4311 53142 4321
rect 52174 3511 52184 4311
rect 52484 3511 53142 4311
rect 52174 3501 53142 3511
rect 5529 1305 5783 1397
rect 5529 1249 5541 1305
rect 5597 1249 5783 1305
rect 5529 1237 5783 1249
rect 15001 1305 15255 1397
rect 15001 1249 15013 1305
rect 15069 1249 15255 1305
rect 15001 1237 15255 1249
rect 24473 1306 24727 1398
rect 24473 1250 24485 1306
rect 24541 1250 24727 1306
rect 24473 1238 24727 1250
rect 33945 1306 34199 1398
rect 33945 1250 33957 1306
rect 34013 1250 34199 1306
rect 33945 1238 34199 1250
rect 43417 1306 43671 1398
rect 43417 1250 43429 1306
rect 43485 1250 43671 1306
rect 43417 1238 43671 1250
rect 52889 1306 53143 1398
rect 52889 1250 52901 1306
rect 52957 1250 53143 1306
rect 52889 1238 53143 1250
use 2inmux  2inmux_0
timestamp 1758084968
transform 1 0 1034 0 1 2370
box -1024 -2340 4350 2140
use 2inmux  2inmux_1
timestamp 1758084968
transform 1 0 48394 0 1 2371
box -1024 -2340 4350 2140
use 2inmux  2inmux_2
timestamp 1758084968
transform 1 0 10506 0 1 2370
box -1024 -2340 4350 2140
use 2inmux  2inmux_3
timestamp 1758084968
transform 1 0 19978 0 1 2371
box -1024 -2340 4350 2140
use 2inmux  2inmux_4
timestamp 1758084968
transform 1 0 29450 0 1 2371
box -1024 -2340 4350 2140
use 2inmux  2inmux_5
timestamp 1758084968
transform 1 0 38922 0 1 2371
box -1024 -2340 4350 2140
use dffrs  dffrs_0
timestamp 1758085300
transform 1 0 6492 0 1 7135
box -848 -5898 2620 2881
use dffrs  dffrs_1
timestamp 1758085300
transform 1 0 15964 0 1 7135
box -848 -5898 2620 2881
use dffrs  dffrs_2
timestamp 1758085300
transform 1 0 25436 0 1 7136
box -848 -5898 2620 2881
use dffrs  dffrs_3
timestamp 1758085300
transform 1 0 34908 0 1 7136
box -848 -5898 2620 2881
use dffrs  dffrs_4
timestamp 1758085300
transform 1 0 44380 0 1 7136
box -848 -5898 2620 2881
use dffrs  dffrs_5
timestamp 1758085300
transform 1 0 53852 0 1 7136
box -848 -5898 2620 2881
<< labels >>
rlabel metal3 -689 -113 -689 -113 7 load
port 0 w
rlabel metal2 39 -370 39 -370 5 B6
port 1 s
rlabel metal2 9511 -370 9511 -370 5 B5
port 2 s
rlabel metal2 18983 -370 18983 -370 5 B4
port 3 s
rlabel metal2 56875 9891 56875 9891 1 serial_out
port 4 n
rlabel metal1 230 4493 230 4493 7 avdd
port 5 w
rlabel metal2 28455 -369 28455 -369 5 B3
port 6 s
rlabel metal1 230 54 230 54 7 avss
port 7 w
rlabel metal2 37927 -369 37927 -369 5 B2
port 8 s
rlabel metal2 47398 -369 47398 -369 5 B1
port 9 s
rlabel metal3 3058 5685 3058 5685 7 clk
port 10 w
<< end >>
