magic
tech gf180mcuD
magscale 1 5
timestamp 1755238359
<< checkpaint >>
rect -1030 230 1248 260
rect -1030 200 1496 230
rect -1030 170 1744 200
rect -1030 -2030 1992 170
rect -782 -2060 1992 -2030
rect -534 -2090 1992 -2060
rect -286 -2120 1992 -2090
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use nfet_03v3_5QDTWG  XM1
timestamp 0
transform 1 0 109 0 1 -885
box -139 -145 139 145
use nfet_03v3_5QDTWG  XM2
timestamp 0
transform 1 0 357 0 1 -915
box -139 -145 139 145
use pfet_03v3_YBHBCY  XM3
timestamp 0
transform 1 0 605 0 1 -945
box -139 -145 139 145
use pfet_03v3_YBHBCY  XM4
timestamp 0
transform 1 0 853 0 1 -975
box -139 -145 139 145
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 Vout1
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 Vout2
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 640 0 0 0 Vin1
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 640 0 0 0 Vin2
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 640 0 0 0 VSS
port 5 nsew
<< end >>
