** sch_path: /foss/designs/comparator/final_magic/nand2/osu_sc_nand2_1.sch
.subckt osu_sc_nand2_1 A B Y VDD VSS
*.PININFO A:I B:I Y:O VDD:I VSS:I
XM1 Y A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 Y B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM3 Y A net1 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM4 net1 B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends
.GLOBAL VDD
.GLOBAL VSS
