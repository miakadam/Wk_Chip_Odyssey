* NGSPICE file created from adc_PISO.ext - technology: (null)

.subckt adc_PISO load B6 B5 B4 serial_out avdd B3 avss B2 B1 clk
X0 a_44488_8266 avdd.t378 avss.t100 avss.t99 nfet_03v3
**devattr s=17600,576 d=10400,304
X1 a_50206_2781 a_48650_3501.t4 avdd.t337 avdd.t336 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X2 a_6600_2510.t2 a_6520_1558.t4 avdd.t51 avdd.t50 pfet_03v3
**devattr s=44000,1176 d=26000,604
X3 a_6520_1558.t2 a_6520_3763.t4 avdd.t329 avdd.t328 pfet_03v3
**devattr s=44000,1176 d=26000,604
X4 avdd.t43 dffrs_1.Q.t4 a_20234_3501.t1 avdd.t42 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X5 avdd.t331 a_6520_3763.t5 2inmux_2.Bit.t2 avdd.t330 pfet_03v3
**devattr s=26000,604 d=26000,604
X6 a_2846_2780 a_1290_3500.t4 avdd.t189 avdd.t188 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X7 dffrs_4.Qb avdd.t379 a_46158_3857 avss.t98 nfet_03v3
**devattr s=10400,304 d=17600,576
X8 a_15992_3763.t1 clk.t0 a_16256_6060 avss.t22 nfet_03v3
**devattr s=10400,304 d=17600,576
X9 2inmux_1.Bit.t2 dffrs_4.Qb a_46158_6061 avss.t255 nfet_03v3
**devattr s=10400,304 d=17600,576
X10 a_10950_2780 2inmux_2.Bit.t4 avss.t262 avss.t261 nfet_03v3
**devattr s=17600,576 d=10400,304
X11 a_15992_5968.t0 a_15992_3763.t4 a_16256_8265 avss.t225 nfet_03v3
**devattr s=10400,304 d=17600,576
X12 a_39178_3501.t1 load.t0 avdd.t169 avdd.t168 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X13 avss.t45 dffrs_2.Q.t4 a_29894_2781 avss.t44 nfet_03v3
**devattr s=10400,304 d=17600,576
X14 a_50206_441 a_48650_1161.t4 avss.t218 avss.t217 nfet_03v3
**devattr s=17600,576 d=17600,576
X15 2inmux_1.OUT.t1 a_50878_1605.t4 avss.t285 avss.t284 nfet_03v3
**devattr s=17600,576 d=17600,576
X16 avdd.t53 a_6520_1558.t5 dffrs_0.Qb avdd.t52 pfet_03v3
**devattr s=26000,604 d=26000,604
X17 avss.t189 a_21790_2781 a_22462_1605.t0 avss.t188 nfet_03v3
**devattr s=17600,576 d=17600,576
X18 a_35016_1651 a_34936_1559.t4 avss.t142 avss.t141 nfet_03v3
**devattr s=17600,576 d=10400,304
X19 a_35016_3856 a_34936_3764.t4 avss.t268 avss.t267 nfet_03v3
**devattr s=17600,576 d=10400,304
X20 2inmux_0.OUT.t1 a_3518_1604.t4 avss.t283 avss.t282 nfet_03v3
**devattr s=17600,576 d=17600,576
X21 a_22462_1605.t2 a_21790_441 a_22650_2325 avdd.t373 pfet_03v3
**devattr s=31200,704 d=52800,1376
X22 a_29000_1361 load.t1 avdd.t69 avdd.t68 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X23 avss.t266 a_47944_1361 a_48838_441 avss.t265 nfet_03v3
**devattr s=10400,304 d=17600,576
X24 avdd.t165 avdd.t163 a_44408_3764.t2 avdd.t164 pfet_03v3
**devattr s=26000,604 d=26000,604
X25 a_21790_441 a_20234_1161.t4 avdd.t237 avdd.t236 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X26 a_1478_2780 load.t2 a_1290_3500.t0 avss.t54 nfet_03v3
**devattr s=17600,576 d=10400,304
X27 avdd.t17 a_29000_1361 a_29706_1161.t0 avdd.t16 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X28 a_25464_3764.t0 clk.t1 avdd.t27 avdd.t26 pfet_03v3
**devattr s=26000,604 d=44000,1176
X29 avdd.t162 avdd.t160 a_6600_2510.t0 avdd.t161 pfet_03v3
**devattr s=26000,604 d=26000,604
X30 a_1478_440 B6.t0 a_1290_1160.t3 avss.t181 nfet_03v3
**devattr s=17600,576 d=10400,304
X31 avdd.t321 a_25464_3764.t4 dffrs_2.Q.t3 avdd.t320 pfet_03v3
**devattr s=26000,604 d=26000,604
X32 a_35200_6061 avdd.t380 a_35016_6061 avss.t97 nfet_03v3
**devattr s=10400,304 d=10400,304
X33 avdd.t357 2inmux_2.Bit.t5 a_10762_3500.t3 avdd.t356 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X34 a_1290_1160.t1 B6.t1 avdd.t75 avdd.t74 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X35 2inmux_2.Bit.t1 dffrs_0.Qb avdd.t13 avdd.t12 pfet_03v3
**devattr s=26000,604 d=44000,1176
X36 avdd.t343 clk.t2 a_6520_1558.t3 avdd.t342 pfet_03v3
**devattr s=26000,604 d=26000,604
X37 a_35200_8266 a_35016_2511.t4 a_35016_8266 avss.t208 nfet_03v3
**devattr s=10400,304 d=10400,304
X38 avss.t180 2inmux_1.Bit.t4 a_48838_2781 avss.t179 nfet_03v3
**devattr s=10400,304 d=17600,576
X39 avss.t24 a_40734_2781 a_41406_1605.t0 avss.t23 nfet_03v3
**devattr s=17600,576 d=17600,576
X40 avdd.t289 a_44488_2511.t4 a_44408_5969.t3 avdd.t288 pfet_03v3
**devattr s=26000,604 d=26000,604
X41 avdd.t363 a_25464_1559.t4 dffrs_2.Qb avdd.t362 pfet_03v3
**devattr s=26000,604 d=26000,604
X42 a_31262_2781 a_29706_3501.t4 avss.t131 avss.t130 nfet_03v3
**devattr s=17600,576 d=17600,576
X43 a_47944_1361 load.t3 avdd.t71 avdd.t70 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X44 a_39366_2781 dffrs_3.Q.t4 avss.t196 avss.t195 nfet_03v3
**devattr s=17600,576 d=10400,304
X45 dffrs_0.Qb avdd.t157 avdd.t159 avdd.t158 pfet_03v3
**devattr s=26000,604 d=44000,1176
X46 avdd.t49 a_584_1360 a_1290_1160.t0 avdd.t48 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X47 2inmux_3.OUT.t1 a_22462_1605.t4 avss.t102 avss.t101 nfet_03v3
**devattr s=17600,576 d=17600,576
X48 a_51066_2325 a_50206_441 a_50878_1605.t2 avdd.t317 pfet_03v3
**devattr s=52800,1376 d=31200,704
X49 a_12990_1604.t2 a_12318_440 a_13178_2324 avdd.t1 pfet_03v3
**devattr s=31200,704 d=52800,1376
X50 a_25464_5969.t3 a_25464_3764.t5 avdd.t323 avdd.t322 pfet_03v3
**devattr s=26000,604 d=44000,1176
X51 a_44488_2511.t3 a_44408_1559.t4 avdd.t281 avdd.t280 pfet_03v3
**devattr s=44000,1176 d=26000,604
X52 avdd.t156 avdd.t154 a_15992_3763.t2 avdd.t155 pfet_03v3
**devattr s=26000,604 d=26000,604
X53 a_44408_3764.t0 clk.t3 avdd.t345 avdd.t344 pfet_03v3
**devattr s=26000,604 d=44000,1176
X54 a_44408_1559.t0 a_44408_3764.t4 avdd.t193 avdd.t192 pfet_03v3
**devattr s=44000,1176 d=26000,604
X55 a_20422_2781 load.t4 a_20234_3501.t2 avss.t123 nfet_03v3
**devattr s=17600,576 d=10400,304
X56 avdd.t195 a_44408_3764.t5 2inmux_1.Bit.t1 avdd.t194 pfet_03v3
**devattr s=26000,604 d=26000,604
X57 a_54144_6061 avdd.t381 a_53960_6061 avss.t96 nfet_03v3
**devattr s=10400,304 d=10400,304
X58 a_55630_3857 a_53880_1559.t4 a_55446_3857 avss.t147 nfet_03v3
**devattr s=10400,304 d=10400,304
X59 a_54144_8266 a_53960_2511.t4 a_53960_8266 avss.t166 nfet_03v3
**devattr s=10400,304 d=10400,304
X60 avdd.t263 a_15992_3763.t5 dffrs_1.Q.t3 avdd.t262 pfet_03v3
**devattr s=26000,604 d=26000,604
X61 a_25544_6061 a_25464_5969.t4 avss.t161 avss.t160 nfet_03v3
**devattr s=17600,576 d=10400,304
X62 a_27030_3857 dffrs_2.Q.t5 avss.t220 avss.t219 nfet_03v3
**devattr s=17600,576 d=10400,304
X63 a_25544_8266 avdd.t382 avss.t95 avss.t94 nfet_03v3
**devattr s=17600,576 d=10400,304
X64 dffrs_2.Q.t1 dffrs_2.Qb avdd.t15 avdd.t14 pfet_03v3
**devattr s=26000,604 d=44000,1176
X65 a_55630_6061 a_53880_3764.t4 a_55446_6061 avss.t143 nfet_03v3
**devattr s=10400,304 d=10400,304
X66 a_3518_1604.t0 a_2846_440 avss.t7 avss.t6 nfet_03v3
**devattr s=17600,576 d=17600,576
X67 a_27030_6061 avdd.t383 avss.t93 avss.t92 nfet_03v3
**devattr s=17600,576 d=10400,304
X68 a_34936_3764.t1 clk.t4 a_35200_6061 avss.t245 nfet_03v3
**devattr s=10400,304 d=17600,576
X69 a_31262_2781 a_29706_3501.t5 avdd.t201 avdd.t200 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X70 avdd.t277 dffrs_3.Q.t5 a_39178_3501.t0 avdd.t276 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X71 a_16072_2510.t1 2inmux_2.OUT.t2 avdd.t249 avdd.t248 pfet_03v3
**devattr s=26000,604 d=44000,1176
X72 a_34936_5969.t2 a_34936_3764.t5 a_35200_8266 avss.t269 nfet_03v3
**devattr s=10400,304 d=17600,576
X73 avdd.t283 a_44408_1559.t5 dffrs_4.Qb avdd.t282 pfet_03v3
**devattr s=26000,604 d=26000,604
X74 a_15992_1558.t1 a_16072_2510.t4 avdd.t241 avdd.t240 pfet_03v3
**devattr s=26000,604 d=44000,1176
X75 a_39366_441 a_38472_1361 avss.t30 avss.t29 nfet_03v3
**devattr s=17600,576 d=10400,304
X76 a_21790_441 a_20234_1161.t5 avss.t151 avss.t150 nfet_03v3
**devattr s=17600,576 d=17600,576
X77 a_1290_1160.t2 B6.t2 a_1478_440 avss.t252 nfet_03v3
**devattr s=10400,304 d=17600,576
X78 a_44408_5969.t0 a_44408_3764.t6 avdd.t197 avdd.t196 pfet_03v3
**devattr s=26000,604 d=44000,1176
X79 avdd.t285 a_15992_1558.t4 dffrs_1.Qb avdd.t284 pfet_03v3
**devattr s=26000,604 d=26000,604
X80 dffrs_2.Qb avdd.t151 avdd.t153 avdd.t152 pfet_03v3
**devattr s=26000,604 d=44000,1176
X81 avss.t26 a_12318_2780 a_12990_1604.t3 avss.t25 nfet_03v3
**devattr s=17600,576 d=17600,576
X82 avdd.t243 a_16072_2510.t5 a_15992_5968.t3 avdd.t242 pfet_03v3
**devattr s=26000,604 d=26000,604
X83 a_53880_3764.t3 a_53880_5969.t4 avdd.t293 avdd.t292 pfet_03v3
**devattr s=44000,1176 d=26000,604
X84 a_2846_440 a_1290_1160.t4 avss.t135 avss.t134 nfet_03v3
**devattr s=17600,576 d=17600,576
X85 a_44672_1651 avdd.t384 a_44488_1651 avss.t91 nfet_03v3
**devattr s=10400,304 d=10400,304
X86 2inmux_4.OUT.t1 a_31934_1605.t4 avss.t201 avss.t200 nfet_03v3
**devattr s=17600,576 d=17600,576
X87 a_44672_3856 clk.t5 a_44488_3856 avss.t249 nfet_03v3
**devattr s=10400,304 d=10400,304
X88 dffrs_3.Q.t3 avdd.t148 avdd.t150 avdd.t149 pfet_03v3
**devattr s=44000,1176 d=26000,604
X89 a_45974_3857 2inmux_1.Bit.t5 avss.t117 avss.t116 nfet_03v3
**devattr s=17600,576 d=10400,304
X90 a_10950_2780 load.t5 a_10762_3500.t2 avss.t124 nfet_03v3
**devattr s=17600,576 d=10400,304
X91 a_25544_2511.t2 2inmux_3.OUT.t2 a_25728_1651 avss.t279 nfet_03v3
**devattr s=10400,304 d=17600,576
X92 a_1478_440 a_584_1360 avss.t38 avss.t37 nfet_03v3
**devattr s=17600,576 d=10400,304
X93 a_16072_6060 a_15992_5968.t4 avss.t271 avss.t270 nfet_03v3
**devattr s=17600,576 d=10400,304
X94 a_25464_1559.t1 a_25544_2511.t4 a_25728_3856 avss.t41 nfet_03v3
**devattr s=10400,304 d=17600,576
X95 a_25728_6061 avdd.t385 a_25544_6061 avss.t90 nfet_03v3
**devattr s=10400,304 d=10400,304
X96 a_45974_6061 avdd.t386 avss.t89 avss.t88 nfet_03v3
**devattr s=17600,576 d=10400,304
X97 a_53880_3764.t0 clk.t6 a_54144_6061 avss.t250 nfet_03v3
**devattr s=10400,304 d=17600,576
X98 dffrs_5.Qb avdd.t387 a_55630_3857 avss.t87 nfet_03v3
**devattr s=10400,304 d=17600,576
X99 a_10762_1160.t0 B5.t0 avdd.t219 avdd.t218 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X100 a_19528_1361 load.t6 avss.t127 avss.t126 nfet_03v3
**devattr s=17600,576 d=17600,576
X101 a_39366_2781 load.t7 a_39178_3501.t3 avss.t128 nfet_03v3
**devattr s=17600,576 d=10400,304
X102 avdd.t147 avdd.t145 a_35016_2511.t1 avdd.t146 pfet_03v3
**devattr s=26000,604 d=26000,604
X103 a_16072_8265 avdd.t388 avss.t86 avss.t85 nfet_03v3
**devattr s=17600,576 d=10400,304
X104 a_25728_8266 a_25544_2511.t5 a_25544_8266 avss.t42 nfet_03v3
**devattr s=10400,304 d=10400,304
X105 a_53880_5969.t2 a_53880_3764.t5 a_54144_8266 avss.t144 nfet_03v3
**devattr s=10400,304 d=17600,576
X106 dffrs_1.Q.t1 dffrs_1.Qb avdd.t199 avdd.t198 pfet_03v3
**devattr s=26000,604 d=44000,1176
X107 a_6520_3763.t3 clk.t7 a_6784_6060 avss.t251 nfet_03v3
**devattr s=10400,304 d=17600,576
X108 avdd.t7 clk.t8 a_34936_1559.t0 avdd.t6 pfet_03v3
**devattr s=26000,604 d=26000,604
X109 avdd.t35 a_12318_2780 a_13178_2324 avdd.t34 pfet_03v3
**devattr s=31200,704 d=52800,1376
X110 a_22462_1605.t3 a_21790_441 avss.t287 avss.t286 nfet_03v3
**devattr s=17600,576 d=17600,576
X111 a_53880_5969.t0 avdd.t142 avdd.t144 avdd.t143 pfet_03v3
**devattr s=44000,1176 d=26000,604
X112 a_6520_5968.t2 a_6520_3763.t6 a_6784_8265 avss.t238 nfet_03v3
**devattr s=10400,304 d=17600,576
X113 serial_out.t3 dffrs_5.Qb a_55630_6061 avss.t242 nfet_03v3
**devattr s=10400,304 d=17600,576
X114 dffrs_3.Qb dffrs_3.Q.t6 avdd.t279 avdd.t278 pfet_03v3
**devattr s=44000,1176 d=26000,604
X115 avss.t28 a_38472_1361 a_39366_441 avss.t27 nfet_03v3
**devattr s=10400,304 d=17600,576
X116 a_39366_441 B2.t0 a_39178_1161.t2 avss.t120 nfet_03v3
**devattr s=17600,576 d=10400,304
X117 dffrs_1.Qb avdd.t139 avdd.t141 avdd.t140 pfet_03v3
**devattr s=26000,604 d=44000,1176
X118 serial_out.t0 avdd.t136 avdd.t138 avdd.t137 pfet_03v3
**devattr s=44000,1176 d=26000,604
X119 a_16256_1650 avdd.t389 a_16072_1650 avss.t84 nfet_03v3
**devattr s=10400,304 d=10400,304
X120 a_44488_2511.t1 2inmux_5.OUT.t2 a_44672_1651 avss.t168 nfet_03v3
**devattr s=10400,304 d=17600,576
X121 a_6520_3763.t1 a_6520_5968.t4 avdd.t187 avdd.t186 pfet_03v3
**devattr s=44000,1176 d=26000,604
X122 a_16256_3855 clk.t9 a_16072_3855 avss.t5 nfet_03v3
**devattr s=10400,304 d=10400,304
X123 a_44408_1559.t2 a_44488_2511.t5 a_44672_3856 avss.t173 nfet_03v3
**devattr s=10400,304 d=17600,576
X124 avss.t36 a_584_1360 a_1478_440 avss.t35 nfet_03v3
**devattr s=10400,304 d=17600,576
X125 a_17558_3856 dffrs_1.Q.t5 avss.t15 avss.t14 nfet_03v3
**devattr s=17600,576 d=10400,304
X126 avdd.t135 avdd.t133 a_53960_2511.t1 avdd.t134 pfet_03v3
**devattr s=26000,604 d=26000,604
X127 a_48650_3501.t1 load.t8 a_48838_2781 avss.t136 nfet_03v3
**devattr s=10400,304 d=17600,576
X128 a_41406_1605.t3 a_40734_441 avss.t47 avss.t46 nfet_03v3
**devattr s=17600,576 d=17600,576
X129 avdd.t361 a_34936_3764.t6 dffrs_3.Q.t0 avdd.t360 pfet_03v3
**devattr s=26000,604 d=26000,604
X130 avdd.t9 clk.t10 a_53880_1559.t0 avdd.t8 pfet_03v3
**devattr s=26000,604 d=26000,604
X131 a_25544_2511.t0 a_25464_1559.t5 avdd.t365 avdd.t364 pfet_03v3
**devattr s=44000,1176 d=26000,604
X132 a_25464_1559.t3 a_25464_3764.t6 avdd.t325 avdd.t324 pfet_03v3
**devattr s=44000,1176 d=26000,604
X133 dffrs_5.Qb serial_out.t4 avdd.t177 avdd.t176 pfet_03v3
**devattr s=44000,1176 d=26000,604
X134 a_12990_1604.t0 a_12318_440 avss.t3 avss.t2 nfet_03v3
**devattr s=17600,576 d=17600,576
X135 2inmux_1.OUT.t0 a_50878_1605.t5 avdd.t215 avdd.t214 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X136 a_17558_6060 avdd.t390 avss.t83 avss.t82 nfet_03v3
**devattr s=17600,576 d=10400,304
X137 avss.t216 avss.t214 a_1478_2780 avss.t215 nfet_03v3
**devattr s=10400,304 d=17600,576
X138 a_22650_2325 a_21790_2781 avdd.t275 avdd.t274 pfet_03v3
**devattr s=52800,1376 d=31200,704
X139 a_35016_2511.t2 2inmux_4.OUT.t2 avdd.t297 avdd.t296 pfet_03v3
**devattr s=26000,604 d=44000,1176
X140 a_34936_1559.t3 a_35016_2511.t5 avdd.t301 avdd.t300 pfet_03v3
**devattr s=26000,604 d=44000,1176
X141 2inmux_0.OUT.t0 a_3518_1604.t5 avdd.t235 avdd.t234 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X142 avss.t115 a_50206_2781 a_50878_1605.t0 avss.t114 nfet_03v3
**devattr s=17600,576 d=17600,576
X143 a_40734_2781 a_39178_3501.t4 avss.t260 avss.t259 nfet_03v3
**devattr s=17600,576 d=17600,576
X144 avdd.t225 a_34936_1559.t5 dffrs_3.Qb avdd.t224 pfet_03v3
**devattr s=26000,604 d=26000,604
X145 a_20422_441 B4.t0 a_20234_1161.t0 avss.t43 nfet_03v3
**devattr s=17600,576 d=10400,304
X146 a_48838_2781 2inmux_1.Bit.t6 avss.t119 avss.t118 nfet_03v3
**devattr s=17600,576 d=10400,304
X147 a_6520_5968.t3 avdd.t130 avdd.t132 avdd.t131 pfet_03v3
**devattr s=44000,1176 d=26000,604
X148 a_53960_1651 a_53880_1559.t5 avss.t149 avss.t148 nfet_03v3
**devattr s=17600,576 d=10400,304
X149 a_53960_3856 a_53880_3764.t6 avss.t146 avss.t145 nfet_03v3
**devattr s=17600,576 d=10400,304
X150 a_12318_440 a_10762_1160.t4 avss.t140 avss.t139 nfet_03v3
**devattr s=17600,576 d=17600,576
X151 a_41406_1605.t2 a_40734_441 a_41594_2325 avdd.t59 pfet_03v3
**devattr s=31200,704 d=52800,1376
X152 a_48650_3501.t2 load.t9 avdd.t213 avdd.t212 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X153 a_29706_3501.t2 load.t10 a_29894_2781 avss.t104 nfet_03v3
**devattr s=10400,304 d=17600,576
X154 avdd.t129 avdd.t127 a_6520_3763.t0 avdd.t128 pfet_03v3
**devattr s=26000,604 d=26000,604
X155 a_35016_6061 a_34936_5969.t4 avss.t172 avss.t171 nfet_03v3
**devattr s=17600,576 d=10400,304
X156 2inmux_2.Bit.t3 avdd.t124 avdd.t126 avdd.t125 pfet_03v3
**devattr s=44000,1176 d=26000,604
X157 a_16072_2510.t3 a_15992_1558.t5 avdd.t287 avdd.t286 pfet_03v3
**devattr s=44000,1176 d=26000,604
X158 a_10056_1360 load.t11 avss.t106 avss.t105 nfet_03v3
**devattr s=17600,576 d=17600,576
X159 a_53960_2511.t3 2inmux_1.OUT.t2 avdd.t309 avdd.t308 pfet_03v3
**devattr s=26000,604 d=44000,1176
X160 a_35016_8266 avdd.t391 avss.t81 avss.t80 nfet_03v3
**devattr s=17600,576 d=10400,304
X161 a_15992_1558.t3 a_15992_3763.t6 avdd.t265 avdd.t264 pfet_03v3
**devattr s=44000,1176 d=26000,604
X162 a_40734_2781 a_39178_3501.t5 avdd.t355 avdd.t354 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X163 avdd.t123 avdd.t121 a_25544_2511.t3 avdd.t122 pfet_03v3
**devattr s=26000,604 d=26000,604
X164 a_41594_2325 a_40734_2781 avdd.t31 avdd.t30 pfet_03v3
**devattr s=52800,1376 d=31200,704
X165 avdd.t205 a_31262_2781 a_32122_2325 avdd.t204 pfet_03v3
**devattr s=31200,704 d=52800,1376
X166 avdd.t23 clk.t11 a_25464_1559.t0 avdd.t22 pfet_03v3
**devattr s=26000,604 d=26000,604
X167 a_53880_1559.t2 a_53960_2511.t5 avdd.t251 avdd.t250 pfet_03v3
**devattr s=26000,604 d=44000,1176
X168 avdd.t185 2inmux_1.Bit.t7 a_48650_3501.t0 avdd.t184 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X169 a_6600_2510.t3 2inmux_0.OUT.t2 avdd.t371 avdd.t370 pfet_03v3
**devattr s=26000,604 d=44000,1176
X170 a_584_1360 load.t12 avss.t183 avss.t182 nfet_03v3
**devattr s=17600,576 d=17600,576
X171 a_6520_1558.t0 a_6600_2510.t4 avdd.t5 avdd.t4 pfet_03v3
**devattr s=26000,604 d=44000,1176
X172 dffrs_3.Qb avdd.t392 a_36686_3857 avss.t79 nfet_03v3
**devattr s=10400,304 d=17600,576
X173 avss.t17 dffrs_1.Q.t6 a_20422_2781 avss.t16 nfet_03v3
**devattr s=10400,304 d=17600,576
X174 2inmux_3.OUT.t0 a_22462_1605.t5 avdd.t167 avdd.t166 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X175 a_20234_1161.t2 B4.t1 avdd.t221 avdd.t220 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X176 dffrs_0.Qb 2inmux_2.Bit.t6 avdd.t369 avdd.t368 pfet_03v3
**devattr s=44000,1176 d=26000,604
X177 a_20234_1161.t3 B4.t2 a_20422_441 avss.t138 nfet_03v3
**devattr s=10400,304 d=17600,576
X178 dffrs_3.Q.t1 dffrs_3.Qb a_36686_6061 avss.t48 nfet_03v3
**devattr s=10400,304 d=17600,576
X179 a_12318_2780 a_10762_3500.t4 avss.t203 avss.t202 nfet_03v3
**devattr s=17600,576 d=17600,576
X180 avdd.t21 a_6600_2510.t5 a_6520_5968.t0 avdd.t20 pfet_03v3
**devattr s=26000,604 d=26000,604
X181 a_29706_3501.t3 load.t13 avdd.t269 avdd.t268 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X182 avss.t289 a_2846_2780 a_3518_1604.t3 avss.t288 nfet_03v3
**devattr s=17600,576 d=17600,576
X183 2inmux_5.OUT.t1 a_41406_1605.t4 avss.t154 avss.t153 nfet_03v3
**devattr s=17600,576 d=17600,576
X184 a_44408_3764.t3 a_44408_5969.t4 avdd.t319 avdd.t318 pfet_03v3
**devattr s=44000,1176 d=26000,604
X185 a_6600_1650 a_6520_1558.t6 avss.t40 avss.t39 nfet_03v3
**devattr s=17600,576 d=10400,304
X186 a_50206_441 a_48650_1161.t5 avdd.t259 avdd.t258 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X187 a_2846_440 a_1290_1160.t5 avdd.t211 avdd.t210 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X188 avdd.t67 a_19528_1361 a_20234_1161.t1 avdd.t66 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X189 a_6600_3855 a_6520_3763.t7 avss.t240 avss.t239 nfet_03v3
**devattr s=17600,576 d=10400,304
X190 a_3706_2324 a_2846_440 a_3518_1604.t2 avdd.t11 pfet_03v3
**devattr s=52800,1376 d=31200,704
X191 avss.t235 a_10056_1360 a_10950_440 avss.t234 nfet_03v3
**devattr s=10400,304 d=17600,576
X192 a_39178_1161.t1 B2.t1 a_39366_441 avss.t165 nfet_03v3
**devattr s=10400,304 d=17600,576
X193 a_20422_441 a_19528_1361 avss.t53 avss.t52 nfet_03v3
**devattr s=17600,576 d=10400,304
X194 a_10950_440 B5.t1 a_10762_1160.t2 avss.t274 nfet_03v3
**devattr s=17600,576 d=10400,304
X195 a_31934_1605.t3 a_31262_441 avss.t224 avss.t223 nfet_03v3
**devattr s=17600,576 d=17600,576
X196 a_15992_3763.t0 clk.t12 avdd.t25 avdd.t24 pfet_03v3
**devattr s=26000,604 d=44000,1176
X197 2inmux_1.Bit.t3 dffrs_4.Qb avdd.t353 avdd.t352 pfet_03v3
**devattr s=26000,604 d=44000,1176
X198 avdd.t377 a_2846_2780 a_3706_2324 avdd.t376 pfet_03v3
**devattr s=31200,704 d=52800,1376
X199 a_40734_441 a_39178_1161.t4 avss.t170 avss.t169 nfet_03v3
**devattr s=17600,576 d=17600,576
X200 a_39178_1161.t3 B2.t2 avdd.t233 avdd.t232 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X201 a_8270_3856 a_6520_1558.t7 a_8086_3856 avss.t20 nfet_03v3
**devattr s=10400,304 d=10400,304
X202 a_12318_2780 a_10762_3500.t5 avdd.t307 avdd.t306 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X203 a_13178_2324 a_12318_2780 avdd.t33 avdd.t32 pfet_03v3
**devattr s=52800,1376 d=31200,704
X204 a_44408_5969.t2 avdd.t118 avdd.t120 avdd.t119 pfet_03v3
**devattr s=44000,1176 d=26000,604
X205 a_8270_6060 a_6520_3763.t8 a_8086_6060 avss.t241 nfet_03v3
**devattr s=10400,304 d=10400,304
X206 2inmux_4.OUT.t0 a_31934_1605.t5 avdd.t295 avdd.t294 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X207 dffrs_4.Qb avdd.t115 avdd.t117 avdd.t116 pfet_03v3
**devattr s=26000,604 d=44000,1176
X208 a_21790_2781 a_20234_3501.t4 avss.t113 avss.t112 nfet_03v3
**devattr s=17600,576 d=17600,576
X209 a_29894_2781 dffrs_2.Q.t6 avss.t222 avss.t221 nfet_03v3
**devattr s=17600,576 d=10400,304
X210 avdd.t327 a_10056_1360 a_10762_1160.t3 avdd.t326 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X211 2inmux_2.OUT.t1 a_12990_1604.t4 avss.t273 avss.t272 nfet_03v3
**devattr s=17600,576 d=17600,576
X212 a_31934_1605.t2 a_31262_441 a_32122_2325 avdd.t315 pfet_03v3
**devattr s=31200,704 d=52800,1376
X213 a_15992_5968.t1 a_15992_3763.t7 avdd.t267 avdd.t266 pfet_03v3
**devattr s=26000,604 d=44000,1176
X214 a_6784_1650 avdd.t393 a_6600_1650 avss.t78 nfet_03v3
**devattr s=10400,304 d=10400,304
X215 a_19528_1361 load.t14 avdd.t171 avdd.t170 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X216 a_22650_2325 a_21790_441 a_22462_1605.t1 avdd.t372 pfet_03v3
**devattr s=52800,1376 d=31200,704
X217 a_6784_3855 clk.t13 a_6600_3855 avss.t21 nfet_03v3
**devattr s=10400,304 d=10400,304
X218 a_1290_3500.t1 load.t15 a_1478_2780 avss.t103 nfet_03v3
**devattr s=10400,304 d=17600,576
X219 a_35016_2511.t0 a_34936_1559.t6 avdd.t217 avdd.t216 pfet_03v3
**devattr s=44000,1176 d=26000,604
X220 avdd.t114 avdd.t112 a_34936_3764.t2 avdd.t113 pfet_03v3
**devattr s=26000,604 d=26000,604
X221 a_34936_1559.t1 a_34936_3764.t7 avdd.t63 avdd.t62 pfet_03v3
**devattr s=44000,1176 d=26000,604
X222 a_44672_6061 avdd.t394 a_44488_6061 avss.t77 nfet_03v3
**devattr s=10400,304 d=10400,304
X223 a_38472_1361 load.t16 avss.t109 avss.t108 nfet_03v3
**devattr s=17600,576 d=17600,576
X224 a_44672_8266 a_44488_2511.t6 a_44488_8266 avss.t174 nfet_03v3
**devattr s=10400,304 d=10400,304
X225 dffrs_0.Qb avdd.t395 a_8270_3856 avss.t76 nfet_03v3
**devattr s=10400,304 d=17600,576
X226 a_27214_3857 a_25464_1559.t6 a_27030_3857 avss.t56 nfet_03v3
**devattr s=10400,304 d=10400,304
X227 a_1478_2780 avss.t211 avss.t213 avss.t212 nfet_03v3
**devattr s=17600,576 d=10400,304
X228 avss.t51 a_19528_1361 a_20422_441 avss.t50 nfet_03v3
**devattr s=10400,304 d=17600,576
X229 a_25464_3764.t1 clk.t14 a_25728_6061 avss.t247 nfet_03v3
**devattr s=10400,304 d=17600,576
X230 a_21790_2781 a_20234_3501.t5 avdd.t261 avdd.t260 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X231 avdd.t313 dffrs_2.Q.t7 a_29706_3501.t0 avdd.t312 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X232 a_25464_5969.t2 a_25464_3764.t7 a_25728_8266 avss.t204 nfet_03v3
**devattr s=10400,304 d=17600,576
X233 a_27214_6061 a_25464_3764.t8 a_27030_6061 avss.t205 nfet_03v3
**devattr s=10400,304 d=10400,304
X234 a_10762_1160.t1 B5.t2 a_10950_440 avss.t209 nfet_03v3
**devattr s=10400,304 d=17600,576
X235 a_10950_440 a_10056_1360 avss.t233 avss.t232 nfet_03v3
**devattr s=17600,576 d=10400,304
X236 2inmux_2.Bit.t0 dffrs_0.Qb a_8270_6060 avss.t8 nfet_03v3
**devattr s=10400,304 d=17600,576
X237 a_50878_1605.t1 a_50206_441 a_51066_2325 avdd.t316 pfet_03v3
**devattr s=31200,704 d=52800,1376
X238 a_44488_1651 a_44408_1559.t6 avss.t158 avss.t157 nfet_03v3
**devattr s=17600,576 d=10400,304
X239 avss.t133 a_31262_2781 a_31934_1605.t0 avss.t132 nfet_03v3
**devattr s=17600,576 d=17600,576
X240 avdd.t303 a_35016_2511.t6 a_34936_5969.t0 avdd.t302 pfet_03v3
**devattr s=26000,604 d=26000,604
X241 a_1290_3500.t2 load.t17 avdd.t175 avdd.t174 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X242 a_44488_3856 a_44408_3764.t7 avss.t176 avss.t175 nfet_03v3
**devattr s=17600,576 d=10400,304
X243 a_41594_2325 a_40734_441 a_41406_1605.t1 avdd.t58 pfet_03v3
**devattr s=52800,1376 d=31200,704
X244 avdd.t111 avdd.t109 a_53880_3764.t2 avdd.t110 pfet_03v3
**devattr s=26000,604 d=26000,604
X245 a_25464_3764.t3 a_25464_5969.t5 avdd.t245 avdd.t244 pfet_03v3
**devattr s=44000,1176 d=26000,604
X246 a_13178_2324 a_12318_440 a_12990_1604.t1 avdd.t0 pfet_03v3
**devattr s=52800,1376 d=31200,704
X247 a_29894_2781 load.t18 a_29706_3501.t1 avss.t187 nfet_03v3
**devattr s=17600,576 d=10400,304
X248 a_31262_441 a_29706_1161.t4 avdd.t57 avdd.t56 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X249 avdd.t37 a_38472_1361 a_39178_1161.t0 avdd.t36 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X250 dffrs_2.Q.t2 avdd.t106 avdd.t108 avdd.t107 pfet_03v3
**devattr s=44000,1176 d=26000,604
X251 a_34936_3764.t0 clk.t15 avdd.t351 avdd.t350 pfet_03v3
**devattr s=26000,604 d=44000,1176
X252 avdd.t227 a_53880_3764.t7 serial_out.t1 avdd.t226 pfet_03v3
**devattr s=26000,604 d=26000,604
X253 a_46158_3857 a_44408_1559.t7 a_45974_3857 avss.t159 nfet_03v3
**devattr s=10400,304 d=10400,304
X254 a_16072_2510.t0 2inmux_2.OUT.t3 a_16256_1650 avss.t162 nfet_03v3
**devattr s=10400,304 d=17600,576
X255 a_51066_2325 a_50206_2781 avdd.t183 avdd.t182 pfet_03v3
**devattr s=52800,1376 d=31200,704
X256 avdd.t55 avss.t290 a_1290_3500.t3 avdd.t54 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X257 a_15992_1558.t0 a_16072_2510.t6 a_16256_3855 avss.t164 nfet_03v3
**devattr s=10400,304 d=17600,576
X258 a_29894_441 a_29000_1361 avss.t13 avss.t12 nfet_03v3
**devattr s=17600,576 d=10400,304
X259 a_16256_6060 avdd.t396 a_16072_6060 avss.t75 nfet_03v3
**devattr s=10400,304 d=10400,304
X260 a_44408_3764.t1 clk.t16 a_44672_6061 avss.t248 nfet_03v3
**devattr s=10400,304 d=17600,576
X261 a_17742_3856 a_15992_1558.t6 a_17558_3856 avss.t192 nfet_03v3
**devattr s=10400,304 d=10400,304
X262 a_16256_8265 a_16072_2510.t7 a_16072_8265 avss.t163 nfet_03v3
**devattr s=10400,304 d=10400,304
X263 a_44408_5969.t1 a_44408_3764.t8 a_44672_8266 avss.t177 nfet_03v3
**devattr s=10400,304 d=17600,576
X264 a_46158_6061 a_44408_3764.t9 a_45974_6061 avss.t178 nfet_03v3
**devattr s=10400,304 d=10400,304
X265 dffrs_2.Qb avdd.t397 a_27214_3857 avss.t74 nfet_03v3
**devattr s=10400,304 d=17600,576
X266 a_17742_6060 a_15992_3763.t8 a_17558_6060 avss.t256 nfet_03v3
**devattr s=10400,304 d=10400,304
X267 dffrs_2.Qb dffrs_2.Q.t8 avdd.t311 avdd.t310 pfet_03v3
**devattr s=44000,1176 d=26000,604
X268 avdd.t39 a_53880_1559.t6 dffrs_5.Qb avdd.t38 pfet_03v3
**devattr s=26000,604 d=26000,604
X269 avdd.t291 a_53960_2511.t6 a_53880_5969.t1 avdd.t290 pfet_03v3
**devattr s=26000,604 d=26000,604
X270 dffrs_2.Q.t0 dffrs_2.Qb a_27214_6061 avss.t9 nfet_03v3
**devattr s=10400,304 d=17600,576
X271 a_25464_5969.t0 avdd.t103 avdd.t105 avdd.t104 pfet_03v3
**devattr s=44000,1176 d=26000,604
X272 a_10056_1360 load.t19 avdd.t271 avdd.t270 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X273 a_34936_5969.t1 a_34936_3764.t8 avdd.t65 avdd.t64 pfet_03v3
**devattr s=26000,604 d=44000,1176
X274 a_31262_441 a_29706_1161.t5 avss.t237 avss.t236 nfet_03v3
**devattr s=17600,576 d=17600,576
X275 a_15992_3763.t3 a_15992_5968.t5 avdd.t299 avdd.t298 pfet_03v3
**devattr s=44000,1176 d=26000,604
X276 a_35200_1651 avdd.t398 a_35016_1651 avss.t73 nfet_03v3
**devattr s=10400,304 d=10400,304
X277 a_10762_3500.t1 load.t21 a_10950_2780 avss.t107 nfet_03v3
**devattr s=10400,304 d=17600,576
X278 a_584_1360 load.t20 avdd.t173 avdd.t172 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X279 a_53880_3764.t1 clk.t17 avdd.t339 avdd.t338 pfet_03v3
**devattr s=26000,604 d=44000,1176
X280 2inmux_1.Bit.t0 avdd.t79 avdd.t81 avdd.t80 pfet_03v3
**devattr s=44000,1176 d=26000,604
X281 avdd.t102 avdd.t100 a_25464_3764.t2 avdd.t101 pfet_03v3
**devattr s=26000,604 d=26000,604
X282 a_35200_3856 clk.t19 a_35016_3856 avss.t244 nfet_03v3
**devattr s=10400,304 d=10400,304
X283 a_53960_6061 a_53880_5969.t5 avss.t199 avss.t198 nfet_03v3
**devattr s=17600,576 d=10400,304
X284 a_6520_3763.t2 clk.t18 avdd.t341 avdd.t340 pfet_03v3
**devattr s=26000,604 d=44000,1176
X285 a_29000_1361 load.t22 avss.t33 avss.t32 nfet_03v3
**devattr s=17600,576 d=17600,576
X286 avdd.t99 avdd.t97 a_44488_2511.t0 avdd.t98 pfet_03v3
**devattr s=26000,604 d=26000,604
X287 avdd.t181 a_50206_2781 a_51066_2325 avdd.t180 pfet_03v3
**devattr s=31200,704 d=52800,1376
X288 a_36502_3857 dffrs_3.Q.t7 avss.t191 avss.t190 nfet_03v3
**devattr s=17600,576 d=10400,304
X289 serial_out.t2 dffrs_5.Qb avdd.t335 avdd.t334 pfet_03v3
**devattr s=26000,604 d=44000,1176
X290 a_53960_8266 avdd.t399 avss.t72 avss.t71 nfet_03v3
**devattr s=17600,576 d=10400,304
X291 a_3706_2324 a_2846_2780 avdd.t375 avdd.t374 pfet_03v3
**devattr s=52800,1376 d=31200,704
X292 avdd.t347 clk.t20 a_44408_1559.t1 avdd.t346 pfet_03v3
**devattr s=26000,604 d=26000,604
X293 2inmux_5.OUT.t0 a_41406_1605.t5 avdd.t239 avdd.t238 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X294 a_25544_2511.t1 2inmux_3.OUT.t3 avdd.t179 avdd.t178 pfet_03v3
**devattr s=26000,604 d=44000,1176
X295 dffrs_1.Qb avdd.t401 a_17742_3856 avss.t68 nfet_03v3
**devattr s=10400,304 d=17600,576
X296 dffrs_4.Qb 2inmux_1.Bit.t8 avdd.t305 avdd.t304 pfet_03v3
**devattr s=44000,1176 d=26000,604
X297 a_36502_6061 avdd.t400 avss.t70 avss.t69 nfet_03v3
**devattr s=17600,576 d=10400,304
X298 dffrs_5.Qb avdd.t94 avdd.t96 avdd.t95 pfet_03v3
**devattr s=26000,604 d=44000,1176
X299 a_25464_1559.t2 a_25544_2511.t6 avdd.t207 avdd.t206 pfet_03v3
**devattr s=26000,604 d=44000,1176
X300 avss.t11 a_29000_1361 a_29894_441 avss.t10 nfet_03v3
**devattr s=10400,304 d=17600,576
X301 dffrs_1.Q.t2 dffrs_1.Qb a_17742_6060 avss.t129 nfet_03v3
**devattr s=10400,304 d=17600,576
X302 a_53880_5969.t3 a_53880_3764.t8 avdd.t229 avdd.t228 pfet_03v3
**devattr s=26000,604 d=44000,1176
X303 a_15992_5968.t2 avdd.t91 avdd.t93 avdd.t92 pfet_03v3
**devattr s=44000,1176 d=26000,604
X304 a_54144_1651 avdd.t402 a_53960_1651 avss.t67 nfet_03v3
**devattr s=10400,304 d=10400,304
X305 a_10762_3500.t0 load.t23 avdd.t45 avdd.t44 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X306 avdd.t209 a_25544_2511.t7 a_25464_5969.t1 avdd.t208 pfet_03v3
**devattr s=26000,604 d=26000,604
X307 a_32122_2325 a_31262_441 a_31934_1605.t1 avdd.t314 pfet_03v3
**devattr s=52800,1376 d=31200,704
X308 a_25544_1651 a_25464_1559.t7 avss.t58 avss.t57 nfet_03v3
**devattr s=17600,576 d=10400,304
X309 a_6520_5968.t1 a_6520_3763.t9 avdd.t333 avdd.t332 pfet_03v3
**devattr s=26000,604 d=44000,1176
X310 a_54144_3856 clk.t21 a_53960_3856 avss.t246 nfet_03v3
**devattr s=10400,304 d=10400,304
X311 a_25544_3856 a_25464_3764.t9 avss.t207 avss.t206 nfet_03v3
**devattr s=17600,576 d=10400,304
X312 a_35016_2511.t3 2inmux_4.OUT.t3 a_35200_1651 avss.t231 nfet_03v3
**devattr s=10400,304 d=17600,576
X313 a_47944_1361 load.t24 avss.t185 avss.t184 nfet_03v3
**devattr s=17600,576 d=17600,576
X314 a_48838_441 B1.t0 a_48650_1161.t0 avss.t4 nfet_03v3
**devattr s=17600,576 d=10400,304
X315 a_55446_3857 serial_out.t5 avss.t111 avss.t110 nfet_03v3
**devattr s=17600,576 d=10400,304
X316 a_50878_1605.t3 a_50206_441 avss.t227 avss.t226 nfet_03v3
**devattr s=17600,576 d=17600,576
X317 a_34936_1559.t2 a_35016_2511.t7 a_35200_3856 avss.t152 nfet_03v3
**devattr s=10400,304 d=17600,576
X318 dffrs_1.Q.t0 avdd.t88 avdd.t90 avdd.t89 pfet_03v3
**devattr s=44000,1176 d=26000,604
X319 a_44488_2511.t2 2inmux_5.OUT.t3 avdd.t253 avdd.t252 pfet_03v3
**devattr s=26000,604 d=44000,1176
X320 a_48838_2781 load.t25 a_48650_3501.t3 avss.t186 nfet_03v3
**devattr s=17600,576 d=10400,304
X321 a_36686_3857 a_34936_1559.t7 a_36502_3857 avss.t137 nfet_03v3
**devattr s=10400,304 d=10400,304
X322 a_55446_6061 avdd.t403 avss.t66 avss.t65 nfet_03v3
**devattr s=17600,576 d=10400,304
X323 a_6600_6060 a_6520_5968.t5 avss.t122 avss.t121 nfet_03v3
**devattr s=17600,576 d=10400,304
X324 avdd.t273 a_21790_2781 a_22650_2325 avdd.t272 pfet_03v3
**devattr s=31200,704 d=52800,1376
X325 avdd.t87 avdd.t85 a_16072_2510.t2 avdd.t86 pfet_03v3
**devattr s=26000,604 d=26000,604
X326 a_44408_1559.t3 a_44488_2511.t7 avdd.t257 avdd.t256 pfet_03v3
**devattr s=26000,604 d=44000,1176
X327 avdd.t349 clk.t22 a_15992_1558.t2 avdd.t348 pfet_03v3
**devattr s=26000,604 d=26000,604
X328 a_36686_6061 a_34936_3764.t9 a_36502_6061 avss.t49 nfet_03v3
**devattr s=10400,304 d=10400,304
X329 a_6600_8265 avdd.t404 avss.t64 avss.t63 nfet_03v3
**devattr s=17600,576 d=10400,304
X330 a_48650_1161.t1 B1.t1 avdd.t3 avdd.t2 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X331 2inmux_2.OUT.t0 a_12990_1604.t5 avdd.t367 avdd.t366 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X332 avss.t276 2inmux_2.Bit.t7 a_10950_2780 avss.t275 nfet_03v3
**devattr s=10400,304 d=17600,576
X333 dffrs_1.Qb dffrs_1.Q.t7 avdd.t19 avdd.t18 pfet_03v3
**devattr s=44000,1176 d=26000,604
X334 avss.t156 dffrs_3.Q.t8 a_39366_2781 avss.t155 nfet_03v3
**devattr s=10400,304 d=17600,576
X335 a_16072_1650 a_15992_1558.t7 avss.t194 avss.t193 nfet_03v3
**devattr s=17600,576 d=10400,304
X336 a_38472_1361 load.t26 avdd.t73 avdd.t72 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X337 a_40734_441 a_39178_1161.t5 avdd.t255 avdd.t254 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X338 a_53960_2511.t2 2inmux_1.OUT.t3 a_54144_1651 avss.t210 nfet_03v3
**devattr s=10400,304 d=17600,576
X339 a_29894_441 B3.t0 a_29706_1161.t2 avss.t34 nfet_03v3
**devattr s=17600,576 d=10400,304
X340 a_25728_1651 avdd.t405 a_25544_1651 avss.t62 nfet_03v3
**devattr s=10400,304 d=10400,304
X341 a_34936_3764.t3 a_34936_5969.t5 avdd.t247 avdd.t246 pfet_03v3
**devattr s=44000,1176 d=26000,604
X342 a_53960_2511.t0 a_53880_1559.t7 avdd.t41 avdd.t40 pfet_03v3
**devattr s=44000,1176 d=26000,604
X343 avdd.t359 a_47944_1361 a_48650_1161.t3 avdd.t358 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X344 a_6600_2510.t1 2inmux_0.OUT.t3 a_6784_1650 avss.t167 nfet_03v3
**devattr s=10400,304 d=17600,576
X345 a_53880_1559.t3 a_53960_2511.t7 a_54144_3856 avss.t197 nfet_03v3
**devattr s=10400,304 d=17600,576
X346 a_16072_3855 a_15992_3763.t9 avss.t258 avss.t257 nfet_03v3
**devattr s=17600,576 d=10400,304
X347 a_20234_3501.t0 load.t27 a_20422_2781 avss.t55 nfet_03v3
**devattr s=10400,304 d=17600,576
X348 a_25728_3856 clk.t23 a_25544_3856 avss.t243 nfet_03v3
**devattr s=10400,304 d=10400,304
X349 a_53880_1559.t1 a_53880_3764.t9 avdd.t231 avdd.t230 pfet_03v3
**devattr s=44000,1176 d=26000,604
X350 avdd.t29 a_40734_2781 a_41594_2325 avdd.t28 pfet_03v3
**devattr s=31200,704 d=52800,1376
X351 a_8086_3856 2inmux_2.Bit.t8 avss.t278 avss.t277 nfet_03v3
**devattr s=17600,576 d=10400,304
X352 a_6520_1558.t1 a_6600_2510.t6 a_6784_3855 avss.t18 nfet_03v3
**devattr s=10400,304 d=17600,576
X353 a_32122_2325 a_31262_2781 avdd.t203 avdd.t202 pfet_03v3
**devattr s=52800,1376 d=31200,704
X354 a_29706_1161.t3 B3.t1 avdd.t47 avdd.t46 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X355 a_6784_6060 avdd.t406 a_6600_6060 avss.t61 nfet_03v3
**devattr s=10400,304 d=10400,304
X356 dffrs_3.Q.t2 dffrs_3.Qb avdd.t61 avdd.t60 pfet_03v3
**devattr s=26000,604 d=44000,1176
X357 a_50206_2781 a_48650_3501.t5 avss.t254 avss.t253 nfet_03v3
**devattr s=17600,576 d=17600,576
X358 a_48650_1161.t2 B1.t2 a_48838_441 avss.t228 nfet_03v3
**devattr s=10400,304 d=17600,576
X359 a_8086_6060 avdd.t407 avss.t60 avss.t59 nfet_03v3
**devattr s=17600,576 d=10400,304
X360 a_6784_8265 a_6600_2510.t7 a_6600_8265 avss.t19 nfet_03v3
**devattr s=10400,304 d=10400,304
X361 a_20422_2781 dffrs_1.Q.t8 avss.t1 avss.t0 nfet_03v3
**devattr s=17600,576 d=10400,304
X362 a_34936_5969.t3 avdd.t82 avdd.t84 avdd.t83 pfet_03v3
**devattr s=44000,1176 d=26000,604
X363 a_2846_2780 a_1290_3500.t5 avss.t281 avss.t280 nfet_03v3
**devattr s=17600,576 d=17600,576
X364 a_29706_1161.t1 B3.t2 a_29894_441 avss.t31 nfet_03v3
**devattr s=10400,304 d=17600,576
X365 dffrs_3.Qb avdd.t76 avdd.t78 avdd.t77 pfet_03v3
**devattr s=26000,604 d=44000,1176
X366 a_20234_3501.t3 load.t28 avdd.t191 avdd.t190 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X367 a_39178_3501.t2 load.t29 a_39366_2781 avss.t125 nfet_03v3
**devattr s=10400,304 d=17600,576
X368 a_48838_441 a_47944_1361 avss.t264 avss.t263 nfet_03v3
**devattr s=17600,576 d=10400,304
X369 a_3518_1604.t1 a_2846_440 a_3706_2324 avdd.t10 pfet_03v3
**devattr s=31200,704 d=52800,1376
X370 a_12318_440 a_10762_1160.t5 avdd.t223 avdd.t222 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X371 a_44488_6061 a_44408_5969.t5 avss.t230 avss.t229 nfet_03v3
**devattr s=17600,576 d=10400,304
R0 avdd.t266 avdd.n390 250.9
R1 avdd.n391 avdd.t92 250.9
R2 avdd.t24 avdd.n401 250.9
R3 avdd.n402 avdd.t298 250.9
R4 avdd.t198 avdd.n396 250.9
R5 avdd.n397 avdd.t89 250.9
R6 avdd.t240 avdd.n413 250.9
R7 avdd.n414 avdd.t264 250.9
R8 avdd.t140 avdd.n407 250.9
R9 avdd.n408 avdd.t18 250.9
R10 avdd.t248 avdd.n425 250.9
R11 avdd.n426 avdd.t286 250.9
R12 avdd.t228 avdd.n98 250.9
R13 avdd.n99 avdd.t143 250.9
R14 avdd.t338 avdd.n109 250.9
R15 avdd.n110 avdd.t292 250.9
R16 avdd.t334 avdd.n104 250.9
R17 avdd.n105 avdd.t137 250.9
R18 avdd.t250 avdd.n121 250.9
R19 avdd.n122 avdd.t230 250.9
R20 avdd.t95 avdd.n115 250.9
R21 avdd.n116 avdd.t176 250.9
R22 avdd.t308 avdd.n132 250.9
R23 avdd.n133 avdd.t40 250.9
R24 avdd.t196 avdd.n171 250.9
R25 avdd.n172 avdd.t119 250.9
R26 avdd.t344 avdd.n182 250.9
R27 avdd.n183 avdd.t318 250.9
R28 avdd.t352 avdd.n177 250.9
R29 avdd.n178 avdd.t80 250.9
R30 avdd.t256 avdd.n194 250.9
R31 avdd.n195 avdd.t192 250.9
R32 avdd.t116 avdd.n188 250.9
R33 avdd.n189 avdd.t304 250.9
R34 avdd.t252 avdd.n205 250.9
R35 avdd.n206 avdd.t280 250.9
R36 avdd.t64 avdd.n244 250.9
R37 avdd.n245 avdd.t83 250.9
R38 avdd.t350 avdd.n255 250.9
R39 avdd.n256 avdd.t246 250.9
R40 avdd.t60 avdd.n250 250.9
R41 avdd.n251 avdd.t149 250.9
R42 avdd.t300 avdd.n267 250.9
R43 avdd.n268 avdd.t62 250.9
R44 avdd.t77 avdd.n261 250.9
R45 avdd.n262 avdd.t278 250.9
R46 avdd.t296 avdd.n278 250.9
R47 avdd.n279 avdd.t216 250.9
R48 avdd.t322 avdd.n317 250.9
R49 avdd.n318 avdd.t104 250.9
R50 avdd.t26 avdd.n328 250.9
R51 avdd.n329 avdd.t244 250.9
R52 avdd.t14 avdd.n323 250.9
R53 avdd.n324 avdd.t107 250.9
R54 avdd.t206 avdd.n340 250.9
R55 avdd.n341 avdd.t324 250.9
R56 avdd.t152 avdd.n334 250.9
R57 avdd.n335 avdd.t310 250.9
R58 avdd.t178 avdd.n351 250.9
R59 avdd.n352 avdd.t364 250.9
R60 avdd.t332 avdd.n4 250.9
R61 avdd.n5 avdd.t131 250.9
R62 avdd.t340 avdd.n528 250.9
R63 avdd.n529 avdd.t186 250.9
R64 avdd.t12 avdd.n9 250.9
R65 avdd.n10 avdd.t125 250.9
R66 avdd.t4 avdd.n516 250.9
R67 avdd.n517 avdd.t328 250.9
R68 avdd.t158 avdd.n522 250.9
R69 avdd.n523 avdd.t368 250.9
R70 avdd.t370 avdd.n465 250.9
R71 avdd.n466 avdd.t50 250.9
R72 avdd.n495 avdd.t188 236.083
R73 avdd.t174 avdd.n491 236.083
R74 avdd.t210 avdd.n499 236.083
R75 avdd.n505 avdd.t74 236.083
R76 avdd.n453 avdd.t306 236.083
R77 avdd.t44 avdd.n450 236.083
R78 avdd.t222 avdd.n433 236.083
R79 avdd.n439 avdd.t218 236.083
R80 avdd.n379 avdd.t260 236.083
R81 avdd.t190 avdd.n376 236.083
R82 avdd.t236 avdd.n359 236.083
R83 avdd.n365 avdd.t220 236.083
R84 avdd.n306 avdd.t200 236.083
R85 avdd.t268 avdd.n303 236.083
R86 avdd.t56 avdd.n286 236.083
R87 avdd.n292 avdd.t46 236.083
R88 avdd.n233 avdd.t354 236.083
R89 avdd.t168 avdd.n230 236.083
R90 avdd.t254 avdd.n213 236.083
R91 avdd.n219 avdd.t232 236.083
R92 avdd.n160 avdd.t336 236.083
R93 avdd.t212 avdd.n157 236.083
R94 avdd.t258 avdd.n140 236.083
R95 avdd.n146 avdd.t2 236.083
R96 avdd.n92 avdd.t214 236.083
R97 avdd.n86 avdd.t182 236.083
R98 avdd.n76 avdd.t238 236.083
R99 avdd.n70 avdd.t30 236.083
R100 avdd.n60 avdd.t294 236.083
R101 avdd.n54 avdd.t202 236.083
R102 avdd.n44 avdd.t166 236.083
R103 avdd.n38 avdd.t274 236.083
R104 avdd.n28 avdd.t366 236.083
R105 avdd.n22 avdd.t32 236.083
R106 avdd.t234 avdd.n470 236.083
R107 avdd.n481 avdd.t374 236.083
R108 avdd.t188 avdd.n494 235.294
R109 avdd.n494 avdd.t174 235.294
R110 avdd.n504 avdd.t210 235.294
R111 avdd.t74 avdd.n504 235.294
R112 avdd.t306 avdd.n452 235.294
R113 avdd.n452 avdd.t44 235.294
R114 avdd.n438 avdd.t222 235.294
R115 avdd.t218 avdd.n438 235.294
R116 avdd.t260 avdd.n378 235.294
R117 avdd.n378 avdd.t190 235.294
R118 avdd.n364 avdd.t236 235.294
R119 avdd.t220 avdd.n364 235.294
R120 avdd.t200 avdd.n305 235.294
R121 avdd.n305 avdd.t268 235.294
R122 avdd.n291 avdd.t56 235.294
R123 avdd.t46 avdd.n291 235.294
R124 avdd.t354 avdd.n232 235.294
R125 avdd.n232 avdd.t168 235.294
R126 avdd.n218 avdd.t254 235.294
R127 avdd.t232 avdd.n218 235.294
R128 avdd.t336 avdd.n159 235.294
R129 avdd.n159 avdd.t212 235.294
R130 avdd.n145 avdd.t258 235.294
R131 avdd.t2 avdd.n145 235.294
R132 avdd.t214 avdd.n91 235.294
R133 avdd.n91 avdd.t316 235.294
R134 avdd.t317 avdd.n89 235.294
R135 avdd.n89 avdd.t180 235.294
R136 avdd.t238 avdd.n75 235.294
R137 avdd.n75 avdd.t59 235.294
R138 avdd.t58 avdd.n73 235.294
R139 avdd.n73 avdd.t28 235.294
R140 avdd.t294 avdd.n59 235.294
R141 avdd.n59 avdd.t315 235.294
R142 avdd.t314 avdd.n57 235.294
R143 avdd.n57 avdd.t204 235.294
R144 avdd.t166 avdd.n43 235.294
R145 avdd.n43 avdd.t373 235.294
R146 avdd.t372 avdd.n41 235.294
R147 avdd.n41 avdd.t272 235.294
R148 avdd.t366 avdd.n27 235.294
R149 avdd.n27 avdd.t1 235.294
R150 avdd.t0 avdd.n25 235.294
R151 avdd.n25 avdd.t34 235.294
R152 avdd.n478 avdd.t234 235.294
R153 avdd.t10 avdd.n478 235.294
R154 avdd.n480 avdd.t11 235.294
R155 avdd.t376 avdd.n480 235.294
R156 avdd.t242 avdd.t266 200
R157 avdd.t92 avdd.t242 200
R158 avdd.t155 avdd.t24 200
R159 avdd.t298 avdd.t155 200
R160 avdd.t262 avdd.t198 200
R161 avdd.t89 avdd.t262 200
R162 avdd.t348 avdd.t240 200
R163 avdd.t264 avdd.t348 200
R164 avdd.t284 avdd.t140 200
R165 avdd.t18 avdd.t284 200
R166 avdd.t86 avdd.t248 200
R167 avdd.t286 avdd.t86 200
R168 avdd.t290 avdd.t228 200
R169 avdd.t143 avdd.t290 200
R170 avdd.t110 avdd.t338 200
R171 avdd.t292 avdd.t110 200
R172 avdd.t226 avdd.t334 200
R173 avdd.t137 avdd.t226 200
R174 avdd.t8 avdd.t250 200
R175 avdd.t230 avdd.t8 200
R176 avdd.t38 avdd.t95 200
R177 avdd.t176 avdd.t38 200
R178 avdd.t134 avdd.t308 200
R179 avdd.t40 avdd.t134 200
R180 avdd.t316 avdd.t317 200
R181 avdd.t182 avdd.t180 200
R182 avdd.t288 avdd.t196 200
R183 avdd.t119 avdd.t288 200
R184 avdd.t164 avdd.t344 200
R185 avdd.t318 avdd.t164 200
R186 avdd.t194 avdd.t352 200
R187 avdd.t80 avdd.t194 200
R188 avdd.t346 avdd.t256 200
R189 avdd.t192 avdd.t346 200
R190 avdd.t282 avdd.t116 200
R191 avdd.t304 avdd.t282 200
R192 avdd.t98 avdd.t252 200
R193 avdd.t280 avdd.t98 200
R194 avdd.t59 avdd.t58 200
R195 avdd.t30 avdd.t28 200
R196 avdd.t302 avdd.t64 200
R197 avdd.t83 avdd.t302 200
R198 avdd.t113 avdd.t350 200
R199 avdd.t246 avdd.t113 200
R200 avdd.t360 avdd.t60 200
R201 avdd.t149 avdd.t360 200
R202 avdd.t6 avdd.t300 200
R203 avdd.t62 avdd.t6 200
R204 avdd.t224 avdd.t77 200
R205 avdd.t278 avdd.t224 200
R206 avdd.t146 avdd.t296 200
R207 avdd.t216 avdd.t146 200
R208 avdd.t315 avdd.t314 200
R209 avdd.t202 avdd.t204 200
R210 avdd.t208 avdd.t322 200
R211 avdd.t104 avdd.t208 200
R212 avdd.t101 avdd.t26 200
R213 avdd.t244 avdd.t101 200
R214 avdd.t320 avdd.t14 200
R215 avdd.t107 avdd.t320 200
R216 avdd.t22 avdd.t206 200
R217 avdd.t324 avdd.t22 200
R218 avdd.t362 avdd.t152 200
R219 avdd.t310 avdd.t362 200
R220 avdd.t122 avdd.t178 200
R221 avdd.t364 avdd.t122 200
R222 avdd.t373 avdd.t372 200
R223 avdd.t274 avdd.t272 200
R224 avdd.t1 avdd.t0 200
R225 avdd.t32 avdd.t34 200
R226 avdd.t20 avdd.t332 200
R227 avdd.t131 avdd.t20 200
R228 avdd.t128 avdd.t340 200
R229 avdd.t186 avdd.t128 200
R230 avdd.t330 avdd.t12 200
R231 avdd.t125 avdd.t330 200
R232 avdd.t342 avdd.t4 200
R233 avdd.t328 avdd.t342 200
R234 avdd.t52 avdd.t158 200
R235 avdd.t368 avdd.t52 200
R236 avdd.t161 avdd.t370 200
R237 avdd.t50 avdd.t161 200
R238 avdd.t11 avdd.t10 200
R239 avdd.t374 avdd.t376 200
R240 avdd.n486 avdd.t54 131.589
R241 avdd.n507 avdd.t48 131.589
R242 avdd.n14 avdd.t356 131.589
R243 avdd.n441 avdd.t326 131.589
R244 avdd.n30 avdd.t42 131.589
R245 avdd.n367 avdd.t66 131.589
R246 avdd.n46 avdd.t312 131.589
R247 avdd.n294 avdd.t16 131.589
R248 avdd.n62 avdd.t276 131.589
R249 avdd.n221 avdd.t36 131.589
R250 avdd.n78 avdd.t184 131.589
R251 avdd.n148 avdd.t358 131.589
R252 avdd.n164 avdd.t70 118.543
R253 avdd.n237 avdd.t72 118.543
R254 avdd.n310 avdd.t68 118.543
R255 avdd.n383 avdd.t170 118.543
R256 avdd.n457 avdd.t270 118.543
R257 avdd.n487 avdd.t172 118.543
R258 avdd.n86 avdd.n85 96.0755
R259 avdd.n87 avdd.n86 96.0755
R260 avdd.n70 avdd.n69 96.0755
R261 avdd.n71 avdd.n70 96.0755
R262 avdd.n54 avdd.n53 96.0755
R263 avdd.n55 avdd.n54 96.0755
R264 avdd.n38 avdd.n37 96.0755
R265 avdd.n39 avdd.n38 96.0755
R266 avdd.n22 avdd.n21 96.0755
R267 avdd.n23 avdd.n22 96.0755
R268 avdd.n481 avdd.n473 96.0755
R269 avdd.n481 avdd.n474 96.0755
R270 avdd.n501 avdd.n499 78.2255
R271 avdd.n505 avdd.n501 78.2255
R272 avdd.n505 avdd.n502 78.2255
R273 avdd.n502 avdd.n499 78.2255
R274 avdd.n435 avdd.n433 78.2255
R275 avdd.n439 avdd.n435 78.2255
R276 avdd.n439 avdd.n436 78.2255
R277 avdd.n436 avdd.n433 78.2255
R278 avdd.n361 avdd.n359 78.2255
R279 avdd.n365 avdd.n361 78.2255
R280 avdd.n365 avdd.n362 78.2255
R281 avdd.n362 avdd.n359 78.2255
R282 avdd.n288 avdd.n286 78.2255
R283 avdd.n292 avdd.n288 78.2255
R284 avdd.n292 avdd.n289 78.2255
R285 avdd.n289 avdd.n286 78.2255
R286 avdd.n215 avdd.n213 78.2255
R287 avdd.n219 avdd.n215 78.2255
R288 avdd.n219 avdd.n216 78.2255
R289 avdd.n216 avdd.n213 78.2255
R290 avdd.n142 avdd.n140 78.2255
R291 avdd.n146 avdd.n142 78.2255
R292 avdd.n146 avdd.n143 78.2255
R293 avdd.n143 avdd.n140 78.2255
R294 avdd.n92 avdd.n83 78.2255
R295 avdd.n92 avdd.n84 78.2255
R296 avdd.n160 avdd.n155 78.2255
R297 avdd.n160 avdd.n156 78.2255
R298 avdd.n157 avdd.n155 78.2255
R299 avdd.n157 avdd.n156 78.2255
R300 avdd.n76 avdd.n67 78.2255
R301 avdd.n76 avdd.n68 78.2255
R302 avdd.n233 avdd.n228 78.2255
R303 avdd.n233 avdd.n229 78.2255
R304 avdd.n230 avdd.n228 78.2255
R305 avdd.n230 avdd.n229 78.2255
R306 avdd.n60 avdd.n51 78.2255
R307 avdd.n60 avdd.n52 78.2255
R308 avdd.n306 avdd.n301 78.2255
R309 avdd.n306 avdd.n302 78.2255
R310 avdd.n303 avdd.n301 78.2255
R311 avdd.n303 avdd.n302 78.2255
R312 avdd.n44 avdd.n35 78.2255
R313 avdd.n44 avdd.n36 78.2255
R314 avdd.n379 avdd.n374 78.2255
R315 avdd.n379 avdd.n375 78.2255
R316 avdd.n376 avdd.n374 78.2255
R317 avdd.n376 avdd.n375 78.2255
R318 avdd.n28 avdd.n19 78.2255
R319 avdd.n28 avdd.n20 78.2255
R320 avdd.n453 avdd.n448 78.2255
R321 avdd.n453 avdd.n449 78.2255
R322 avdd.n450 avdd.n448 78.2255
R323 avdd.n450 avdd.n449 78.2255
R324 avdd.n475 avdd.n470 78.2255
R325 avdd.n476 avdd.n470 78.2255
R326 avdd.n495 avdd.n484 78.2255
R327 avdd.n495 avdd.n485 78.2255
R328 avdd.n491 avdd.n484 78.2255
R329 avdd.n491 avdd.n485 78.2255
R330 avdd.n391 avdd.n390 68.0765
R331 avdd.n402 avdd.n401 68.0765
R332 avdd.n397 avdd.n396 68.0765
R333 avdd.n414 avdd.n413 68.0765
R334 avdd.n408 avdd.n407 68.0765
R335 avdd.n426 avdd.n425 68.0765
R336 avdd.n99 avdd.n98 68.0765
R337 avdd.n110 avdd.n109 68.0765
R338 avdd.n105 avdd.n104 68.0765
R339 avdd.n122 avdd.n121 68.0765
R340 avdd.n116 avdd.n115 68.0765
R341 avdd.n133 avdd.n132 68.0765
R342 avdd.n172 avdd.n171 68.0765
R343 avdd.n183 avdd.n182 68.0765
R344 avdd.n178 avdd.n177 68.0765
R345 avdd.n195 avdd.n194 68.0765
R346 avdd.n189 avdd.n188 68.0765
R347 avdd.n206 avdd.n205 68.0765
R348 avdd.n245 avdd.n244 68.0765
R349 avdd.n256 avdd.n255 68.0765
R350 avdd.n251 avdd.n250 68.0765
R351 avdd.n268 avdd.n267 68.0765
R352 avdd.n262 avdd.n261 68.0765
R353 avdd.n279 avdd.n278 68.0765
R354 avdd.n318 avdd.n317 68.0765
R355 avdd.n329 avdd.n328 68.0765
R356 avdd.n324 avdd.n323 68.0765
R357 avdd.n341 avdd.n340 68.0765
R358 avdd.n335 avdd.n334 68.0765
R359 avdd.n352 avdd.n351 68.0765
R360 avdd.n5 avdd.n4 68.0765
R361 avdd.n529 avdd.n528 68.0765
R362 avdd.n10 avdd.n9 68.0765
R363 avdd.n517 avdd.n516 68.0765
R364 avdd.n523 avdd.n522 68.0765
R365 avdd.n466 avdd.n465 68.0765
R366 avdd.n85 avdd.n83 59.8505
R367 avdd.n87 avdd.n84 59.8505
R368 avdd.n69 avdd.n67 59.8505
R369 avdd.n71 avdd.n68 59.8505
R370 avdd.n53 avdd.n51 59.8505
R371 avdd.n55 avdd.n52 59.8505
R372 avdd.n37 avdd.n35 59.8505
R373 avdd.n39 avdd.n36 59.8505
R374 avdd.n21 avdd.n19 59.8505
R375 avdd.n23 avdd.n20 59.8505
R376 avdd.n475 avdd.n473 59.8505
R377 avdd.n476 avdd.n474 59.8505
R378 avdd.n419 avdd.t139 41.0041
R379 avdd.n126 avdd.t94 41.0041
R380 avdd.n199 avdd.t115 41.0041
R381 avdd.n272 avdd.t76 41.0041
R382 avdd.n345 avdd.t151 41.0041
R383 avdd.n459 avdd.t157 41.0041
R384 avdd.n421 avdd.t85 40.8177
R385 avdd.n420 avdd.t154 40.8177
R386 avdd.n128 avdd.t133 40.8177
R387 avdd.n127 avdd.t109 40.8177
R388 avdd.n201 avdd.t97 40.8177
R389 avdd.n200 avdd.t163 40.8177
R390 avdd.n274 avdd.t145 40.8177
R391 avdd.n273 avdd.t112 40.8177
R392 avdd.n347 avdd.t121 40.8177
R393 avdd.n346 avdd.t100 40.8177
R394 avdd.n461 avdd.t160 40.8177
R395 avdd.n460 avdd.t127 40.8177
R396 avdd.n386 avdd.t91 40.6313
R397 avdd.n385 avdd.t88 40.6313
R398 avdd.n94 avdd.t142 40.6313
R399 avdd.n93 avdd.t136 40.6313
R400 avdd.n167 avdd.t118 40.6313
R401 avdd.n166 avdd.t79 40.6313
R402 avdd.n240 avdd.t82 40.6313
R403 avdd.n239 avdd.t148 40.6313
R404 avdd.n313 avdd.t103 40.6313
R405 avdd.n312 avdd.t106 40.6313
R406 avdd.n1 avdd.t130 40.6313
R407 avdd.n0 avdd.t124 40.6313
R408 avdd.n503 avdd.n501 36.2255
R409 avdd.n503 avdd.n502 36.2255
R410 avdd.n437 avdd.n435 36.2255
R411 avdd.n437 avdd.n436 36.2255
R412 avdd.n363 avdd.n361 36.2255
R413 avdd.n363 avdd.n362 36.2255
R414 avdd.n290 avdd.n288 36.2255
R415 avdd.n290 avdd.n289 36.2255
R416 avdd.n217 avdd.n215 36.2255
R417 avdd.n217 avdd.n216 36.2255
R418 avdd.n144 avdd.n142 36.2255
R419 avdd.n144 avdd.n143 36.2255
R420 avdd.n88 avdd.n85 36.2255
R421 avdd.n88 avdd.n87 36.2255
R422 avdd.n90 avdd.n83 36.2255
R423 avdd.n90 avdd.n84 36.2255
R424 avdd.n158 avdd.n155 36.2255
R425 avdd.n158 avdd.n156 36.2255
R426 avdd.n72 avdd.n69 36.2255
R427 avdd.n72 avdd.n71 36.2255
R428 avdd.n74 avdd.n67 36.2255
R429 avdd.n74 avdd.n68 36.2255
R430 avdd.n231 avdd.n228 36.2255
R431 avdd.n231 avdd.n229 36.2255
R432 avdd.n56 avdd.n53 36.2255
R433 avdd.n56 avdd.n55 36.2255
R434 avdd.n58 avdd.n51 36.2255
R435 avdd.n58 avdd.n52 36.2255
R436 avdd.n304 avdd.n301 36.2255
R437 avdd.n304 avdd.n302 36.2255
R438 avdd.n40 avdd.n37 36.2255
R439 avdd.n40 avdd.n39 36.2255
R440 avdd.n42 avdd.n35 36.2255
R441 avdd.n42 avdd.n36 36.2255
R442 avdd.n377 avdd.n374 36.2255
R443 avdd.n377 avdd.n375 36.2255
R444 avdd.n24 avdd.n21 36.2255
R445 avdd.n24 avdd.n23 36.2255
R446 avdd.n26 avdd.n19 36.2255
R447 avdd.n26 avdd.n20 36.2255
R448 avdd.n451 avdd.n448 36.2255
R449 avdd.n451 avdd.n449 36.2255
R450 avdd.n479 avdd.n473 36.2255
R451 avdd.n479 avdd.n474 36.2255
R452 avdd.n477 avdd.n475 36.2255
R453 avdd.n477 avdd.n476 36.2255
R454 avdd.n493 avdd.n484 36.2255
R455 avdd.n493 avdd.n485 36.2255
R456 avdd.n386 avdd.t388 27.3166
R457 avdd.n385 avdd.t390 27.3166
R458 avdd.n94 avdd.t399 27.3166
R459 avdd.n93 avdd.t403 27.3166
R460 avdd.n167 avdd.t378 27.3166
R461 avdd.n166 avdd.t386 27.3166
R462 avdd.n240 avdd.t391 27.3166
R463 avdd.n239 avdd.t400 27.3166
R464 avdd.n313 avdd.t382 27.3166
R465 avdd.n312 avdd.t383 27.3166
R466 avdd.n1 avdd.t404 27.3166
R467 avdd.n0 avdd.t407 27.3166
R468 avdd.n421 avdd.t389 27.1302
R469 avdd.n420 avdd.t396 27.1302
R470 avdd.n128 avdd.t402 27.1302
R471 avdd.n127 avdd.t381 27.1302
R472 avdd.n201 avdd.t384 27.1302
R473 avdd.n200 avdd.t394 27.1302
R474 avdd.n274 avdd.t398 27.1302
R475 avdd.n273 avdd.t380 27.1302
R476 avdd.n347 avdd.t405 27.1302
R477 avdd.n346 avdd.t385 27.1302
R478 avdd.n461 avdd.t393 27.1302
R479 avdd.n460 avdd.t406 27.1302
R480 avdd.n419 avdd.t401 26.9438
R481 avdd.n126 avdd.t387 26.9438
R482 avdd.n199 avdd.t379 26.9438
R483 avdd.n272 avdd.t392 26.9438
R484 avdd.n345 avdd.t397 26.9438
R485 avdd.n459 avdd.t395 26.9438
R486 avdd.n429 dffrs_1.resetb 18.2415
R487 avdd.n136 dffrs_5.resetb 18.2415
R488 avdd.n209 dffrs_4.resetb 18.2415
R489 avdd.n282 dffrs_3.resetb 18.2415
R490 avdd.n355 dffrs_2.resetb 18.2415
R491 avdd.n469 dffrs_0.resetb 18.2415
R492 avdd.n394 avdd.n388 18.0418
R493 avdd.n102 avdd.n96 18.0418
R494 avdd.n175 avdd.n169 18.0418
R495 avdd.n248 avdd.n242 18.0418
R496 avdd.n321 avdd.n315 18.0418
R497 avdd.n534 avdd.n533 18.0418
R498 avdd.n422 avdd.n420 17.6364
R499 avdd.n129 avdd.n127 17.6364
R500 avdd.n202 avdd.n200 17.6364
R501 avdd.n275 avdd.n273 17.6364
R502 avdd.n348 avdd.n346 17.6364
R503 avdd.n462 avdd.n460 17.6364
R504 avdd.n387 avdd.n385 14.3609
R505 avdd.n95 avdd.n93 14.3609
R506 avdd.n168 avdd.n166 14.3609
R507 avdd.n241 avdd.n239 14.3609
R508 avdd.n314 avdd.n312 14.3609
R509 avdd.n2 avdd.n0 14.3609
R510 avdd.n394 avdd.n393 13.5174
R511 avdd.n102 avdd.n101 13.5174
R512 avdd.n175 avdd.n174 13.5174
R513 avdd.n248 avdd.n247 13.5174
R514 avdd.n321 avdd.n320 13.5174
R515 avdd.n533 avdd.n7 13.5174
R516 avdd.n405 avdd.n404 13.5005
R517 avdd.n405 avdd.n399 13.5005
R518 avdd.n417 avdd.n416 13.5005
R519 avdd.n411 avdd.n410 13.5005
R520 avdd.n429 avdd.n428 13.5005
R521 avdd.n113 avdd.n112 13.5005
R522 avdd.n113 avdd.n107 13.5005
R523 avdd.n125 avdd.n124 13.5005
R524 avdd.n119 avdd.n118 13.5005
R525 avdd.n136 avdd.n135 13.5005
R526 avdd.n186 avdd.n185 13.5005
R527 avdd.n186 avdd.n180 13.5005
R528 avdd.n198 avdd.n197 13.5005
R529 avdd.n192 avdd.n191 13.5005
R530 avdd.n209 avdd.n208 13.5005
R531 avdd.n259 avdd.n258 13.5005
R532 avdd.n259 avdd.n253 13.5005
R533 avdd.n271 avdd.n270 13.5005
R534 avdd.n265 avdd.n264 13.5005
R535 avdd.n282 avdd.n281 13.5005
R536 avdd.n332 avdd.n331 13.5005
R537 avdd.n332 avdd.n326 13.5005
R538 avdd.n344 avdd.n343 13.5005
R539 avdd.n338 avdd.n337 13.5005
R540 avdd.n355 avdd.n354 13.5005
R541 avdd.n532 avdd.n531 13.5005
R542 avdd.n532 avdd.n12 13.5005
R543 avdd.n520 avdd.n519 13.5005
R544 avdd.n526 avdd.n525 13.5005
R545 avdd.n469 avdd.n468 13.5005
R546 avdd.n423 avdd.n419 13.4839
R547 avdd.n130 avdd.n126 13.4839
R548 avdd.n203 avdd.n199 13.4839
R549 avdd.n276 avdd.n272 13.4839
R550 avdd.n349 avdd.n345 13.4839
R551 avdd.n463 avdd.n459 13.4839
R552 avdd.n422 avdd.n421 10.5752
R553 avdd.n129 avdd.n128 10.5752
R554 avdd.n202 avdd.n201 10.5752
R555 avdd.n275 avdd.n274 10.5752
R556 avdd.n348 avdd.n347 10.5752
R557 avdd.n462 avdd.n461 10.5752
R558 avdd.n393 avdd.n390 6.4802
R559 avdd.n404 avdd.n401 6.4802
R560 avdd.n399 avdd.n396 6.4802
R561 avdd.n416 avdd.n413 6.4802
R562 avdd.n410 avdd.n407 6.4802
R563 avdd.n428 avdd.n425 6.4802
R564 avdd.n101 avdd.n98 6.4802
R565 avdd.n112 avdd.n109 6.4802
R566 avdd.n107 avdd.n104 6.4802
R567 avdd.n124 avdd.n121 6.4802
R568 avdd.n118 avdd.n115 6.4802
R569 avdd.n135 avdd.n132 6.4802
R570 avdd.n174 avdd.n171 6.4802
R571 avdd.n185 avdd.n182 6.4802
R572 avdd.n180 avdd.n177 6.4802
R573 avdd.n197 avdd.n194 6.4802
R574 avdd.n191 avdd.n188 6.4802
R575 avdd.n208 avdd.n205 6.4802
R576 avdd.n247 avdd.n244 6.4802
R577 avdd.n258 avdd.n255 6.4802
R578 avdd.n253 avdd.n250 6.4802
R579 avdd.n270 avdd.n267 6.4802
R580 avdd.n264 avdd.n261 6.4802
R581 avdd.n281 avdd.n278 6.4802
R582 avdd.n320 avdd.n317 6.4802
R583 avdd.n331 avdd.n328 6.4802
R584 avdd.n326 avdd.n323 6.4802
R585 avdd.n343 avdd.n340 6.4802
R586 avdd.n337 avdd.n334 6.4802
R587 avdd.n354 avdd.n351 6.4802
R588 avdd.n7 avdd.n4 6.4802
R589 avdd.n531 avdd.n528 6.4802
R590 avdd.n12 avdd.n9 6.4802
R591 avdd.n519 avdd.n516 6.4802
R592 avdd.n525 avdd.n522 6.4802
R593 avdd.n468 avdd.n465 6.4802
R594 avdd.n393 avdd.n389 6.25878
R595 avdd.n404 avdd.n400 6.25878
R596 avdd.n399 avdd.n395 6.25878
R597 avdd.n416 avdd.n412 6.25878
R598 avdd.n410 avdd.n406 6.25878
R599 avdd.n428 avdd.n424 6.25878
R600 avdd.n101 avdd.n97 6.25878
R601 avdd.n112 avdd.n108 6.25878
R602 avdd.n107 avdd.n103 6.25878
R603 avdd.n124 avdd.n120 6.25878
R604 avdd.n118 avdd.n114 6.25878
R605 avdd.n135 avdd.n131 6.25878
R606 avdd.n174 avdd.n170 6.25878
R607 avdd.n185 avdd.n181 6.25878
R608 avdd.n180 avdd.n176 6.25878
R609 avdd.n197 avdd.n193 6.25878
R610 avdd.n191 avdd.n187 6.25878
R611 avdd.n208 avdd.n204 6.25878
R612 avdd.n247 avdd.n243 6.25878
R613 avdd.n258 avdd.n254 6.25878
R614 avdd.n253 avdd.n249 6.25878
R615 avdd.n270 avdd.n266 6.25878
R616 avdd.n264 avdd.n260 6.25878
R617 avdd.n281 avdd.n277 6.25878
R618 avdd.n320 avdd.n316 6.25878
R619 avdd.n331 avdd.n327 6.25878
R620 avdd.n326 avdd.n322 6.25878
R621 avdd.n343 avdd.n339 6.25878
R622 avdd.n337 avdd.n333 6.25878
R623 avdd.n354 avdd.n350 6.25878
R624 avdd.n7 avdd.n3 6.25878
R625 avdd.n531 avdd.n527 6.25878
R626 avdd.n12 avdd.n8 6.25878
R627 avdd.n519 avdd.n515 6.25878
R628 avdd.n525 avdd.n521 6.25878
R629 avdd.n468 avdd.n464 6.25878
R630 avdd.n423 avdd.n422 5.93546
R631 avdd.n130 avdd.n129 5.93546
R632 avdd.n203 avdd.n202 5.93546
R633 avdd.n276 avdd.n275 5.93546
R634 avdd.n349 avdd.n348 5.93546
R635 avdd.n463 avdd.n462 5.93546
R636 avdd.n393 avdd.n392 5.44497
R637 avdd.n404 avdd.n403 5.44497
R638 avdd.n399 avdd.n398 5.44497
R639 avdd.n416 avdd.n415 5.44497
R640 avdd.n410 avdd.n409 5.44497
R641 avdd.n428 avdd.n427 5.44497
R642 avdd.n101 avdd.n100 5.44497
R643 avdd.n112 avdd.n111 5.44497
R644 avdd.n107 avdd.n106 5.44497
R645 avdd.n124 avdd.n123 5.44497
R646 avdd.n118 avdd.n117 5.44497
R647 avdd.n135 avdd.n134 5.44497
R648 avdd.n174 avdd.n173 5.44497
R649 avdd.n185 avdd.n184 5.44497
R650 avdd.n180 avdd.n179 5.44497
R651 avdd.n197 avdd.n196 5.44497
R652 avdd.n191 avdd.n190 5.44497
R653 avdd.n208 avdd.n207 5.44497
R654 avdd.n247 avdd.n246 5.44497
R655 avdd.n258 avdd.n257 5.44497
R656 avdd.n253 avdd.n252 5.44497
R657 avdd.n270 avdd.n269 5.44497
R658 avdd.n264 avdd.n263 5.44497
R659 avdd.n281 avdd.n280 5.44497
R660 avdd.n320 avdd.n319 5.44497
R661 avdd.n331 avdd.n330 5.44497
R662 avdd.n326 avdd.n325 5.44497
R663 avdd.n343 avdd.n342 5.44497
R664 avdd.n337 avdd.n336 5.44497
R665 avdd.n354 avdd.n353 5.44497
R666 avdd.n7 avdd.n6 5.44497
R667 avdd.n531 avdd.n530 5.44497
R668 avdd.n12 avdd.n11 5.44497
R669 avdd.n519 avdd.n518 5.44497
R670 avdd.n525 avdd.n524 5.44497
R671 avdd.n468 avdd.n467 5.44497
R672 avdd.n387 avdd.n386 5.14711
R673 avdd.n95 avdd.n94 5.14711
R674 avdd.n168 avdd.n167 5.14711
R675 avdd.n241 avdd.n240 5.14711
R676 avdd.n314 avdd.n313 5.14711
R677 avdd.n2 avdd.n1 5.14711
R678 avdd.n511 avdd.n510 2.49936
R679 avdd.n445 avdd.n444 2.49936
R680 avdd.n371 avdd.n370 2.49936
R681 avdd.n298 avdd.n297 2.49936
R682 avdd.n225 avdd.n224 2.49936
R683 avdd.n152 avdd.n151 2.49936
R684 avdd.n510 avdd.n499 1.93883
R685 avdd.n444 avdd.n433 1.93883
R686 avdd.n370 avdd.n359 1.93883
R687 avdd.n297 avdd.n286 1.93883
R688 avdd.n224 avdd.n213 1.93883
R689 avdd.n151 avdd.n140 1.93883
R690 avdd.n392 avdd.t93 1.85637
R691 avdd.n403 avdd.t299 1.85637
R692 avdd.n398 avdd.t90 1.85637
R693 avdd.n415 avdd.t265 1.85637
R694 avdd.n409 avdd.t19 1.85637
R695 avdd.n427 avdd.t287 1.85637
R696 avdd.n100 avdd.t144 1.85637
R697 avdd.n111 avdd.t293 1.85637
R698 avdd.n106 avdd.t138 1.85637
R699 avdd.n123 avdd.t231 1.85637
R700 avdd.n117 avdd.t177 1.85637
R701 avdd.n134 avdd.t41 1.85637
R702 avdd.n173 avdd.t120 1.85637
R703 avdd.n184 avdd.t319 1.85637
R704 avdd.n179 avdd.t81 1.85637
R705 avdd.n196 avdd.t193 1.85637
R706 avdd.n190 avdd.t305 1.85637
R707 avdd.n207 avdd.t281 1.85637
R708 avdd.n246 avdd.t84 1.85637
R709 avdd.n257 avdd.t247 1.85637
R710 avdd.n252 avdd.t150 1.85637
R711 avdd.n269 avdd.t63 1.85637
R712 avdd.n263 avdd.t279 1.85637
R713 avdd.n280 avdd.t217 1.85637
R714 avdd.n319 avdd.t105 1.85637
R715 avdd.n330 avdd.t245 1.85637
R716 avdd.n325 avdd.t108 1.85637
R717 avdd.n342 avdd.t325 1.85637
R718 avdd.n336 avdd.t311 1.85637
R719 avdd.n353 avdd.t365 1.85637
R720 avdd.n6 avdd.t132 1.85637
R721 avdd.n530 avdd.t187 1.85637
R722 avdd.n11 avdd.t126 1.85637
R723 avdd.n518 avdd.t329 1.85637
R724 avdd.n524 avdd.t369 1.85637
R725 avdd.n467 avdd.t51 1.85637
R726 avdd.n138 avdd.n92 1.80479
R727 avdd.n211 avdd.n76 1.80479
R728 avdd.n284 avdd.n60 1.80479
R729 avdd.n357 avdd.n44 1.80479
R730 avdd.n431 avdd.n28 1.80479
R731 avdd.n513 avdd.n470 1.80479
R732 avdd.n161 avdd.n160 1.78583
R733 avdd.n234 avdd.n233 1.78583
R734 avdd.n307 avdd.n306 1.78583
R735 avdd.n380 avdd.n379 1.78583
R736 avdd.n454 avdd.n453 1.78583
R737 avdd.n496 avdd.n495 1.78583
R738 avdd.n164 avdd.t71 1.74654
R739 avdd.n237 avdd.t73 1.74654
R740 avdd.n310 avdd.t69 1.74654
R741 avdd.n383 avdd.t171 1.74654
R742 avdd.n457 avdd.t271 1.74654
R743 avdd.n487 avdd.t173 1.74654
R744 avdd.n486 avdd.t55 1.49467
R745 avdd.n507 avdd.t49 1.49467
R746 avdd.n506 avdd.t75 1.49467
R747 avdd.n14 avdd.t357 1.49467
R748 avdd.n441 avdd.t327 1.49467
R749 avdd.n440 avdd.t219 1.49467
R750 avdd.n30 avdd.t43 1.49467
R751 avdd.n367 avdd.t67 1.49467
R752 avdd.n366 avdd.t221 1.49467
R753 avdd.n46 avdd.t313 1.49467
R754 avdd.n294 avdd.t17 1.49467
R755 avdd.n293 avdd.t47 1.49467
R756 avdd.n62 avdd.t277 1.49467
R757 avdd.n221 avdd.t37 1.49467
R758 avdd.n220 avdd.t233 1.49467
R759 avdd.n78 avdd.t185 1.49467
R760 avdd.n148 avdd.t359 1.49467
R761 avdd.n147 avdd.t3 1.49467
R762 avdd.n77 avdd.t213 1.49467
R763 avdd.n61 avdd.t169 1.49467
R764 avdd.n45 avdd.t269 1.49467
R765 avdd.n29 avdd.t191 1.49467
R766 avdd.n13 avdd.t45 1.49467
R767 avdd.n490 avdd.t175 1.49467
R768 avdd.n500 avdd.t211 1.47383
R769 avdd.n434 avdd.t223 1.47383
R770 avdd.n360 avdd.t237 1.47383
R771 avdd.n287 avdd.t57 1.47383
R772 avdd.n214 avdd.t255 1.47383
R773 avdd.n141 avdd.t259 1.47383
R774 avdd.n80 avdd.t183 1.47383
R775 avdd.n81 avdd.t181 1.47383
R776 avdd.n82 avdd.t215 1.47383
R777 avdd.n79 avdd.t337 1.47383
R778 avdd.n64 avdd.t31 1.47383
R779 avdd.n65 avdd.t29 1.47383
R780 avdd.n66 avdd.t239 1.47383
R781 avdd.n63 avdd.t355 1.47383
R782 avdd.n48 avdd.t203 1.47383
R783 avdd.n49 avdd.t205 1.47383
R784 avdd.n50 avdd.t295 1.47383
R785 avdd.n47 avdd.t201 1.47383
R786 avdd.n32 avdd.t275 1.47383
R787 avdd.n33 avdd.t273 1.47383
R788 avdd.n34 avdd.t167 1.47383
R789 avdd.n31 avdd.t261 1.47383
R790 avdd.n16 avdd.t33 1.47383
R791 avdd.n17 avdd.t35 1.47383
R792 avdd.n18 avdd.t367 1.47383
R793 avdd.n15 avdd.t307 1.47383
R794 avdd.n482 avdd.t375 1.47383
R795 avdd.n472 avdd.t377 1.47383
R796 avdd.n471 avdd.t235 1.47383
R797 avdd.n492 avdd.t189 1.47383
R798 avdd.n210 avdd.n165 1.19311
R799 avdd.n283 avdd.n238 1.19311
R800 avdd.n356 avdd.n311 1.19311
R801 avdd.n418 avdd.n384 1.19311
R802 avdd.n514 avdd.n458 1.19311
R803 avdd.n392 avdd.n391 1.04105
R804 avdd.n403 avdd.n402 1.04105
R805 avdd.n398 avdd.n397 1.04105
R806 avdd.n415 avdd.n414 1.04105
R807 avdd.n409 avdd.n408 1.04105
R808 avdd.n427 avdd.n426 1.04105
R809 avdd.n100 avdd.n99 1.04105
R810 avdd.n111 avdd.n110 1.04105
R811 avdd.n106 avdd.n105 1.04105
R812 avdd.n123 avdd.n122 1.04105
R813 avdd.n117 avdd.n116 1.04105
R814 avdd.n134 avdd.n133 1.04105
R815 avdd.n173 avdd.n172 1.04105
R816 avdd.n184 avdd.n183 1.04105
R817 avdd.n179 avdd.n178 1.04105
R818 avdd.n196 avdd.n195 1.04105
R819 avdd.n190 avdd.n189 1.04105
R820 avdd.n207 avdd.n206 1.04105
R821 avdd.n246 avdd.n245 1.04105
R822 avdd.n257 avdd.n256 1.04105
R823 avdd.n252 avdd.n251 1.04105
R824 avdd.n269 avdd.n268 1.04105
R825 avdd.n263 avdd.n262 1.04105
R826 avdd.n280 avdd.n279 1.04105
R827 avdd.n319 avdd.n318 1.04105
R828 avdd.n330 avdd.n329 1.04105
R829 avdd.n325 avdd.n324 1.04105
R830 avdd.n342 avdd.n341 1.04105
R831 avdd.n336 avdd.n335 1.04105
R832 avdd.n353 avdd.n352 1.04105
R833 avdd.n6 avdd.n5 1.04105
R834 avdd.n530 avdd.n529 1.04105
R835 avdd.n11 avdd.n10 1.04105
R836 avdd.n518 avdd.n517 1.04105
R837 avdd.n524 avdd.n523 1.04105
R838 avdd.n467 avdd.n466 1.04105
R839 avdd.n138 avdd.n137 0.809622
R840 avdd.n211 avdd.n210 0.809622
R841 avdd.n284 avdd.n283 0.809622
R842 avdd.n357 avdd.n356 0.809622
R843 avdd.n431 avdd.n430 0.809622
R844 avdd.n514 avdd.n513 0.809622
R845 avdd.n503 avdd.n500 0.788
R846 avdd.n504 avdd.n503 0.788
R847 avdd.n506 avdd.n505 0.788
R848 avdd.n437 avdd.n434 0.788
R849 avdd.n438 avdd.n437 0.788
R850 avdd.n440 avdd.n439 0.788
R851 avdd.n363 avdd.n360 0.788
R852 avdd.n364 avdd.n363 0.788
R853 avdd.n366 avdd.n365 0.788
R854 avdd.n290 avdd.n287 0.788
R855 avdd.n291 avdd.n290 0.788
R856 avdd.n293 avdd.n292 0.788
R857 avdd.n217 avdd.n214 0.788
R858 avdd.n218 avdd.n217 0.788
R859 avdd.n220 avdd.n219 0.788
R860 avdd.n144 avdd.n141 0.788
R861 avdd.n145 avdd.n144 0.788
R862 avdd.n147 avdd.n146 0.788
R863 avdd.n88 avdd.n81 0.788
R864 avdd.n89 avdd.n88 0.788
R865 avdd.n90 avdd.n82 0.788
R866 avdd.n91 avdd.n90 0.788
R867 avdd.n86 avdd.n80 0.788
R868 avdd.n158 avdd.n79 0.788
R869 avdd.n159 avdd.n158 0.788
R870 avdd.n157 avdd.n77 0.788
R871 avdd.n72 avdd.n65 0.788
R872 avdd.n73 avdd.n72 0.788
R873 avdd.n74 avdd.n66 0.788
R874 avdd.n75 avdd.n74 0.788
R875 avdd.n70 avdd.n64 0.788
R876 avdd.n231 avdd.n63 0.788
R877 avdd.n232 avdd.n231 0.788
R878 avdd.n230 avdd.n61 0.788
R879 avdd.n56 avdd.n49 0.788
R880 avdd.n57 avdd.n56 0.788
R881 avdd.n58 avdd.n50 0.788
R882 avdd.n59 avdd.n58 0.788
R883 avdd.n54 avdd.n48 0.788
R884 avdd.n304 avdd.n47 0.788
R885 avdd.n305 avdd.n304 0.788
R886 avdd.n303 avdd.n45 0.788
R887 avdd.n40 avdd.n33 0.788
R888 avdd.n41 avdd.n40 0.788
R889 avdd.n42 avdd.n34 0.788
R890 avdd.n43 avdd.n42 0.788
R891 avdd.n38 avdd.n32 0.788
R892 avdd.n377 avdd.n31 0.788
R893 avdd.n378 avdd.n377 0.788
R894 avdd.n376 avdd.n29 0.788
R895 avdd.n24 avdd.n17 0.788
R896 avdd.n25 avdd.n24 0.788
R897 avdd.n26 avdd.n18 0.788
R898 avdd.n27 avdd.n26 0.788
R899 avdd.n22 avdd.n16 0.788
R900 avdd.n451 avdd.n15 0.788
R901 avdd.n452 avdd.n451 0.788
R902 avdd.n450 avdd.n13 0.788
R903 avdd.n479 avdd.n472 0.788
R904 avdd.n480 avdd.n479 0.788
R905 avdd.n477 avdd.n471 0.788
R906 avdd.n478 avdd.n477 0.788
R907 avdd.n482 avdd.n481 0.788
R908 avdd.n493 avdd.n492 0.788
R909 avdd.n494 avdd.n493 0.788
R910 avdd.n491 avdd.n490 0.788
R911 avdd.n388 avdd.n387 0.754571
R912 avdd.n96 avdd.n95 0.754571
R913 avdd.n169 avdd.n168 0.754571
R914 avdd.n242 avdd.n241 0.754571
R915 avdd.n315 avdd.n314 0.754571
R916 avdd.n534 avdd.n2 0.754571
R917 avdd.n389 avdd.t267 0.7285
R918 avdd.n389 avdd.t243 0.7285
R919 avdd.n400 avdd.t25 0.7285
R920 avdd.n400 avdd.t156 0.7285
R921 avdd.n395 avdd.t199 0.7285
R922 avdd.n395 avdd.t263 0.7285
R923 avdd.n412 avdd.t241 0.7285
R924 avdd.n412 avdd.t349 0.7285
R925 avdd.n406 avdd.t141 0.7285
R926 avdd.n406 avdd.t285 0.7285
R927 avdd.n424 avdd.t249 0.7285
R928 avdd.n424 avdd.t87 0.7285
R929 avdd.n97 avdd.t229 0.7285
R930 avdd.n97 avdd.t291 0.7285
R931 avdd.n108 avdd.t339 0.7285
R932 avdd.n108 avdd.t111 0.7285
R933 avdd.n103 avdd.t335 0.7285
R934 avdd.n103 avdd.t227 0.7285
R935 avdd.n120 avdd.t251 0.7285
R936 avdd.n120 avdd.t9 0.7285
R937 avdd.n114 avdd.t96 0.7285
R938 avdd.n114 avdd.t39 0.7285
R939 avdd.n131 avdd.t309 0.7285
R940 avdd.n131 avdd.t135 0.7285
R941 avdd.n170 avdd.t197 0.7285
R942 avdd.n170 avdd.t289 0.7285
R943 avdd.n181 avdd.t345 0.7285
R944 avdd.n181 avdd.t165 0.7285
R945 avdd.n176 avdd.t353 0.7285
R946 avdd.n176 avdd.t195 0.7285
R947 avdd.n193 avdd.t257 0.7285
R948 avdd.n193 avdd.t347 0.7285
R949 avdd.n187 avdd.t117 0.7285
R950 avdd.n187 avdd.t283 0.7285
R951 avdd.n204 avdd.t253 0.7285
R952 avdd.n204 avdd.t99 0.7285
R953 avdd.n243 avdd.t65 0.7285
R954 avdd.n243 avdd.t303 0.7285
R955 avdd.n254 avdd.t351 0.7285
R956 avdd.n254 avdd.t114 0.7285
R957 avdd.n249 avdd.t61 0.7285
R958 avdd.n249 avdd.t361 0.7285
R959 avdd.n266 avdd.t301 0.7285
R960 avdd.n266 avdd.t7 0.7285
R961 avdd.n260 avdd.t78 0.7285
R962 avdd.n260 avdd.t225 0.7285
R963 avdd.n277 avdd.t297 0.7285
R964 avdd.n277 avdd.t147 0.7285
R965 avdd.n316 avdd.t323 0.7285
R966 avdd.n316 avdd.t209 0.7285
R967 avdd.n327 avdd.t27 0.7285
R968 avdd.n327 avdd.t102 0.7285
R969 avdd.n322 avdd.t15 0.7285
R970 avdd.n322 avdd.t321 0.7285
R971 avdd.n339 avdd.t207 0.7285
R972 avdd.n339 avdd.t23 0.7285
R973 avdd.n333 avdd.t153 0.7285
R974 avdd.n333 avdd.t363 0.7285
R975 avdd.n350 avdd.t179 0.7285
R976 avdd.n350 avdd.t123 0.7285
R977 avdd.n3 avdd.t333 0.7285
R978 avdd.n3 avdd.t21 0.7285
R979 avdd.n527 avdd.t341 0.7285
R980 avdd.n527 avdd.t129 0.7285
R981 avdd.n8 avdd.t13 0.7285
R982 avdd.n8 avdd.t331 0.7285
R983 avdd.n515 avdd.t5 0.7285
R984 avdd.n515 avdd.t343 0.7285
R985 avdd.n521 avdd.t159 0.7285
R986 avdd.n521 avdd.t53 0.7285
R987 avdd.n464 avdd.t371 0.7285
R988 avdd.n464 avdd.t162 0.7285
R989 avdd.n509 avdd.n500 0.561043
R990 avdd.n443 avdd.n434 0.561043
R991 avdd.n369 avdd.n360 0.561043
R992 avdd.n296 avdd.n287 0.561043
R993 avdd.n223 avdd.n214 0.561043
R994 avdd.n150 avdd.n141 0.561043
R995 avdd.n154 avdd.n80 0.561043
R996 avdd.n153 avdd.n81 0.561043
R997 avdd.n139 avdd.n82 0.561043
R998 avdd.n162 avdd.n79 0.561043
R999 avdd.n227 avdd.n64 0.561043
R1000 avdd.n226 avdd.n65 0.561043
R1001 avdd.n212 avdd.n66 0.561043
R1002 avdd.n235 avdd.n63 0.561043
R1003 avdd.n300 avdd.n48 0.561043
R1004 avdd.n299 avdd.n49 0.561043
R1005 avdd.n285 avdd.n50 0.561043
R1006 avdd.n308 avdd.n47 0.561043
R1007 avdd.n373 avdd.n32 0.561043
R1008 avdd.n372 avdd.n33 0.561043
R1009 avdd.n358 avdd.n34 0.561043
R1010 avdd.n381 avdd.n31 0.561043
R1011 avdd.n447 avdd.n16 0.561043
R1012 avdd.n446 avdd.n17 0.561043
R1013 avdd.n432 avdd.n18 0.561043
R1014 avdd.n455 avdd.n15 0.561043
R1015 avdd.n497 avdd.n482 0.561043
R1016 avdd.n498 avdd.n472 0.561043
R1017 avdd.n512 avdd.n471 0.561043
R1018 avdd.n492 avdd.n483 0.561043
R1019 avdd.n488 avdd.n487 0.510024
R1020 avdd.n165 avdd.n163 0.490037
R1021 avdd.n238 avdd.n236 0.490037
R1022 avdd.n311 avdd.n309 0.490037
R1023 avdd.n384 avdd.n382 0.490037
R1024 avdd.n458 avdd.n456 0.490037
R1025 avdd.n165 avdd.n164 0.436534
R1026 avdd.n238 avdd.n237 0.436534
R1027 avdd.n311 avdd.n310 0.436534
R1028 avdd.n384 avdd.n383 0.436534
R1029 avdd.n458 avdd.n457 0.436534
R1030 avdd.n489 avdd.n488 0.415037
R1031 avdd.n509 avdd.n508 0.255737
R1032 avdd.n443 avdd.n442 0.255737
R1033 avdd.n369 avdd.n368 0.255737
R1034 avdd.n296 avdd.n295 0.255737
R1035 avdd.n223 avdd.n222 0.255737
R1036 avdd.n150 avdd.n149 0.255737
R1037 avdd.n163 avdd.n162 0.255737
R1038 avdd.n236 avdd.n235 0.255737
R1039 avdd.n309 avdd.n308 0.255737
R1040 avdd.n382 avdd.n381 0.255737
R1041 avdd.n456 avdd.n455 0.255737
R1042 avdd.n489 avdd.n483 0.255737
R1043 avdd.n162 avdd.n161 0.2165
R1044 avdd.n235 avdd.n234 0.2165
R1045 avdd.n308 avdd.n307 0.2165
R1046 avdd.n381 avdd.n380 0.2165
R1047 avdd.n455 avdd.n454 0.2165
R1048 avdd.n496 avdd.n483 0.2165
R1049 avdd.n161 avdd.n154 0.148424
R1050 avdd.n234 avdd.n227 0.148424
R1051 avdd.n307 avdd.n300 0.148424
R1052 avdd.n380 avdd.n373 0.148424
R1053 avdd.n454 avdd.n447 0.148424
R1054 avdd.n497 avdd.n496 0.148424
R1055 dffrs_1.resetb avdd.n423 0.136036
R1056 dffrs_5.resetb avdd.n130 0.136036
R1057 dffrs_4.resetb avdd.n203 0.136036
R1058 dffrs_3.resetb avdd.n276 0.136036
R1059 dffrs_2.resetb avdd.n349 0.136036
R1060 dffrs_0.resetb avdd.n463 0.136036
R1061 avdd.n510 avdd.n509 0.0635
R1062 avdd.n444 avdd.n443 0.0635
R1063 avdd.n370 avdd.n369 0.0635
R1064 avdd.n297 avdd.n296 0.0635
R1065 avdd.n224 avdd.n223 0.0635
R1066 avdd.n151 avdd.n150 0.0635
R1067 avdd.n154 avdd.n153 0.0452384
R1068 avdd.n227 avdd.n226 0.0452384
R1069 avdd.n300 avdd.n299 0.0452384
R1070 avdd.n373 avdd.n372 0.0452384
R1071 avdd.n447 avdd.n446 0.0452384
R1072 avdd.n498 avdd.n497 0.0452384
R1073 avdd.n119 avdd.n113 0.0405727
R1074 avdd.n192 avdd.n186 0.0405727
R1075 avdd.n265 avdd.n259 0.0405727
R1076 avdd.n338 avdd.n332 0.0405727
R1077 avdd.n411 avdd.n405 0.0405727
R1078 avdd.n532 avdd.n526 0.0405727
R1079 avdd.n388 dffrs_1.setb 0.032
R1080 avdd.n96 dffrs_5.setb 0.032
R1081 avdd.n169 dffrs_4.setb 0.032
R1082 avdd.n242 dffrs_3.setb 0.032
R1083 avdd.n315 dffrs_2.setb 0.032
R1084 dffrs_0.setb avdd.n534 0.032
R1085 avdd.n508 avdd.n506 0.0313054
R1086 avdd.n508 avdd.n507 0.0313054
R1087 avdd.n442 avdd.n440 0.0313054
R1088 avdd.n442 avdd.n441 0.0313054
R1089 avdd.n368 avdd.n366 0.0313054
R1090 avdd.n368 avdd.n367 0.0313054
R1091 avdd.n295 avdd.n293 0.0313054
R1092 avdd.n295 avdd.n294 0.0313054
R1093 avdd.n222 avdd.n220 0.0313054
R1094 avdd.n222 avdd.n221 0.0313054
R1095 avdd.n149 avdd.n147 0.0313054
R1096 avdd.n149 avdd.n148 0.0313054
R1097 avdd.n163 avdd.n77 0.0313054
R1098 avdd.n163 avdd.n78 0.0313054
R1099 avdd.n236 avdd.n61 0.0313054
R1100 avdd.n236 avdd.n62 0.0313054
R1101 avdd.n309 avdd.n45 0.0313054
R1102 avdd.n309 avdd.n46 0.0313054
R1103 avdd.n382 avdd.n29 0.0313054
R1104 avdd.n382 avdd.n30 0.0313054
R1105 avdd.n456 avdd.n13 0.0313054
R1106 avdd.n456 avdd.n14 0.0313054
R1107 avdd.n490 avdd.n489 0.0313054
R1108 avdd.n489 avdd.n486 0.0313054
R1109 avdd.n152 avdd.n139 0.0295407
R1110 avdd.n225 avdd.n212 0.0295407
R1111 avdd.n298 avdd.n285 0.0295407
R1112 avdd.n371 avdd.n358 0.0295407
R1113 avdd.n445 avdd.n432 0.0295407
R1114 avdd.n512 avdd.n511 0.0295407
R1115 avdd.n137 avdd.n125 0.0288636
R1116 avdd.n210 avdd.n198 0.0288636
R1117 avdd.n283 avdd.n271 0.0288636
R1118 avdd.n356 avdd.n344 0.0288636
R1119 avdd.n520 avdd.n514 0.0288636
R1120 avdd.n418 avdd.n417 0.0288455
R1121 avdd.n113 avdd.n102 0.0237
R1122 avdd.n186 avdd.n175 0.0237
R1123 avdd.n259 avdd.n248 0.0237
R1124 avdd.n332 avdd.n321 0.0237
R1125 avdd.n405 avdd.n394 0.0237
R1126 avdd.n533 avdd.n532 0.0237
R1127 avdd.n153 avdd.n152 0.0161977
R1128 avdd.n226 avdd.n225 0.0161977
R1129 avdd.n299 avdd.n298 0.0161977
R1130 avdd.n372 avdd.n371 0.0161977
R1131 avdd.n446 avdd.n445 0.0161977
R1132 avdd.n511 avdd.n498 0.0161977
R1133 avdd.n139 avdd.n138 0.0129273
R1134 avdd.n212 avdd.n211 0.0129273
R1135 avdd.n285 avdd.n284 0.0129273
R1136 avdd.n358 avdd.n357 0.0129273
R1137 avdd.n432 avdd.n431 0.0129273
R1138 avdd.n513 avdd.n512 0.0129273
R1139 avdd.n488 avdd 0.0128676
R1140 avdd.n137 avdd.n136 0.0122273
R1141 avdd.n210 avdd.n209 0.0122273
R1142 avdd.n283 avdd.n282 0.0122273
R1143 avdd.n356 avdd.n355 0.0122273
R1144 avdd.n430 avdd.n429 0.0122273
R1145 avdd.n514 avdd.n469 0.0122273
R1146 avdd.n125 avdd.n119 0.000518182
R1147 avdd.n198 avdd.n192 0.000518182
R1148 avdd.n271 avdd.n265 0.000518182
R1149 avdd.n344 avdd.n338 0.000518182
R1150 avdd.n417 avdd.n411 0.000518182
R1151 avdd.n430 avdd.n418 0.000518182
R1152 avdd.n526 avdd.n520 0.000518182
R1153 avss.n259 avss.n258 21124.8
R1154 avss.n216 avss.n215 21124.8
R1155 avss.n173 avss.n172 21124.8
R1156 avss.n124 avss.n51 21034.5
R1157 avss.n787 avss.n786 21034.5
R1158 avss.n321 avss.n301 21026.3
R1159 avss.n374 avss.n373 21012.5
R1160 avss.n474 avss.n473 21012.5
R1161 avss.n574 avss.n573 21012.5
R1162 avss.n674 avss.n673 21012.5
R1163 avss.n757 avss.n756 21000
R1164 avss.n825 avss.n824 21000
R1165 avss.n381 avss.n267 16221.9
R1166 avss.n481 avss.n224 16221.9
R1167 avss.n581 avss.n181 16221.9
R1168 avss.n681 avss.n132 16221.9
R1169 avss.n785 avss.n53 16221.9
R1170 avss.n836 avss.n833 11510.4
R1171 avss.n382 avss.n381 11510.4
R1172 avss.n482 avss.n481 11510.4
R1173 avss.n582 avss.n581 11510.4
R1174 avss.n682 avss.n681 11510.4
R1175 avss.n764 avss.n53 11510.4
R1176 avss.n836 avss.n6 11510.4
R1177 avss.n826 avss.n825 7422.73
R1178 avss.n758 avss.n757 7422.73
R1179 avss.n373 avss.n372 7422.62
R1180 avss.n473 avss.n472 7422.62
R1181 avss.n573 avss.n572 7422.62
R1182 avss.n673 avss.n672 7422.62
R1183 avss.n423 avss.n422 6961.73
R1184 avss.n523 avss.n522 6961.73
R1185 avss.n623 avss.n622 6961.73
R1186 avss.n716 avss.n715 6961.73
R1187 avss.n55 avss.n50 6961.73
R1188 avss.n854 avss.n5 6190.48
R1189 avss.n781 avss.n81 6190.48
R1190 avss.n699 avss.n139 6190.48
R1191 avss.n606 avss.n182 6190.48
R1192 avss.n506 avss.n225 6190.48
R1193 avss.n406 avss.n268 6190.48
R1194 avss.n323 avss.n322 5557.62
R1195 avss.n323 avss.n291 5551.58
R1196 avss.n423 avss.n250 5551.58
R1197 avss.n523 avss.n207 5551.58
R1198 avss.n623 avss.n164 5551.58
R1199 avss.n716 avss.n116 5551.58
R1200 avss.n55 avss.n42 5551.58
R1201 avss.n408 avss.n249 5290.17
R1202 avss.n508 avss.n206 5290.17
R1203 avss.n608 avss.n163 5290.17
R1204 avss.n701 avss.n115 5286.93
R1205 avss.n783 avss.n41 5286.93
R1206 avss.n854 avss.n853 4683.14
R1207 avss.n300 avss.n299 4273.71
R1208 avss.n409 avss.n408 4062.5
R1209 avss.n509 avss.n508 4062.5
R1210 avss.n609 avss.n608 4062.5
R1211 avss.n702 avss.n701 4062.5
R1212 avss.n784 avss.n783 4062.5
R1213 avss.n322 avss.n300 3568.02
R1214 avss.n854 avss.n6 3123.51
R1215 avss.n374 avss.n284 2944.22
R1216 avss.n474 avss.n241 2944.22
R1217 avss.n574 avss.n198 2944.22
R1218 avss.n674 avss.n155 2944.22
R1219 avss.n756 avss.n750 2944.22
R1220 avss.n824 avss.n822 2944.22
R1221 avss.n267 avss.n258 2845.46
R1222 avss.n224 avss.n215 2845.46
R1223 avss.n181 avss.n172 2845.46
R1224 avss.n786 avss.n785 2845.46
R1225 avss.n132 avss.n124 2843.75
R1226 avss.n325 avss.n283 2257.8
R1227 avss.n425 avss.n240 2257.8
R1228 avss.n525 avss.n197 2257.8
R1229 avss.n625 avss.n154 2257.8
R1230 avss.n97 avss.n52 2257.8
R1231 avss.n789 avss.n23 2257.8
R1232 avss.n702 avss.n132 1878.69
R1233 avss.n409 avss.n267 1876.98
R1234 avss.n509 avss.n224 1876.98
R1235 avss.n609 avss.n181 1876.98
R1236 avss.n785 avss.n784 1876.98
R1237 avss.n347 avss.n346 1486.9
R1238 avss.n309 avss.n300 1212.42
R1239 avss.n422 avss.n258 1205.08
R1240 avss.n522 avss.n215 1205.08
R1241 avss.n622 avss.n172 1205.08
R1242 avss.n715 avss.n124 1205.08
R1243 avss.n786 avss.n50 1205.08
R1244 avss.n301 avss.n267 1135.55
R1245 avss.n259 avss.n224 1135.55
R1246 avss.n216 avss.n181 1135.55
R1247 avss.n173 avss.n132 1135.55
R1248 avss.n785 avss.n51 1135.55
R1249 avss.n788 avss.n787 1135.55
R1250 avss.n325 avss.n267 1122.24
R1251 avss.n425 avss.n224 1122.24
R1252 avss.n525 avss.n181 1122.24
R1253 avss.n625 avss.n132 1122.24
R1254 avss.n785 avss.n52 1122.24
R1255 avss.n789 avss.n788 1122.24
R1256 avss.n739 avss.n738 977.434
R1257 avss.n811 avss.n810 977.434
R1258 avss.n447 avss.n446 977.068
R1259 avss.n547 avss.n546 977.068
R1260 avss.n647 avss.n646 977.068
R1261 avss.n738 avss.n115 904.402
R1262 avss.n810 avss.n41 904.402
R1263 avss.n446 avss.n249 904.062
R1264 avss.n546 avss.n206 904.062
R1265 avss.n646 avss.n163 904.062
R1266 avss.n322 avss.n321 897.806
R1267 avss.n323 avss.n298 832.22
R1268 avss.n423 avss.n257 832.22
R1269 avss.n523 avss.n214 832.22
R1270 avss.n623 avss.n171 832.22
R1271 avss.n716 avss.n123 832.22
R1272 avss.n56 avss.n55 832.22
R1273 avss.n324 avss.n323 832.101
R1274 avss.n424 avss.n423 832.101
R1275 avss.n524 avss.n523 832.101
R1276 avss.n624 avss.n623 832.101
R1277 avss.n717 avss.n716 832.101
R1278 avss.n55 avss.n54 832.101
R1279 avss.n75 avss.n41 784.409
R1280 avss.n133 avss.n115 784.37
R1281 avss.n588 avss.n163 784.37
R1282 avss.n488 avss.n206 784.37
R1283 avss.n388 avss.n249 784.37
R1284 avss.n788 avss.n6 697.039
R1285 avss.n374 avss.n283 665.564
R1286 avss.n474 avss.n240 665.564
R1287 avss.n574 avss.n197 665.564
R1288 avss.n674 avss.n154 665.564
R1289 avss.n756 avss.n97 665.564
R1290 avss.n824 avss.n23 665.564
R1291 avss.n822 avss.n821 654.253
R1292 avss.n750 avss.n749 654.253
R1293 avss.n156 avss.n155 654.005
R1294 avss.n199 avss.n198 654.005
R1295 avss.n242 avss.n241 654.005
R1296 avss.n285 avss.n284 654.005
R1297 avss.n750 avss.n98 648.784
R1298 avss.n822 avss.n24 648.784
R1299 avss.n348 avss.n284 648.54
R1300 avss.n448 avss.n241 648.54
R1301 avss.n548 avss.n198 648.54
R1302 avss.n648 avss.n155 648.54
R1303 avss.t134 avss.n826 590.909
R1304 avss.n827 avss.t134 590.909
R1305 avss.n827 avss.t252 590.909
R1306 avss.n833 avss.t181 590.909
R1307 avss.n833 avss.t35 590.909
R1308 avss.t37 avss.n832 590.909
R1309 avss.t253 avss.n375 590.909
R1310 avss.n379 avss.t253 590.909
R1311 avss.t136 avss.n379 590.909
R1312 avss.n381 avss.t186 590.909
R1313 avss.n381 avss.t179 590.909
R1314 avss.n405 avss.t118 590.909
R1315 avss.t259 avss.n475 590.909
R1316 avss.n479 avss.t259 590.909
R1317 avss.t125 avss.n479 590.909
R1318 avss.n481 avss.t128 590.909
R1319 avss.n481 avss.t155 590.909
R1320 avss.n505 avss.t195 590.909
R1321 avss.t130 avss.n575 590.909
R1322 avss.n579 avss.t130 590.909
R1323 avss.t104 avss.n579 590.909
R1324 avss.n581 avss.t187 590.909
R1325 avss.n581 avss.t44 590.909
R1326 avss.n605 avss.t221 590.909
R1327 avss.t112 avss.n675 590.909
R1328 avss.n679 avss.t112 590.909
R1329 avss.t55 avss.n679 590.909
R1330 avss.n681 avss.t123 590.909
R1331 avss.n681 avss.t16 590.909
R1332 avss.n698 avss.t0 590.909
R1333 avss.t139 avss.n758 590.909
R1334 avss.n762 avss.t139 590.909
R1335 avss.t209 avss.n762 590.909
R1336 avss.n764 avss.t274 590.909
R1337 avss.t234 avss.n764 590.909
R1338 avss.n765 avss.t232 590.909
R1339 avss.n755 avss.t202 590.909
R1340 avss.t202 avss.n754 590.909
R1341 avss.n754 avss.t107 590.909
R1342 avss.t124 avss.n53 590.909
R1343 avss.t275 avss.n53 590.909
R1344 avss.n780 avss.t261 590.909
R1345 avss.n823 avss.t280 590.909
R1346 avss.n837 avss.t280 590.909
R1347 avss.n837 avss.t103 590.909
R1348 avss.t54 avss.n836 590.909
R1349 avss.n836 avss.t215 590.909
R1350 avss.n855 avss.t212 590.909
R1351 avss.n372 avss.t217 590.462
R1352 avss.t217 avss.n371 590.462
R1353 avss.n371 avss.t228 590.462
R1354 avss.n382 avss.t4 590.462
R1355 avss.t265 avss.n382 590.462
R1356 avss.n383 avss.t263 590.462
R1357 avss.n472 avss.t169 590.462
R1358 avss.t169 avss.n471 590.462
R1359 avss.n471 avss.t165 590.462
R1360 avss.n482 avss.t120 590.462
R1361 avss.t27 avss.n482 590.462
R1362 avss.n483 avss.t29 590.462
R1363 avss.n572 avss.t236 590.462
R1364 avss.t236 avss.n571 590.462
R1365 avss.n571 avss.t31 590.462
R1366 avss.n582 avss.t34 590.462
R1367 avss.t10 avss.n582 590.462
R1368 avss.n583 avss.t12 590.462
R1369 avss.n672 avss.t150 590.462
R1370 avss.t150 avss.n671 590.462
R1371 avss.n671 avss.t138 590.462
R1372 avss.n682 avss.t43 590.462
R1373 avss.t50 avss.n682 590.462
R1374 avss.n683 avss.t52 590.462
R1375 avss.n309 avss.t242 582.165
R1376 avss.t65 avss.n298 582.165
R1377 avss.n410 avss.t255 582.165
R1378 avss.t88 avss.n257 582.165
R1379 avss.n510 avss.t48 582.165
R1380 avss.t69 avss.n214 582.165
R1381 avss.n610 avss.t9 582.165
R1382 avss.t92 avss.n171 582.165
R1383 avss.n703 avss.t129 582.165
R1384 avss.t82 avss.n123 582.165
R1385 avss.n74 avss.t8 582.165
R1386 avss.n56 avss.t59 582.165
R1387 avss.t250 avss.n324 581.712
R1388 avss.n326 avss.t198 581.712
R1389 avss.n320 avss.t144 581.712
R1390 avss.n302 avss.t71 581.712
R1391 avss.t248 avss.n424 581.712
R1392 avss.n426 avss.t229 581.712
R1393 avss.n421 avss.t177 581.712
R1394 avss.n260 avss.t99 581.712
R1395 avss.t245 avss.n524 581.712
R1396 avss.n526 avss.t171 581.712
R1397 avss.n521 avss.t269 581.712
R1398 avss.n217 avss.t80 581.712
R1399 avss.t247 avss.n624 581.712
R1400 avss.n626 avss.t160 581.712
R1401 avss.n621 avss.t204 581.712
R1402 avss.n174 avss.t94 581.712
R1403 avss.t22 avss.n717 581.712
R1404 avss.n718 avss.t270 581.712
R1405 avss.n714 avss.t225 581.712
R1406 avss.n125 avss.t85 581.712
R1407 avss.n54 avss.t251 581.712
R1408 avss.n790 avss.t121 581.712
R1409 avss.n60 avss.t238 581.712
R1410 avss.t63 avss.n49 581.712
R1411 avss.t197 avss.n334 581.712
R1412 avss.n335 avss.t145 581.712
R1413 avss.t173 avss.n434 581.712
R1414 avss.n435 avss.t175 581.712
R1415 avss.t152 avss.n534 581.712
R1416 avss.n535 avss.t267 581.712
R1417 avss.t41 avss.n634 581.712
R1418 avss.n635 avss.t206 581.712
R1419 avss.t164 avss.n726 581.712
R1420 avss.n727 avss.t257 581.712
R1421 avss.t18 avss.n798 581.712
R1422 avss.n799 avss.t239 581.712
R1423 avss.n701 avss.n699 574.192
R1424 avss.n408 avss.n406 574.061
R1425 avss.n508 avss.n506 574.061
R1426 avss.n608 avss.n606 574.061
R1427 avss.n783 avss.n781 574.061
R1428 avss.n334 avss.n291 548.058
R1429 avss.n434 avss.n250 548.058
R1430 avss.n534 avss.n207 548.058
R1431 avss.n634 avss.n164 548.058
R1432 avss.n726 avss.n116 548.058
R1433 avss.n798 avss.n42 548.058
R1434 avss.t252 avss.t181 502.274
R1435 avss.t35 avss.t37 502.274
R1436 avss.t186 avss.t136 502.274
R1437 avss.t179 avss.t118 502.274
R1438 avss.t128 avss.t125 502.274
R1439 avss.t155 avss.t195 502.274
R1440 avss.t187 avss.t104 502.274
R1441 avss.t44 avss.t221 502.274
R1442 avss.t123 avss.t55 502.274
R1443 avss.t16 avss.t0 502.274
R1444 avss.t274 avss.t209 502.274
R1445 avss.t232 avss.t234 502.274
R1446 avss.t107 avss.t124 502.274
R1447 avss.t261 avss.t275 502.274
R1448 avss.t103 avss.t54 502.274
R1449 avss.t215 avss.t212 502.274
R1450 avss.t228 avss.t4 501.892
R1451 avss.t263 avss.t265 501.892
R1452 avss.t165 avss.t120 501.892
R1453 avss.t29 avss.t27 501.892
R1454 avss.t31 avss.t34 501.892
R1455 avss.t12 avss.t10 501.892
R1456 avss.t138 avss.t43 501.892
R1457 avss.t52 avss.t50 501.892
R1458 avss.n345 avss.n291 484.702
R1459 avss.n445 avss.n250 484.702
R1460 avss.n545 avss.n207 484.702
R1461 avss.n645 avss.n164 484.702
R1462 avss.n737 avss.n116 484.702
R1463 avss.n809 avss.n42 484.702
R1464 avss.t242 avss.t143 465.733
R1465 avss.t143 avss.t65 465.733
R1466 avss.t255 avss.t178 465.733
R1467 avss.t178 avss.t88 465.733
R1468 avss.t48 avss.t49 465.733
R1469 avss.t49 avss.t69 465.733
R1470 avss.t9 avss.t205 465.733
R1471 avss.t205 avss.t92 465.733
R1472 avss.t129 avss.t256 465.733
R1473 avss.t256 avss.t82 465.733
R1474 avss.t241 avss.t8 465.733
R1475 avss.t59 avss.t241 465.733
R1476 avss.t96 avss.t250 465.37
R1477 avss.t198 avss.t96 465.37
R1478 avss.t166 avss.t144 465.37
R1479 avss.t71 avss.t166 465.37
R1480 avss.t77 avss.t248 465.37
R1481 avss.t229 avss.t77 465.37
R1482 avss.t174 avss.t177 465.37
R1483 avss.t99 avss.t174 465.37
R1484 avss.t97 avss.t245 465.37
R1485 avss.t171 avss.t97 465.37
R1486 avss.t208 avss.t269 465.37
R1487 avss.t80 avss.t208 465.37
R1488 avss.t90 avss.t247 465.37
R1489 avss.t160 avss.t90 465.37
R1490 avss.t42 avss.t204 465.37
R1491 avss.t94 avss.t42 465.37
R1492 avss.t75 avss.t22 465.37
R1493 avss.t270 avss.t75 465.37
R1494 avss.t163 avss.t225 465.37
R1495 avss.t85 avss.t163 465.37
R1496 avss.t251 avss.t61 465.37
R1497 avss.t61 avss.t121 465.37
R1498 avss.t238 avss.t19 465.37
R1499 avss.t19 avss.t63 465.37
R1500 avss.t246 avss.t197 465.37
R1501 avss.t145 avss.t246 465.37
R1502 avss.t249 avss.t173 465.37
R1503 avss.t175 avss.t249 465.37
R1504 avss.t244 avss.t152 465.37
R1505 avss.t267 avss.t244 465.37
R1506 avss.t243 avss.t41 465.37
R1507 avss.t206 avss.t243 465.37
R1508 avss.t5 avss.t164 465.37
R1509 avss.t257 avss.t5 465.37
R1510 avss.t21 avss.t18 465.37
R1511 avss.t239 avss.t21 465.37
R1512 avss.n832 avss.n5 361.01
R1513 avss.n765 avss.n81 361.01
R1514 avss.n683 avss.n139 360.803
R1515 avss.n583 avss.n182 360.803
R1516 avss.n483 avss.n225 360.803
R1517 avss.n383 avss.n268 360.803
R1518 avss.n80 avss.t105 348.214
R1519 avss.n75 avss.t105 348.214
R1520 avss.n7 avss.t182 348.214
R1521 avss.n853 avss.t182 348.214
R1522 avss.n138 avss.t126 348.06
R1523 avss.n133 avss.t126 348.06
R1524 avss.t32 avss.n587 348.06
R1525 avss.n588 avss.t32 348.06
R1526 avss.t108 avss.n487 348.06
R1527 avss.n488 avss.t108 348.06
R1528 avss.t184 avss.n387 348.06
R1529 avss.n388 avss.t184 348.06
R1530 avss.n299 avss.t87 338.849
R1531 avss.t110 avss.n345 338.849
R1532 avss.n407 avss.t98 338.849
R1533 avss.n507 avss.t79 338.849
R1534 avss.n607 avss.t74 338.849
R1535 avss.n700 avss.t68 338.849
R1536 avss.n782 avss.t76 338.849
R1537 avss.n821 avss.t282 314.01
R1538 avss.n33 avss.t282 314.01
R1539 avss.n32 avss.t6 314.01
R1540 avss.n29 avss.t6 314.01
R1541 avss.n28 avss.t288 314.01
R1542 avss.t288 avss.n22 314.01
R1543 avss.n749 avss.t272 314.01
R1544 avss.n107 avss.t272 314.01
R1545 avss.n106 avss.t2 314.01
R1546 avss.n103 avss.t2 314.01
R1547 avss.n102 avss.t25 314.01
R1548 avss.t25 avss.n96 314.01
R1549 avss.n156 avss.t101 313.884
R1550 avss.n658 avss.t101 313.884
R1551 avss.n659 avss.t286 313.884
R1552 avss.n663 avss.t286 313.884
R1553 avss.t188 avss.n666 313.884
R1554 avss.n667 avss.t188 313.884
R1555 avss.n199 avss.t200 313.884
R1556 avss.n558 avss.t200 313.884
R1557 avss.n559 avss.t223 313.884
R1558 avss.n563 avss.t223 313.884
R1559 avss.t132 avss.n566 313.884
R1560 avss.n567 avss.t132 313.884
R1561 avss.n242 avss.t153 313.884
R1562 avss.n458 avss.t153 313.884
R1563 avss.n459 avss.t46 313.884
R1564 avss.n463 avss.t46 313.884
R1565 avss.t23 avss.n466 313.884
R1566 avss.n467 avss.t23 313.884
R1567 avss.n285 avss.t284 313.884
R1568 avss.n358 avss.t284 313.884
R1569 avss.n359 avss.t226 313.884
R1570 avss.n363 avss.t226 313.884
R1571 avss.t114 avss.n366 313.884
R1572 avss.n367 avss.t114 313.884
R1573 avss.n81 avss.n80 300.336
R1574 avss.n7 avss.n5 300.336
R1575 avss.n139 avss.n138 300.202
R1576 avss.n587 avss.n182 300.202
R1577 avss.n487 avss.n225 300.202
R1578 avss.n387 avss.n268 300.202
R1579 avss.n739 avss.t162 279.964
R1580 avss.t193 avss.n98 279.964
R1581 avss.n811 avss.t167 279.964
R1582 avss.t39 avss.n24 279.964
R1583 avss.t210 avss.n347 279.858
R1584 avss.n348 avss.t148 279.858
R1585 avss.t168 avss.n447 279.858
R1586 avss.n448 avss.t157 279.858
R1587 avss.t231 avss.n547 279.858
R1588 avss.n548 avss.t141 279.858
R1589 avss.t279 avss.n647 279.858
R1590 avss.n648 avss.t57 279.858
R1591 avss.t147 avss.t110 271.079
R1592 avss.t98 avss.t159 271.079
R1593 avss.t159 avss.t116 271.079
R1594 avss.t79 avss.t137 271.079
R1595 avss.t137 avss.t190 271.079
R1596 avss.t74 avss.t56 271.079
R1597 avss.t56 avss.t219 271.079
R1598 avss.t68 avss.t192 271.079
R1599 avss.t192 avss.t14 271.079
R1600 avss.t76 avss.t20 271.079
R1601 avss.t20 avss.t277 271.079
R1602 avss.n33 avss.n32 266.909
R1603 avss.n29 avss.n28 266.909
R1604 avss.n107 avss.n106 266.909
R1605 avss.n103 avss.n102 266.909
R1606 avss.n659 avss.n658 266.801
R1607 avss.n666 avss.n663 266.801
R1608 avss.n559 avss.n558 266.801
R1609 avss.n566 avss.n563 266.801
R1610 avss.n459 avss.n458 266.801
R1611 avss.n466 avss.n463 266.801
R1612 avss.n359 avss.n358 266.801
R1613 avss.n366 avss.n363 266.801
R1614 avss.t162 avss.t84 223.97
R1615 avss.t84 avss.t193 223.97
R1616 avss.t167 avss.t78 223.97
R1617 avss.t78 avss.t39 223.97
R1618 avss.t67 avss.t210 223.887
R1619 avss.t148 avss.t67 223.887
R1620 avss.t91 avss.t168 223.887
R1621 avss.t157 avss.t91 223.887
R1622 avss.t73 avss.t231 223.887
R1623 avss.t141 avss.t73 223.887
R1624 avss.t62 avss.t279 223.887
R1625 avss.t57 avss.t62 223.887
R1626 avss.n346 avss.t147 220.988
R1627 avss.n446 avss.n445 213.623
R1628 avss.n546 avss.n545 213.623
R1629 avss.n646 avss.n645 213.623
R1630 avss.n738 avss.n737 213.623
R1631 avss.n810 avss.n809 213.623
R1632 avss.n410 avss.n409 151.869
R1633 avss.n510 avss.n509 151.869
R1634 avss.n610 avss.n609 151.869
R1635 avss.n703 avss.n702 151.869
R1636 avss.n784 avss.n74 151.869
R1637 avss.n326 avss.n325 151.751
R1638 avss.n321 avss.n320 151.751
R1639 avss.n302 avss.n301 151.751
R1640 avss.n426 avss.n425 151.751
R1641 avss.n422 avss.n421 151.751
R1642 avss.n260 avss.n259 151.751
R1643 avss.n526 avss.n525 151.751
R1644 avss.n522 avss.n521 151.751
R1645 avss.n217 avss.n216 151.751
R1646 avss.n626 avss.n625 151.751
R1647 avss.n622 avss.n621 151.751
R1648 avss.n174 avss.n173 151.751
R1649 avss.n718 avss.n52 151.751
R1650 avss.n715 avss.n714 151.751
R1651 avss.n125 avss.n51 151.751
R1652 avss.n790 avss.n789 151.751
R1653 avss.n60 avss.n50 151.751
R1654 avss.n787 avss.n49 151.751
R1655 avss.n335 avss.n283 151.751
R1656 avss.n435 avss.n240 151.751
R1657 avss.n535 avss.n197 151.751
R1658 avss.n635 avss.n154 151.751
R1659 avss.n727 avss.n97 151.751
R1660 avss.n799 avss.n23 151.751
R1661 avss.n375 avss.n374 147.727
R1662 avss.n406 avss.n405 147.727
R1663 avss.n475 avss.n474 147.727
R1664 avss.n506 avss.n505 147.727
R1665 avss.n575 avss.n574 147.727
R1666 avss.n606 avss.n605 147.727
R1667 avss.n675 avss.n674 147.727
R1668 avss.n699 avss.n698 147.727
R1669 avss.n756 avss.n755 147.727
R1670 avss.n781 avss.n780 147.727
R1671 avss.n824 avss.n823 147.727
R1672 avss.n855 avss.n854 147.727
R1673 avss.n446 avss.t116 125.228
R1674 avss.n546 avss.t190 125.228
R1675 avss.n646 avss.t219 125.228
R1676 avss.n738 avss.t14 125.228
R1677 avss.n810 avss.t277 125.228
R1678 avss.n408 avss.n407 88.3958
R1679 avss.n508 avss.n507 88.3958
R1680 avss.n608 avss.n607 88.3958
R1681 avss.n701 avss.n700 88.3958
R1682 avss.n783 avss.n782 88.3958
R1683 avss.n856 avss.n3 87.3061
R1684 avss.n856 avss.n4 87.3061
R1685 avss.n779 avss.n82 87.3061
R1686 avss.n779 avss.n83 87.3061
R1687 avss.n766 avss.n94 87.3061
R1688 avss.n766 avss.n95 87.3061
R1689 avss.n697 avss.n140 87.3061
R1690 avss.n697 avss.n141 87.3061
R1691 avss.n684 avss.n151 87.3061
R1692 avss.n684 avss.n152 87.3061
R1693 avss.n604 avss.n183 87.3061
R1694 avss.n604 avss.n184 87.3061
R1695 avss.n584 avss.n194 87.3061
R1696 avss.n584 avss.n195 87.3061
R1697 avss.n504 avss.n226 87.3061
R1698 avss.n504 avss.n227 87.3061
R1699 avss.n484 avss.n237 87.3061
R1700 avss.n484 avss.n238 87.3061
R1701 avss.n404 avss.n269 87.3061
R1702 avss.n404 avss.n270 87.3061
R1703 avss.n384 avss.n280 87.3061
R1704 avss.n384 avss.n281 87.3061
R1705 avss.n831 avss.n20 87.3061
R1706 avss.n831 avss.n830 87.3061
R1707 avss.n825 avss.n22 78.5029
R1708 avss.n757 avss.n96 78.5029
R1709 avss.n673 avss.n667 78.4713
R1710 avss.n573 avss.n567 78.4713
R1711 avss.n473 avss.n467 78.4713
R1712 avss.n373 avss.n367 78.4713
R1713 avss.n17 avss.n16 67.4727
R1714 avss.n18 avss.n16 67.4727
R1715 avss.n751 avss.n87 67.4727
R1716 avss.n752 avss.n87 67.4727
R1717 avss.n759 avss.n91 67.4727
R1718 avss.n760 avss.n91 67.4727
R1719 avss.n676 avss.n144 67.4727
R1720 avss.n677 avss.n144 67.4727
R1721 avss.n668 avss.n148 67.4727
R1722 avss.n669 avss.n148 67.4727
R1723 avss.n576 avss.n187 67.4727
R1724 avss.n577 avss.n187 67.4727
R1725 avss.n568 avss.n191 67.4727
R1726 avss.n569 avss.n191 67.4727
R1727 avss.n476 avss.n230 67.4727
R1728 avss.n477 avss.n230 67.4727
R1729 avss.n468 avss.n234 67.4727
R1730 avss.n469 avss.n234 67.4727
R1731 avss.n376 avss.n273 67.4727
R1732 avss.n377 avss.n273 67.4727
R1733 avss.n368 avss.n277 67.4727
R1734 avss.n369 avss.n277 67.4727
R1735 avss.n21 avss.n12 67.4727
R1736 avss.n829 avss.n12 67.4727
R1737 avss.n17 avss.n3 66.5005
R1738 avss.n18 avss.n4 66.5005
R1739 avss.n751 avss.n82 66.5005
R1740 avss.n752 avss.n83 66.5005
R1741 avss.n759 avss.n94 66.5005
R1742 avss.n760 avss.n95 66.5005
R1743 avss.n676 avss.n140 66.5005
R1744 avss.n677 avss.n141 66.5005
R1745 avss.n668 avss.n151 66.5005
R1746 avss.n669 avss.n152 66.5005
R1747 avss.n576 avss.n183 66.5005
R1748 avss.n577 avss.n184 66.5005
R1749 avss.n568 avss.n194 66.5005
R1750 avss.n569 avss.n195 66.5005
R1751 avss.n476 avss.n226 66.5005
R1752 avss.n477 avss.n227 66.5005
R1753 avss.n468 avss.n237 66.5005
R1754 avss.n469 avss.n238 66.5005
R1755 avss.n376 avss.n269 66.5005
R1756 avss.n377 avss.n270 66.5005
R1757 avss.n368 avss.n280 66.5005
R1758 avss.n369 avss.n281 66.5005
R1759 avss.n21 avss.n20 66.5005
R1760 avss.n830 avss.n829 66.5005
R1761 avss.n319 avss.n303 61.0571
R1762 avss.n420 avss.n261 61.0571
R1763 avss.n520 avss.n218 61.0571
R1764 avss.n620 avss.n175 61.0571
R1765 avss.n713 avss.n126 61.0571
R1766 avss.n62 avss.n61 61.0571
R1767 avss.n800 avss.n797 61.0561
R1768 avss.n808 avss.n43 61.0561
R1769 avss.n813 avss.n812 61.0561
R1770 avss.n728 avss.n725 61.0561
R1771 avss.n736 avss.n117 61.0561
R1772 avss.n741 avss.n740 61.0561
R1773 avss.n636 avss.n633 61.0561
R1774 avss.n644 avss.n165 61.0561
R1775 avss.n649 avss.n162 61.0561
R1776 avss.n536 avss.n533 61.0561
R1777 avss.n544 avss.n208 61.0561
R1778 avss.n549 avss.n205 61.0561
R1779 avss.n436 avss.n433 61.0561
R1780 avss.n444 avss.n251 61.0561
R1781 avss.n449 avss.n248 61.0561
R1782 avss.n336 avss.n333 61.0561
R1783 avss.n344 avss.n292 61.0561
R1784 avss.n349 avss.n290 61.0561
R1785 avss.n327 avss.n297 61.0561
R1786 avss.n311 avss.n310 61.0561
R1787 avss.n427 avss.n256 61.0561
R1788 avss.n412 avss.n411 61.0561
R1789 avss.n527 avss.n213 61.0561
R1790 avss.n512 avss.n511 61.0561
R1791 avss.n627 avss.n170 61.0561
R1792 avss.n612 avss.n611 61.0561
R1793 avss.n719 avss.n122 61.0561
R1794 avss.n705 avss.n704 61.0561
R1795 avss.n791 avss.n48 61.0561
R1796 avss.n73 avss.n57 61.0561
R1797 avss.n346 avss.t87 50.0912
R1798 avss.n31 avss.n30 44.1404
R1799 avss.n27 avss.n13 44.1404
R1800 avss.n79 avss.n76 44.1404
R1801 avss.n105 avss.n104 44.1404
R1802 avss.n101 avss.n90 44.1404
R1803 avss.n137 avss.n134 44.1404
R1804 avss.n662 avss.n660 44.1404
R1805 avss.n665 avss.n147 44.1404
R1806 avss.n589 avss.n586 44.1404
R1807 avss.n562 avss.n560 44.1404
R1808 avss.n565 avss.n190 44.1404
R1809 avss.n489 avss.n486 44.1404
R1810 avss.n462 avss.n460 44.1404
R1811 avss.n465 avss.n233 44.1404
R1812 avss.n389 avss.n386 44.1404
R1813 avss.n852 avss.n8 44.1404
R1814 avss.n365 avss.n276 44.1394
R1815 avss.n362 avss.n360 44.1394
R1816 avss.n357 avss.n286 44.1394
R1817 avss.n820 avss.n34 44.1394
R1818 avss.n748 avss.n108 44.1394
R1819 avss.n657 avss.n157 44.1394
R1820 avss.n557 avss.n200 44.1394
R1821 avss.n457 avss.n243 44.1394
R1822 avss.n1 avss.t290 34.1066
R1823 avss.n835 avss.n3 20.8061
R1824 avss.n835 avss.n4 20.8061
R1825 avss.n838 avss.n17 20.8061
R1826 avss.n838 avss.n18 20.8061
R1827 avss.n84 avss.n82 20.8061
R1828 avss.n84 avss.n83 20.8061
R1829 avss.n753 avss.n751 20.8061
R1830 avss.n753 avss.n752 20.8061
R1831 avss.n763 avss.n94 20.8061
R1832 avss.n763 avss.n95 20.8061
R1833 avss.n761 avss.n759 20.8061
R1834 avss.n761 avss.n760 20.8061
R1835 avss.n680 avss.n140 20.8061
R1836 avss.n680 avss.n141 20.8061
R1837 avss.n678 avss.n676 20.8061
R1838 avss.n678 avss.n677 20.8061
R1839 avss.n153 avss.n151 20.8061
R1840 avss.n153 avss.n152 20.8061
R1841 avss.n670 avss.n668 20.8061
R1842 avss.n670 avss.n669 20.8061
R1843 avss.n580 avss.n183 20.8061
R1844 avss.n580 avss.n184 20.8061
R1845 avss.n578 avss.n576 20.8061
R1846 avss.n578 avss.n577 20.8061
R1847 avss.n196 avss.n194 20.8061
R1848 avss.n196 avss.n195 20.8061
R1849 avss.n570 avss.n568 20.8061
R1850 avss.n570 avss.n569 20.8061
R1851 avss.n480 avss.n226 20.8061
R1852 avss.n480 avss.n227 20.8061
R1853 avss.n478 avss.n476 20.8061
R1854 avss.n478 avss.n477 20.8061
R1855 avss.n239 avss.n237 20.8061
R1856 avss.n239 avss.n238 20.8061
R1857 avss.n470 avss.n468 20.8061
R1858 avss.n470 avss.n469 20.8061
R1859 avss.n380 avss.n269 20.8061
R1860 avss.n380 avss.n270 20.8061
R1861 avss.n378 avss.n376 20.8061
R1862 avss.n378 avss.n377 20.8061
R1863 avss.n282 avss.n280 20.8061
R1864 avss.n282 avss.n281 20.8061
R1865 avss.n370 avss.n368 20.8061
R1866 avss.n370 avss.n369 20.8061
R1867 avss.n828 avss.n21 20.8061
R1868 avss.n829 avss.n828 20.8061
R1869 avss.n20 avss.n19 20.8061
R1870 avss.n830 avss.n19 20.8061
R1871 avss.n0 avss.t214 19.673
R1872 avss.n0 avss.t211 19.4007
R1873 avss.n859 avss.n858 14.6135
R1874 avss.n289 avss.n287 9.0005
R1875 avss.n340 avss.n339 9.0005
R1876 avss.n318 avss.n317 9.0005
R1877 avss.n305 avss.n294 9.0005
R1878 avss.n308 avss.n307 9.0005
R1879 avss.n314 avss.n313 9.0005
R1880 avss.n296 avss.n295 9.0005
R1881 avss.n330 avss.n329 9.0005
R1882 avss.n338 avss.n288 9.0005
R1883 avss.n352 avss.n351 9.0005
R1884 avss.n247 avss.n245 9.0005
R1885 avss.n440 avss.n439 9.0005
R1886 avss.n419 avss.n418 9.0005
R1887 avss.n263 avss.n253 9.0005
R1888 avss.n266 avss.n265 9.0005
R1889 avss.n415 avss.n414 9.0005
R1890 avss.n255 avss.n254 9.0005
R1891 avss.n430 avss.n429 9.0005
R1892 avss.n438 avss.n246 9.0005
R1893 avss.n452 avss.n451 9.0005
R1894 avss.n204 avss.n202 9.0005
R1895 avss.n540 avss.n539 9.0005
R1896 avss.n519 avss.n518 9.0005
R1897 avss.n220 avss.n210 9.0005
R1898 avss.n223 avss.n222 9.0005
R1899 avss.n515 avss.n514 9.0005
R1900 avss.n212 avss.n211 9.0005
R1901 avss.n530 avss.n529 9.0005
R1902 avss.n538 avss.n203 9.0005
R1903 avss.n552 avss.n551 9.0005
R1904 avss.n161 avss.n159 9.0005
R1905 avss.n640 avss.n639 9.0005
R1906 avss.n619 avss.n618 9.0005
R1907 avss.n177 avss.n167 9.0005
R1908 avss.n180 avss.n179 9.0005
R1909 avss.n615 avss.n614 9.0005
R1910 avss.n169 avss.n168 9.0005
R1911 avss.n630 avss.n629 9.0005
R1912 avss.n638 avss.n160 9.0005
R1913 avss.n652 avss.n651 9.0005
R1914 avss.n114 avss.n112 9.0005
R1915 avss.n732 avss.n731 9.0005
R1916 avss.n712 avss.n711 9.0005
R1917 avss.n128 avss.n119 9.0005
R1918 avss.n131 avss.n130 9.0005
R1919 avss.n708 avss.n707 9.0005
R1920 avss.n121 avss.n120 9.0005
R1921 avss.n722 avss.n721 9.0005
R1922 avss.n730 avss.n113 9.0005
R1923 avss.n744 avss.n743 9.0005
R1924 avss.n40 avss.n38 9.0005
R1925 avss.n804 avss.n803 9.0005
R1926 avss.n66 avss.n65 9.0005
R1927 avss.n64 avss.n45 9.0005
R1928 avss.n72 avss.n58 9.0005
R1929 avss.n71 avss.n69 9.0005
R1930 avss.n47 avss.n46 9.0005
R1931 avss.n794 avss.n793 9.0005
R1932 avss.n802 avss.n39 9.0005
R1933 avss.n816 avss.n815 9.0005
R1934 avss.n342 avss.n292 6.9012
R1935 avss.n442 avss.n251 6.9012
R1936 avss.n542 avss.n208 6.9012
R1937 avss.n642 avss.n165 6.9012
R1938 avss.n734 avss.n117 6.9012
R1939 avss.n806 avss.n43 6.9012
R1940 avss.n339 avss.n333 6.46296
R1941 avss.n297 avss.n296 6.46296
R1942 avss.n310 avss.n308 6.46296
R1943 avss.n439 avss.n433 6.46296
R1944 avss.n256 avss.n255 6.46296
R1945 avss.n411 avss.n266 6.46296
R1946 avss.n539 avss.n533 6.46296
R1947 avss.n213 avss.n212 6.46296
R1948 avss.n511 avss.n223 6.46296
R1949 avss.n639 avss.n633 6.46296
R1950 avss.n170 avss.n169 6.46296
R1951 avss.n611 avss.n180 6.46296
R1952 avss.n731 avss.n725 6.46296
R1953 avss.n122 avss.n121 6.46296
R1954 avss.n704 avss.n131 6.46296
R1955 avss.n803 avss.n797 6.46296
R1956 avss.n48 avss.n47 6.46296
R1957 avss.n73 avss.n72 6.46296
R1958 avss.n290 avss.n289 6.4618
R1959 avss.n319 avss.n318 6.4618
R1960 avss.n248 avss.n247 6.4618
R1961 avss.n420 avss.n419 6.4618
R1962 avss.n205 avss.n204 6.4618
R1963 avss.n520 avss.n519 6.4618
R1964 avss.n162 avss.n161 6.4618
R1965 avss.n620 avss.n619 6.4618
R1966 avss.n740 avss.n114 6.4618
R1967 avss.n713 avss.n712 6.4618
R1968 avss.n812 avss.n40 6.4618
R1969 avss.n65 avss.n61 6.4618
R1970 avss.n343 avss.n342 5.47239
R1971 avss.n443 avss.n442 5.47239
R1972 avss.n543 avss.n542 5.47239
R1973 avss.n643 avss.n642 5.47239
R1974 avss.n735 avss.n734 5.47239
R1975 avss.n807 avss.n806 5.47239
R1976 avss.n859 avss.n1 5.18044
R1977 avss.n351 avss.n350 5.03414
R1978 avss.n338 avss.n337 5.03414
R1979 avss.n329 avss.n328 5.03414
R1980 avss.n313 avss.n312 5.03414
R1981 avss.n305 avss.n304 5.03414
R1982 avss.n451 avss.n450 5.03414
R1983 avss.n438 avss.n437 5.03414
R1984 avss.n429 avss.n428 5.03414
R1985 avss.n414 avss.n413 5.03414
R1986 avss.n263 avss.n262 5.03414
R1987 avss.n551 avss.n550 5.03414
R1988 avss.n538 avss.n537 5.03414
R1989 avss.n529 avss.n528 5.03414
R1990 avss.n514 avss.n513 5.03414
R1991 avss.n220 avss.n219 5.03414
R1992 avss.n651 avss.n650 5.03414
R1993 avss.n638 avss.n637 5.03414
R1994 avss.n629 avss.n628 5.03414
R1995 avss.n614 avss.n613 5.03414
R1996 avss.n177 avss.n176 5.03414
R1997 avss.n743 avss.n742 5.03414
R1998 avss.n730 avss.n729 5.03414
R1999 avss.n721 avss.n720 5.03414
R2000 avss.n707 avss.n706 5.03414
R2001 avss.n128 avss.n127 5.03414
R2002 avss.n815 avss.n814 5.03414
R2003 avss.n802 avss.n801 5.03414
R2004 avss.n793 avss.n792 5.03414
R2005 avss.n71 avss.n70 5.03414
R2006 avss.n64 avss.n63 5.03414
R2007 avss.n26 avss.t289 4.84702
R2008 avss.n25 avss.t7 4.84702
R2009 avss.n100 avss.t26 4.84702
R2010 avss.n99 avss.t3 4.84702
R2011 avss.n664 avss.t189 4.84702
R2012 avss.n661 avss.t287 4.84702
R2013 avss.n564 avss.t133 4.84702
R2014 avss.n561 avss.t224 4.84702
R2015 avss.n464 avss.t24 4.84702
R2016 avss.n461 avss.t47 4.84702
R2017 avss.n364 avss.t115 4.84702
R2018 avss.n361 avss.t227 4.84702
R2019 avss.n272 avss.t254 4.7885
R2020 avss.n271 avss.t180 4.7885
R2021 avss.n403 avss.t119 4.7885
R2022 avss.n350 avss.t149 4.7885
R2023 avss.n337 avss.t146 4.7885
R2024 avss.n343 avss.t111 4.7885
R2025 avss.n328 avss.t199 4.7885
R2026 avss.n312 avss.t66 4.7885
R2027 avss.n304 avss.t72 4.7885
R2028 avss.n229 avss.t260 4.7885
R2029 avss.n228 avss.t156 4.7885
R2030 avss.n503 avss.t196 4.7885
R2031 avss.n450 avss.t158 4.7885
R2032 avss.n437 avss.t176 4.7885
R2033 avss.n443 avss.t117 4.7885
R2034 avss.n428 avss.t230 4.7885
R2035 avss.n413 avss.t89 4.7885
R2036 avss.n262 avss.t100 4.7885
R2037 avss.n186 avss.t131 4.7885
R2038 avss.n185 avss.t45 4.7885
R2039 avss.n603 avss.t222 4.7885
R2040 avss.n550 avss.t142 4.7885
R2041 avss.n537 avss.t268 4.7885
R2042 avss.n543 avss.t191 4.7885
R2043 avss.n528 avss.t172 4.7885
R2044 avss.n513 avss.t70 4.7885
R2045 avss.n219 avss.t81 4.7885
R2046 avss.n143 avss.t113 4.7885
R2047 avss.n142 avss.t17 4.7885
R2048 avss.n696 avss.t1 4.7885
R2049 avss.n650 avss.t58 4.7885
R2050 avss.n637 avss.t207 4.7885
R2051 avss.n643 avss.t220 4.7885
R2052 avss.n628 avss.t161 4.7885
R2053 avss.n613 avss.t93 4.7885
R2054 avss.n176 avss.t95 4.7885
R2055 avss.n86 avss.t203 4.7885
R2056 avss.n85 avss.t276 4.7885
R2057 avss.n778 avss.t262 4.7885
R2058 avss.n742 avss.t194 4.7885
R2059 avss.n729 avss.t258 4.7885
R2060 avss.n735 avss.t15 4.7885
R2061 avss.n720 avss.t271 4.7885
R2062 avss.n706 avss.t83 4.7885
R2063 avss.n127 avss.t86 4.7885
R2064 avss.n814 avss.t40 4.7885
R2065 avss.n801 avss.t240 4.7885
R2066 avss.n807 avss.t278 4.7885
R2067 avss.n792 avss.t122 4.7885
R2068 avss.n70 avss.t60 4.7885
R2069 avss.n63 avss.t64 4.7885
R2070 avss.n839 avss.t281 4.7885
R2071 avss.n834 avss.t216 4.7885
R2072 avss.n857 avss.t213 4.7885
R2073 avss.n10 avss.t36 4.7885
R2074 avss.n11 avss.t135 4.7885
R2075 avss.n9 avss.t38 4.7885
R2076 avss.n36 avss.t283 4.7885
R2077 avss.n77 avss.t106 4.7885
R2078 avss.n92 avss.t140 4.7885
R2079 avss.n93 avss.t235 4.7885
R2080 avss.n767 avss.t233 4.7885
R2081 avss.n110 avss.t273 4.7885
R2082 avss.n135 avss.t127 4.7885
R2083 avss.n149 avss.t151 4.7885
R2084 avss.n150 avss.t51 4.7885
R2085 avss.n685 avss.t53 4.7885
R2086 avss.n656 avss.t102 4.7885
R2087 avss.n590 avss.t33 4.7885
R2088 avss.n192 avss.t237 4.7885
R2089 avss.n193 avss.t11 4.7885
R2090 avss.n585 avss.t13 4.7885
R2091 avss.n556 avss.t201 4.7885
R2092 avss.n490 avss.t109 4.7885
R2093 avss.n235 avss.t170 4.7885
R2094 avss.n236 avss.t28 4.7885
R2095 avss.n485 avss.t30 4.7885
R2096 avss.n456 avss.t154 4.7885
R2097 avss.n390 avss.t185 4.7885
R2098 avss.n278 avss.t218 4.7885
R2099 avss.n279 avss.t266 4.7885
R2100 avss.n385 avss.t264 4.7885
R2101 avss.n356 avss.t285 4.7885
R2102 avss.n851 avss.t183 4.7885
R2103 avss.n342 avss.n341 4.28213
R2104 avss.n442 avss.n441 4.28213
R2105 avss.n542 avss.n541 4.28213
R2106 avss.n642 avss.n641 4.28213
R2107 avss.n734 avss.n733 4.28213
R2108 avss.n806 avss.n805 4.28213
R2109 avss.n400 avss.n399 3.51467
R2110 avss.n500 avss.n499 3.51467
R2111 avss.n600 avss.n599 3.51467
R2112 avss.n693 avss.n692 3.51467
R2113 avss.n775 avss.n774 3.51467
R2114 avss.n842 avss.n841 3.51467
R2115 avss.n400 avss.n273 2.06002
R2116 avss.n500 avss.n230 2.06002
R2117 avss.n600 avss.n187 2.06002
R2118 avss.n693 avss.n144 2.06002
R2119 avss.n775 avss.n87 2.06002
R2120 avss.n841 avss.n16 2.06002
R2121 avss.n354 avss.n286 1.92616
R2122 avss.n845 avss.n12 1.90702
R2123 avss.n820 avss.n819 1.90702
R2124 avss.n31 avss.n15 1.90702
R2125 avss.n844 avss.n13 1.90702
R2126 avss.n79 avss.n78 1.90702
R2127 avss.n771 avss.n91 1.90702
R2128 avss.n748 avss.n747 1.90702
R2129 avss.n105 avss.n88 1.90702
R2130 avss.n772 avss.n90 1.90702
R2131 avss.n137 avss.n136 1.90702
R2132 avss.n689 avss.n148 1.90702
R2133 avss.n158 avss.n157 1.90702
R2134 avss.n660 avss.n145 1.90702
R2135 avss.n690 avss.n147 1.90702
R2136 avss.n591 avss.n586 1.90702
R2137 avss.n596 avss.n191 1.90702
R2138 avss.n201 avss.n200 1.90702
R2139 avss.n560 avss.n188 1.90702
R2140 avss.n597 avss.n190 1.90702
R2141 avss.n491 avss.n486 1.90702
R2142 avss.n496 avss.n234 1.90702
R2143 avss.n244 avss.n243 1.90702
R2144 avss.n460 avss.n231 1.90702
R2145 avss.n497 avss.n233 1.90702
R2146 avss.n391 avss.n386 1.90702
R2147 avss.n396 avss.n277 1.90702
R2148 avss.n360 avss.n274 1.90702
R2149 avss.n397 avss.n276 1.90702
R2150 avss.n850 avss.n8 1.90702
R2151 2inmux_0.Bit avss.n859 1.54251
R2152 avss.n310 avss.n309 1.3005
R2153 avss.n312 avss.n311 1.3005
R2154 avss.n311 avss.n298 1.3005
R2155 avss.n324 avss.n297 1.3005
R2156 avss.n328 avss.n327 1.3005
R2157 avss.n327 avss.n326 1.3005
R2158 avss.n304 avss.n303 1.3005
R2159 avss.n303 avss.n302 1.3005
R2160 avss.n320 avss.n319 1.3005
R2161 avss.n411 avss.n410 1.3005
R2162 avss.n413 avss.n412 1.3005
R2163 avss.n412 avss.n257 1.3005
R2164 avss.n424 avss.n256 1.3005
R2165 avss.n428 avss.n427 1.3005
R2166 avss.n427 avss.n426 1.3005
R2167 avss.n262 avss.n261 1.3005
R2168 avss.n261 avss.n260 1.3005
R2169 avss.n421 avss.n420 1.3005
R2170 avss.n511 avss.n510 1.3005
R2171 avss.n513 avss.n512 1.3005
R2172 avss.n512 avss.n214 1.3005
R2173 avss.n524 avss.n213 1.3005
R2174 avss.n528 avss.n527 1.3005
R2175 avss.n527 avss.n526 1.3005
R2176 avss.n219 avss.n218 1.3005
R2177 avss.n218 avss.n217 1.3005
R2178 avss.n521 avss.n520 1.3005
R2179 avss.n611 avss.n610 1.3005
R2180 avss.n613 avss.n612 1.3005
R2181 avss.n612 avss.n171 1.3005
R2182 avss.n624 avss.n170 1.3005
R2183 avss.n628 avss.n627 1.3005
R2184 avss.n627 avss.n626 1.3005
R2185 avss.n176 avss.n175 1.3005
R2186 avss.n175 avss.n174 1.3005
R2187 avss.n621 avss.n620 1.3005
R2188 avss.n704 avss.n703 1.3005
R2189 avss.n706 avss.n705 1.3005
R2190 avss.n705 avss.n123 1.3005
R2191 avss.n717 avss.n122 1.3005
R2192 avss.n720 avss.n719 1.3005
R2193 avss.n719 avss.n718 1.3005
R2194 avss.n127 avss.n126 1.3005
R2195 avss.n126 avss.n125 1.3005
R2196 avss.n714 avss.n713 1.3005
R2197 avss.n74 avss.n73 1.3005
R2198 avss.n70 avss.n57 1.3005
R2199 avss.n57 avss.n56 1.3005
R2200 avss.n54 avss.n48 1.3005
R2201 avss.n792 avss.n791 1.3005
R2202 avss.n791 avss.n790 1.3005
R2203 avss.n63 avss.n62 1.3005
R2204 avss.n62 avss.n49 1.3005
R2205 avss.n61 avss.n60 1.3005
R2206 avss.n828 avss.n11 1.3005
R2207 avss.n828 avss.n827 1.3005
R2208 avss.n826 avss.n12 1.3005
R2209 avss.n19 avss.n10 1.3005
R2210 avss.n833 avss.n19 1.3005
R2211 avss.n831 avss.n9 1.3005
R2212 avss.n832 avss.n831 1.3005
R2213 avss.n821 avss.n820 1.3005
R2214 avss.n36 avss.n34 1.3005
R2215 avss.n34 avss.n33 1.3005
R2216 avss.n32 avss.n31 1.3005
R2217 avss.n30 avss.n25 1.3005
R2218 avss.n30 avss.n29 1.3005
R2219 avss.n27 avss.n26 1.3005
R2220 avss.n28 avss.n27 1.3005
R2221 avss.n22 avss.n13 1.3005
R2222 avss.n77 avss.n76 1.3005
R2223 avss.n76 avss.n75 1.3005
R2224 avss.n80 avss.n79 1.3005
R2225 avss.n749 avss.n748 1.3005
R2226 avss.n110 avss.n108 1.3005
R2227 avss.n108 avss.n107 1.3005
R2228 avss.n106 avss.n105 1.3005
R2229 avss.n104 avss.n99 1.3005
R2230 avss.n104 avss.n103 1.3005
R2231 avss.n101 avss.n100 1.3005
R2232 avss.n102 avss.n101 1.3005
R2233 avss.n96 avss.n90 1.3005
R2234 avss.n135 avss.n134 1.3005
R2235 avss.n134 avss.n133 1.3005
R2236 avss.n138 avss.n137 1.3005
R2237 avss.n157 avss.n156 1.3005
R2238 avss.n657 avss.n656 1.3005
R2239 avss.n658 avss.n657 1.3005
R2240 avss.n660 avss.n659 1.3005
R2241 avss.n662 avss.n661 1.3005
R2242 avss.n663 avss.n662 1.3005
R2243 avss.n665 avss.n664 1.3005
R2244 avss.n666 avss.n665 1.3005
R2245 avss.n667 avss.n147 1.3005
R2246 avss.n590 avss.n589 1.3005
R2247 avss.n589 avss.n588 1.3005
R2248 avss.n587 avss.n586 1.3005
R2249 avss.n200 avss.n199 1.3005
R2250 avss.n557 avss.n556 1.3005
R2251 avss.n558 avss.n557 1.3005
R2252 avss.n560 avss.n559 1.3005
R2253 avss.n562 avss.n561 1.3005
R2254 avss.n563 avss.n562 1.3005
R2255 avss.n565 avss.n564 1.3005
R2256 avss.n566 avss.n565 1.3005
R2257 avss.n567 avss.n190 1.3005
R2258 avss.n490 avss.n489 1.3005
R2259 avss.n489 avss.n488 1.3005
R2260 avss.n487 avss.n486 1.3005
R2261 avss.n243 avss.n242 1.3005
R2262 avss.n457 avss.n456 1.3005
R2263 avss.n458 avss.n457 1.3005
R2264 avss.n460 avss.n459 1.3005
R2265 avss.n462 avss.n461 1.3005
R2266 avss.n463 avss.n462 1.3005
R2267 avss.n465 avss.n464 1.3005
R2268 avss.n466 avss.n465 1.3005
R2269 avss.n467 avss.n233 1.3005
R2270 avss.n390 avss.n389 1.3005
R2271 avss.n389 avss.n388 1.3005
R2272 avss.n387 avss.n386 1.3005
R2273 avss.n286 avss.n285 1.3005
R2274 avss.n357 avss.n356 1.3005
R2275 avss.n358 avss.n357 1.3005
R2276 avss.n360 avss.n359 1.3005
R2277 avss.n362 avss.n361 1.3005
R2278 avss.n363 avss.n362 1.3005
R2279 avss.n365 avss.n364 1.3005
R2280 avss.n366 avss.n365 1.3005
R2281 avss.n367 avss.n276 1.3005
R2282 avss.n347 avss.n290 1.3005
R2283 avss.n350 avss.n349 1.3005
R2284 avss.n349 avss.n348 1.3005
R2285 avss.n299 avss.n292 1.3005
R2286 avss.n344 avss.n343 1.3005
R2287 avss.n345 avss.n344 1.3005
R2288 avss.n334 avss.n333 1.3005
R2289 avss.n337 avss.n336 1.3005
R2290 avss.n336 avss.n335 1.3005
R2291 avss.n372 avss.n277 1.3005
R2292 avss.n370 avss.n278 1.3005
R2293 avss.n371 avss.n370 1.3005
R2294 avss.n282 avss.n279 1.3005
R2295 avss.n382 avss.n282 1.3005
R2296 avss.n385 avss.n384 1.3005
R2297 avss.n384 avss.n383 1.3005
R2298 avss.n375 avss.n273 1.3005
R2299 avss.n378 avss.n272 1.3005
R2300 avss.n379 avss.n378 1.3005
R2301 avss.n380 avss.n271 1.3005
R2302 avss.n381 avss.n380 1.3005
R2303 avss.n404 avss.n403 1.3005
R2304 avss.n405 avss.n404 1.3005
R2305 avss.n447 avss.n248 1.3005
R2306 avss.n450 avss.n449 1.3005
R2307 avss.n449 avss.n448 1.3005
R2308 avss.n407 avss.n251 1.3005
R2309 avss.n444 avss.n443 1.3005
R2310 avss.n445 avss.n444 1.3005
R2311 avss.n434 avss.n433 1.3005
R2312 avss.n437 avss.n436 1.3005
R2313 avss.n436 avss.n435 1.3005
R2314 avss.n472 avss.n234 1.3005
R2315 avss.n470 avss.n235 1.3005
R2316 avss.n471 avss.n470 1.3005
R2317 avss.n239 avss.n236 1.3005
R2318 avss.n482 avss.n239 1.3005
R2319 avss.n485 avss.n484 1.3005
R2320 avss.n484 avss.n483 1.3005
R2321 avss.n475 avss.n230 1.3005
R2322 avss.n478 avss.n229 1.3005
R2323 avss.n479 avss.n478 1.3005
R2324 avss.n480 avss.n228 1.3005
R2325 avss.n481 avss.n480 1.3005
R2326 avss.n504 avss.n503 1.3005
R2327 avss.n505 avss.n504 1.3005
R2328 avss.n547 avss.n205 1.3005
R2329 avss.n550 avss.n549 1.3005
R2330 avss.n549 avss.n548 1.3005
R2331 avss.n507 avss.n208 1.3005
R2332 avss.n544 avss.n543 1.3005
R2333 avss.n545 avss.n544 1.3005
R2334 avss.n534 avss.n533 1.3005
R2335 avss.n537 avss.n536 1.3005
R2336 avss.n536 avss.n535 1.3005
R2337 avss.n572 avss.n191 1.3005
R2338 avss.n570 avss.n192 1.3005
R2339 avss.n571 avss.n570 1.3005
R2340 avss.n196 avss.n193 1.3005
R2341 avss.n582 avss.n196 1.3005
R2342 avss.n585 avss.n584 1.3005
R2343 avss.n584 avss.n583 1.3005
R2344 avss.n575 avss.n187 1.3005
R2345 avss.n578 avss.n186 1.3005
R2346 avss.n579 avss.n578 1.3005
R2347 avss.n580 avss.n185 1.3005
R2348 avss.n581 avss.n580 1.3005
R2349 avss.n604 avss.n603 1.3005
R2350 avss.n605 avss.n604 1.3005
R2351 avss.n647 avss.n162 1.3005
R2352 avss.n650 avss.n649 1.3005
R2353 avss.n649 avss.n648 1.3005
R2354 avss.n607 avss.n165 1.3005
R2355 avss.n644 avss.n643 1.3005
R2356 avss.n645 avss.n644 1.3005
R2357 avss.n634 avss.n633 1.3005
R2358 avss.n637 avss.n636 1.3005
R2359 avss.n636 avss.n635 1.3005
R2360 avss.n672 avss.n148 1.3005
R2361 avss.n670 avss.n149 1.3005
R2362 avss.n671 avss.n670 1.3005
R2363 avss.n153 avss.n150 1.3005
R2364 avss.n682 avss.n153 1.3005
R2365 avss.n685 avss.n684 1.3005
R2366 avss.n684 avss.n683 1.3005
R2367 avss.n675 avss.n144 1.3005
R2368 avss.n678 avss.n143 1.3005
R2369 avss.n679 avss.n678 1.3005
R2370 avss.n680 avss.n142 1.3005
R2371 avss.n681 avss.n680 1.3005
R2372 avss.n697 avss.n696 1.3005
R2373 avss.n698 avss.n697 1.3005
R2374 avss.n740 avss.n739 1.3005
R2375 avss.n742 avss.n741 1.3005
R2376 avss.n741 avss.n98 1.3005
R2377 avss.n700 avss.n117 1.3005
R2378 avss.n736 avss.n735 1.3005
R2379 avss.n737 avss.n736 1.3005
R2380 avss.n726 avss.n725 1.3005
R2381 avss.n729 avss.n728 1.3005
R2382 avss.n728 avss.n727 1.3005
R2383 avss.n758 avss.n91 1.3005
R2384 avss.n761 avss.n92 1.3005
R2385 avss.n762 avss.n761 1.3005
R2386 avss.n763 avss.n93 1.3005
R2387 avss.n764 avss.n763 1.3005
R2388 avss.n767 avss.n766 1.3005
R2389 avss.n766 avss.n765 1.3005
R2390 avss.n755 avss.n87 1.3005
R2391 avss.n753 avss.n86 1.3005
R2392 avss.n754 avss.n753 1.3005
R2393 avss.n85 avss.n84 1.3005
R2394 avss.n84 avss.n53 1.3005
R2395 avss.n779 avss.n778 1.3005
R2396 avss.n780 avss.n779 1.3005
R2397 avss.n812 avss.n811 1.3005
R2398 avss.n814 avss.n813 1.3005
R2399 avss.n813 avss.n24 1.3005
R2400 avss.n782 avss.n43 1.3005
R2401 avss.n808 avss.n807 1.3005
R2402 avss.n809 avss.n808 1.3005
R2403 avss.n798 avss.n797 1.3005
R2404 avss.n801 avss.n800 1.3005
R2405 avss.n800 avss.n799 1.3005
R2406 avss.n823 avss.n16 1.3005
R2407 avss.n839 avss.n838 1.3005
R2408 avss.n838 avss.n837 1.3005
R2409 avss.n835 avss.n834 1.3005
R2410 avss.n836 avss.n835 1.3005
R2411 avss.n857 avss.n856 1.3005
R2412 avss.n856 avss.n855 1.3005
R2413 avss.n852 avss.n851 1.3005
R2414 avss.n853 avss.n852 1.3005
R2415 avss.n8 avss.n7 1.3005
R2416 avss.n819 avss.n35 0.990409
R2417 avss.n747 avss.n109 0.990409
R2418 avss.n592 avss.n158 0.990409
R2419 avss.n492 avss.n201 0.990409
R2420 avss.n392 avss.n244 0.990409
R2421 avss.n351 avss.n289 0.92075
R2422 avss.n339 avss.n338 0.92075
R2423 avss.n329 avss.n296 0.92075
R2424 avss.n313 avss.n308 0.92075
R2425 avss.n318 avss.n305 0.92075
R2426 avss.n451 avss.n247 0.92075
R2427 avss.n439 avss.n438 0.92075
R2428 avss.n429 avss.n255 0.92075
R2429 avss.n414 avss.n266 0.92075
R2430 avss.n419 avss.n263 0.92075
R2431 avss.n551 avss.n204 0.92075
R2432 avss.n539 avss.n538 0.92075
R2433 avss.n529 avss.n212 0.92075
R2434 avss.n514 avss.n223 0.92075
R2435 avss.n519 avss.n220 0.92075
R2436 avss.n651 avss.n161 0.92075
R2437 avss.n639 avss.n638 0.92075
R2438 avss.n629 avss.n169 0.92075
R2439 avss.n614 avss.n180 0.92075
R2440 avss.n619 avss.n177 0.92075
R2441 avss.n743 avss.n114 0.92075
R2442 avss.n731 avss.n730 0.92075
R2443 avss.n721 avss.n121 0.92075
R2444 avss.n707 avss.n131 0.92075
R2445 avss.n712 avss.n128 0.92075
R2446 avss.n815 avss.n40 0.92075
R2447 avss.n803 avss.n802 0.92075
R2448 avss.n793 avss.n47 0.92075
R2449 avss.n72 avss.n71 0.92075
R2450 avss.n65 avss.n64 0.92075
R2451 avss.n403 avss.n402 0.771017
R2452 avss.n503 avss.n502 0.771017
R2453 avss.n603 avss.n602 0.771017
R2454 avss.n696 avss.n695 0.771017
R2455 avss.n778 avss.n777 0.771017
R2456 avss.n354 avss.n353 0.709028
R2457 avss.n454 avss.n453 0.709028
R2458 avss.n554 avss.n553 0.709028
R2459 avss.n654 avss.n653 0.709028
R2460 avss.n746 avss.n745 0.709028
R2461 avss.n818 avss.n817 0.709028
R2462 avss.n858 avss.n857 0.471317
R2463 avss.n401 avss.n272 0.463217
R2464 avss.n402 avss.n271 0.463217
R2465 avss.n501 avss.n229 0.463217
R2466 avss.n502 avss.n228 0.463217
R2467 avss.n601 avss.n186 0.463217
R2468 avss.n602 avss.n185 0.463217
R2469 avss.n694 avss.n143 0.463217
R2470 avss.n695 avss.n142 0.463217
R2471 avss.n776 avss.n86 0.463217
R2472 avss.n777 avss.n85 0.463217
R2473 avss.n840 avss.n839 0.463217
R2474 avss.n834 avss.n2 0.463217
R2475 avss.n847 avss.n10 0.463217
R2476 avss.n846 avss.n11 0.463217
R2477 avss.n848 avss.n9 0.463217
R2478 avss.n37 avss.n36 0.463217
R2479 avss.n78 avss.n77 0.463217
R2480 avss.n770 avss.n92 0.463217
R2481 avss.n769 avss.n93 0.463217
R2482 avss.n768 avss.n767 0.463217
R2483 avss.n111 avss.n110 0.463217
R2484 avss.n136 avss.n135 0.463217
R2485 avss.n688 avss.n149 0.463217
R2486 avss.n687 avss.n150 0.463217
R2487 avss.n686 avss.n685 0.463217
R2488 avss.n656 avss.n655 0.463217
R2489 avss.n591 avss.n590 0.463217
R2490 avss.n595 avss.n192 0.463217
R2491 avss.n594 avss.n193 0.463217
R2492 avss.n593 avss.n585 0.463217
R2493 avss.n556 avss.n555 0.463217
R2494 avss.n491 avss.n490 0.463217
R2495 avss.n495 avss.n235 0.463217
R2496 avss.n494 avss.n236 0.463217
R2497 avss.n493 avss.n485 0.463217
R2498 avss.n456 avss.n455 0.463217
R2499 avss.n391 avss.n390 0.463217
R2500 avss.n395 avss.n278 0.463217
R2501 avss.n394 avss.n279 0.463217
R2502 avss.n393 avss.n385 0.463217
R2503 avss.n356 avss.n355 0.463217
R2504 avss.n851 avss.n850 0.463217
R2505 avss.n402 avss.n401 0.3083
R2506 avss.n502 avss.n501 0.3083
R2507 avss.n602 avss.n601 0.3083
R2508 avss.n695 avss.n694 0.3083
R2509 avss.n777 avss.n776 0.3083
R2510 avss.n840 avss.n2 0.3083
R2511 avss.n847 avss.n846 0.3083
R2512 avss.n848 avss.n847 0.3083
R2513 avss.n770 avss.n769 0.3083
R2514 avss.n769 avss.n768 0.3083
R2515 avss.n688 avss.n687 0.3083
R2516 avss.n687 avss.n686 0.3083
R2517 avss.n595 avss.n594 0.3083
R2518 avss.n594 avss.n593 0.3083
R2519 avss.n495 avss.n494 0.3083
R2520 avss.n494 avss.n493 0.3083
R2521 avss.n395 avss.n394 0.3083
R2522 avss.n394 avss.n393 0.3083
R2523 avss.n858 avss.n2 0.3002
R2524 avss.n1 avss.n0 0.252687
R2525 avss.n846 avss.n845 0.2165
R2526 avss.n771 avss.n770 0.2165
R2527 avss.n689 avss.n688 0.2165
R2528 avss.n596 avss.n595 0.2165
R2529 avss.n496 avss.n495 0.2165
R2530 avss.n396 avss.n395 0.2165
R2531 avss.n768 avss.n35 0.1748
R2532 avss.n593 avss.n592 0.1748
R2533 avss.n493 avss.n492 0.1748
R2534 avss.n393 avss.n392 0.1748
R2535 avss.n686 avss.n109 0.17465
R2536 avss.n849 avss.n848 0.1598
R2537 avss.n850 avss.n849 0.152487
R2538 avss.n845 avss.n844 0.148459
R2539 avss.n772 avss.n771 0.148459
R2540 avss.n690 avss.n689 0.148459
R2541 avss.n597 avss.n596 0.148459
R2542 avss.n497 avss.n496 0.148459
R2543 avss.n397 avss.n396 0.148459
R2544 avss.n136 avss.n109 0.13865
R2545 avss.n78 avss.n35 0.1385
R2546 avss.n592 avss.n591 0.1385
R2547 avss.n492 avss.n491 0.1385
R2548 avss.n392 avss.n391 0.1385
R2549 avss.n316 avss.n306 0.122607
R2550 avss.n417 avss.n264 0.122607
R2551 avss.n517 avss.n221 0.122607
R2552 avss.n617 avss.n178 0.122607
R2553 avss.n710 avss.n129 0.122607
R2554 avss.n67 avss.n59 0.122607
R2555 avss.n332 avss.n331 0.10457
R2556 avss.n432 avss.n431 0.10457
R2557 avss.n532 avss.n531 0.10457
R2558 avss.n632 avss.n631 0.10457
R2559 avss.n724 avss.n723 0.10457
R2560 avss.n796 avss.n795 0.10457
R2561 avss.n843 avss.n14 0.073981
R2562 avss.n773 avss.n89 0.073981
R2563 avss.n691 avss.n146 0.073981
R2564 avss.n598 avss.n189 0.073981
R2565 avss.n498 avss.n232 0.073981
R2566 avss.n398 avss.n275 0.073981
R2567 avss.n340 avss.n287 0.0679983
R2568 avss.n440 avss.n245 0.0679983
R2569 avss.n540 avss.n202 0.0679983
R2570 avss.n640 avss.n159 0.0679983
R2571 avss.n732 avss.n112 0.0679983
R2572 avss.n804 avss.n38 0.0679983
R2573 avss.n401 avss.n400 0.0635
R2574 avss.n501 avss.n500 0.0635
R2575 avss.n601 avss.n600 0.0635
R2576 avss.n694 avss.n693 0.0635
R2577 avss.n776 avss.n775 0.0635
R2578 avss.n841 avss.n840 0.0635
R2579 avss.n306 avss.n293 0.0622481
R2580 avss.n264 avss.n252 0.0622481
R2581 avss.n221 avss.n209 0.0622481
R2582 avss.n178 avss.n166 0.0622481
R2583 avss.n129 avss.n118 0.0622481
R2584 avss.n59 avss.n44 0.0622481
R2585 avss.n352 avss.n288 0.0568904
R2586 avss.n452 avss.n246 0.0568904
R2587 avss.n552 avss.n203 0.0568904
R2588 avss.n652 avss.n160 0.0568904
R2589 avss.n744 avss.n113 0.0568904
R2590 avss.n816 avss.n39 0.0568904
R2591 avss.n332 avss.n288 0.054837
R2592 avss.n432 avss.n246 0.054837
R2593 avss.n532 avss.n203 0.054837
R2594 avss.n632 avss.n160 0.054837
R2595 avss.n724 avss.n113 0.054837
R2596 avss.n796 avss.n39 0.054837
R2597 avss.n331 avss.n294 0.0466843
R2598 avss.n431 avss.n253 0.0466843
R2599 avss.n531 avss.n210 0.0466843
R2600 avss.n631 avss.n167 0.0466843
R2601 avss.n723 avss.n119 0.0466843
R2602 avss.n795 avss.n45 0.0466843
R2603 avss.n332 avss.n293 0.0415307
R2604 avss.n432 avss.n252 0.0415307
R2605 avss.n532 avss.n209 0.0415307
R2606 avss.n632 avss.n166 0.0415307
R2607 avss.n724 avss.n118 0.0415307
R2608 avss.n796 avss.n44 0.0415307
R2609 avss.n317 avss.n294 0.0405109
R2610 avss.n314 avss.n307 0.0405109
R2611 avss.n330 avss.n295 0.0405109
R2612 avss.n418 avss.n253 0.0405109
R2613 avss.n415 avss.n265 0.0405109
R2614 avss.n430 avss.n254 0.0405109
R2615 avss.n518 avss.n210 0.0405109
R2616 avss.n515 avss.n222 0.0405109
R2617 avss.n530 avss.n211 0.0405109
R2618 avss.n618 avss.n167 0.0405109
R2619 avss.n615 avss.n179 0.0405109
R2620 avss.n630 avss.n168 0.0405109
R2621 avss.n711 avss.n119 0.0405109
R2622 avss.n708 avss.n130 0.0405109
R2623 avss.n722 avss.n120 0.0405109
R2624 avss.n66 avss.n45 0.0405109
R2625 avss.n69 avss.n58 0.0405109
R2626 avss.n794 avss.n46 0.0405109
R2627 avss.n844 avss.n843 0.0389018
R2628 avss.n773 avss.n772 0.0389018
R2629 avss.n691 avss.n690 0.0389018
R2630 avss.n598 avss.n597 0.0389018
R2631 avss.n498 avss.n497 0.0389018
R2632 avss.n398 avss.n397 0.0389018
R2633 avss.n353 avss.n287 0.035635
R2634 avss.n453 avss.n245 0.035635
R2635 avss.n553 avss.n202 0.035635
R2636 avss.n653 avss.n159 0.035635
R2637 avss.n745 avss.n112 0.035635
R2638 avss.n817 avss.n38 0.035635
R2639 avss.n341 avss.n332 0.0349747
R2640 avss.n441 avss.n432 0.0349747
R2641 avss.n541 avss.n532 0.0349747
R2642 avss.n641 avss.n632 0.0349747
R2643 avss.n733 avss.n724 0.0349747
R2644 avss.n805 avss.n796 0.0349747
R2645 avss.n316 avss.n315 0.0322085
R2646 avss.n315 avss.n293 0.0322085
R2647 avss.n417 avss.n416 0.0322085
R2648 avss.n416 avss.n252 0.0322085
R2649 avss.n517 avss.n516 0.0322085
R2650 avss.n516 avss.n209 0.0322085
R2651 avss.n617 avss.n616 0.0322085
R2652 avss.n616 avss.n166 0.0322085
R2653 avss.n710 avss.n709 0.0322085
R2654 avss.n709 avss.n118 0.0322085
R2655 avss.n68 avss.n67 0.0322085
R2656 avss.n68 avss.n44 0.0322085
R2657 avss.n25 avss.n14 0.0258591
R2658 avss.n26 avss.n14 0.0258591
R2659 avss.n99 avss.n89 0.0258591
R2660 avss.n100 avss.n89 0.0258591
R2661 avss.n661 avss.n146 0.0258591
R2662 avss.n664 avss.n146 0.0258591
R2663 avss.n561 avss.n189 0.0258591
R2664 avss.n564 avss.n189 0.0258591
R2665 avss.n461 avss.n232 0.0258591
R2666 avss.n464 avss.n232 0.0258591
R2667 avss.n361 avss.n275 0.0258591
R2668 avss.n364 avss.n275 0.0258591
R2669 avss.n843 avss.n842 0.023066
R2670 avss.n774 avss.n773 0.023066
R2671 avss.n692 avss.n691 0.023066
R2672 avss.n599 avss.n598 0.023066
R2673 avss.n499 avss.n498 0.023066
R2674 avss.n399 avss.n398 0.023066
R2675 avss.n317 avss.n316 0.0214837
R2676 avss.n315 avss.n295 0.0214837
R2677 avss.n418 avss.n417 0.0214837
R2678 avss.n416 avss.n254 0.0214837
R2679 avss.n518 avss.n517 0.0214837
R2680 avss.n516 avss.n211 0.0214837
R2681 avss.n618 avss.n617 0.0214837
R2682 avss.n616 avss.n168 0.0214837
R2683 avss.n711 avss.n710 0.0214837
R2684 avss.n709 avss.n120 0.0214837
R2685 avss.n67 avss.n66 0.0214837
R2686 avss.n68 avss.n46 0.0214837
R2687 avss.n819 avss.n818 0.0196349
R2688 avss.n747 avss.n746 0.0196349
R2689 avss.n654 avss.n158 0.0196349
R2690 avss.n554 avss.n201 0.0196349
R2691 avss.n454 avss.n244 0.0196349
R2692 avss.n842 avss.n15 0.0163358
R2693 avss.n774 avss.n88 0.0163358
R2694 avss.n692 avss.n145 0.0163358
R2695 avss.n599 avss.n188 0.0163358
R2696 avss.n499 avss.n231 0.0163358
R2697 avss.n399 avss.n274 0.0163358
R2698 avss.n37 avss.n15 0.0139604
R2699 avss.n111 avss.n88 0.0139604
R2700 avss.n655 avss.n145 0.0139604
R2701 avss.n555 avss.n188 0.0139604
R2702 avss.n455 avss.n231 0.0139604
R2703 avss.n355 avss.n274 0.0139604
R2704 avss.n818 avss.n37 0.0130367
R2705 avss.n746 avss.n111 0.0130367
R2706 avss.n655 avss.n654 0.0130367
R2707 avss.n555 avss.n554 0.0130367
R2708 avss.n455 avss.n454 0.0130367
R2709 avss.n355 avss.n354 0.0130367
R2710 avss.n315 avss.n314 0.0121902
R2711 avss.n416 avss.n415 0.0121902
R2712 avss.n516 avss.n515 0.0121902
R2713 avss.n616 avss.n615 0.0121902
R2714 avss.n709 avss.n708 0.0121902
R2715 avss.n69 avss.n68 0.0121902
R2716 avss.n849 avss 0.0118245
R2717 avss.n307 avss.n306 0.00915761
R2718 avss.n265 avss.n264 0.00915761
R2719 avss.n222 avss.n221 0.00915761
R2720 avss.n179 avss.n178 0.00915761
R2721 avss.n130 avss.n129 0.00915761
R2722 avss.n59 avss.n58 0.00915761
R2723 avss.n331 avss.n330 0.00720109
R2724 avss.n431 avss.n430 0.00720109
R2725 avss.n531 avss.n530 0.00720109
R2726 avss.n631 avss.n630 0.00720109
R2727 avss.n723 avss.n722 0.00720109
R2728 avss.n795 avss.n794 0.00720109
R2729 avss.n353 avss.n352 0.00511663
R2730 avss.n453 avss.n452 0.00511663
R2731 avss.n553 avss.n552 0.00511663
R2732 avss.n653 avss.n652 0.00511663
R2733 avss.n745 avss.n744 0.00511663
R2734 avss.n817 avss.n816 0.00511663
R2735 avss.n341 avss.n340 0.000544599
R2736 avss.n441 avss.n440 0.000544599
R2737 avss.n541 avss.n540 0.000544599
R2738 avss.n641 avss.n640 0.000544599
R2739 avss.n733 avss.n732 0.000544599
R2740 avss.n805 avss.n804 0.000544599
R2741 a_48650_3501.n0 a_48650_3501.t4 34.1797
R2742 a_48650_3501.n0 a_48650_3501.t5 19.5798
R2743 a_48650_3501.n1 a_48650_3501.t3 18.7717
R2744 a_48650_3501.n1 a_48650_3501.t1 9.2885
R2745 a_48650_3501.n2 a_48650_3501.n0 4.93379
R2746 a_48650_3501.t0 a_48650_3501.n3 4.23346
R2747 a_48650_3501.n3 a_48650_3501.t2 3.85546
R2748 a_48650_3501.n2 a_48650_3501.n1 0.4055
R2749 a_48650_3501.n3 a_48650_3501.n2 0.352625
R2750 a_6520_1558.n0 a_6520_1558.t5 40.8177
R2751 a_6520_1558.n1 a_6520_1558.t4 40.6313
R2752 a_6520_1558.n1 a_6520_1558.t6 27.3166
R2753 a_6520_1558.n0 a_6520_1558.t7 27.1302
R2754 a_6520_1558.n2 a_6520_1558.n1 19.2576
R2755 a_6520_1558.n3 a_6520_1558.t1 10.0473
R2756 a_6520_1558.t0 a_6520_1558.n5 6.51042
R2757 a_6520_1558.n5 a_6520_1558.n4 6.04952
R2758 a_6520_1558.n2 a_6520_1558.n0 5.91752
R2759 a_6520_1558.n3 a_6520_1558.n2 4.89565
R2760 a_6520_1558.n5 a_6520_1558.n3 0.732092
R2761 a_6520_1558.n4 a_6520_1558.t3 0.7285
R2762 a_6520_1558.n4 a_6520_1558.t2 0.7285
R2763 a_6600_2510.n0 a_6600_2510.t4 41.0041
R2764 a_6600_2510.n1 a_6600_2510.t5 40.8177
R2765 a_6600_2510.n1 a_6600_2510.t7 27.1302
R2766 a_6600_2510.n0 a_6600_2510.t6 26.9438
R2767 a_6600_2510.n2 a_6600_2510.n1 22.5284
R2768 a_6600_2510.n3 a_6600_2510.n2 19.5781
R2769 a_6600_2510.n3 a_6600_2510.t1 10.0473
R2770 a_6600_2510.n4 a_6600_2510.t3 6.51042
R2771 a_6600_2510.n5 a_6600_2510.n4 6.04952
R2772 a_6600_2510.n2 a_6600_2510.n0 5.7305
R2773 a_6600_2510.n4 a_6600_2510.n3 0.732092
R2774 a_6600_2510.t0 a_6600_2510.n5 0.7285
R2775 a_6600_2510.n5 a_6600_2510.t2 0.7285
R2776 a_6520_3763.n1 a_6520_3763.t9 41.0041
R2777 a_6520_3763.n0 a_6520_3763.t5 40.8177
R2778 a_6520_3763.n2 a_6520_3763.t4 40.6313
R2779 a_6520_3763.n2 a_6520_3763.t7 27.3166
R2780 a_6520_3763.n0 a_6520_3763.t8 27.1302
R2781 a_6520_3763.n1 a_6520_3763.t6 26.9438
R2782 a_6520_3763.n3 a_6520_3763.n1 15.6312
R2783 a_6520_3763.n3 a_6520_3763.n2 15.046
R2784 a_6520_3763.n5 a_6520_3763.t3 10.0473
R2785 a_6520_3763.n6 a_6520_3763.t2 6.51042
R2786 a_6520_3763.n7 a_6520_3763.n6 6.04952
R2787 a_6520_3763.n4 a_6520_3763.n0 5.64619
R2788 a_6520_3763.n5 a_6520_3763.n4 5.17851
R2789 a_6520_3763.n4 a_6520_3763.n3 4.5005
R2790 a_6520_3763.n6 a_6520_3763.n5 0.732092
R2791 a_6520_3763.t0 a_6520_3763.n7 0.7285
R2792 a_6520_3763.n7 a_6520_3763.t1 0.7285
R2793 dffrs_1.Q.n3 dffrs_1.Q.t7 40.6313
R2794 dffrs_1.Q.n1 dffrs_1.Q.t4 34.1066
R2795 dffrs_1.Q.n3 dffrs_1.Q.t5 27.3166
R2796 dffrs_1.Q.n0 dffrs_1.Q.t6 19.673
R2797 dffrs_1.Q.n0 dffrs_1.Q.t8 19.4007
R2798 dffrs_1.Q.n7 dffrs_1.Q.n3 14.6967
R2799 dffrs_1.Q.n6 dffrs_1.Q.t2 10.0473
R2800 dffrs_1.Q.n7 dffrs_1.Q.n6 9.39565
R2801 dffrs_1.Q.n2 dffrs_1.Q.n1 6.70486
R2802 dffrs_1.Q.n5 dffrs_1.Q.t1 6.51042
R2803 dffrs_1.Q.n5 dffrs_1.Q.n4 6.04952
R2804 dffrs_1.Q dffrs_1.Q.n2 5.81354
R2805 dffrs_1.Q.n6 dffrs_1.Q.n5 0.732092
R2806 dffrs_1.Q.n4 dffrs_1.Q.t3 0.7285
R2807 dffrs_1.Q.n4 dffrs_1.Q.t0 0.7285
R2808 dffrs_1.Q dffrs_1.Q.n7 0.458082
R2809 dffrs_1.Q.n1 dffrs_1.Q.n0 0.252687
R2810 dffrs_1.Q.n2 2inmux_3.Bit 0.0519286
R2811 a_20234_3501.n0 a_20234_3501.t5 34.1797
R2812 a_20234_3501.n0 a_20234_3501.t4 19.5798
R2813 a_20234_3501.n3 a_20234_3501.t2 18.7717
R2814 a_20234_3501.t0 a_20234_3501.n3 9.2885
R2815 a_20234_3501.n2 a_20234_3501.n0 4.93379
R2816 a_20234_3501.n1 a_20234_3501.t1 4.23346
R2817 a_20234_3501.n1 a_20234_3501.t3 3.85546
R2818 a_20234_3501.n3 a_20234_3501.n2 0.4055
R2819 a_20234_3501.n2 a_20234_3501.n1 0.352625
R2820 2inmux_2.Bit.n3 2inmux_2.Bit.t6 40.6313
R2821 2inmux_2.Bit.n1 2inmux_2.Bit.t5 34.1066
R2822 2inmux_2.Bit.n3 2inmux_2.Bit.t8 27.3166
R2823 2inmux_2.Bit.n0 2inmux_2.Bit.t7 19.673
R2824 2inmux_2.Bit.n0 2inmux_2.Bit.t4 19.4007
R2825 2inmux_2.Bit.n7 2inmux_2.Bit.n3 14.6967
R2826 2inmux_2.Bit.n6 2inmux_2.Bit.t0 10.0473
R2827 2inmux_2.Bit.n7 2inmux_2.Bit.n6 9.39565
R2828 2inmux_2.Bit.n2 2inmux_2.Bit.n1 6.70486
R2829 2inmux_2.Bit.n5 2inmux_2.Bit.t1 6.51042
R2830 2inmux_2.Bit.n5 2inmux_2.Bit.n4 6.04952
R2831 dffrs_0.Q 2inmux_2.Bit.n2 5.81514
R2832 2inmux_2.Bit.n6 2inmux_2.Bit.n5 0.732092
R2833 2inmux_2.Bit.n4 2inmux_2.Bit.t2 0.7285
R2834 2inmux_2.Bit.n4 2inmux_2.Bit.t3 0.7285
R2835 dffrs_0.Q 2inmux_2.Bit.n7 0.458082
R2836 2inmux_2.Bit.n1 2inmux_2.Bit.n0 0.252687
R2837 2inmux_2.Bit.n2 2inmux_2.Bit 0.0519286
R2838 a_1290_3500.n0 a_1290_3500.t4 34.1797
R2839 a_1290_3500.n0 a_1290_3500.t5 19.5798
R2840 a_1290_3500.t0 a_1290_3500.n3 18.7717
R2841 a_1290_3500.n3 a_1290_3500.t1 9.2885
R2842 a_1290_3500.n2 a_1290_3500.n0 4.93379
R2843 a_1290_3500.n1 a_1290_3500.t3 4.23346
R2844 a_1290_3500.n1 a_1290_3500.t2 3.85546
R2845 a_1290_3500.n3 a_1290_3500.n2 0.4055
R2846 a_1290_3500.n2 a_1290_3500.n1 0.352625
R2847 clk.n3 clk.t18 41.0041
R2848 clk.n7 clk.t12 41.0041
R2849 clk.n11 clk.t1 41.0041
R2850 clk.n15 clk.t15 41.0041
R2851 clk.n19 clk.t3 41.0041
R2852 clk.n0 clk.t17 41.0041
R2853 clk.n4 clk.t2 40.8177
R2854 clk.n8 clk.t22 40.8177
R2855 clk.n12 clk.t11 40.8177
R2856 clk.n16 clk.t8 40.8177
R2857 clk.n20 clk.t20 40.8177
R2858 clk.n1 clk.t10 40.8177
R2859 clk.n4 clk.t13 27.1302
R2860 clk.n8 clk.t9 27.1302
R2861 clk.n12 clk.t23 27.1302
R2862 clk.n16 clk.t19 27.1302
R2863 clk.n20 clk.t5 27.1302
R2864 clk.n1 clk.t21 27.1302
R2865 clk.n3 clk.t7 26.9438
R2866 clk.n7 clk.t0 26.9438
R2867 clk.n11 clk.t14 26.9438
R2868 clk.n15 clk.t4 26.9438
R2869 clk.n19 clk.t16 26.9438
R2870 clk.n0 clk.t6 26.9438
R2871 dffrs_5.clk clk.n22 23.2034
R2872 clk.n10 clk.n6 13.9468
R2873 clk.n14 clk.n10 13.9463
R2874 clk.n22 clk.n18 13.9457
R2875 clk.n18 clk.n14 13.9457
R2876 clk.n6 dffrs_0.clk 9.25764
R2877 clk.n10 dffrs_1.clk 9.25764
R2878 clk.n14 dffrs_2.clk 9.25764
R2879 clk.n18 dffrs_3.clk 9.25764
R2880 clk.n22 dffrs_4.clk 9.25764
R2881 clk.n5 clk.n4 7.65746
R2882 clk.n9 clk.n8 7.65746
R2883 clk.n13 clk.n12 7.65746
R2884 clk.n17 clk.n16 7.65746
R2885 clk.n21 clk.n20 7.65746
R2886 clk.n2 clk.n1 7.65746
R2887 clk.n5 clk.n3 7.12229
R2888 clk.n9 clk.n7 7.12229
R2889 clk.n13 clk.n11 7.12229
R2890 clk.n17 clk.n15 7.12229
R2891 clk.n21 clk.n19 7.12229
R2892 clk.n2 clk.n0 7.12229
R2893 clk.n6 clk 3.54742
R2894 dffrs_0.clk clk.n5 0.611214
R2895 dffrs_1.clk clk.n9 0.611214
R2896 dffrs_2.clk clk.n13 0.611214
R2897 dffrs_3.clk clk.n17 0.611214
R2898 dffrs_4.clk clk.n21 0.611214
R2899 dffrs_5.clk clk.n2 0.611214
R2900 a_15992_3763.n1 a_15992_3763.t7 41.0041
R2901 a_15992_3763.n0 a_15992_3763.t5 40.8177
R2902 a_15992_3763.n2 a_15992_3763.t6 40.6313
R2903 a_15992_3763.n2 a_15992_3763.t9 27.3166
R2904 a_15992_3763.n0 a_15992_3763.t8 27.1302
R2905 a_15992_3763.n1 a_15992_3763.t4 26.9438
R2906 a_15992_3763.n3 a_15992_3763.n1 15.6312
R2907 a_15992_3763.n3 a_15992_3763.n2 15.046
R2908 a_15992_3763.n5 a_15992_3763.t1 10.0473
R2909 a_15992_3763.t0 a_15992_3763.n7 6.51042
R2910 a_15992_3763.n7 a_15992_3763.n6 6.04952
R2911 a_15992_3763.n4 a_15992_3763.n0 5.64619
R2912 a_15992_3763.n5 a_15992_3763.n4 5.17851
R2913 a_15992_3763.n4 a_15992_3763.n3 4.5005
R2914 a_15992_3763.n7 a_15992_3763.n5 0.732092
R2915 a_15992_3763.n6 a_15992_3763.t2 0.7285
R2916 a_15992_3763.n6 a_15992_3763.t3 0.7285
R2917 2inmux_1.Bit.n3 2inmux_1.Bit.t8 40.6313
R2918 2inmux_1.Bit.n1 2inmux_1.Bit.t7 34.1066
R2919 2inmux_1.Bit.n3 2inmux_1.Bit.t5 27.3166
R2920 2inmux_1.Bit.n0 2inmux_1.Bit.t4 19.673
R2921 2inmux_1.Bit.n0 2inmux_1.Bit.t6 19.4007
R2922 2inmux_1.Bit.n7 2inmux_1.Bit.n3 14.6967
R2923 2inmux_1.Bit.n6 2inmux_1.Bit.t2 10.0473
R2924 2inmux_1.Bit.n7 2inmux_1.Bit.n6 9.39565
R2925 2inmux_1.Bit.n2 2inmux_1.Bit.n1 6.70486
R2926 2inmux_1.Bit.n5 2inmux_1.Bit.t3 6.51042
R2927 2inmux_1.Bit.n5 2inmux_1.Bit.n4 6.04952
R2928 dffrs_4.Q 2inmux_1.Bit.n2 5.81514
R2929 2inmux_1.Bit.n6 2inmux_1.Bit.n5 0.732092
R2930 2inmux_1.Bit.n4 2inmux_1.Bit.t1 0.7285
R2931 2inmux_1.Bit.n4 2inmux_1.Bit.t0 0.7285
R2932 dffrs_4.Q 2inmux_1.Bit.n7 0.458082
R2933 2inmux_1.Bit.n1 2inmux_1.Bit.n0 0.252687
R2934 2inmux_1.Bit.n2 2inmux_1.Bit 0.0519286
R2935 a_15992_5968.n2 a_15992_5968.t5 40.6313
R2936 a_15992_5968.n2 a_15992_5968.t4 27.3166
R2937 a_15992_5968.n3 a_15992_5968.n2 24.1527
R2938 a_15992_5968.t0 a_15992_5968.n3 10.0473
R2939 a_15992_5968.n1 a_15992_5968.t1 6.51042
R2940 a_15992_5968.n1 a_15992_5968.n0 6.04952
R2941 a_15992_5968.n3 a_15992_5968.n1 0.732092
R2942 a_15992_5968.n0 a_15992_5968.t3 0.7285
R2943 a_15992_5968.n0 a_15992_5968.t2 0.7285
R2944 load.n4 load.t17 34.2529
R2945 load.n10 load.t23 34.2529
R2946 load.n16 load.t28 34.2529
R2947 load.n22 load.t13 34.2529
R2948 load.n28 load.t0 34.2529
R2949 load.n1 load.t9 34.2529
R2950 load.n6 load.t20 34.1797
R2951 load.n12 load.t19 34.1797
R2952 load.n18 load.t14 34.1797
R2953 load.n24 load.t1 34.1797
R2954 load.n30 load.t26 34.1797
R2955 load.n2 load.t3 34.1797
R2956 load.n3 load.t2 19.673
R2957 load.n9 load.t5 19.673
R2958 load.n15 load.t4 19.673
R2959 load.n21 load.t18 19.673
R2960 load.n27 load.t7 19.673
R2961 load.n0 load.t25 19.673
R2962 load.n6 load.t12 19.5798
R2963 load.n12 load.t11 19.5798
R2964 load.n18 load.t6 19.5798
R2965 load.n24 load.t22 19.5798
R2966 load.n30 load.t16 19.5798
R2967 load.n2 load.t24 19.5798
R2968 load.n3 load.t15 19.4007
R2969 load.n9 load.t21 19.4007
R2970 load.n15 load.t27 19.4007
R2971 load.n21 load.t10 19.4007
R2972 load.n27 load.t29 19.4007
R2973 load.n0 load.t8 19.4007
R2974 load.n33 load.n32 15.5531
R2975 load.n8 load.n7 8.46371
R2976 load.n20 load.n19 8.37371
R2977 load.n14 load.n13 8.32871
R2978 load.n26 load.n25 8.32871
R2979 load.n32 load.n31 8.32871
R2980 load.n5 load.n4 7.87164
R2981 load.n11 load.n10 7.87164
R2982 load.n17 load.n16 7.87164
R2983 load.n23 load.n22 7.87164
R2984 load.n29 load.n28 7.87164
R2985 load.n34 load.n1 7.87164
R2986 load.n14 load.n8 7.26762
R2987 load.n32 load.n26 7.22491
R2988 load.n26 load.n20 7.22491
R2989 load.n20 load.n14 7.22491
R2990 load.n7 load.n6 5.00771
R2991 load.n19 load.n18 5.00771
R2992 load.n13 load.n12 4.96432
R2993 load.n25 load.n24 4.96432
R2994 load.n31 load.n30 4.96432
R2995 load.n33 load.n2 4.96432
R2996 load.n13 load.n11 2.11068
R2997 load.n25 load.n23 2.11068
R2998 load.n31 load.n29 2.11068
R2999 load.n34 load.n33 2.11068
R3000 load.n7 load.n5 2.06729
R3001 load.n19 load.n17 2.06729
R3002 load.n5 2inmux_0.Load 0.2255
R3003 load.n11 2inmux_2.Load 0.2255
R3004 load.n17 2inmux_3.Load 0.2255
R3005 load.n23 2inmux_4.Load 0.2255
R3006 load.n29 2inmux_5.Load 0.2255
R3007 2inmux_1.Load load.n34 0.2255
R3008 load.n8 load 0.211008
R3009 load.n4 load.n3 0.106438
R3010 load.n10 load.n9 0.106438
R3011 load.n16 load.n15 0.106438
R3012 load.n22 load.n21 0.106438
R3013 load.n28 load.n27 0.106438
R3014 load.n1 load.n0 0.106438
R3015 a_39178_3501.n0 a_39178_3501.t5 34.1797
R3016 a_39178_3501.n0 a_39178_3501.t4 19.5798
R3017 a_39178_3501.n1 a_39178_3501.t3 18.7717
R3018 a_39178_3501.n1 a_39178_3501.t2 9.2885
R3019 a_39178_3501.n2 a_39178_3501.n0 4.93379
R3020 a_39178_3501.t0 a_39178_3501.n3 4.23346
R3021 a_39178_3501.n3 a_39178_3501.t1 3.85546
R3022 a_39178_3501.n2 a_39178_3501.n1 0.4055
R3023 a_39178_3501.n3 a_39178_3501.n2 0.352625
R3024 dffrs_2.Q.n3 dffrs_2.Q.t8 40.6313
R3025 dffrs_2.Q.n1 dffrs_2.Q.t7 34.1066
R3026 dffrs_2.Q.n3 dffrs_2.Q.t5 27.3166
R3027 dffrs_2.Q.n0 dffrs_2.Q.t4 19.673
R3028 dffrs_2.Q.n0 dffrs_2.Q.t6 19.4007
R3029 dffrs_2.Q.n7 dffrs_2.Q.n3 14.6967
R3030 dffrs_2.Q.n6 dffrs_2.Q.t0 10.0473
R3031 dffrs_2.Q.n7 dffrs_2.Q.n6 9.39565
R3032 dffrs_2.Q.n2 dffrs_2.Q.n1 6.70486
R3033 dffrs_2.Q.n5 dffrs_2.Q.t1 6.51042
R3034 dffrs_2.Q.n5 dffrs_2.Q.n4 6.04952
R3035 dffrs_2.Q dffrs_2.Q.n2 5.81514
R3036 dffrs_2.Q.n6 dffrs_2.Q.n5 0.732092
R3037 dffrs_2.Q.n4 dffrs_2.Q.t3 0.7285
R3038 dffrs_2.Q.n4 dffrs_2.Q.t2 0.7285
R3039 dffrs_2.Q dffrs_2.Q.n7 0.458082
R3040 dffrs_2.Q.n1 dffrs_2.Q.n0 0.252687
R3041 dffrs_2.Q.n2 2inmux_4.Bit 0.0519286
R3042 a_48650_1161.n0 a_48650_1161.t5 34.1797
R3043 a_48650_1161.n0 a_48650_1161.t4 19.5798
R3044 a_48650_1161.t0 a_48650_1161.n3 18.7717
R3045 a_48650_1161.n3 a_48650_1161.t2 9.2885
R3046 a_48650_1161.n2 a_48650_1161.n0 4.93379
R3047 a_48650_1161.n1 a_48650_1161.t3 4.23346
R3048 a_48650_1161.n1 a_48650_1161.t1 3.85546
R3049 a_48650_1161.n3 a_48650_1161.n2 0.4055
R3050 a_48650_1161.n2 a_48650_1161.n1 0.352625
R3051 a_50878_1605.n0 a_50878_1605.t5 34.1797
R3052 a_50878_1605.n0 a_50878_1605.t4 19.5798
R3053 a_50878_1605.t0 a_50878_1605.n3 10.3401
R3054 a_50878_1605.n3 a_50878_1605.t3 9.2885
R3055 a_50878_1605.n2 a_50878_1605.n0 4.93379
R3056 a_50878_1605.n1 a_50878_1605.t2 4.09202
R3057 a_50878_1605.n1 a_50878_1605.t1 3.95079
R3058 a_50878_1605.n3 a_50878_1605.n2 0.599711
R3059 a_50878_1605.n2 a_50878_1605.n1 0.296375
R3060 2inmux_1.OUT.n0 2inmux_1.OUT.t2 41.0041
R3061 2inmux_1.OUT.n0 2inmux_1.OUT.t3 26.9438
R3062 2inmux_1.OUT.n1 2inmux_1.OUT.t1 9.6935
R3063 dffrs_5.d 2inmux_1.OUT.n0 6.55979
R3064 2inmux_1.OUT dffrs_5.d 4.883
R3065 2inmux_1.OUT.n1 2inmux_1.OUT.t0 4.35383
R3066 2inmux_1.OUT 2inmux_1.OUT.n1 0.350857
R3067 a_22462_1605.n0 a_22462_1605.t5 34.1797
R3068 a_22462_1605.n0 a_22462_1605.t4 19.5798
R3069 a_22462_1605.t0 a_22462_1605.n3 10.3401
R3070 a_22462_1605.n3 a_22462_1605.t3 9.2885
R3071 a_22462_1605.n2 a_22462_1605.n0 4.93379
R3072 a_22462_1605.n1 a_22462_1605.t1 4.09202
R3073 a_22462_1605.n1 a_22462_1605.t2 3.95079
R3074 a_22462_1605.n3 a_22462_1605.n2 0.599711
R3075 a_22462_1605.n2 a_22462_1605.n1 0.296375
R3076 a_34936_1559.n0 a_34936_1559.t5 40.8177
R3077 a_34936_1559.n1 a_34936_1559.t6 40.6313
R3078 a_34936_1559.n1 a_34936_1559.t4 27.3166
R3079 a_34936_1559.n0 a_34936_1559.t7 27.1302
R3080 a_34936_1559.n2 a_34936_1559.n1 19.2576
R3081 a_34936_1559.n3 a_34936_1559.t2 10.0473
R3082 a_34936_1559.n4 a_34936_1559.t3 6.51042
R3083 a_34936_1559.n5 a_34936_1559.n4 6.04952
R3084 a_34936_1559.n2 a_34936_1559.n0 5.91752
R3085 a_34936_1559.n3 a_34936_1559.n2 4.89565
R3086 a_34936_1559.n4 a_34936_1559.n3 0.732092
R3087 a_34936_1559.t0 a_34936_1559.n5 0.7285
R3088 a_34936_1559.n5 a_34936_1559.t1 0.7285
R3089 a_34936_3764.n1 a_34936_3764.t8 41.0041
R3090 a_34936_3764.n0 a_34936_3764.t6 40.8177
R3091 a_34936_3764.n2 a_34936_3764.t7 40.6313
R3092 a_34936_3764.n2 a_34936_3764.t4 27.3166
R3093 a_34936_3764.n0 a_34936_3764.t9 27.1302
R3094 a_34936_3764.n1 a_34936_3764.t5 26.9438
R3095 a_34936_3764.n3 a_34936_3764.n1 15.6312
R3096 a_34936_3764.n3 a_34936_3764.n2 15.046
R3097 a_34936_3764.n5 a_34936_3764.t1 10.0473
R3098 a_34936_3764.t0 a_34936_3764.n7 6.51042
R3099 a_34936_3764.n7 a_34936_3764.n6 6.04952
R3100 a_34936_3764.n4 a_34936_3764.n0 5.64619
R3101 a_34936_3764.n5 a_34936_3764.n4 5.17851
R3102 a_34936_3764.n4 a_34936_3764.n3 4.5005
R3103 a_34936_3764.n7 a_34936_3764.n5 0.732092
R3104 a_34936_3764.n6 a_34936_3764.t2 0.7285
R3105 a_34936_3764.n6 a_34936_3764.t3 0.7285
R3106 a_3518_1604.n0 a_3518_1604.t5 34.1797
R3107 a_3518_1604.n0 a_3518_1604.t4 19.5798
R3108 a_3518_1604.n3 a_3518_1604.t3 10.3401
R3109 a_3518_1604.t0 a_3518_1604.n3 9.2885
R3110 a_3518_1604.n2 a_3518_1604.n0 4.93379
R3111 a_3518_1604.n1 a_3518_1604.t2 4.09202
R3112 a_3518_1604.n1 a_3518_1604.t1 3.95079
R3113 a_3518_1604.n3 a_3518_1604.n2 0.599711
R3114 a_3518_1604.n2 a_3518_1604.n1 0.296375
R3115 2inmux_0.OUT.n0 2inmux_0.OUT.t2 41.0041
R3116 2inmux_0.OUT.n0 2inmux_0.OUT.t3 26.9438
R3117 2inmux_0.OUT.n1 2inmux_0.OUT.t1 9.6935
R3118 dffrs_0.d 2inmux_0.OUT.n0 6.55979
R3119 2inmux_0.OUT dffrs_0.d 4.883
R3120 2inmux_0.OUT.n1 2inmux_0.OUT.t0 4.35383
R3121 2inmux_0.OUT 2inmux_0.OUT.n1 0.350857
R3122 a_44408_3764.n1 a_44408_3764.t6 41.0041
R3123 a_44408_3764.n0 a_44408_3764.t5 40.8177
R3124 a_44408_3764.n2 a_44408_3764.t4 40.6313
R3125 a_44408_3764.n2 a_44408_3764.t7 27.3166
R3126 a_44408_3764.n0 a_44408_3764.t9 27.1302
R3127 a_44408_3764.n1 a_44408_3764.t8 26.9438
R3128 a_44408_3764.n3 a_44408_3764.n1 15.6312
R3129 a_44408_3764.n3 a_44408_3764.n2 15.046
R3130 a_44408_3764.n5 a_44408_3764.t1 10.0473
R3131 a_44408_3764.t0 a_44408_3764.n7 6.51042
R3132 a_44408_3764.n7 a_44408_3764.n6 6.04952
R3133 a_44408_3764.n4 a_44408_3764.n0 5.64619
R3134 a_44408_3764.n5 a_44408_3764.n4 5.17851
R3135 a_44408_3764.n4 a_44408_3764.n3 4.5005
R3136 a_44408_3764.n7 a_44408_3764.n5 0.732092
R3137 a_44408_3764.n6 a_44408_3764.t2 0.7285
R3138 a_44408_3764.n6 a_44408_3764.t3 0.7285
R3139 a_20234_1161.n0 a_20234_1161.t4 34.1797
R3140 a_20234_1161.n0 a_20234_1161.t5 19.5798
R3141 a_20234_1161.t0 a_20234_1161.n3 18.7717
R3142 a_20234_1161.n3 a_20234_1161.t3 9.2885
R3143 a_20234_1161.n2 a_20234_1161.n0 4.93379
R3144 a_20234_1161.n1 a_20234_1161.t1 4.23346
R3145 a_20234_1161.n1 a_20234_1161.t2 3.85546
R3146 a_20234_1161.n3 a_20234_1161.n2 0.4055
R3147 a_20234_1161.n2 a_20234_1161.n1 0.352625
R3148 a_29706_1161.n0 a_29706_1161.t4 34.1797
R3149 a_29706_1161.n0 a_29706_1161.t5 19.5798
R3150 a_29706_1161.n1 a_29706_1161.t2 18.7717
R3151 a_29706_1161.n1 a_29706_1161.t1 9.2885
R3152 a_29706_1161.n2 a_29706_1161.n0 4.93379
R3153 a_29706_1161.t0 a_29706_1161.n3 4.23346
R3154 a_29706_1161.n3 a_29706_1161.t3 3.85546
R3155 a_29706_1161.n2 a_29706_1161.n1 0.4055
R3156 a_29706_1161.n3 a_29706_1161.n2 0.352625
R3157 a_25464_3764.n1 a_25464_3764.t5 41.0041
R3158 a_25464_3764.n0 a_25464_3764.t4 40.8177
R3159 a_25464_3764.n2 a_25464_3764.t6 40.6313
R3160 a_25464_3764.n2 a_25464_3764.t9 27.3166
R3161 a_25464_3764.n0 a_25464_3764.t8 27.1302
R3162 a_25464_3764.n1 a_25464_3764.t7 26.9438
R3163 a_25464_3764.n3 a_25464_3764.n1 15.6312
R3164 a_25464_3764.n3 a_25464_3764.n2 15.046
R3165 a_25464_3764.n5 a_25464_3764.t1 10.0473
R3166 a_25464_3764.t0 a_25464_3764.n7 6.51042
R3167 a_25464_3764.n7 a_25464_3764.n6 6.04952
R3168 a_25464_3764.n4 a_25464_3764.n0 5.64619
R3169 a_25464_3764.n5 a_25464_3764.n4 5.17851
R3170 a_25464_3764.n4 a_25464_3764.n3 4.5005
R3171 a_25464_3764.n7 a_25464_3764.n5 0.732092
R3172 a_25464_3764.n6 a_25464_3764.t2 0.7285
R3173 a_25464_3764.n6 a_25464_3764.t3 0.7285
R3174 B6.n1 B6.t1 34.2529
R3175 B6.n0 B6.t0 19.673
R3176 B6.n0 B6.t2 19.4007
R3177 B6.n2 B6.n1 8.05164
R3178 B6.n2 B6 1.87121
R3179 B6.n1 B6.n0 0.106438
R3180 2inmux_0.In B6.n2 0.0455
R3181 a_1290_1160.n0 a_1290_1160.t5 34.1797
R3182 a_1290_1160.n0 a_1290_1160.t4 19.5798
R3183 a_1290_1160.n1 a_1290_1160.t3 18.7717
R3184 a_1290_1160.n1 a_1290_1160.t2 9.2885
R3185 a_1290_1160.n2 a_1290_1160.n0 4.93379
R3186 a_1290_1160.t0 a_1290_1160.n3 4.23346
R3187 a_1290_1160.n3 a_1290_1160.t1 3.85546
R3188 a_1290_1160.n2 a_1290_1160.n1 0.4055
R3189 a_1290_1160.n3 a_1290_1160.n2 0.352625
R3190 a_10762_3500.n0 a_10762_3500.t5 34.1797
R3191 a_10762_3500.n0 a_10762_3500.t4 19.5798
R3192 a_10762_3500.n1 a_10762_3500.t2 18.7717
R3193 a_10762_3500.n1 a_10762_3500.t1 9.2885
R3194 a_10762_3500.n2 a_10762_3500.n0 4.93379
R3195 a_10762_3500.n3 a_10762_3500.t3 4.23346
R3196 a_10762_3500.t0 a_10762_3500.n3 3.85546
R3197 a_10762_3500.n2 a_10762_3500.n1 0.4055
R3198 a_10762_3500.n3 a_10762_3500.n2 0.352625
R3199 a_35016_2511.n0 a_35016_2511.t5 41.0041
R3200 a_35016_2511.n1 a_35016_2511.t6 40.8177
R3201 a_35016_2511.n1 a_35016_2511.t4 27.1302
R3202 a_35016_2511.n0 a_35016_2511.t7 26.9438
R3203 a_35016_2511.n2 a_35016_2511.n1 22.5284
R3204 a_35016_2511.n3 a_35016_2511.n2 19.5781
R3205 a_35016_2511.n3 a_35016_2511.t3 10.0473
R3206 a_35016_2511.n4 a_35016_2511.t2 6.51042
R3207 a_35016_2511.n5 a_35016_2511.n4 6.04952
R3208 a_35016_2511.n2 a_35016_2511.n0 5.7305
R3209 a_35016_2511.n4 a_35016_2511.n3 0.732092
R3210 a_35016_2511.n5 a_35016_2511.t1 0.7285
R3211 a_35016_2511.t0 a_35016_2511.n5 0.7285
R3212 a_41406_1605.n0 a_41406_1605.t5 34.1797
R3213 a_41406_1605.n0 a_41406_1605.t4 19.5798
R3214 a_41406_1605.t0 a_41406_1605.n3 10.3401
R3215 a_41406_1605.n3 a_41406_1605.t3 9.2885
R3216 a_41406_1605.n2 a_41406_1605.n0 4.93379
R3217 a_41406_1605.n1 a_41406_1605.t1 4.09202
R3218 a_41406_1605.n1 a_41406_1605.t2 3.95079
R3219 a_41406_1605.n3 a_41406_1605.n2 0.599711
R3220 a_41406_1605.n2 a_41406_1605.n1 0.296375
R3221 a_44488_2511.n0 a_44488_2511.t7 41.0041
R3222 a_44488_2511.n1 a_44488_2511.t4 40.8177
R3223 a_44488_2511.n1 a_44488_2511.t6 27.1302
R3224 a_44488_2511.n0 a_44488_2511.t5 26.9438
R3225 a_44488_2511.n2 a_44488_2511.n1 22.5284
R3226 a_44488_2511.n3 a_44488_2511.n2 19.5781
R3227 a_44488_2511.n3 a_44488_2511.t1 10.0473
R3228 a_44488_2511.n4 a_44488_2511.t2 6.51042
R3229 a_44488_2511.n5 a_44488_2511.n4 6.04952
R3230 a_44488_2511.n2 a_44488_2511.n0 5.7305
R3231 a_44488_2511.n4 a_44488_2511.n3 0.732092
R3232 a_44488_2511.t0 a_44488_2511.n5 0.7285
R3233 a_44488_2511.n5 a_44488_2511.t3 0.7285
R3234 a_44408_5969.n0 a_44408_5969.t4 40.6313
R3235 a_44408_5969.n0 a_44408_5969.t5 27.3166
R3236 a_44408_5969.n1 a_44408_5969.n0 24.1527
R3237 a_44408_5969.n1 a_44408_5969.t1 10.0473
R3238 a_44408_5969.t0 a_44408_5969.n3 6.51042
R3239 a_44408_5969.n3 a_44408_5969.n2 6.04952
R3240 a_44408_5969.n3 a_44408_5969.n1 0.732092
R3241 a_44408_5969.n2 a_44408_5969.t3 0.7285
R3242 a_44408_5969.n2 a_44408_5969.t2 0.7285
R3243 a_25464_1559.n0 a_25464_1559.t4 40.8177
R3244 a_25464_1559.n1 a_25464_1559.t5 40.6313
R3245 a_25464_1559.n1 a_25464_1559.t7 27.3166
R3246 a_25464_1559.n0 a_25464_1559.t6 27.1302
R3247 a_25464_1559.n2 a_25464_1559.n1 19.2576
R3248 a_25464_1559.n3 a_25464_1559.t1 10.0473
R3249 a_25464_1559.n4 a_25464_1559.t2 6.51042
R3250 a_25464_1559.n5 a_25464_1559.n4 6.04952
R3251 a_25464_1559.n2 a_25464_1559.n0 5.91752
R3252 a_25464_1559.n3 a_25464_1559.n2 4.89565
R3253 a_25464_1559.n4 a_25464_1559.n3 0.732092
R3254 a_25464_1559.t0 a_25464_1559.n5 0.7285
R3255 a_25464_1559.n5 a_25464_1559.t3 0.7285
R3256 a_29706_3501.n0 a_29706_3501.t5 34.1797
R3257 a_29706_3501.n0 a_29706_3501.t4 19.5798
R3258 a_29706_3501.n1 a_29706_3501.t1 18.7717
R3259 a_29706_3501.n1 a_29706_3501.t2 9.2885
R3260 a_29706_3501.n2 a_29706_3501.n0 4.93379
R3261 a_29706_3501.t0 a_29706_3501.n3 4.23346
R3262 a_29706_3501.n3 a_29706_3501.t3 3.85546
R3263 a_29706_3501.n2 a_29706_3501.n1 0.4055
R3264 a_29706_3501.n3 a_29706_3501.n2 0.352625
R3265 dffrs_3.Q.n3 dffrs_3.Q.t6 40.6313
R3266 dffrs_3.Q.n1 dffrs_3.Q.t5 34.1066
R3267 dffrs_3.Q.n3 dffrs_3.Q.t7 27.3166
R3268 dffrs_3.Q.n0 dffrs_3.Q.t8 19.673
R3269 dffrs_3.Q.n0 dffrs_3.Q.t4 19.4007
R3270 dffrs_3.Q.n7 dffrs_3.Q.n3 14.6967
R3271 dffrs_3.Q.n6 dffrs_3.Q.t1 10.0473
R3272 dffrs_3.Q.n7 dffrs_3.Q.n6 9.39565
R3273 dffrs_3.Q.n2 dffrs_3.Q.n1 6.70486
R3274 dffrs_3.Q.n5 dffrs_3.Q.t2 6.51042
R3275 dffrs_3.Q.n5 dffrs_3.Q.n4 6.04952
R3276 dffrs_3.Q dffrs_3.Q.n2 5.81514
R3277 dffrs_3.Q.n6 dffrs_3.Q.n5 0.732092
R3278 dffrs_3.Q.n4 dffrs_3.Q.t0 0.7285
R3279 dffrs_3.Q.n4 dffrs_3.Q.t3 0.7285
R3280 dffrs_3.Q dffrs_3.Q.n7 0.458082
R3281 dffrs_3.Q.n1 dffrs_3.Q.n0 0.252687
R3282 dffrs_3.Q.n2 2inmux_5.Bit 0.0519286
R3283 2inmux_3.OUT.n0 2inmux_3.OUT.t3 41.0041
R3284 2inmux_3.OUT.n0 2inmux_3.OUT.t2 26.9438
R3285 2inmux_3.OUT.n1 2inmux_3.OUT.t1 9.6935
R3286 dffrs_2.d 2inmux_3.OUT.n0 6.55979
R3287 2inmux_3.OUT dffrs_2.d 4.883
R3288 2inmux_3.OUT.n1 2inmux_3.OUT.t0 4.35383
R3289 2inmux_3.OUT 2inmux_3.OUT.n1 0.350857
R3290 a_12990_1604.n0 a_12990_1604.t5 34.1797
R3291 a_12990_1604.n0 a_12990_1604.t4 19.5798
R3292 a_12990_1604.n3 a_12990_1604.t3 10.3401
R3293 a_12990_1604.t0 a_12990_1604.n3 9.2885
R3294 a_12990_1604.n2 a_12990_1604.n0 4.93379
R3295 a_12990_1604.n1 a_12990_1604.t1 4.09202
R3296 a_12990_1604.n1 a_12990_1604.t2 3.95079
R3297 a_12990_1604.n3 a_12990_1604.n2 0.599711
R3298 a_12990_1604.n2 a_12990_1604.n1 0.296375
R3299 a_25464_5969.n0 a_25464_5969.t5 40.6313
R3300 a_25464_5969.n0 a_25464_5969.t4 27.3166
R3301 a_25464_5969.n1 a_25464_5969.n0 24.1527
R3302 a_25464_5969.n1 a_25464_5969.t2 10.0473
R3303 a_25464_5969.n2 a_25464_5969.t3 6.51042
R3304 a_25464_5969.n3 a_25464_5969.n2 6.04952
R3305 a_25464_5969.n2 a_25464_5969.n1 0.732092
R3306 a_25464_5969.n3 a_25464_5969.t1 0.7285
R3307 a_25464_5969.t0 a_25464_5969.n3 0.7285
R3308 a_44408_1559.n0 a_44408_1559.t5 40.8177
R3309 a_44408_1559.n1 a_44408_1559.t4 40.6313
R3310 a_44408_1559.n1 a_44408_1559.t6 27.3166
R3311 a_44408_1559.n0 a_44408_1559.t7 27.1302
R3312 a_44408_1559.n2 a_44408_1559.n1 19.2576
R3313 a_44408_1559.n3 a_44408_1559.t2 10.0473
R3314 a_44408_1559.n4 a_44408_1559.t3 6.51042
R3315 a_44408_1559.n5 a_44408_1559.n4 6.04952
R3316 a_44408_1559.n2 a_44408_1559.n0 5.91752
R3317 a_44408_1559.n3 a_44408_1559.n2 4.89565
R3318 a_44408_1559.n4 a_44408_1559.n3 0.732092
R3319 a_44408_1559.n5 a_44408_1559.t1 0.7285
R3320 a_44408_1559.t0 a_44408_1559.n5 0.7285
R3321 a_53880_1559.n0 a_53880_1559.t6 40.8177
R3322 a_53880_1559.n1 a_53880_1559.t7 40.6313
R3323 a_53880_1559.n1 a_53880_1559.t5 27.3166
R3324 a_53880_1559.n0 a_53880_1559.t4 27.1302
R3325 a_53880_1559.n2 a_53880_1559.n1 19.2576
R3326 a_53880_1559.n3 a_53880_1559.t3 10.0473
R3327 a_53880_1559.n4 a_53880_1559.t2 6.51042
R3328 a_53880_1559.n5 a_53880_1559.n4 6.04952
R3329 a_53880_1559.n2 a_53880_1559.n0 5.91752
R3330 a_53880_1559.n3 a_53880_1559.n2 4.89565
R3331 a_53880_1559.n4 a_53880_1559.n3 0.732092
R3332 a_53880_1559.t0 a_53880_1559.n5 0.7285
R3333 a_53880_1559.n5 a_53880_1559.t1 0.7285
R3334 a_53960_2511.n0 a_53960_2511.t5 41.0041
R3335 a_53960_2511.n1 a_53960_2511.t6 40.8177
R3336 a_53960_2511.n1 a_53960_2511.t4 27.1302
R3337 a_53960_2511.n0 a_53960_2511.t7 26.9438
R3338 a_53960_2511.n2 a_53960_2511.n1 22.5284
R3339 a_53960_2511.n3 a_53960_2511.n2 19.5781
R3340 a_53960_2511.n3 a_53960_2511.t2 10.0473
R3341 a_53960_2511.n4 a_53960_2511.t3 6.51042
R3342 a_53960_2511.n5 a_53960_2511.n4 6.04952
R3343 a_53960_2511.n2 a_53960_2511.n0 5.7305
R3344 a_53960_2511.n4 a_53960_2511.n3 0.732092
R3345 a_53960_2511.n5 a_53960_2511.t1 0.7285
R3346 a_53960_2511.t0 a_53960_2511.n5 0.7285
R3347 a_53880_3764.n3 a_53880_3764.t8 41.0041
R3348 a_53880_3764.n2 a_53880_3764.t7 40.8177
R3349 a_53880_3764.n4 a_53880_3764.t9 40.6313
R3350 a_53880_3764.n4 a_53880_3764.t6 27.3166
R3351 a_53880_3764.n2 a_53880_3764.t4 27.1302
R3352 a_53880_3764.n3 a_53880_3764.t5 26.9438
R3353 a_53880_3764.n5 a_53880_3764.n3 15.6312
R3354 a_53880_3764.n5 a_53880_3764.n4 15.046
R3355 a_53880_3764.t0 a_53880_3764.n7 10.0473
R3356 a_53880_3764.n1 a_53880_3764.t1 6.51042
R3357 a_53880_3764.n1 a_53880_3764.n0 6.04952
R3358 a_53880_3764.n6 a_53880_3764.n2 5.64619
R3359 a_53880_3764.n7 a_53880_3764.n6 5.17851
R3360 a_53880_3764.n6 a_53880_3764.n5 4.5005
R3361 a_53880_3764.n7 a_53880_3764.n1 0.732092
R3362 a_53880_3764.n0 a_53880_3764.t2 0.7285
R3363 a_53880_3764.n0 a_53880_3764.t3 0.7285
R3364 2inmux_2.OUT.n0 2inmux_2.OUT.t2 41.0041
R3365 2inmux_2.OUT.n0 2inmux_2.OUT.t3 26.9438
R3366 2inmux_2.OUT.n1 2inmux_2.OUT.t1 9.6935
R3367 dffrs_1.d 2inmux_2.OUT.n0 6.55979
R3368 2inmux_2.OUT dffrs_1.d 4.883
R3369 2inmux_2.OUT.n1 2inmux_2.OUT.t0 4.35383
R3370 2inmux_2.OUT 2inmux_2.OUT.n1 0.350857
R3371 a_16072_2510.n2 a_16072_2510.t4 41.0041
R3372 a_16072_2510.n3 a_16072_2510.t5 40.8177
R3373 a_16072_2510.n3 a_16072_2510.t7 27.1302
R3374 a_16072_2510.n2 a_16072_2510.t6 26.9438
R3375 a_16072_2510.n4 a_16072_2510.n3 22.5284
R3376 a_16072_2510.n5 a_16072_2510.n4 19.5781
R3377 a_16072_2510.t0 a_16072_2510.n5 10.0473
R3378 a_16072_2510.n1 a_16072_2510.t1 6.51042
R3379 a_16072_2510.n1 a_16072_2510.n0 6.04952
R3380 a_16072_2510.n4 a_16072_2510.n2 5.7305
R3381 a_16072_2510.n5 a_16072_2510.n1 0.732092
R3382 a_16072_2510.n0 a_16072_2510.t2 0.7285
R3383 a_16072_2510.n0 a_16072_2510.t3 0.7285
R3384 a_34936_5969.n0 a_34936_5969.t5 40.6313
R3385 a_34936_5969.n0 a_34936_5969.t4 27.3166
R3386 a_34936_5969.n1 a_34936_5969.n0 24.1527
R3387 a_34936_5969.n1 a_34936_5969.t2 10.0473
R3388 a_34936_5969.n2 a_34936_5969.t1 6.51042
R3389 a_34936_5969.n3 a_34936_5969.n2 6.04952
R3390 a_34936_5969.n2 a_34936_5969.n1 0.732092
R3391 a_34936_5969.t0 a_34936_5969.n3 0.7285
R3392 a_34936_5969.n3 a_34936_5969.t3 0.7285
R3393 a_15992_1558.n2 a_15992_1558.t4 40.8177
R3394 a_15992_1558.n3 a_15992_1558.t5 40.6313
R3395 a_15992_1558.n3 a_15992_1558.t7 27.3166
R3396 a_15992_1558.n2 a_15992_1558.t6 27.1302
R3397 a_15992_1558.n4 a_15992_1558.n3 19.2576
R3398 a_15992_1558.t0 a_15992_1558.n5 10.0473
R3399 a_15992_1558.n1 a_15992_1558.t1 6.51042
R3400 a_15992_1558.n1 a_15992_1558.n0 6.04952
R3401 a_15992_1558.n4 a_15992_1558.n2 5.91752
R3402 a_15992_1558.n5 a_15992_1558.n4 4.89565
R3403 a_15992_1558.n5 a_15992_1558.n1 0.732092
R3404 a_15992_1558.n0 a_15992_1558.t2 0.7285
R3405 a_15992_1558.n0 a_15992_1558.t3 0.7285
R3406 a_53880_5969.n0 a_53880_5969.t4 40.6313
R3407 a_53880_5969.n0 a_53880_5969.t5 27.3166
R3408 a_53880_5969.n1 a_53880_5969.n0 24.1527
R3409 a_53880_5969.n1 a_53880_5969.t2 10.0473
R3410 a_53880_5969.n2 a_53880_5969.t3 6.51042
R3411 a_53880_5969.n3 a_53880_5969.n2 6.04952
R3412 a_53880_5969.n2 a_53880_5969.n1 0.732092
R3413 a_53880_5969.n3 a_53880_5969.t1 0.7285
R3414 a_53880_5969.t0 a_53880_5969.n3 0.7285
R3415 a_31934_1605.n0 a_31934_1605.t5 34.1797
R3416 a_31934_1605.n0 a_31934_1605.t4 19.5798
R3417 a_31934_1605.t0 a_31934_1605.n3 10.3401
R3418 a_31934_1605.n3 a_31934_1605.t3 9.2885
R3419 a_31934_1605.n2 a_31934_1605.n0 4.93379
R3420 a_31934_1605.n1 a_31934_1605.t1 4.09202
R3421 a_31934_1605.n1 a_31934_1605.t2 3.95079
R3422 a_31934_1605.n3 a_31934_1605.n2 0.599711
R3423 a_31934_1605.n2 a_31934_1605.n1 0.296375
R3424 2inmux_4.OUT.n0 2inmux_4.OUT.t2 41.0041
R3425 2inmux_4.OUT.n0 2inmux_4.OUT.t3 26.9438
R3426 2inmux_4.OUT.n1 2inmux_4.OUT.t1 9.6935
R3427 dffrs_3.d 2inmux_4.OUT.n0 6.55979
R3428 2inmux_4.OUT dffrs_3.d 4.883
R3429 2inmux_4.OUT.n1 2inmux_4.OUT.t0 4.35383
R3430 2inmux_4.OUT 2inmux_4.OUT.n1 0.350857
R3431 a_25544_2511.n0 a_25544_2511.t6 41.0041
R3432 a_25544_2511.n1 a_25544_2511.t7 40.8177
R3433 a_25544_2511.n1 a_25544_2511.t5 27.1302
R3434 a_25544_2511.n0 a_25544_2511.t4 26.9438
R3435 a_25544_2511.n2 a_25544_2511.n1 22.5284
R3436 a_25544_2511.n3 a_25544_2511.n2 19.5781
R3437 a_25544_2511.n3 a_25544_2511.t2 10.0473
R3438 a_25544_2511.n4 a_25544_2511.t1 6.51042
R3439 a_25544_2511.n5 a_25544_2511.n4 6.04952
R3440 a_25544_2511.n2 a_25544_2511.n0 5.7305
R3441 a_25544_2511.n4 a_25544_2511.n3 0.732092
R3442 a_25544_2511.n5 a_25544_2511.t3 0.7285
R3443 a_25544_2511.t0 a_25544_2511.n5 0.7285
R3444 B5.n1 B5.t0 34.2529
R3445 B5.n0 B5.t1 19.673
R3446 B5.n0 B5.t2 19.4007
R3447 B5.n2 B5.n1 8.05164
R3448 B5.n2 B5 1.87121
R3449 B5.n1 B5.n0 0.106438
R3450 2inmux_2.In B5.n2 0.0455
R3451 a_10762_1160.n0 a_10762_1160.t5 34.1797
R3452 a_10762_1160.n0 a_10762_1160.t4 19.5798
R3453 a_10762_1160.n1 a_10762_1160.t2 18.7717
R3454 a_10762_1160.n1 a_10762_1160.t1 9.2885
R3455 a_10762_1160.n2 a_10762_1160.n0 4.93379
R3456 a_10762_1160.n3 a_10762_1160.t3 4.23346
R3457 a_10762_1160.t0 a_10762_1160.n3 3.85546
R3458 a_10762_1160.n2 a_10762_1160.n1 0.4055
R3459 a_10762_1160.n3 a_10762_1160.n2 0.352625
R3460 a_6520_5968.n0 a_6520_5968.t4 40.6313
R3461 a_6520_5968.n0 a_6520_5968.t5 27.3166
R3462 a_6520_5968.n1 a_6520_5968.n0 24.1527
R3463 a_6520_5968.n1 a_6520_5968.t2 10.0473
R3464 a_6520_5968.n2 a_6520_5968.t1 6.51042
R3465 a_6520_5968.n3 a_6520_5968.n2 6.04952
R3466 a_6520_5968.n2 a_6520_5968.n1 0.732092
R3467 a_6520_5968.t0 a_6520_5968.n3 0.7285
R3468 a_6520_5968.n3 a_6520_5968.t3 0.7285
R3469 serial_out.n0 serial_out.t4 40.6313
R3470 serial_out.n0 serial_out.t5 27.3166
R3471 serial_out.n4 serial_out.n0 14.6967
R3472 serial_out.n3 serial_out.t3 10.0473
R3473 serial_out.n4 serial_out.n3 9.39565
R3474 serial_out.n2 serial_out.t2 6.51042
R3475 serial_out.n2 serial_out.n1 6.04952
R3476 dffrs_5.Q serial_out 5.90514
R3477 serial_out.n3 serial_out.n2 0.732092
R3478 serial_out.n1 serial_out.t1 0.7285
R3479 serial_out.n1 serial_out.t0 0.7285
R3480 dffrs_5.Q serial_out.n4 0.458082
R3481 B2.n1 B2.t2 34.2529
R3482 B2.n0 B2.t0 19.673
R3483 B2.n0 B2.t1 19.4007
R3484 B2.n2 B2.n1 8.05164
R3485 B2.n2 B2 1.87121
R3486 B2.n1 B2.n0 0.106438
R3487 2inmux_5.In B2.n2 0.0455
R3488 a_39178_1161.n0 a_39178_1161.t5 34.1797
R3489 a_39178_1161.n0 a_39178_1161.t4 19.5798
R3490 a_39178_1161.n1 a_39178_1161.t2 18.7717
R3491 a_39178_1161.n1 a_39178_1161.t1 9.2885
R3492 a_39178_1161.n2 a_39178_1161.n0 4.93379
R3493 a_39178_1161.t0 a_39178_1161.n3 4.23346
R3494 a_39178_1161.n3 a_39178_1161.t3 3.85546
R3495 a_39178_1161.n2 a_39178_1161.n1 0.4055
R3496 a_39178_1161.n3 a_39178_1161.n2 0.352625
R3497 2inmux_5.OUT.n0 2inmux_5.OUT.t3 41.0041
R3498 2inmux_5.OUT.n0 2inmux_5.OUT.t2 26.9438
R3499 2inmux_5.OUT.n1 2inmux_5.OUT.t1 9.6935
R3500 dffrs_4.d 2inmux_5.OUT.n0 6.55979
R3501 2inmux_5.OUT dffrs_4.d 4.883
R3502 2inmux_5.OUT.n1 2inmux_5.OUT.t0 4.35383
R3503 2inmux_5.OUT 2inmux_5.OUT.n1 0.350857
R3504 B4.n1 B4.t1 34.2529
R3505 B4.n0 B4.t0 19.673
R3506 B4.n0 B4.t2 19.4007
R3507 B4.n2 B4.n1 8.05164
R3508 B4.n2 B4 1.87282
R3509 B4.n1 B4.n0 0.106438
R3510 2inmux_3.In B4.n2 0.0455
R3511 B1.n1 B1.t1 34.2529
R3512 B1.n0 B1.t0 19.673
R3513 B1.n0 B1.t2 19.4007
R3514 B1.n2 B1.n1 8.05164
R3515 B1.n2 B1 1.87121
R3516 B1.n1 B1.n0 0.106438
R3517 2inmux_1.In B1.n2 0.0455
R3518 B3.n1 B3.t1 34.2529
R3519 B3.n0 B3.t0 19.673
R3520 B3.n0 B3.t2 19.4007
R3521 B3.n2 B3.n1 8.05164
R3522 B3.n2 B3 1.87121
R3523 B3.n1 B3.n0 0.106438
R3524 2inmux_4.In B3.n2 0.0455
R3525 avdd.t266 avdd.n390 250.9
R3526 avdd.n391 avdd.t92 250.9
R3527 avdd.t24 avdd.n401 250.9
R3528 avdd.n402 avdd.t298 250.9
R3529 avdd.t198 avdd.n396 250.9
R3530 avdd.n397 avdd.t89 250.9
R3531 avdd.t240 avdd.n413 250.9
R3532 avdd.n414 avdd.t264 250.9
R3533 avdd.t140 avdd.n407 250.9
R3534 avdd.n408 avdd.t18 250.9
R3535 avdd.t248 avdd.n425 250.9
R3536 avdd.n426 avdd.t286 250.9
R3537 avdd.t228 avdd.n98 250.9
R3538 avdd.n99 avdd.t143 250.9
R3539 avdd.t338 avdd.n109 250.9
R3540 avdd.n110 avdd.t292 250.9
R3541 avdd.t334 avdd.n104 250.9
R3542 avdd.n105 avdd.t137 250.9
R3543 avdd.t250 avdd.n121 250.9
R3544 avdd.n122 avdd.t230 250.9
R3545 avdd.t95 avdd.n115 250.9
R3546 avdd.n116 avdd.t176 250.9
R3547 avdd.t308 avdd.n132 250.9
R3548 avdd.n133 avdd.t40 250.9
R3549 avdd.t196 avdd.n171 250.9
R3550 avdd.n172 avdd.t119 250.9
R3551 avdd.t344 avdd.n182 250.9
R3552 avdd.n183 avdd.t318 250.9
R3553 avdd.t352 avdd.n177 250.9
R3554 avdd.n178 avdd.t80 250.9
R3555 avdd.t256 avdd.n194 250.9
R3556 avdd.n195 avdd.t192 250.9
R3557 avdd.t116 avdd.n188 250.9
R3558 avdd.n189 avdd.t304 250.9
R3559 avdd.t252 avdd.n205 250.9
R3560 avdd.n206 avdd.t280 250.9
R3561 avdd.t64 avdd.n244 250.9
R3562 avdd.n245 avdd.t83 250.9
R3563 avdd.t350 avdd.n255 250.9
R3564 avdd.n256 avdd.t246 250.9
R3565 avdd.t60 avdd.n250 250.9
R3566 avdd.n251 avdd.t149 250.9
R3567 avdd.t300 avdd.n267 250.9
R3568 avdd.n268 avdd.t62 250.9
R3569 avdd.t77 avdd.n261 250.9
R3570 avdd.n262 avdd.t278 250.9
R3571 avdd.t296 avdd.n278 250.9
R3572 avdd.n279 avdd.t216 250.9
R3573 avdd.t322 avdd.n317 250.9
R3574 avdd.n318 avdd.t104 250.9
R3575 avdd.t26 avdd.n328 250.9
R3576 avdd.n329 avdd.t244 250.9
R3577 avdd.t14 avdd.n323 250.9
R3578 avdd.n324 avdd.t107 250.9
R3579 avdd.t206 avdd.n340 250.9
R3580 avdd.n341 avdd.t324 250.9
R3581 avdd.t152 avdd.n334 250.9
R3582 avdd.n335 avdd.t310 250.9
R3583 avdd.t178 avdd.n351 250.9
R3584 avdd.n352 avdd.t364 250.9
R3585 avdd.t332 avdd.n4 250.9
R3586 avdd.n5 avdd.t131 250.9
R3587 avdd.t340 avdd.n528 250.9
R3588 avdd.n529 avdd.t186 250.9
R3589 avdd.t12 avdd.n9 250.9
R3590 avdd.n10 avdd.t125 250.9
R3591 avdd.t4 avdd.n516 250.9
R3592 avdd.n517 avdd.t328 250.9
R3593 avdd.t158 avdd.n522 250.9
R3594 avdd.n523 avdd.t368 250.9
R3595 avdd.t370 avdd.n465 250.9
R3596 avdd.n466 avdd.t50 250.9
R3597 avdd.n495 avdd.t188 236.083
R3598 avdd.t174 avdd.n491 236.083
R3599 avdd.t210 avdd.n499 236.083
R3600 avdd.n505 avdd.t74 236.083
R3601 avdd.n453 avdd.t306 236.083
R3602 avdd.t44 avdd.n450 236.083
R3603 avdd.t222 avdd.n433 236.083
R3604 avdd.n439 avdd.t218 236.083
R3605 avdd.n379 avdd.t260 236.083
R3606 avdd.t190 avdd.n376 236.083
R3607 avdd.t236 avdd.n359 236.083
R3608 avdd.n365 avdd.t220 236.083
R3609 avdd.n306 avdd.t200 236.083
R3610 avdd.t268 avdd.n303 236.083
R3611 avdd.t56 avdd.n286 236.083
R3612 avdd.n292 avdd.t46 236.083
R3613 avdd.n233 avdd.t354 236.083
R3614 avdd.t168 avdd.n230 236.083
R3615 avdd.t254 avdd.n213 236.083
R3616 avdd.n219 avdd.t232 236.083
R3617 avdd.n160 avdd.t336 236.083
R3618 avdd.t212 avdd.n157 236.083
R3619 avdd.t258 avdd.n140 236.083
R3620 avdd.n146 avdd.t2 236.083
R3621 avdd.n92 avdd.t214 236.083
R3622 avdd.n86 avdd.t182 236.083
R3623 avdd.n76 avdd.t238 236.083
R3624 avdd.n70 avdd.t30 236.083
R3625 avdd.n60 avdd.t294 236.083
R3626 avdd.n54 avdd.t202 236.083
R3627 avdd.n44 avdd.t166 236.083
R3628 avdd.n38 avdd.t274 236.083
R3629 avdd.n28 avdd.t366 236.083
R3630 avdd.n22 avdd.t32 236.083
R3631 avdd.t234 avdd.n470 236.083
R3632 avdd.n481 avdd.t374 236.083
R3633 avdd.t188 avdd.n494 235.294
R3634 avdd.n494 avdd.t174 235.294
R3635 avdd.n504 avdd.t210 235.294
R3636 avdd.t74 avdd.n504 235.294
R3637 avdd.t306 avdd.n452 235.294
R3638 avdd.n452 avdd.t44 235.294
R3639 avdd.n438 avdd.t222 235.294
R3640 avdd.t218 avdd.n438 235.294
R3641 avdd.t260 avdd.n378 235.294
R3642 avdd.n378 avdd.t190 235.294
R3643 avdd.n364 avdd.t236 235.294
R3644 avdd.t220 avdd.n364 235.294
R3645 avdd.t200 avdd.n305 235.294
R3646 avdd.n305 avdd.t268 235.294
R3647 avdd.n291 avdd.t56 235.294
R3648 avdd.t46 avdd.n291 235.294
R3649 avdd.t354 avdd.n232 235.294
R3650 avdd.n232 avdd.t168 235.294
R3651 avdd.n218 avdd.t254 235.294
R3652 avdd.t232 avdd.n218 235.294
R3653 avdd.t336 avdd.n159 235.294
R3654 avdd.n159 avdd.t212 235.294
R3655 avdd.n145 avdd.t258 235.294
R3656 avdd.t2 avdd.n145 235.294
R3657 avdd.t214 avdd.n91 235.294
R3658 avdd.n91 avdd.t316 235.294
R3659 avdd.t317 avdd.n89 235.294
R3660 avdd.n89 avdd.t180 235.294
R3661 avdd.t238 avdd.n75 235.294
R3662 avdd.n75 avdd.t59 235.294
R3663 avdd.t58 avdd.n73 235.294
R3664 avdd.n73 avdd.t28 235.294
R3665 avdd.t294 avdd.n59 235.294
R3666 avdd.n59 avdd.t315 235.294
R3667 avdd.t314 avdd.n57 235.294
R3668 avdd.n57 avdd.t204 235.294
R3669 avdd.t166 avdd.n43 235.294
R3670 avdd.n43 avdd.t373 235.294
R3671 avdd.t372 avdd.n41 235.294
R3672 avdd.n41 avdd.t272 235.294
R3673 avdd.t366 avdd.n27 235.294
R3674 avdd.n27 avdd.t1 235.294
R3675 avdd.t0 avdd.n25 235.294
R3676 avdd.n25 avdd.t34 235.294
R3677 avdd.n478 avdd.t234 235.294
R3678 avdd.t10 avdd.n478 235.294
R3679 avdd.n480 avdd.t11 235.294
R3680 avdd.t376 avdd.n480 235.294
R3681 avdd.t242 avdd.t266 200
R3682 avdd.t92 avdd.t242 200
R3683 avdd.t155 avdd.t24 200
R3684 avdd.t298 avdd.t155 200
R3685 avdd.t262 avdd.t198 200
R3686 avdd.t89 avdd.t262 200
R3687 avdd.t348 avdd.t240 200
R3688 avdd.t264 avdd.t348 200
R3689 avdd.t284 avdd.t140 200
R3690 avdd.t18 avdd.t284 200
R3691 avdd.t86 avdd.t248 200
R3692 avdd.t286 avdd.t86 200
R3693 avdd.t290 avdd.t228 200
R3694 avdd.t143 avdd.t290 200
R3695 avdd.t110 avdd.t338 200
R3696 avdd.t292 avdd.t110 200
R3697 avdd.t226 avdd.t334 200
R3698 avdd.t137 avdd.t226 200
R3699 avdd.t8 avdd.t250 200
R3700 avdd.t230 avdd.t8 200
R3701 avdd.t38 avdd.t95 200
R3702 avdd.t176 avdd.t38 200
R3703 avdd.t134 avdd.t308 200
R3704 avdd.t40 avdd.t134 200
R3705 avdd.t316 avdd.t317 200
R3706 avdd.t182 avdd.t180 200
R3707 avdd.t288 avdd.t196 200
R3708 avdd.t119 avdd.t288 200
R3709 avdd.t164 avdd.t344 200
R3710 avdd.t318 avdd.t164 200
R3711 avdd.t194 avdd.t352 200
R3712 avdd.t80 avdd.t194 200
R3713 avdd.t346 avdd.t256 200
R3714 avdd.t192 avdd.t346 200
R3715 avdd.t282 avdd.t116 200
R3716 avdd.t304 avdd.t282 200
R3717 avdd.t98 avdd.t252 200
R3718 avdd.t280 avdd.t98 200
R3719 avdd.t59 avdd.t58 200
R3720 avdd.t30 avdd.t28 200
R3721 avdd.t302 avdd.t64 200
R3722 avdd.t83 avdd.t302 200
R3723 avdd.t113 avdd.t350 200
R3724 avdd.t246 avdd.t113 200
R3725 avdd.t360 avdd.t60 200
R3726 avdd.t149 avdd.t360 200
R3727 avdd.t6 avdd.t300 200
R3728 avdd.t62 avdd.t6 200
R3729 avdd.t224 avdd.t77 200
R3730 avdd.t278 avdd.t224 200
R3731 avdd.t146 avdd.t296 200
R3732 avdd.t216 avdd.t146 200
R3733 avdd.t315 avdd.t314 200
R3734 avdd.t202 avdd.t204 200
R3735 avdd.t208 avdd.t322 200
R3736 avdd.t104 avdd.t208 200
R3737 avdd.t101 avdd.t26 200
R3738 avdd.t244 avdd.t101 200
R3739 avdd.t320 avdd.t14 200
R3740 avdd.t107 avdd.t320 200
R3741 avdd.t22 avdd.t206 200
R3742 avdd.t324 avdd.t22 200
R3743 avdd.t362 avdd.t152 200
R3744 avdd.t310 avdd.t362 200
R3745 avdd.t122 avdd.t178 200
R3746 avdd.t364 avdd.t122 200
R3747 avdd.t373 avdd.t372 200
R3748 avdd.t274 avdd.t272 200
R3749 avdd.t1 avdd.t0 200
R3750 avdd.t32 avdd.t34 200
R3751 avdd.t20 avdd.t332 200
R3752 avdd.t131 avdd.t20 200
R3753 avdd.t128 avdd.t340 200
R3754 avdd.t186 avdd.t128 200
R3755 avdd.t330 avdd.t12 200
R3756 avdd.t125 avdd.t330 200
R3757 avdd.t342 avdd.t4 200
R3758 avdd.t328 avdd.t342 200
R3759 avdd.t52 avdd.t158 200
R3760 avdd.t368 avdd.t52 200
R3761 avdd.t161 avdd.t370 200
R3762 avdd.t50 avdd.t161 200
R3763 avdd.t11 avdd.t10 200
R3764 avdd.t374 avdd.t376 200
R3765 avdd.n486 avdd.t54 131.589
R3766 avdd.n507 avdd.t48 131.589
R3767 avdd.n14 avdd.t356 131.589
R3768 avdd.n441 avdd.t326 131.589
R3769 avdd.n30 avdd.t42 131.589
R3770 avdd.n367 avdd.t66 131.589
R3771 avdd.n46 avdd.t312 131.589
R3772 avdd.n294 avdd.t16 131.589
R3773 avdd.n62 avdd.t276 131.589
R3774 avdd.n221 avdd.t36 131.589
R3775 avdd.n78 avdd.t184 131.589
R3776 avdd.n148 avdd.t358 131.589
R3777 avdd.n164 avdd.t70 118.543
R3778 avdd.n237 avdd.t72 118.543
R3779 avdd.n310 avdd.t68 118.543
R3780 avdd.n383 avdd.t170 118.543
R3781 avdd.n457 avdd.t270 118.543
R3782 avdd.n487 avdd.t172 118.543
R3783 avdd.n86 avdd.n85 96.0755
R3784 avdd.n87 avdd.n86 96.0755
R3785 avdd.n70 avdd.n69 96.0755
R3786 avdd.n71 avdd.n70 96.0755
R3787 avdd.n54 avdd.n53 96.0755
R3788 avdd.n55 avdd.n54 96.0755
R3789 avdd.n38 avdd.n37 96.0755
R3790 avdd.n39 avdd.n38 96.0755
R3791 avdd.n22 avdd.n21 96.0755
R3792 avdd.n23 avdd.n22 96.0755
R3793 avdd.n481 avdd.n473 96.0755
R3794 avdd.n481 avdd.n474 96.0755
R3795 avdd.n501 avdd.n499 78.2255
R3796 avdd.n505 avdd.n501 78.2255
R3797 avdd.n505 avdd.n502 78.2255
R3798 avdd.n502 avdd.n499 78.2255
R3799 avdd.n435 avdd.n433 78.2255
R3800 avdd.n439 avdd.n435 78.2255
R3801 avdd.n439 avdd.n436 78.2255
R3802 avdd.n436 avdd.n433 78.2255
R3803 avdd.n361 avdd.n359 78.2255
R3804 avdd.n365 avdd.n361 78.2255
R3805 avdd.n365 avdd.n362 78.2255
R3806 avdd.n362 avdd.n359 78.2255
R3807 avdd.n288 avdd.n286 78.2255
R3808 avdd.n292 avdd.n288 78.2255
R3809 avdd.n292 avdd.n289 78.2255
R3810 avdd.n289 avdd.n286 78.2255
R3811 avdd.n215 avdd.n213 78.2255
R3812 avdd.n219 avdd.n215 78.2255
R3813 avdd.n219 avdd.n216 78.2255
R3814 avdd.n216 avdd.n213 78.2255
R3815 avdd.n142 avdd.n140 78.2255
R3816 avdd.n146 avdd.n142 78.2255
R3817 avdd.n146 avdd.n143 78.2255
R3818 avdd.n143 avdd.n140 78.2255
R3819 avdd.n92 avdd.n83 78.2255
R3820 avdd.n92 avdd.n84 78.2255
R3821 avdd.n160 avdd.n155 78.2255
R3822 avdd.n160 avdd.n156 78.2255
R3823 avdd.n157 avdd.n155 78.2255
R3824 avdd.n157 avdd.n156 78.2255
R3825 avdd.n76 avdd.n67 78.2255
R3826 avdd.n76 avdd.n68 78.2255
R3827 avdd.n233 avdd.n228 78.2255
R3828 avdd.n233 avdd.n229 78.2255
R3829 avdd.n230 avdd.n228 78.2255
R3830 avdd.n230 avdd.n229 78.2255
R3831 avdd.n60 avdd.n51 78.2255
R3832 avdd.n60 avdd.n52 78.2255
R3833 avdd.n306 avdd.n301 78.2255
R3834 avdd.n306 avdd.n302 78.2255
R3835 avdd.n303 avdd.n301 78.2255
R3836 avdd.n303 avdd.n302 78.2255
R3837 avdd.n44 avdd.n35 78.2255
R3838 avdd.n44 avdd.n36 78.2255
R3839 avdd.n379 avdd.n374 78.2255
R3840 avdd.n379 avdd.n375 78.2255
R3841 avdd.n376 avdd.n374 78.2255
R3842 avdd.n376 avdd.n375 78.2255
R3843 avdd.n28 avdd.n19 78.2255
R3844 avdd.n28 avdd.n20 78.2255
R3845 avdd.n453 avdd.n448 78.2255
R3846 avdd.n453 avdd.n449 78.2255
R3847 avdd.n450 avdd.n448 78.2255
R3848 avdd.n450 avdd.n449 78.2255
R3849 avdd.n475 avdd.n470 78.2255
R3850 avdd.n476 avdd.n470 78.2255
R3851 avdd.n495 avdd.n484 78.2255
R3852 avdd.n495 avdd.n485 78.2255
R3853 avdd.n491 avdd.n484 78.2255
R3854 avdd.n491 avdd.n485 78.2255
R3855 avdd.n391 avdd.n390 68.0765
R3856 avdd.n402 avdd.n401 68.0765
R3857 avdd.n397 avdd.n396 68.0765
R3858 avdd.n414 avdd.n413 68.0765
R3859 avdd.n408 avdd.n407 68.0765
R3860 avdd.n426 avdd.n425 68.0765
R3861 avdd.n99 avdd.n98 68.0765
R3862 avdd.n110 avdd.n109 68.0765
R3863 avdd.n105 avdd.n104 68.0765
R3864 avdd.n122 avdd.n121 68.0765
R3865 avdd.n116 avdd.n115 68.0765
R3866 avdd.n133 avdd.n132 68.0765
R3867 avdd.n172 avdd.n171 68.0765
R3868 avdd.n183 avdd.n182 68.0765
R3869 avdd.n178 avdd.n177 68.0765
R3870 avdd.n195 avdd.n194 68.0765
R3871 avdd.n189 avdd.n188 68.0765
R3872 avdd.n206 avdd.n205 68.0765
R3873 avdd.n245 avdd.n244 68.0765
R3874 avdd.n256 avdd.n255 68.0765
R3875 avdd.n251 avdd.n250 68.0765
R3876 avdd.n268 avdd.n267 68.0765
R3877 avdd.n262 avdd.n261 68.0765
R3878 avdd.n279 avdd.n278 68.0765
R3879 avdd.n318 avdd.n317 68.0765
R3880 avdd.n329 avdd.n328 68.0765
R3881 avdd.n324 avdd.n323 68.0765
R3882 avdd.n341 avdd.n340 68.0765
R3883 avdd.n335 avdd.n334 68.0765
R3884 avdd.n352 avdd.n351 68.0765
R3885 avdd.n5 avdd.n4 68.0765
R3886 avdd.n529 avdd.n528 68.0765
R3887 avdd.n10 avdd.n9 68.0765
R3888 avdd.n517 avdd.n516 68.0765
R3889 avdd.n523 avdd.n522 68.0765
R3890 avdd.n466 avdd.n465 68.0765
R3891 avdd.n85 avdd.n83 59.8505
R3892 avdd.n87 avdd.n84 59.8505
R3893 avdd.n69 avdd.n67 59.8505
R3894 avdd.n71 avdd.n68 59.8505
R3895 avdd.n53 avdd.n51 59.8505
R3896 avdd.n55 avdd.n52 59.8505
R3897 avdd.n37 avdd.n35 59.8505
R3898 avdd.n39 avdd.n36 59.8505
R3899 avdd.n21 avdd.n19 59.8505
R3900 avdd.n23 avdd.n20 59.8505
R3901 avdd.n475 avdd.n473 59.8505
R3902 avdd.n476 avdd.n474 59.8505
R3903 avdd.n419 avdd.t139 41.0041
R3904 avdd.n126 avdd.t94 41.0041
R3905 avdd.n199 avdd.t115 41.0041
R3906 avdd.n272 avdd.t76 41.0041
R3907 avdd.n345 avdd.t151 41.0041
R3908 avdd.n459 avdd.t157 41.0041
R3909 avdd.n421 avdd.t85 40.8177
R3910 avdd.n420 avdd.t154 40.8177
R3911 avdd.n128 avdd.t133 40.8177
R3912 avdd.n127 avdd.t109 40.8177
R3913 avdd.n201 avdd.t97 40.8177
R3914 avdd.n200 avdd.t163 40.8177
R3915 avdd.n274 avdd.t145 40.8177
R3916 avdd.n273 avdd.t112 40.8177
R3917 avdd.n347 avdd.t121 40.8177
R3918 avdd.n346 avdd.t100 40.8177
R3919 avdd.n461 avdd.t160 40.8177
R3920 avdd.n460 avdd.t127 40.8177
R3921 avdd.n386 avdd.t91 40.6313
R3922 avdd.n385 avdd.t88 40.6313
R3923 avdd.n94 avdd.t142 40.6313
R3924 avdd.n93 avdd.t136 40.6313
R3925 avdd.n167 avdd.t118 40.6313
R3926 avdd.n166 avdd.t79 40.6313
R3927 avdd.n240 avdd.t82 40.6313
R3928 avdd.n239 avdd.t148 40.6313
R3929 avdd.n313 avdd.t103 40.6313
R3930 avdd.n312 avdd.t106 40.6313
R3931 avdd.n1 avdd.t130 40.6313
R3932 avdd.n0 avdd.t124 40.6313
R3933 avdd.n503 avdd.n501 36.2255
R3934 avdd.n503 avdd.n502 36.2255
R3935 avdd.n437 avdd.n435 36.2255
R3936 avdd.n437 avdd.n436 36.2255
R3937 avdd.n363 avdd.n361 36.2255
R3938 avdd.n363 avdd.n362 36.2255
R3939 avdd.n290 avdd.n288 36.2255
R3940 avdd.n290 avdd.n289 36.2255
R3941 avdd.n217 avdd.n215 36.2255
R3942 avdd.n217 avdd.n216 36.2255
R3943 avdd.n144 avdd.n142 36.2255
R3944 avdd.n144 avdd.n143 36.2255
R3945 avdd.n88 avdd.n85 36.2255
R3946 avdd.n88 avdd.n87 36.2255
R3947 avdd.n90 avdd.n83 36.2255
R3948 avdd.n90 avdd.n84 36.2255
R3949 avdd.n158 avdd.n155 36.2255
R3950 avdd.n158 avdd.n156 36.2255
R3951 avdd.n72 avdd.n69 36.2255
R3952 avdd.n72 avdd.n71 36.2255
R3953 avdd.n74 avdd.n67 36.2255
R3954 avdd.n74 avdd.n68 36.2255
R3955 avdd.n231 avdd.n228 36.2255
R3956 avdd.n231 avdd.n229 36.2255
R3957 avdd.n56 avdd.n53 36.2255
R3958 avdd.n56 avdd.n55 36.2255
R3959 avdd.n58 avdd.n51 36.2255
R3960 avdd.n58 avdd.n52 36.2255
R3961 avdd.n304 avdd.n301 36.2255
R3962 avdd.n304 avdd.n302 36.2255
R3963 avdd.n40 avdd.n37 36.2255
R3964 avdd.n40 avdd.n39 36.2255
R3965 avdd.n42 avdd.n35 36.2255
R3966 avdd.n42 avdd.n36 36.2255
R3967 avdd.n377 avdd.n374 36.2255
R3968 avdd.n377 avdd.n375 36.2255
R3969 avdd.n24 avdd.n21 36.2255
R3970 avdd.n24 avdd.n23 36.2255
R3971 avdd.n26 avdd.n19 36.2255
R3972 avdd.n26 avdd.n20 36.2255
R3973 avdd.n451 avdd.n448 36.2255
R3974 avdd.n451 avdd.n449 36.2255
R3975 avdd.n479 avdd.n473 36.2255
R3976 avdd.n479 avdd.n474 36.2255
R3977 avdd.n477 avdd.n475 36.2255
R3978 avdd.n477 avdd.n476 36.2255
R3979 avdd.n493 avdd.n484 36.2255
R3980 avdd.n493 avdd.n485 36.2255
R3981 avdd.n386 avdd.t388 27.3166
R3982 avdd.n385 avdd.t390 27.3166
R3983 avdd.n94 avdd.t399 27.3166
R3984 avdd.n93 avdd.t403 27.3166
R3985 avdd.n167 avdd.t378 27.3166
R3986 avdd.n166 avdd.t386 27.3166
R3987 avdd.n240 avdd.t391 27.3166
R3988 avdd.n239 avdd.t400 27.3166
R3989 avdd.n313 avdd.t382 27.3166
R3990 avdd.n312 avdd.t383 27.3166
R3991 avdd.n1 avdd.t404 27.3166
R3992 avdd.n0 avdd.t407 27.3166
R3993 avdd.n421 avdd.t389 27.1302
R3994 avdd.n420 avdd.t396 27.1302
R3995 avdd.n128 avdd.t402 27.1302
R3996 avdd.n127 avdd.t381 27.1302
R3997 avdd.n201 avdd.t384 27.1302
R3998 avdd.n200 avdd.t394 27.1302
R3999 avdd.n274 avdd.t398 27.1302
R4000 avdd.n273 avdd.t380 27.1302
R4001 avdd.n347 avdd.t405 27.1302
R4002 avdd.n346 avdd.t385 27.1302
R4003 avdd.n461 avdd.t393 27.1302
R4004 avdd.n460 avdd.t406 27.1302
R4005 avdd.n419 avdd.t401 26.9438
R4006 avdd.n126 avdd.t387 26.9438
R4007 avdd.n199 avdd.t379 26.9438
R4008 avdd.n272 avdd.t392 26.9438
R4009 avdd.n345 avdd.t397 26.9438
R4010 avdd.n459 avdd.t395 26.9438
R4011 avdd.n429 dffrs_1.resetb 18.2415
R4012 avdd.n136 dffrs_5.resetb 18.2415
R4013 avdd.n209 dffrs_4.resetb 18.2415
R4014 avdd.n282 dffrs_3.resetb 18.2415
R4015 avdd.n355 dffrs_2.resetb 18.2415
R4016 avdd.n469 dffrs_0.resetb 18.2415
R4017 avdd.n394 avdd.n388 18.0418
R4018 avdd.n102 avdd.n96 18.0418
R4019 avdd.n175 avdd.n169 18.0418
R4020 avdd.n248 avdd.n242 18.0418
R4021 avdd.n321 avdd.n315 18.0418
R4022 avdd.n534 avdd.n533 18.0418
R4023 avdd.n422 avdd.n420 17.6364
R4024 avdd.n129 avdd.n127 17.6364
R4025 avdd.n202 avdd.n200 17.6364
R4026 avdd.n275 avdd.n273 17.6364
R4027 avdd.n348 avdd.n346 17.6364
R4028 avdd.n462 avdd.n460 17.6364
R4029 avdd.n387 avdd.n385 14.3609
R4030 avdd.n95 avdd.n93 14.3609
R4031 avdd.n168 avdd.n166 14.3609
R4032 avdd.n241 avdd.n239 14.3609
R4033 avdd.n314 avdd.n312 14.3609
R4034 avdd.n2 avdd.n0 14.3609
R4035 avdd.n394 avdd.n393 13.5174
R4036 avdd.n102 avdd.n101 13.5174
R4037 avdd.n175 avdd.n174 13.5174
R4038 avdd.n248 avdd.n247 13.5174
R4039 avdd.n321 avdd.n320 13.5174
R4040 avdd.n533 avdd.n7 13.5174
R4041 avdd.n405 avdd.n404 13.5005
R4042 avdd.n405 avdd.n399 13.5005
R4043 avdd.n417 avdd.n416 13.5005
R4044 avdd.n411 avdd.n410 13.5005
R4045 avdd.n429 avdd.n428 13.5005
R4046 avdd.n113 avdd.n112 13.5005
R4047 avdd.n113 avdd.n107 13.5005
R4048 avdd.n125 avdd.n124 13.5005
R4049 avdd.n119 avdd.n118 13.5005
R4050 avdd.n136 avdd.n135 13.5005
R4051 avdd.n186 avdd.n185 13.5005
R4052 avdd.n186 avdd.n180 13.5005
R4053 avdd.n198 avdd.n197 13.5005
R4054 avdd.n192 avdd.n191 13.5005
R4055 avdd.n209 avdd.n208 13.5005
R4056 avdd.n259 avdd.n258 13.5005
R4057 avdd.n259 avdd.n253 13.5005
R4058 avdd.n271 avdd.n270 13.5005
R4059 avdd.n265 avdd.n264 13.5005
R4060 avdd.n282 avdd.n281 13.5005
R4061 avdd.n332 avdd.n331 13.5005
R4062 avdd.n332 avdd.n326 13.5005
R4063 avdd.n344 avdd.n343 13.5005
R4064 avdd.n338 avdd.n337 13.5005
R4065 avdd.n355 avdd.n354 13.5005
R4066 avdd.n532 avdd.n531 13.5005
R4067 avdd.n532 avdd.n12 13.5005
R4068 avdd.n520 avdd.n519 13.5005
R4069 avdd.n526 avdd.n525 13.5005
R4070 avdd.n469 avdd.n468 13.5005
R4071 avdd.n423 avdd.n419 13.4839
R4072 avdd.n130 avdd.n126 13.4839
R4073 avdd.n203 avdd.n199 13.4839
R4074 avdd.n276 avdd.n272 13.4839
R4075 avdd.n349 avdd.n345 13.4839
R4076 avdd.n463 avdd.n459 13.4839
R4077 avdd.n422 avdd.n421 10.5752
R4078 avdd.n129 avdd.n128 10.5752
R4079 avdd.n202 avdd.n201 10.5752
R4080 avdd.n275 avdd.n274 10.5752
R4081 avdd.n348 avdd.n347 10.5752
R4082 avdd.n462 avdd.n461 10.5752
R4083 avdd.n393 avdd.n390 6.4802
R4084 avdd.n404 avdd.n401 6.4802
R4085 avdd.n399 avdd.n396 6.4802
R4086 avdd.n416 avdd.n413 6.4802
R4087 avdd.n410 avdd.n407 6.4802
R4088 avdd.n428 avdd.n425 6.4802
R4089 avdd.n101 avdd.n98 6.4802
R4090 avdd.n112 avdd.n109 6.4802
R4091 avdd.n107 avdd.n104 6.4802
R4092 avdd.n124 avdd.n121 6.4802
R4093 avdd.n118 avdd.n115 6.4802
R4094 avdd.n135 avdd.n132 6.4802
R4095 avdd.n174 avdd.n171 6.4802
R4096 avdd.n185 avdd.n182 6.4802
R4097 avdd.n180 avdd.n177 6.4802
R4098 avdd.n197 avdd.n194 6.4802
R4099 avdd.n191 avdd.n188 6.4802
R4100 avdd.n208 avdd.n205 6.4802
R4101 avdd.n247 avdd.n244 6.4802
R4102 avdd.n258 avdd.n255 6.4802
R4103 avdd.n253 avdd.n250 6.4802
R4104 avdd.n270 avdd.n267 6.4802
R4105 avdd.n264 avdd.n261 6.4802
R4106 avdd.n281 avdd.n278 6.4802
R4107 avdd.n320 avdd.n317 6.4802
R4108 avdd.n331 avdd.n328 6.4802
R4109 avdd.n326 avdd.n323 6.4802
R4110 avdd.n343 avdd.n340 6.4802
R4111 avdd.n337 avdd.n334 6.4802
R4112 avdd.n354 avdd.n351 6.4802
R4113 avdd.n7 avdd.n4 6.4802
R4114 avdd.n531 avdd.n528 6.4802
R4115 avdd.n12 avdd.n9 6.4802
R4116 avdd.n519 avdd.n516 6.4802
R4117 avdd.n525 avdd.n522 6.4802
R4118 avdd.n468 avdd.n465 6.4802
R4119 avdd.n393 avdd.n389 6.25878
R4120 avdd.n404 avdd.n400 6.25878
R4121 avdd.n399 avdd.n395 6.25878
R4122 avdd.n416 avdd.n412 6.25878
R4123 avdd.n410 avdd.n406 6.25878
R4124 avdd.n428 avdd.n424 6.25878
R4125 avdd.n101 avdd.n97 6.25878
R4126 avdd.n112 avdd.n108 6.25878
R4127 avdd.n107 avdd.n103 6.25878
R4128 avdd.n124 avdd.n120 6.25878
R4129 avdd.n118 avdd.n114 6.25878
R4130 avdd.n135 avdd.n131 6.25878
R4131 avdd.n174 avdd.n170 6.25878
R4132 avdd.n185 avdd.n181 6.25878
R4133 avdd.n180 avdd.n176 6.25878
R4134 avdd.n197 avdd.n193 6.25878
R4135 avdd.n191 avdd.n187 6.25878
R4136 avdd.n208 avdd.n204 6.25878
R4137 avdd.n247 avdd.n243 6.25878
R4138 avdd.n258 avdd.n254 6.25878
R4139 avdd.n253 avdd.n249 6.25878
R4140 avdd.n270 avdd.n266 6.25878
R4141 avdd.n264 avdd.n260 6.25878
R4142 avdd.n281 avdd.n277 6.25878
R4143 avdd.n320 avdd.n316 6.25878
R4144 avdd.n331 avdd.n327 6.25878
R4145 avdd.n326 avdd.n322 6.25878
R4146 avdd.n343 avdd.n339 6.25878
R4147 avdd.n337 avdd.n333 6.25878
R4148 avdd.n354 avdd.n350 6.25878
R4149 avdd.n7 avdd.n3 6.25878
R4150 avdd.n531 avdd.n527 6.25878
R4151 avdd.n12 avdd.n8 6.25878
R4152 avdd.n519 avdd.n515 6.25878
R4153 avdd.n525 avdd.n521 6.25878
R4154 avdd.n468 avdd.n464 6.25878
R4155 avdd.n423 avdd.n422 5.93546
R4156 avdd.n130 avdd.n129 5.93546
R4157 avdd.n203 avdd.n202 5.93546
R4158 avdd.n276 avdd.n275 5.93546
R4159 avdd.n349 avdd.n348 5.93546
R4160 avdd.n463 avdd.n462 5.93546
R4161 avdd.n393 avdd.n392 5.44497
R4162 avdd.n404 avdd.n403 5.44497
R4163 avdd.n399 avdd.n398 5.44497
R4164 avdd.n416 avdd.n415 5.44497
R4165 avdd.n410 avdd.n409 5.44497
R4166 avdd.n428 avdd.n427 5.44497
R4167 avdd.n101 avdd.n100 5.44497
R4168 avdd.n112 avdd.n111 5.44497
R4169 avdd.n107 avdd.n106 5.44497
R4170 avdd.n124 avdd.n123 5.44497
R4171 avdd.n118 avdd.n117 5.44497
R4172 avdd.n135 avdd.n134 5.44497
R4173 avdd.n174 avdd.n173 5.44497
R4174 avdd.n185 avdd.n184 5.44497
R4175 avdd.n180 avdd.n179 5.44497
R4176 avdd.n197 avdd.n196 5.44497
R4177 avdd.n191 avdd.n190 5.44497
R4178 avdd.n208 avdd.n207 5.44497
R4179 avdd.n247 avdd.n246 5.44497
R4180 avdd.n258 avdd.n257 5.44497
R4181 avdd.n253 avdd.n252 5.44497
R4182 avdd.n270 avdd.n269 5.44497
R4183 avdd.n264 avdd.n263 5.44497
R4184 avdd.n281 avdd.n280 5.44497
R4185 avdd.n320 avdd.n319 5.44497
R4186 avdd.n331 avdd.n330 5.44497
R4187 avdd.n326 avdd.n325 5.44497
R4188 avdd.n343 avdd.n342 5.44497
R4189 avdd.n337 avdd.n336 5.44497
R4190 avdd.n354 avdd.n353 5.44497
R4191 avdd.n7 avdd.n6 5.44497
R4192 avdd.n531 avdd.n530 5.44497
R4193 avdd.n12 avdd.n11 5.44497
R4194 avdd.n519 avdd.n518 5.44497
R4195 avdd.n525 avdd.n524 5.44497
R4196 avdd.n468 avdd.n467 5.44497
R4197 avdd.n387 avdd.n386 5.14711
R4198 avdd.n95 avdd.n94 5.14711
R4199 avdd.n168 avdd.n167 5.14711
R4200 avdd.n241 avdd.n240 5.14711
R4201 avdd.n314 avdd.n313 5.14711
R4202 avdd.n2 avdd.n1 5.14711
R4203 avdd.n511 avdd.n510 2.49936
R4204 avdd.n445 avdd.n444 2.49936
R4205 avdd.n371 avdd.n370 2.49936
R4206 avdd.n298 avdd.n297 2.49936
R4207 avdd.n225 avdd.n224 2.49936
R4208 avdd.n152 avdd.n151 2.49936
R4209 avdd.n510 avdd.n499 1.93883
R4210 avdd.n444 avdd.n433 1.93883
R4211 avdd.n370 avdd.n359 1.93883
R4212 avdd.n297 avdd.n286 1.93883
R4213 avdd.n224 avdd.n213 1.93883
R4214 avdd.n151 avdd.n140 1.93883
R4215 avdd.n392 avdd.t93 1.85637
R4216 avdd.n403 avdd.t299 1.85637
R4217 avdd.n398 avdd.t90 1.85637
R4218 avdd.n415 avdd.t265 1.85637
R4219 avdd.n409 avdd.t19 1.85637
R4220 avdd.n427 avdd.t287 1.85637
R4221 avdd.n100 avdd.t144 1.85637
R4222 avdd.n111 avdd.t293 1.85637
R4223 avdd.n106 avdd.t138 1.85637
R4224 avdd.n123 avdd.t231 1.85637
R4225 avdd.n117 avdd.t177 1.85637
R4226 avdd.n134 avdd.t41 1.85637
R4227 avdd.n173 avdd.t120 1.85637
R4228 avdd.n184 avdd.t319 1.85637
R4229 avdd.n179 avdd.t81 1.85637
R4230 avdd.n196 avdd.t193 1.85637
R4231 avdd.n190 avdd.t305 1.85637
R4232 avdd.n207 avdd.t281 1.85637
R4233 avdd.n246 avdd.t84 1.85637
R4234 avdd.n257 avdd.t247 1.85637
R4235 avdd.n252 avdd.t150 1.85637
R4236 avdd.n269 avdd.t63 1.85637
R4237 avdd.n263 avdd.t279 1.85637
R4238 avdd.n280 avdd.t217 1.85637
R4239 avdd.n319 avdd.t105 1.85637
R4240 avdd.n330 avdd.t245 1.85637
R4241 avdd.n325 avdd.t108 1.85637
R4242 avdd.n342 avdd.t325 1.85637
R4243 avdd.n336 avdd.t311 1.85637
R4244 avdd.n353 avdd.t365 1.85637
R4245 avdd.n6 avdd.t132 1.85637
R4246 avdd.n530 avdd.t187 1.85637
R4247 avdd.n11 avdd.t126 1.85637
R4248 avdd.n518 avdd.t329 1.85637
R4249 avdd.n524 avdd.t369 1.85637
R4250 avdd.n467 avdd.t51 1.85637
R4251 avdd.n138 avdd.n92 1.80479
R4252 avdd.n211 avdd.n76 1.80479
R4253 avdd.n284 avdd.n60 1.80479
R4254 avdd.n357 avdd.n44 1.80479
R4255 avdd.n431 avdd.n28 1.80479
R4256 avdd.n513 avdd.n470 1.80479
R4257 avdd.n161 avdd.n160 1.78583
R4258 avdd.n234 avdd.n233 1.78583
R4259 avdd.n307 avdd.n306 1.78583
R4260 avdd.n380 avdd.n379 1.78583
R4261 avdd.n454 avdd.n453 1.78583
R4262 avdd.n496 avdd.n495 1.78583
R4263 avdd.n164 avdd.t71 1.74654
R4264 avdd.n237 avdd.t73 1.74654
R4265 avdd.n310 avdd.t69 1.74654
R4266 avdd.n383 avdd.t171 1.74654
R4267 avdd.n457 avdd.t271 1.74654
R4268 avdd.n487 avdd.t173 1.74654
R4269 avdd.n486 avdd.t55 1.49467
R4270 avdd.n507 avdd.t49 1.49467
R4271 avdd.n506 avdd.t75 1.49467
R4272 avdd.n14 avdd.t357 1.49467
R4273 avdd.n441 avdd.t327 1.49467
R4274 avdd.n440 avdd.t219 1.49467
R4275 avdd.n30 avdd.t43 1.49467
R4276 avdd.n367 avdd.t67 1.49467
R4277 avdd.n366 avdd.t221 1.49467
R4278 avdd.n46 avdd.t313 1.49467
R4279 avdd.n294 avdd.t17 1.49467
R4280 avdd.n293 avdd.t47 1.49467
R4281 avdd.n62 avdd.t277 1.49467
R4282 avdd.n221 avdd.t37 1.49467
R4283 avdd.n220 avdd.t233 1.49467
R4284 avdd.n78 avdd.t185 1.49467
R4285 avdd.n148 avdd.t359 1.49467
R4286 avdd.n147 avdd.t3 1.49467
R4287 avdd.n77 avdd.t213 1.49467
R4288 avdd.n61 avdd.t169 1.49467
R4289 avdd.n45 avdd.t269 1.49467
R4290 avdd.n29 avdd.t191 1.49467
R4291 avdd.n13 avdd.t45 1.49467
R4292 avdd.n490 avdd.t175 1.49467
R4293 avdd.n500 avdd.t211 1.47383
R4294 avdd.n434 avdd.t223 1.47383
R4295 avdd.n360 avdd.t237 1.47383
R4296 avdd.n287 avdd.t57 1.47383
R4297 avdd.n214 avdd.t255 1.47383
R4298 avdd.n141 avdd.t259 1.47383
R4299 avdd.n80 avdd.t183 1.47383
R4300 avdd.n81 avdd.t181 1.47383
R4301 avdd.n82 avdd.t215 1.47383
R4302 avdd.n79 avdd.t337 1.47383
R4303 avdd.n64 avdd.t31 1.47383
R4304 avdd.n65 avdd.t29 1.47383
R4305 avdd.n66 avdd.t239 1.47383
R4306 avdd.n63 avdd.t355 1.47383
R4307 avdd.n48 avdd.t203 1.47383
R4308 avdd.n49 avdd.t205 1.47383
R4309 avdd.n50 avdd.t295 1.47383
R4310 avdd.n47 avdd.t201 1.47383
R4311 avdd.n32 avdd.t275 1.47383
R4312 avdd.n33 avdd.t273 1.47383
R4313 avdd.n34 avdd.t167 1.47383
R4314 avdd.n31 avdd.t261 1.47383
R4315 avdd.n16 avdd.t33 1.47383
R4316 avdd.n17 avdd.t35 1.47383
R4317 avdd.n18 avdd.t367 1.47383
R4318 avdd.n15 avdd.t307 1.47383
R4319 avdd.n482 avdd.t375 1.47383
R4320 avdd.n472 avdd.t377 1.47383
R4321 avdd.n471 avdd.t235 1.47383
R4322 avdd.n492 avdd.t189 1.47383
R4323 avdd.n210 avdd.n165 1.19311
R4324 avdd.n283 avdd.n238 1.19311
R4325 avdd.n356 avdd.n311 1.19311
R4326 avdd.n418 avdd.n384 1.19311
R4327 avdd.n514 avdd.n458 1.19311
R4328 avdd.n392 avdd.n391 1.04105
R4329 avdd.n403 avdd.n402 1.04105
R4330 avdd.n398 avdd.n397 1.04105
R4331 avdd.n415 avdd.n414 1.04105
R4332 avdd.n409 avdd.n408 1.04105
R4333 avdd.n427 avdd.n426 1.04105
R4334 avdd.n100 avdd.n99 1.04105
R4335 avdd.n111 avdd.n110 1.04105
R4336 avdd.n106 avdd.n105 1.04105
R4337 avdd.n123 avdd.n122 1.04105
R4338 avdd.n117 avdd.n116 1.04105
R4339 avdd.n134 avdd.n133 1.04105
R4340 avdd.n173 avdd.n172 1.04105
R4341 avdd.n184 avdd.n183 1.04105
R4342 avdd.n179 avdd.n178 1.04105
R4343 avdd.n196 avdd.n195 1.04105
R4344 avdd.n190 avdd.n189 1.04105
R4345 avdd.n207 avdd.n206 1.04105
R4346 avdd.n246 avdd.n245 1.04105
R4347 avdd.n257 avdd.n256 1.04105
R4348 avdd.n252 avdd.n251 1.04105
R4349 avdd.n269 avdd.n268 1.04105
R4350 avdd.n263 avdd.n262 1.04105
R4351 avdd.n280 avdd.n279 1.04105
R4352 avdd.n319 avdd.n318 1.04105
R4353 avdd.n330 avdd.n329 1.04105
R4354 avdd.n325 avdd.n324 1.04105
R4355 avdd.n342 avdd.n341 1.04105
R4356 avdd.n336 avdd.n335 1.04105
R4357 avdd.n353 avdd.n352 1.04105
R4358 avdd.n6 avdd.n5 1.04105
R4359 avdd.n530 avdd.n529 1.04105
R4360 avdd.n11 avdd.n10 1.04105
R4361 avdd.n518 avdd.n517 1.04105
R4362 avdd.n524 avdd.n523 1.04105
R4363 avdd.n467 avdd.n466 1.04105
R4364 avdd.n138 avdd.n137 0.809622
R4365 avdd.n211 avdd.n210 0.809622
R4366 avdd.n284 avdd.n283 0.809622
R4367 avdd.n357 avdd.n356 0.809622
R4368 avdd.n431 avdd.n430 0.809622
R4369 avdd.n514 avdd.n513 0.809622
R4370 avdd.n503 avdd.n500 0.788
R4371 avdd.n504 avdd.n503 0.788
R4372 avdd.n506 avdd.n505 0.788
R4373 avdd.n437 avdd.n434 0.788
R4374 avdd.n438 avdd.n437 0.788
R4375 avdd.n440 avdd.n439 0.788
R4376 avdd.n363 avdd.n360 0.788
R4377 avdd.n364 avdd.n363 0.788
R4378 avdd.n366 avdd.n365 0.788
R4379 avdd.n290 avdd.n287 0.788
R4380 avdd.n291 avdd.n290 0.788
R4381 avdd.n293 avdd.n292 0.788
R4382 avdd.n217 avdd.n214 0.788
R4383 avdd.n218 avdd.n217 0.788
R4384 avdd.n220 avdd.n219 0.788
R4385 avdd.n144 avdd.n141 0.788
R4386 avdd.n145 avdd.n144 0.788
R4387 avdd.n147 avdd.n146 0.788
R4388 avdd.n88 avdd.n81 0.788
R4389 avdd.n89 avdd.n88 0.788
R4390 avdd.n90 avdd.n82 0.788
R4391 avdd.n91 avdd.n90 0.788
R4392 avdd.n86 avdd.n80 0.788
R4393 avdd.n158 avdd.n79 0.788
R4394 avdd.n159 avdd.n158 0.788
R4395 avdd.n157 avdd.n77 0.788
R4396 avdd.n72 avdd.n65 0.788
R4397 avdd.n73 avdd.n72 0.788
R4398 avdd.n74 avdd.n66 0.788
R4399 avdd.n75 avdd.n74 0.788
R4400 avdd.n70 avdd.n64 0.788
R4401 avdd.n231 avdd.n63 0.788
R4402 avdd.n232 avdd.n231 0.788
R4403 avdd.n230 avdd.n61 0.788
R4404 avdd.n56 avdd.n49 0.788
R4405 avdd.n57 avdd.n56 0.788
R4406 avdd.n58 avdd.n50 0.788
R4407 avdd.n59 avdd.n58 0.788
R4408 avdd.n54 avdd.n48 0.788
R4409 avdd.n304 avdd.n47 0.788
R4410 avdd.n305 avdd.n304 0.788
R4411 avdd.n303 avdd.n45 0.788
R4412 avdd.n40 avdd.n33 0.788
R4413 avdd.n41 avdd.n40 0.788
R4414 avdd.n42 avdd.n34 0.788
R4415 avdd.n43 avdd.n42 0.788
R4416 avdd.n38 avdd.n32 0.788
R4417 avdd.n377 avdd.n31 0.788
R4418 avdd.n378 avdd.n377 0.788
R4419 avdd.n376 avdd.n29 0.788
R4420 avdd.n24 avdd.n17 0.788
R4421 avdd.n25 avdd.n24 0.788
R4422 avdd.n26 avdd.n18 0.788
R4423 avdd.n27 avdd.n26 0.788
R4424 avdd.n22 avdd.n16 0.788
R4425 avdd.n451 avdd.n15 0.788
R4426 avdd.n452 avdd.n451 0.788
R4427 avdd.n450 avdd.n13 0.788
R4428 avdd.n479 avdd.n472 0.788
R4429 avdd.n480 avdd.n479 0.788
R4430 avdd.n477 avdd.n471 0.788
R4431 avdd.n478 avdd.n477 0.788
R4432 avdd.n482 avdd.n481 0.788
R4433 avdd.n493 avdd.n492 0.788
R4434 avdd.n494 avdd.n493 0.788
R4435 avdd.n491 avdd.n490 0.788
R4436 avdd.n388 avdd.n387 0.754571
R4437 avdd.n96 avdd.n95 0.754571
R4438 avdd.n169 avdd.n168 0.754571
R4439 avdd.n242 avdd.n241 0.754571
R4440 avdd.n315 avdd.n314 0.754571
R4441 avdd.n534 avdd.n2 0.754571
R4442 avdd.n389 avdd.t267 0.7285
R4443 avdd.n389 avdd.t243 0.7285
R4444 avdd.n400 avdd.t25 0.7285
R4445 avdd.n400 avdd.t156 0.7285
R4446 avdd.n395 avdd.t199 0.7285
R4447 avdd.n395 avdd.t263 0.7285
R4448 avdd.n412 avdd.t241 0.7285
R4449 avdd.n412 avdd.t349 0.7285
R4450 avdd.n406 avdd.t141 0.7285
R4451 avdd.n406 avdd.t285 0.7285
R4452 avdd.n424 avdd.t249 0.7285
R4453 avdd.n424 avdd.t87 0.7285
R4454 avdd.n97 avdd.t229 0.7285
R4455 avdd.n97 avdd.t291 0.7285
R4456 avdd.n108 avdd.t339 0.7285
R4457 avdd.n108 avdd.t111 0.7285
R4458 avdd.n103 avdd.t335 0.7285
R4459 avdd.n103 avdd.t227 0.7285
R4460 avdd.n120 avdd.t251 0.7285
R4461 avdd.n120 avdd.t9 0.7285
R4462 avdd.n114 avdd.t96 0.7285
R4463 avdd.n114 avdd.t39 0.7285
R4464 avdd.n131 avdd.t309 0.7285
R4465 avdd.n131 avdd.t135 0.7285
R4466 avdd.n170 avdd.t197 0.7285
R4467 avdd.n170 avdd.t289 0.7285
R4468 avdd.n181 avdd.t345 0.7285
R4469 avdd.n181 avdd.t165 0.7285
R4470 avdd.n176 avdd.t353 0.7285
R4471 avdd.n176 avdd.t195 0.7285
R4472 avdd.n193 avdd.t257 0.7285
R4473 avdd.n193 avdd.t347 0.7285
R4474 avdd.n187 avdd.t117 0.7285
R4475 avdd.n187 avdd.t283 0.7285
R4476 avdd.n204 avdd.t253 0.7285
R4477 avdd.n204 avdd.t99 0.7285
R4478 avdd.n243 avdd.t65 0.7285
R4479 avdd.n243 avdd.t303 0.7285
R4480 avdd.n254 avdd.t351 0.7285
R4481 avdd.n254 avdd.t114 0.7285
R4482 avdd.n249 avdd.t61 0.7285
R4483 avdd.n249 avdd.t361 0.7285
R4484 avdd.n266 avdd.t301 0.7285
R4485 avdd.n266 avdd.t7 0.7285
R4486 avdd.n260 avdd.t78 0.7285
R4487 avdd.n260 avdd.t225 0.7285
R4488 avdd.n277 avdd.t297 0.7285
R4489 avdd.n277 avdd.t147 0.7285
R4490 avdd.n316 avdd.t323 0.7285
R4491 avdd.n316 avdd.t209 0.7285
R4492 avdd.n327 avdd.t27 0.7285
R4493 avdd.n327 avdd.t102 0.7285
R4494 avdd.n322 avdd.t15 0.7285
R4495 avdd.n322 avdd.t321 0.7285
R4496 avdd.n339 avdd.t207 0.7285
R4497 avdd.n339 avdd.t23 0.7285
R4498 avdd.n333 avdd.t153 0.7285
R4499 avdd.n333 avdd.t363 0.7285
R4500 avdd.n350 avdd.t179 0.7285
R4501 avdd.n350 avdd.t123 0.7285
R4502 avdd.n3 avdd.t333 0.7285
R4503 avdd.n3 avdd.t21 0.7285
R4504 avdd.n527 avdd.t341 0.7285
R4505 avdd.n527 avdd.t129 0.7285
R4506 avdd.n8 avdd.t13 0.7285
R4507 avdd.n8 avdd.t331 0.7285
R4508 avdd.n515 avdd.t5 0.7285
R4509 avdd.n515 avdd.t343 0.7285
R4510 avdd.n521 avdd.t159 0.7285
R4511 avdd.n521 avdd.t53 0.7285
R4512 avdd.n464 avdd.t371 0.7285
R4513 avdd.n464 avdd.t162 0.7285
R4514 avdd.n509 avdd.n500 0.561043
R4515 avdd.n443 avdd.n434 0.561043
R4516 avdd.n369 avdd.n360 0.561043
R4517 avdd.n296 avdd.n287 0.561043
R4518 avdd.n223 avdd.n214 0.561043
R4519 avdd.n150 avdd.n141 0.561043
R4520 avdd.n154 avdd.n80 0.561043
R4521 avdd.n153 avdd.n81 0.561043
R4522 avdd.n139 avdd.n82 0.561043
R4523 avdd.n162 avdd.n79 0.561043
R4524 avdd.n227 avdd.n64 0.561043
R4525 avdd.n226 avdd.n65 0.561043
R4526 avdd.n212 avdd.n66 0.561043
R4527 avdd.n235 avdd.n63 0.561043
R4528 avdd.n300 avdd.n48 0.561043
R4529 avdd.n299 avdd.n49 0.561043
R4530 avdd.n285 avdd.n50 0.561043
R4531 avdd.n308 avdd.n47 0.561043
R4532 avdd.n373 avdd.n32 0.561043
R4533 avdd.n372 avdd.n33 0.561043
R4534 avdd.n358 avdd.n34 0.561043
R4535 avdd.n381 avdd.n31 0.561043
R4536 avdd.n447 avdd.n16 0.561043
R4537 avdd.n446 avdd.n17 0.561043
R4538 avdd.n432 avdd.n18 0.561043
R4539 avdd.n455 avdd.n15 0.561043
R4540 avdd.n497 avdd.n482 0.561043
R4541 avdd.n498 avdd.n472 0.561043
R4542 avdd.n512 avdd.n471 0.561043
R4543 avdd.n492 avdd.n483 0.561043
R4544 avdd.n488 avdd.n487 0.510024
R4545 avdd.n165 avdd.n163 0.490037
R4546 avdd.n238 avdd.n236 0.490037
R4547 avdd.n311 avdd.n309 0.490037
R4548 avdd.n384 avdd.n382 0.490037
R4549 avdd.n458 avdd.n456 0.490037
R4550 avdd.n165 avdd.n164 0.436534
R4551 avdd.n238 avdd.n237 0.436534
R4552 avdd.n311 avdd.n310 0.436534
R4553 avdd.n384 avdd.n383 0.436534
R4554 avdd.n458 avdd.n457 0.436534
R4555 avdd.n489 avdd.n488 0.415037
R4556 avdd.n509 avdd.n508 0.255737
R4557 avdd.n443 avdd.n442 0.255737
R4558 avdd.n369 avdd.n368 0.255737
R4559 avdd.n296 avdd.n295 0.255737
R4560 avdd.n223 avdd.n222 0.255737
R4561 avdd.n150 avdd.n149 0.255737
R4562 avdd.n163 avdd.n162 0.255737
R4563 avdd.n236 avdd.n235 0.255737
R4564 avdd.n309 avdd.n308 0.255737
R4565 avdd.n382 avdd.n381 0.255737
R4566 avdd.n456 avdd.n455 0.255737
R4567 avdd.n489 avdd.n483 0.255737
R4568 avdd.n162 avdd.n161 0.2165
R4569 avdd.n235 avdd.n234 0.2165
R4570 avdd.n308 avdd.n307 0.2165
R4571 avdd.n381 avdd.n380 0.2165
R4572 avdd.n455 avdd.n454 0.2165
R4573 avdd.n496 avdd.n483 0.2165
R4574 avdd.n161 avdd.n154 0.148424
R4575 avdd.n234 avdd.n227 0.148424
R4576 avdd.n307 avdd.n300 0.148424
R4577 avdd.n380 avdd.n373 0.148424
R4578 avdd.n454 avdd.n447 0.148424
R4579 avdd.n497 avdd.n496 0.148424
R4580 dffrs_1.resetb avdd.n423 0.136036
R4581 dffrs_5.resetb avdd.n130 0.136036
R4582 dffrs_4.resetb avdd.n203 0.136036
R4583 dffrs_3.resetb avdd.n276 0.136036
R4584 dffrs_2.resetb avdd.n349 0.136036
R4585 dffrs_0.resetb avdd.n463 0.136036
R4586 avdd.n510 avdd.n509 0.0635
R4587 avdd.n444 avdd.n443 0.0635
R4588 avdd.n370 avdd.n369 0.0635
R4589 avdd.n297 avdd.n296 0.0635
R4590 avdd.n224 avdd.n223 0.0635
R4591 avdd.n151 avdd.n150 0.0635
R4592 avdd.n154 avdd.n153 0.0452384
R4593 avdd.n227 avdd.n226 0.0452384
R4594 avdd.n300 avdd.n299 0.0452384
R4595 avdd.n373 avdd.n372 0.0452384
R4596 avdd.n447 avdd.n446 0.0452384
R4597 avdd.n498 avdd.n497 0.0452384
R4598 avdd.n119 avdd.n113 0.0405727
R4599 avdd.n192 avdd.n186 0.0405727
R4600 avdd.n265 avdd.n259 0.0405727
R4601 avdd.n338 avdd.n332 0.0405727
R4602 avdd.n411 avdd.n405 0.0405727
R4603 avdd.n532 avdd.n526 0.0405727
R4604 avdd.n388 dffrs_1.setb 0.032
R4605 avdd.n96 dffrs_5.setb 0.032
R4606 avdd.n169 dffrs_4.setb 0.032
R4607 avdd.n242 dffrs_3.setb 0.032
R4608 avdd.n315 dffrs_2.setb 0.032
R4609 dffrs_0.setb avdd.n534 0.032
R4610 avdd.n508 avdd.n506 0.0313054
R4611 avdd.n508 avdd.n507 0.0313054
R4612 avdd.n442 avdd.n440 0.0313054
R4613 avdd.n442 avdd.n441 0.0313054
R4614 avdd.n368 avdd.n366 0.0313054
R4615 avdd.n368 avdd.n367 0.0313054
R4616 avdd.n295 avdd.n293 0.0313054
R4617 avdd.n295 avdd.n294 0.0313054
R4618 avdd.n222 avdd.n220 0.0313054
R4619 avdd.n222 avdd.n221 0.0313054
R4620 avdd.n149 avdd.n147 0.0313054
R4621 avdd.n149 avdd.n148 0.0313054
R4622 avdd.n163 avdd.n77 0.0313054
R4623 avdd.n163 avdd.n78 0.0313054
R4624 avdd.n236 avdd.n61 0.0313054
R4625 avdd.n236 avdd.n62 0.0313054
R4626 avdd.n309 avdd.n45 0.0313054
R4627 avdd.n309 avdd.n46 0.0313054
R4628 avdd.n382 avdd.n29 0.0313054
R4629 avdd.n382 avdd.n30 0.0313054
R4630 avdd.n456 avdd.n13 0.0313054
R4631 avdd.n456 avdd.n14 0.0313054
R4632 avdd.n490 avdd.n489 0.0313054
R4633 avdd.n489 avdd.n486 0.0313054
R4634 avdd.n152 avdd.n139 0.0295407
R4635 avdd.n225 avdd.n212 0.0295407
R4636 avdd.n298 avdd.n285 0.0295407
R4637 avdd.n371 avdd.n358 0.0295407
R4638 avdd.n445 avdd.n432 0.0295407
R4639 avdd.n512 avdd.n511 0.0295407
R4640 avdd.n137 avdd.n125 0.0288636
R4641 avdd.n210 avdd.n198 0.0288636
R4642 avdd.n283 avdd.n271 0.0288636
R4643 avdd.n356 avdd.n344 0.0288636
R4644 avdd.n520 avdd.n514 0.0288636
R4645 avdd.n418 avdd.n417 0.0288455
R4646 avdd.n113 avdd.n102 0.0237
R4647 avdd.n186 avdd.n175 0.0237
R4648 avdd.n259 avdd.n248 0.0237
R4649 avdd.n332 avdd.n321 0.0237
R4650 avdd.n405 avdd.n394 0.0237
R4651 avdd.n533 avdd.n532 0.0237
R4652 avdd.n153 avdd.n152 0.0161977
R4653 avdd.n226 avdd.n225 0.0161977
R4654 avdd.n299 avdd.n298 0.0161977
R4655 avdd.n372 avdd.n371 0.0161977
R4656 avdd.n446 avdd.n445 0.0161977
R4657 avdd.n511 avdd.n498 0.0161977
R4658 avdd.n139 avdd.n138 0.0129273
R4659 avdd.n212 avdd.n211 0.0129273
R4660 avdd.n285 avdd.n284 0.0129273
R4661 avdd.n358 avdd.n357 0.0129273
R4662 avdd.n432 avdd.n431 0.0129273
R4663 avdd.n513 avdd.n512 0.0129273
R4664 avdd.n488 avdd 0.0128676
R4665 avdd.n137 avdd.n136 0.0122273
R4666 avdd.n210 avdd.n209 0.0122273
R4667 avdd.n283 avdd.n282 0.0122273
R4668 avdd.n356 avdd.n355 0.0122273
R4669 avdd.n430 avdd.n429 0.0122273
R4670 avdd.n514 avdd.n469 0.0122273
R4671 avdd.n125 avdd.n119 0.000518182
R4672 avdd.n198 avdd.n192 0.000518182
R4673 avdd.n271 avdd.n265 0.000518182
R4674 avdd.n344 avdd.n338 0.000518182
R4675 avdd.n417 avdd.n411 0.000518182
R4676 avdd.n430 avdd.n418 0.000518182
R4677 avdd.n526 avdd.n520 0.000518182
R4678 avss.n259 avss.n258 21124.8
R4679 avss.n216 avss.n215 21124.8
R4680 avss.n173 avss.n172 21124.8
R4681 avss.n124 avss.n51 21034.5
R4682 avss.n787 avss.n786 21034.5
R4683 avss.n321 avss.n301 21026.3
R4684 avss.n374 avss.n373 21012.5
R4685 avss.n474 avss.n473 21012.5
R4686 avss.n574 avss.n573 21012.5
R4687 avss.n674 avss.n673 21012.5
R4688 avss.n757 avss.n756 21000
R4689 avss.n825 avss.n824 21000
R4690 avss.n381 avss.n267 16221.9
R4691 avss.n481 avss.n224 16221.9
R4692 avss.n581 avss.n181 16221.9
R4693 avss.n681 avss.n132 16221.9
R4694 avss.n785 avss.n53 16221.9
R4695 avss.n836 avss.n833 11510.4
R4696 avss.n382 avss.n381 11510.4
R4697 avss.n482 avss.n481 11510.4
R4698 avss.n582 avss.n581 11510.4
R4699 avss.n682 avss.n681 11510.4
R4700 avss.n764 avss.n53 11510.4
R4701 avss.n836 avss.n6 11510.4
R4702 avss.n826 avss.n825 7422.73
R4703 avss.n758 avss.n757 7422.73
R4704 avss.n373 avss.n372 7422.62
R4705 avss.n473 avss.n472 7422.62
R4706 avss.n573 avss.n572 7422.62
R4707 avss.n673 avss.n672 7422.62
R4708 avss.n423 avss.n422 6961.73
R4709 avss.n523 avss.n522 6961.73
R4710 avss.n623 avss.n622 6961.73
R4711 avss.n716 avss.n715 6961.73
R4712 avss.n55 avss.n50 6961.73
R4713 avss.n854 avss.n5 6190.48
R4714 avss.n781 avss.n81 6190.48
R4715 avss.n699 avss.n139 6190.48
R4716 avss.n606 avss.n182 6190.48
R4717 avss.n506 avss.n225 6190.48
R4718 avss.n406 avss.n268 6190.48
R4719 avss.n323 avss.n322 5557.62
R4720 avss.n323 avss.n291 5551.58
R4721 avss.n423 avss.n250 5551.58
R4722 avss.n523 avss.n207 5551.58
R4723 avss.n623 avss.n164 5551.58
R4724 avss.n716 avss.n116 5551.58
R4725 avss.n55 avss.n42 5551.58
R4726 avss.n408 avss.n249 5290.17
R4727 avss.n508 avss.n206 5290.17
R4728 avss.n608 avss.n163 5290.17
R4729 avss.n701 avss.n115 5286.93
R4730 avss.n783 avss.n41 5286.93
R4731 avss.n854 avss.n853 4683.14
R4732 avss.n300 avss.n299 4273.71
R4733 avss.n409 avss.n408 4062.5
R4734 avss.n509 avss.n508 4062.5
R4735 avss.n609 avss.n608 4062.5
R4736 avss.n702 avss.n701 4062.5
R4737 avss.n784 avss.n783 4062.5
R4738 avss.n322 avss.n300 3568.02
R4739 avss.n854 avss.n6 3123.51
R4740 avss.n374 avss.n284 2944.22
R4741 avss.n474 avss.n241 2944.22
R4742 avss.n574 avss.n198 2944.22
R4743 avss.n674 avss.n155 2944.22
R4744 avss.n756 avss.n750 2944.22
R4745 avss.n824 avss.n822 2944.22
R4746 avss.n267 avss.n258 2845.46
R4747 avss.n224 avss.n215 2845.46
R4748 avss.n181 avss.n172 2845.46
R4749 avss.n786 avss.n785 2845.46
R4750 avss.n132 avss.n124 2843.75
R4751 avss.n325 avss.n283 2257.8
R4752 avss.n425 avss.n240 2257.8
R4753 avss.n525 avss.n197 2257.8
R4754 avss.n625 avss.n154 2257.8
R4755 avss.n97 avss.n52 2257.8
R4756 avss.n789 avss.n23 2257.8
R4757 avss.n702 avss.n132 1878.69
R4758 avss.n409 avss.n267 1876.98
R4759 avss.n509 avss.n224 1876.98
R4760 avss.n609 avss.n181 1876.98
R4761 avss.n785 avss.n784 1876.98
R4762 avss.n347 avss.n346 1486.9
R4763 avss.n309 avss.n300 1212.42
R4764 avss.n422 avss.n258 1205.08
R4765 avss.n522 avss.n215 1205.08
R4766 avss.n622 avss.n172 1205.08
R4767 avss.n715 avss.n124 1205.08
R4768 avss.n786 avss.n50 1205.08
R4769 avss.n301 avss.n267 1135.55
R4770 avss.n259 avss.n224 1135.55
R4771 avss.n216 avss.n181 1135.55
R4772 avss.n173 avss.n132 1135.55
R4773 avss.n785 avss.n51 1135.55
R4774 avss.n788 avss.n787 1135.55
R4775 avss.n325 avss.n267 1122.24
R4776 avss.n425 avss.n224 1122.24
R4777 avss.n525 avss.n181 1122.24
R4778 avss.n625 avss.n132 1122.24
R4779 avss.n785 avss.n52 1122.24
R4780 avss.n789 avss.n788 1122.24
R4781 avss.n739 avss.n738 977.434
R4782 avss.n811 avss.n810 977.434
R4783 avss.n447 avss.n446 977.068
R4784 avss.n547 avss.n546 977.068
R4785 avss.n647 avss.n646 977.068
R4786 avss.n738 avss.n115 904.402
R4787 avss.n810 avss.n41 904.402
R4788 avss.n446 avss.n249 904.062
R4789 avss.n546 avss.n206 904.062
R4790 avss.n646 avss.n163 904.062
R4791 avss.n322 avss.n321 897.806
R4792 avss.n323 avss.n298 832.22
R4793 avss.n423 avss.n257 832.22
R4794 avss.n523 avss.n214 832.22
R4795 avss.n623 avss.n171 832.22
R4796 avss.n716 avss.n123 832.22
R4797 avss.n56 avss.n55 832.22
R4798 avss.n324 avss.n323 832.101
R4799 avss.n424 avss.n423 832.101
R4800 avss.n524 avss.n523 832.101
R4801 avss.n624 avss.n623 832.101
R4802 avss.n717 avss.n716 832.101
R4803 avss.n55 avss.n54 832.101
R4804 avss.n75 avss.n41 784.409
R4805 avss.n133 avss.n115 784.37
R4806 avss.n588 avss.n163 784.37
R4807 avss.n488 avss.n206 784.37
R4808 avss.n388 avss.n249 784.37
R4809 avss.n788 avss.n6 697.039
R4810 avss.n374 avss.n283 665.564
R4811 avss.n474 avss.n240 665.564
R4812 avss.n574 avss.n197 665.564
R4813 avss.n674 avss.n154 665.564
R4814 avss.n756 avss.n97 665.564
R4815 avss.n824 avss.n23 665.564
R4816 avss.n822 avss.n821 654.253
R4817 avss.n750 avss.n749 654.253
R4818 avss.n156 avss.n155 654.005
R4819 avss.n199 avss.n198 654.005
R4820 avss.n242 avss.n241 654.005
R4821 avss.n285 avss.n284 654.005
R4822 avss.n750 avss.n98 648.784
R4823 avss.n822 avss.n24 648.784
R4824 avss.n348 avss.n284 648.54
R4825 avss.n448 avss.n241 648.54
R4826 avss.n548 avss.n198 648.54
R4827 avss.n648 avss.n155 648.54
R4828 avss.t134 avss.n826 590.909
R4829 avss.n827 avss.t134 590.909
R4830 avss.n827 avss.t252 590.909
R4831 avss.n833 avss.t181 590.909
R4832 avss.n833 avss.t35 590.909
R4833 avss.t37 avss.n832 590.909
R4834 avss.t253 avss.n375 590.909
R4835 avss.n379 avss.t253 590.909
R4836 avss.t136 avss.n379 590.909
R4837 avss.n381 avss.t186 590.909
R4838 avss.n381 avss.t179 590.909
R4839 avss.n405 avss.t118 590.909
R4840 avss.t259 avss.n475 590.909
R4841 avss.n479 avss.t259 590.909
R4842 avss.t125 avss.n479 590.909
R4843 avss.n481 avss.t128 590.909
R4844 avss.n481 avss.t155 590.909
R4845 avss.n505 avss.t195 590.909
R4846 avss.t130 avss.n575 590.909
R4847 avss.n579 avss.t130 590.909
R4848 avss.t104 avss.n579 590.909
R4849 avss.n581 avss.t187 590.909
R4850 avss.n581 avss.t44 590.909
R4851 avss.n605 avss.t221 590.909
R4852 avss.t112 avss.n675 590.909
R4853 avss.n679 avss.t112 590.909
R4854 avss.t55 avss.n679 590.909
R4855 avss.n681 avss.t123 590.909
R4856 avss.n681 avss.t16 590.909
R4857 avss.n698 avss.t0 590.909
R4858 avss.t139 avss.n758 590.909
R4859 avss.n762 avss.t139 590.909
R4860 avss.t209 avss.n762 590.909
R4861 avss.n764 avss.t274 590.909
R4862 avss.t234 avss.n764 590.909
R4863 avss.n765 avss.t232 590.909
R4864 avss.n755 avss.t202 590.909
R4865 avss.t202 avss.n754 590.909
R4866 avss.n754 avss.t107 590.909
R4867 avss.t124 avss.n53 590.909
R4868 avss.t275 avss.n53 590.909
R4869 avss.n780 avss.t261 590.909
R4870 avss.n823 avss.t280 590.909
R4871 avss.n837 avss.t280 590.909
R4872 avss.n837 avss.t103 590.909
R4873 avss.t54 avss.n836 590.909
R4874 avss.n836 avss.t215 590.909
R4875 avss.n855 avss.t212 590.909
R4876 avss.n372 avss.t217 590.462
R4877 avss.t217 avss.n371 590.462
R4878 avss.n371 avss.t228 590.462
R4879 avss.n382 avss.t4 590.462
R4880 avss.t265 avss.n382 590.462
R4881 avss.n383 avss.t263 590.462
R4882 avss.n472 avss.t169 590.462
R4883 avss.t169 avss.n471 590.462
R4884 avss.n471 avss.t165 590.462
R4885 avss.n482 avss.t120 590.462
R4886 avss.t27 avss.n482 590.462
R4887 avss.n483 avss.t29 590.462
R4888 avss.n572 avss.t236 590.462
R4889 avss.t236 avss.n571 590.462
R4890 avss.n571 avss.t31 590.462
R4891 avss.n582 avss.t34 590.462
R4892 avss.t10 avss.n582 590.462
R4893 avss.n583 avss.t12 590.462
R4894 avss.n672 avss.t150 590.462
R4895 avss.t150 avss.n671 590.462
R4896 avss.n671 avss.t138 590.462
R4897 avss.n682 avss.t43 590.462
R4898 avss.t50 avss.n682 590.462
R4899 avss.n683 avss.t52 590.462
R4900 avss.n309 avss.t242 582.165
R4901 avss.t65 avss.n298 582.165
R4902 avss.n410 avss.t255 582.165
R4903 avss.t88 avss.n257 582.165
R4904 avss.n510 avss.t48 582.165
R4905 avss.t69 avss.n214 582.165
R4906 avss.n610 avss.t9 582.165
R4907 avss.t92 avss.n171 582.165
R4908 avss.n703 avss.t129 582.165
R4909 avss.t82 avss.n123 582.165
R4910 avss.n74 avss.t8 582.165
R4911 avss.n56 avss.t59 582.165
R4912 avss.t250 avss.n324 581.712
R4913 avss.n326 avss.t198 581.712
R4914 avss.n320 avss.t144 581.712
R4915 avss.n302 avss.t71 581.712
R4916 avss.t248 avss.n424 581.712
R4917 avss.n426 avss.t229 581.712
R4918 avss.n421 avss.t177 581.712
R4919 avss.n260 avss.t99 581.712
R4920 avss.t245 avss.n524 581.712
R4921 avss.n526 avss.t171 581.712
R4922 avss.n521 avss.t269 581.712
R4923 avss.n217 avss.t80 581.712
R4924 avss.t247 avss.n624 581.712
R4925 avss.n626 avss.t160 581.712
R4926 avss.n621 avss.t204 581.712
R4927 avss.n174 avss.t94 581.712
R4928 avss.t22 avss.n717 581.712
R4929 avss.n718 avss.t270 581.712
R4930 avss.n714 avss.t225 581.712
R4931 avss.n125 avss.t85 581.712
R4932 avss.n54 avss.t251 581.712
R4933 avss.n790 avss.t121 581.712
R4934 avss.n60 avss.t238 581.712
R4935 avss.t63 avss.n49 581.712
R4936 avss.t197 avss.n334 581.712
R4937 avss.n335 avss.t145 581.712
R4938 avss.t173 avss.n434 581.712
R4939 avss.n435 avss.t175 581.712
R4940 avss.t152 avss.n534 581.712
R4941 avss.n535 avss.t267 581.712
R4942 avss.t41 avss.n634 581.712
R4943 avss.n635 avss.t206 581.712
R4944 avss.t164 avss.n726 581.712
R4945 avss.n727 avss.t257 581.712
R4946 avss.t18 avss.n798 581.712
R4947 avss.n799 avss.t239 581.712
R4948 avss.n701 avss.n699 574.192
R4949 avss.n408 avss.n406 574.061
R4950 avss.n508 avss.n506 574.061
R4951 avss.n608 avss.n606 574.061
R4952 avss.n783 avss.n781 574.061
R4953 avss.n334 avss.n291 548.058
R4954 avss.n434 avss.n250 548.058
R4955 avss.n534 avss.n207 548.058
R4956 avss.n634 avss.n164 548.058
R4957 avss.n726 avss.n116 548.058
R4958 avss.n798 avss.n42 548.058
R4959 avss.t252 avss.t181 502.274
R4960 avss.t35 avss.t37 502.274
R4961 avss.t186 avss.t136 502.274
R4962 avss.t179 avss.t118 502.274
R4963 avss.t128 avss.t125 502.274
R4964 avss.t155 avss.t195 502.274
R4965 avss.t187 avss.t104 502.274
R4966 avss.t44 avss.t221 502.274
R4967 avss.t123 avss.t55 502.274
R4968 avss.t16 avss.t0 502.274
R4969 avss.t274 avss.t209 502.274
R4970 avss.t232 avss.t234 502.274
R4971 avss.t107 avss.t124 502.274
R4972 avss.t261 avss.t275 502.274
R4973 avss.t103 avss.t54 502.274
R4974 avss.t215 avss.t212 502.274
R4975 avss.t228 avss.t4 501.892
R4976 avss.t263 avss.t265 501.892
R4977 avss.t165 avss.t120 501.892
R4978 avss.t29 avss.t27 501.892
R4979 avss.t31 avss.t34 501.892
R4980 avss.t12 avss.t10 501.892
R4981 avss.t138 avss.t43 501.892
R4982 avss.t52 avss.t50 501.892
R4983 avss.n345 avss.n291 484.702
R4984 avss.n445 avss.n250 484.702
R4985 avss.n545 avss.n207 484.702
R4986 avss.n645 avss.n164 484.702
R4987 avss.n737 avss.n116 484.702
R4988 avss.n809 avss.n42 484.702
R4989 avss.t242 avss.t143 465.733
R4990 avss.t143 avss.t65 465.733
R4991 avss.t255 avss.t178 465.733
R4992 avss.t178 avss.t88 465.733
R4993 avss.t48 avss.t49 465.733
R4994 avss.t49 avss.t69 465.733
R4995 avss.t9 avss.t205 465.733
R4996 avss.t205 avss.t92 465.733
R4997 avss.t129 avss.t256 465.733
R4998 avss.t256 avss.t82 465.733
R4999 avss.t241 avss.t8 465.733
R5000 avss.t59 avss.t241 465.733
R5001 avss.t96 avss.t250 465.37
R5002 avss.t198 avss.t96 465.37
R5003 avss.t166 avss.t144 465.37
R5004 avss.t71 avss.t166 465.37
R5005 avss.t77 avss.t248 465.37
R5006 avss.t229 avss.t77 465.37
R5007 avss.t174 avss.t177 465.37
R5008 avss.t99 avss.t174 465.37
R5009 avss.t97 avss.t245 465.37
R5010 avss.t171 avss.t97 465.37
R5011 avss.t208 avss.t269 465.37
R5012 avss.t80 avss.t208 465.37
R5013 avss.t90 avss.t247 465.37
R5014 avss.t160 avss.t90 465.37
R5015 avss.t42 avss.t204 465.37
R5016 avss.t94 avss.t42 465.37
R5017 avss.t75 avss.t22 465.37
R5018 avss.t270 avss.t75 465.37
R5019 avss.t163 avss.t225 465.37
R5020 avss.t85 avss.t163 465.37
R5021 avss.t251 avss.t61 465.37
R5022 avss.t61 avss.t121 465.37
R5023 avss.t238 avss.t19 465.37
R5024 avss.t19 avss.t63 465.37
R5025 avss.t246 avss.t197 465.37
R5026 avss.t145 avss.t246 465.37
R5027 avss.t249 avss.t173 465.37
R5028 avss.t175 avss.t249 465.37
R5029 avss.t244 avss.t152 465.37
R5030 avss.t267 avss.t244 465.37
R5031 avss.t243 avss.t41 465.37
R5032 avss.t206 avss.t243 465.37
R5033 avss.t5 avss.t164 465.37
R5034 avss.t257 avss.t5 465.37
R5035 avss.t21 avss.t18 465.37
R5036 avss.t239 avss.t21 465.37
R5037 avss.n832 avss.n5 361.01
R5038 avss.n765 avss.n81 361.01
R5039 avss.n683 avss.n139 360.803
R5040 avss.n583 avss.n182 360.803
R5041 avss.n483 avss.n225 360.803
R5042 avss.n383 avss.n268 360.803
R5043 avss.n80 avss.t105 348.214
R5044 avss.n75 avss.t105 348.214
R5045 avss.n7 avss.t182 348.214
R5046 avss.n853 avss.t182 348.214
R5047 avss.n138 avss.t126 348.06
R5048 avss.n133 avss.t126 348.06
R5049 avss.t32 avss.n587 348.06
R5050 avss.n588 avss.t32 348.06
R5051 avss.t108 avss.n487 348.06
R5052 avss.n488 avss.t108 348.06
R5053 avss.t184 avss.n387 348.06
R5054 avss.n388 avss.t184 348.06
R5055 avss.n299 avss.t87 338.849
R5056 avss.t110 avss.n345 338.849
R5057 avss.n407 avss.t98 338.849
R5058 avss.n507 avss.t79 338.849
R5059 avss.n607 avss.t74 338.849
R5060 avss.n700 avss.t68 338.849
R5061 avss.n782 avss.t76 338.849
R5062 avss.n821 avss.t282 314.01
R5063 avss.n33 avss.t282 314.01
R5064 avss.n32 avss.t6 314.01
R5065 avss.n29 avss.t6 314.01
R5066 avss.n28 avss.t288 314.01
R5067 avss.t288 avss.n22 314.01
R5068 avss.n749 avss.t272 314.01
R5069 avss.n107 avss.t272 314.01
R5070 avss.n106 avss.t2 314.01
R5071 avss.n103 avss.t2 314.01
R5072 avss.n102 avss.t25 314.01
R5073 avss.t25 avss.n96 314.01
R5074 avss.n156 avss.t101 313.884
R5075 avss.n658 avss.t101 313.884
R5076 avss.n659 avss.t286 313.884
R5077 avss.n663 avss.t286 313.884
R5078 avss.t188 avss.n666 313.884
R5079 avss.n667 avss.t188 313.884
R5080 avss.n199 avss.t200 313.884
R5081 avss.n558 avss.t200 313.884
R5082 avss.n559 avss.t223 313.884
R5083 avss.n563 avss.t223 313.884
R5084 avss.t132 avss.n566 313.884
R5085 avss.n567 avss.t132 313.884
R5086 avss.n242 avss.t153 313.884
R5087 avss.n458 avss.t153 313.884
R5088 avss.n459 avss.t46 313.884
R5089 avss.n463 avss.t46 313.884
R5090 avss.t23 avss.n466 313.884
R5091 avss.n467 avss.t23 313.884
R5092 avss.n285 avss.t284 313.884
R5093 avss.n358 avss.t284 313.884
R5094 avss.n359 avss.t226 313.884
R5095 avss.n363 avss.t226 313.884
R5096 avss.t114 avss.n366 313.884
R5097 avss.n367 avss.t114 313.884
R5098 avss.n81 avss.n80 300.336
R5099 avss.n7 avss.n5 300.336
R5100 avss.n139 avss.n138 300.202
R5101 avss.n587 avss.n182 300.202
R5102 avss.n487 avss.n225 300.202
R5103 avss.n387 avss.n268 300.202
R5104 avss.n739 avss.t162 279.964
R5105 avss.t193 avss.n98 279.964
R5106 avss.n811 avss.t167 279.964
R5107 avss.t39 avss.n24 279.964
R5108 avss.t210 avss.n347 279.858
R5109 avss.n348 avss.t148 279.858
R5110 avss.t168 avss.n447 279.858
R5111 avss.n448 avss.t157 279.858
R5112 avss.t231 avss.n547 279.858
R5113 avss.n548 avss.t141 279.858
R5114 avss.t279 avss.n647 279.858
R5115 avss.n648 avss.t57 279.858
R5116 avss.t147 avss.t110 271.079
R5117 avss.t98 avss.t159 271.079
R5118 avss.t159 avss.t116 271.079
R5119 avss.t79 avss.t137 271.079
R5120 avss.t137 avss.t190 271.079
R5121 avss.t74 avss.t56 271.079
R5122 avss.t56 avss.t219 271.079
R5123 avss.t68 avss.t192 271.079
R5124 avss.t192 avss.t14 271.079
R5125 avss.t76 avss.t20 271.079
R5126 avss.t20 avss.t277 271.079
R5127 avss.n33 avss.n32 266.909
R5128 avss.n29 avss.n28 266.909
R5129 avss.n107 avss.n106 266.909
R5130 avss.n103 avss.n102 266.909
R5131 avss.n659 avss.n658 266.801
R5132 avss.n666 avss.n663 266.801
R5133 avss.n559 avss.n558 266.801
R5134 avss.n566 avss.n563 266.801
R5135 avss.n459 avss.n458 266.801
R5136 avss.n466 avss.n463 266.801
R5137 avss.n359 avss.n358 266.801
R5138 avss.n366 avss.n363 266.801
R5139 avss.t162 avss.t84 223.97
R5140 avss.t84 avss.t193 223.97
R5141 avss.t167 avss.t78 223.97
R5142 avss.t78 avss.t39 223.97
R5143 avss.t67 avss.t210 223.887
R5144 avss.t148 avss.t67 223.887
R5145 avss.t91 avss.t168 223.887
R5146 avss.t157 avss.t91 223.887
R5147 avss.t73 avss.t231 223.887
R5148 avss.t141 avss.t73 223.887
R5149 avss.t62 avss.t279 223.887
R5150 avss.t57 avss.t62 223.887
R5151 avss.n346 avss.t147 220.988
R5152 avss.n446 avss.n445 213.623
R5153 avss.n546 avss.n545 213.623
R5154 avss.n646 avss.n645 213.623
R5155 avss.n738 avss.n737 213.623
R5156 avss.n810 avss.n809 213.623
R5157 avss.n410 avss.n409 151.869
R5158 avss.n510 avss.n509 151.869
R5159 avss.n610 avss.n609 151.869
R5160 avss.n703 avss.n702 151.869
R5161 avss.n784 avss.n74 151.869
R5162 avss.n326 avss.n325 151.751
R5163 avss.n321 avss.n320 151.751
R5164 avss.n302 avss.n301 151.751
R5165 avss.n426 avss.n425 151.751
R5166 avss.n422 avss.n421 151.751
R5167 avss.n260 avss.n259 151.751
R5168 avss.n526 avss.n525 151.751
R5169 avss.n522 avss.n521 151.751
R5170 avss.n217 avss.n216 151.751
R5171 avss.n626 avss.n625 151.751
R5172 avss.n622 avss.n621 151.751
R5173 avss.n174 avss.n173 151.751
R5174 avss.n718 avss.n52 151.751
R5175 avss.n715 avss.n714 151.751
R5176 avss.n125 avss.n51 151.751
R5177 avss.n790 avss.n789 151.751
R5178 avss.n60 avss.n50 151.751
R5179 avss.n787 avss.n49 151.751
R5180 avss.n335 avss.n283 151.751
R5181 avss.n435 avss.n240 151.751
R5182 avss.n535 avss.n197 151.751
R5183 avss.n635 avss.n154 151.751
R5184 avss.n727 avss.n97 151.751
R5185 avss.n799 avss.n23 151.751
R5186 avss.n375 avss.n374 147.727
R5187 avss.n406 avss.n405 147.727
R5188 avss.n475 avss.n474 147.727
R5189 avss.n506 avss.n505 147.727
R5190 avss.n575 avss.n574 147.727
R5191 avss.n606 avss.n605 147.727
R5192 avss.n675 avss.n674 147.727
R5193 avss.n699 avss.n698 147.727
R5194 avss.n756 avss.n755 147.727
R5195 avss.n781 avss.n780 147.727
R5196 avss.n824 avss.n823 147.727
R5197 avss.n855 avss.n854 147.727
R5198 avss.n446 avss.t116 125.228
R5199 avss.n546 avss.t190 125.228
R5200 avss.n646 avss.t219 125.228
R5201 avss.n738 avss.t14 125.228
R5202 avss.n810 avss.t277 125.228
R5203 avss.n408 avss.n407 88.3958
R5204 avss.n508 avss.n507 88.3958
R5205 avss.n608 avss.n607 88.3958
R5206 avss.n701 avss.n700 88.3958
R5207 avss.n783 avss.n782 88.3958
R5208 avss.n856 avss.n3 87.3061
R5209 avss.n856 avss.n4 87.3061
R5210 avss.n779 avss.n82 87.3061
R5211 avss.n779 avss.n83 87.3061
R5212 avss.n766 avss.n94 87.3061
R5213 avss.n766 avss.n95 87.3061
R5214 avss.n697 avss.n140 87.3061
R5215 avss.n697 avss.n141 87.3061
R5216 avss.n684 avss.n151 87.3061
R5217 avss.n684 avss.n152 87.3061
R5218 avss.n604 avss.n183 87.3061
R5219 avss.n604 avss.n184 87.3061
R5220 avss.n584 avss.n194 87.3061
R5221 avss.n584 avss.n195 87.3061
R5222 avss.n504 avss.n226 87.3061
R5223 avss.n504 avss.n227 87.3061
R5224 avss.n484 avss.n237 87.3061
R5225 avss.n484 avss.n238 87.3061
R5226 avss.n404 avss.n269 87.3061
R5227 avss.n404 avss.n270 87.3061
R5228 avss.n384 avss.n280 87.3061
R5229 avss.n384 avss.n281 87.3061
R5230 avss.n831 avss.n20 87.3061
R5231 avss.n831 avss.n830 87.3061
R5232 avss.n825 avss.n22 78.5029
R5233 avss.n757 avss.n96 78.5029
R5234 avss.n673 avss.n667 78.4713
R5235 avss.n573 avss.n567 78.4713
R5236 avss.n473 avss.n467 78.4713
R5237 avss.n373 avss.n367 78.4713
R5238 avss.n17 avss.n16 67.4727
R5239 avss.n18 avss.n16 67.4727
R5240 avss.n751 avss.n87 67.4727
R5241 avss.n752 avss.n87 67.4727
R5242 avss.n759 avss.n91 67.4727
R5243 avss.n760 avss.n91 67.4727
R5244 avss.n676 avss.n144 67.4727
R5245 avss.n677 avss.n144 67.4727
R5246 avss.n668 avss.n148 67.4727
R5247 avss.n669 avss.n148 67.4727
R5248 avss.n576 avss.n187 67.4727
R5249 avss.n577 avss.n187 67.4727
R5250 avss.n568 avss.n191 67.4727
R5251 avss.n569 avss.n191 67.4727
R5252 avss.n476 avss.n230 67.4727
R5253 avss.n477 avss.n230 67.4727
R5254 avss.n468 avss.n234 67.4727
R5255 avss.n469 avss.n234 67.4727
R5256 avss.n376 avss.n273 67.4727
R5257 avss.n377 avss.n273 67.4727
R5258 avss.n368 avss.n277 67.4727
R5259 avss.n369 avss.n277 67.4727
R5260 avss.n21 avss.n12 67.4727
R5261 avss.n829 avss.n12 67.4727
R5262 avss.n17 avss.n3 66.5005
R5263 avss.n18 avss.n4 66.5005
R5264 avss.n751 avss.n82 66.5005
R5265 avss.n752 avss.n83 66.5005
R5266 avss.n759 avss.n94 66.5005
R5267 avss.n760 avss.n95 66.5005
R5268 avss.n676 avss.n140 66.5005
R5269 avss.n677 avss.n141 66.5005
R5270 avss.n668 avss.n151 66.5005
R5271 avss.n669 avss.n152 66.5005
R5272 avss.n576 avss.n183 66.5005
R5273 avss.n577 avss.n184 66.5005
R5274 avss.n568 avss.n194 66.5005
R5275 avss.n569 avss.n195 66.5005
R5276 avss.n476 avss.n226 66.5005
R5277 avss.n477 avss.n227 66.5005
R5278 avss.n468 avss.n237 66.5005
R5279 avss.n469 avss.n238 66.5005
R5280 avss.n376 avss.n269 66.5005
R5281 avss.n377 avss.n270 66.5005
R5282 avss.n368 avss.n280 66.5005
R5283 avss.n369 avss.n281 66.5005
R5284 avss.n21 avss.n20 66.5005
R5285 avss.n830 avss.n829 66.5005
R5286 avss.n319 avss.n303 61.0571
R5287 avss.n420 avss.n261 61.0571
R5288 avss.n520 avss.n218 61.0571
R5289 avss.n620 avss.n175 61.0571
R5290 avss.n713 avss.n126 61.0571
R5291 avss.n62 avss.n61 61.0571
R5292 avss.n800 avss.n797 61.0561
R5293 avss.n808 avss.n43 61.0561
R5294 avss.n813 avss.n812 61.0561
R5295 avss.n728 avss.n725 61.0561
R5296 avss.n736 avss.n117 61.0561
R5297 avss.n741 avss.n740 61.0561
R5298 avss.n636 avss.n633 61.0561
R5299 avss.n644 avss.n165 61.0561
R5300 avss.n649 avss.n162 61.0561
R5301 avss.n536 avss.n533 61.0561
R5302 avss.n544 avss.n208 61.0561
R5303 avss.n549 avss.n205 61.0561
R5304 avss.n436 avss.n433 61.0561
R5305 avss.n444 avss.n251 61.0561
R5306 avss.n449 avss.n248 61.0561
R5307 avss.n336 avss.n333 61.0561
R5308 avss.n344 avss.n292 61.0561
R5309 avss.n349 avss.n290 61.0561
R5310 avss.n327 avss.n297 61.0561
R5311 avss.n311 avss.n310 61.0561
R5312 avss.n427 avss.n256 61.0561
R5313 avss.n412 avss.n411 61.0561
R5314 avss.n527 avss.n213 61.0561
R5315 avss.n512 avss.n511 61.0561
R5316 avss.n627 avss.n170 61.0561
R5317 avss.n612 avss.n611 61.0561
R5318 avss.n719 avss.n122 61.0561
R5319 avss.n705 avss.n704 61.0561
R5320 avss.n791 avss.n48 61.0561
R5321 avss.n73 avss.n57 61.0561
R5322 avss.n346 avss.t87 50.0912
R5323 avss.n31 avss.n30 44.1404
R5324 avss.n27 avss.n13 44.1404
R5325 avss.n79 avss.n76 44.1404
R5326 avss.n105 avss.n104 44.1404
R5327 avss.n101 avss.n90 44.1404
R5328 avss.n137 avss.n134 44.1404
R5329 avss.n662 avss.n660 44.1404
R5330 avss.n665 avss.n147 44.1404
R5331 avss.n589 avss.n586 44.1404
R5332 avss.n562 avss.n560 44.1404
R5333 avss.n565 avss.n190 44.1404
R5334 avss.n489 avss.n486 44.1404
R5335 avss.n462 avss.n460 44.1404
R5336 avss.n465 avss.n233 44.1404
R5337 avss.n389 avss.n386 44.1404
R5338 avss.n852 avss.n8 44.1404
R5339 avss.n365 avss.n276 44.1394
R5340 avss.n362 avss.n360 44.1394
R5341 avss.n357 avss.n286 44.1394
R5342 avss.n820 avss.n34 44.1394
R5343 avss.n748 avss.n108 44.1394
R5344 avss.n657 avss.n157 44.1394
R5345 avss.n557 avss.n200 44.1394
R5346 avss.n457 avss.n243 44.1394
R5347 avss.n1 avss.t290 34.1066
R5348 avss.n835 avss.n3 20.8061
R5349 avss.n835 avss.n4 20.8061
R5350 avss.n838 avss.n17 20.8061
R5351 avss.n838 avss.n18 20.8061
R5352 avss.n84 avss.n82 20.8061
R5353 avss.n84 avss.n83 20.8061
R5354 avss.n753 avss.n751 20.8061
R5355 avss.n753 avss.n752 20.8061
R5356 avss.n763 avss.n94 20.8061
R5357 avss.n763 avss.n95 20.8061
R5358 avss.n761 avss.n759 20.8061
R5359 avss.n761 avss.n760 20.8061
R5360 avss.n680 avss.n140 20.8061
R5361 avss.n680 avss.n141 20.8061
R5362 avss.n678 avss.n676 20.8061
R5363 avss.n678 avss.n677 20.8061
R5364 avss.n153 avss.n151 20.8061
R5365 avss.n153 avss.n152 20.8061
R5366 avss.n670 avss.n668 20.8061
R5367 avss.n670 avss.n669 20.8061
R5368 avss.n580 avss.n183 20.8061
R5369 avss.n580 avss.n184 20.8061
R5370 avss.n578 avss.n576 20.8061
R5371 avss.n578 avss.n577 20.8061
R5372 avss.n196 avss.n194 20.8061
R5373 avss.n196 avss.n195 20.8061
R5374 avss.n570 avss.n568 20.8061
R5375 avss.n570 avss.n569 20.8061
R5376 avss.n480 avss.n226 20.8061
R5377 avss.n480 avss.n227 20.8061
R5378 avss.n478 avss.n476 20.8061
R5379 avss.n478 avss.n477 20.8061
R5380 avss.n239 avss.n237 20.8061
R5381 avss.n239 avss.n238 20.8061
R5382 avss.n470 avss.n468 20.8061
R5383 avss.n470 avss.n469 20.8061
R5384 avss.n380 avss.n269 20.8061
R5385 avss.n380 avss.n270 20.8061
R5386 avss.n378 avss.n376 20.8061
R5387 avss.n378 avss.n377 20.8061
R5388 avss.n282 avss.n280 20.8061
R5389 avss.n282 avss.n281 20.8061
R5390 avss.n370 avss.n368 20.8061
R5391 avss.n370 avss.n369 20.8061
R5392 avss.n828 avss.n21 20.8061
R5393 avss.n829 avss.n828 20.8061
R5394 avss.n20 avss.n19 20.8061
R5395 avss.n830 avss.n19 20.8061
R5396 avss.n0 avss.t214 19.673
R5397 avss.n0 avss.t211 19.4007
R5398 avss.n859 avss.n858 14.6135
R5399 avss.n289 avss.n287 9.0005
R5400 avss.n340 avss.n339 9.0005
R5401 avss.n318 avss.n317 9.0005
R5402 avss.n305 avss.n294 9.0005
R5403 avss.n308 avss.n307 9.0005
R5404 avss.n314 avss.n313 9.0005
R5405 avss.n296 avss.n295 9.0005
R5406 avss.n330 avss.n329 9.0005
R5407 avss.n338 avss.n288 9.0005
R5408 avss.n352 avss.n351 9.0005
R5409 avss.n247 avss.n245 9.0005
R5410 avss.n440 avss.n439 9.0005
R5411 avss.n419 avss.n418 9.0005
R5412 avss.n263 avss.n253 9.0005
R5413 avss.n266 avss.n265 9.0005
R5414 avss.n415 avss.n414 9.0005
R5415 avss.n255 avss.n254 9.0005
R5416 avss.n430 avss.n429 9.0005
R5417 avss.n438 avss.n246 9.0005
R5418 avss.n452 avss.n451 9.0005
R5419 avss.n204 avss.n202 9.0005
R5420 avss.n540 avss.n539 9.0005
R5421 avss.n519 avss.n518 9.0005
R5422 avss.n220 avss.n210 9.0005
R5423 avss.n223 avss.n222 9.0005
R5424 avss.n515 avss.n514 9.0005
R5425 avss.n212 avss.n211 9.0005
R5426 avss.n530 avss.n529 9.0005
R5427 avss.n538 avss.n203 9.0005
R5428 avss.n552 avss.n551 9.0005
R5429 avss.n161 avss.n159 9.0005
R5430 avss.n640 avss.n639 9.0005
R5431 avss.n619 avss.n618 9.0005
R5432 avss.n177 avss.n167 9.0005
R5433 avss.n180 avss.n179 9.0005
R5434 avss.n615 avss.n614 9.0005
R5435 avss.n169 avss.n168 9.0005
R5436 avss.n630 avss.n629 9.0005
R5437 avss.n638 avss.n160 9.0005
R5438 avss.n652 avss.n651 9.0005
R5439 avss.n114 avss.n112 9.0005
R5440 avss.n732 avss.n731 9.0005
R5441 avss.n712 avss.n711 9.0005
R5442 avss.n128 avss.n119 9.0005
R5443 avss.n131 avss.n130 9.0005
R5444 avss.n708 avss.n707 9.0005
R5445 avss.n121 avss.n120 9.0005
R5446 avss.n722 avss.n721 9.0005
R5447 avss.n730 avss.n113 9.0005
R5448 avss.n744 avss.n743 9.0005
R5449 avss.n40 avss.n38 9.0005
R5450 avss.n804 avss.n803 9.0005
R5451 avss.n66 avss.n65 9.0005
R5452 avss.n64 avss.n45 9.0005
R5453 avss.n72 avss.n58 9.0005
R5454 avss.n71 avss.n69 9.0005
R5455 avss.n47 avss.n46 9.0005
R5456 avss.n794 avss.n793 9.0005
R5457 avss.n802 avss.n39 9.0005
R5458 avss.n816 avss.n815 9.0005
R5459 avss.n342 avss.n292 6.9012
R5460 avss.n442 avss.n251 6.9012
R5461 avss.n542 avss.n208 6.9012
R5462 avss.n642 avss.n165 6.9012
R5463 avss.n734 avss.n117 6.9012
R5464 avss.n806 avss.n43 6.9012
R5465 avss.n339 avss.n333 6.46296
R5466 avss.n297 avss.n296 6.46296
R5467 avss.n310 avss.n308 6.46296
R5468 avss.n439 avss.n433 6.46296
R5469 avss.n256 avss.n255 6.46296
R5470 avss.n411 avss.n266 6.46296
R5471 avss.n539 avss.n533 6.46296
R5472 avss.n213 avss.n212 6.46296
R5473 avss.n511 avss.n223 6.46296
R5474 avss.n639 avss.n633 6.46296
R5475 avss.n170 avss.n169 6.46296
R5476 avss.n611 avss.n180 6.46296
R5477 avss.n731 avss.n725 6.46296
R5478 avss.n122 avss.n121 6.46296
R5479 avss.n704 avss.n131 6.46296
R5480 avss.n803 avss.n797 6.46296
R5481 avss.n48 avss.n47 6.46296
R5482 avss.n73 avss.n72 6.46296
R5483 avss.n290 avss.n289 6.4618
R5484 avss.n319 avss.n318 6.4618
R5485 avss.n248 avss.n247 6.4618
R5486 avss.n420 avss.n419 6.4618
R5487 avss.n205 avss.n204 6.4618
R5488 avss.n520 avss.n519 6.4618
R5489 avss.n162 avss.n161 6.4618
R5490 avss.n620 avss.n619 6.4618
R5491 avss.n740 avss.n114 6.4618
R5492 avss.n713 avss.n712 6.4618
R5493 avss.n812 avss.n40 6.4618
R5494 avss.n65 avss.n61 6.4618
R5495 avss.n343 avss.n342 5.47239
R5496 avss.n443 avss.n442 5.47239
R5497 avss.n543 avss.n542 5.47239
R5498 avss.n643 avss.n642 5.47239
R5499 avss.n735 avss.n734 5.47239
R5500 avss.n807 avss.n806 5.47239
R5501 avss.n859 avss.n1 5.18044
R5502 avss.n351 avss.n350 5.03414
R5503 avss.n338 avss.n337 5.03414
R5504 avss.n329 avss.n328 5.03414
R5505 avss.n313 avss.n312 5.03414
R5506 avss.n305 avss.n304 5.03414
R5507 avss.n451 avss.n450 5.03414
R5508 avss.n438 avss.n437 5.03414
R5509 avss.n429 avss.n428 5.03414
R5510 avss.n414 avss.n413 5.03414
R5511 avss.n263 avss.n262 5.03414
R5512 avss.n551 avss.n550 5.03414
R5513 avss.n538 avss.n537 5.03414
R5514 avss.n529 avss.n528 5.03414
R5515 avss.n514 avss.n513 5.03414
R5516 avss.n220 avss.n219 5.03414
R5517 avss.n651 avss.n650 5.03414
R5518 avss.n638 avss.n637 5.03414
R5519 avss.n629 avss.n628 5.03414
R5520 avss.n614 avss.n613 5.03414
R5521 avss.n177 avss.n176 5.03414
R5522 avss.n743 avss.n742 5.03414
R5523 avss.n730 avss.n729 5.03414
R5524 avss.n721 avss.n720 5.03414
R5525 avss.n707 avss.n706 5.03414
R5526 avss.n128 avss.n127 5.03414
R5527 avss.n815 avss.n814 5.03414
R5528 avss.n802 avss.n801 5.03414
R5529 avss.n793 avss.n792 5.03414
R5530 avss.n71 avss.n70 5.03414
R5531 avss.n64 avss.n63 5.03414
R5532 avss.n26 avss.t289 4.84702
R5533 avss.n25 avss.t7 4.84702
R5534 avss.n100 avss.t26 4.84702
R5535 avss.n99 avss.t3 4.84702
R5536 avss.n664 avss.t189 4.84702
R5537 avss.n661 avss.t287 4.84702
R5538 avss.n564 avss.t133 4.84702
R5539 avss.n561 avss.t224 4.84702
R5540 avss.n464 avss.t24 4.84702
R5541 avss.n461 avss.t47 4.84702
R5542 avss.n364 avss.t115 4.84702
R5543 avss.n361 avss.t227 4.84702
R5544 avss.n272 avss.t254 4.7885
R5545 avss.n271 avss.t180 4.7885
R5546 avss.n403 avss.t119 4.7885
R5547 avss.n350 avss.t149 4.7885
R5548 avss.n337 avss.t146 4.7885
R5549 avss.n343 avss.t111 4.7885
R5550 avss.n328 avss.t199 4.7885
R5551 avss.n312 avss.t66 4.7885
R5552 avss.n304 avss.t72 4.7885
R5553 avss.n229 avss.t260 4.7885
R5554 avss.n228 avss.t156 4.7885
R5555 avss.n503 avss.t196 4.7885
R5556 avss.n450 avss.t158 4.7885
R5557 avss.n437 avss.t176 4.7885
R5558 avss.n443 avss.t117 4.7885
R5559 avss.n428 avss.t230 4.7885
R5560 avss.n413 avss.t89 4.7885
R5561 avss.n262 avss.t100 4.7885
R5562 avss.n186 avss.t131 4.7885
R5563 avss.n185 avss.t45 4.7885
R5564 avss.n603 avss.t222 4.7885
R5565 avss.n550 avss.t142 4.7885
R5566 avss.n537 avss.t268 4.7885
R5567 avss.n543 avss.t191 4.7885
R5568 avss.n528 avss.t172 4.7885
R5569 avss.n513 avss.t70 4.7885
R5570 avss.n219 avss.t81 4.7885
R5571 avss.n143 avss.t113 4.7885
R5572 avss.n142 avss.t17 4.7885
R5573 avss.n696 avss.t1 4.7885
R5574 avss.n650 avss.t58 4.7885
R5575 avss.n637 avss.t207 4.7885
R5576 avss.n643 avss.t220 4.7885
R5577 avss.n628 avss.t161 4.7885
R5578 avss.n613 avss.t93 4.7885
R5579 avss.n176 avss.t95 4.7885
R5580 avss.n86 avss.t203 4.7885
R5581 avss.n85 avss.t276 4.7885
R5582 avss.n778 avss.t262 4.7885
R5583 avss.n742 avss.t194 4.7885
R5584 avss.n729 avss.t258 4.7885
R5585 avss.n735 avss.t15 4.7885
R5586 avss.n720 avss.t271 4.7885
R5587 avss.n706 avss.t83 4.7885
R5588 avss.n127 avss.t86 4.7885
R5589 avss.n814 avss.t40 4.7885
R5590 avss.n801 avss.t240 4.7885
R5591 avss.n807 avss.t278 4.7885
R5592 avss.n792 avss.t122 4.7885
R5593 avss.n70 avss.t60 4.7885
R5594 avss.n63 avss.t64 4.7885
R5595 avss.n839 avss.t281 4.7885
R5596 avss.n834 avss.t216 4.7885
R5597 avss.n857 avss.t213 4.7885
R5598 avss.n10 avss.t36 4.7885
R5599 avss.n11 avss.t135 4.7885
R5600 avss.n9 avss.t38 4.7885
R5601 avss.n36 avss.t283 4.7885
R5602 avss.n77 avss.t106 4.7885
R5603 avss.n92 avss.t140 4.7885
R5604 avss.n93 avss.t235 4.7885
R5605 avss.n767 avss.t233 4.7885
R5606 avss.n110 avss.t273 4.7885
R5607 avss.n135 avss.t127 4.7885
R5608 avss.n149 avss.t151 4.7885
R5609 avss.n150 avss.t51 4.7885
R5610 avss.n685 avss.t53 4.7885
R5611 avss.n656 avss.t102 4.7885
R5612 avss.n590 avss.t33 4.7885
R5613 avss.n192 avss.t237 4.7885
R5614 avss.n193 avss.t11 4.7885
R5615 avss.n585 avss.t13 4.7885
R5616 avss.n556 avss.t201 4.7885
R5617 avss.n490 avss.t109 4.7885
R5618 avss.n235 avss.t170 4.7885
R5619 avss.n236 avss.t28 4.7885
R5620 avss.n485 avss.t30 4.7885
R5621 avss.n456 avss.t154 4.7885
R5622 avss.n390 avss.t185 4.7885
R5623 avss.n278 avss.t218 4.7885
R5624 avss.n279 avss.t266 4.7885
R5625 avss.n385 avss.t264 4.7885
R5626 avss.n356 avss.t285 4.7885
R5627 avss.n851 avss.t183 4.7885
R5628 avss.n342 avss.n341 4.28213
R5629 avss.n442 avss.n441 4.28213
R5630 avss.n542 avss.n541 4.28213
R5631 avss.n642 avss.n641 4.28213
R5632 avss.n734 avss.n733 4.28213
R5633 avss.n806 avss.n805 4.28213
R5634 avss.n400 avss.n399 3.51467
R5635 avss.n500 avss.n499 3.51467
R5636 avss.n600 avss.n599 3.51467
R5637 avss.n693 avss.n692 3.51467
R5638 avss.n775 avss.n774 3.51467
R5639 avss.n842 avss.n841 3.51467
R5640 avss.n400 avss.n273 2.06002
R5641 avss.n500 avss.n230 2.06002
R5642 avss.n600 avss.n187 2.06002
R5643 avss.n693 avss.n144 2.06002
R5644 avss.n775 avss.n87 2.06002
R5645 avss.n841 avss.n16 2.06002
R5646 avss.n354 avss.n286 1.92616
R5647 avss.n845 avss.n12 1.90702
R5648 avss.n820 avss.n819 1.90702
R5649 avss.n31 avss.n15 1.90702
R5650 avss.n844 avss.n13 1.90702
R5651 avss.n79 avss.n78 1.90702
R5652 avss.n771 avss.n91 1.90702
R5653 avss.n748 avss.n747 1.90702
R5654 avss.n105 avss.n88 1.90702
R5655 avss.n772 avss.n90 1.90702
R5656 avss.n137 avss.n136 1.90702
R5657 avss.n689 avss.n148 1.90702
R5658 avss.n158 avss.n157 1.90702
R5659 avss.n660 avss.n145 1.90702
R5660 avss.n690 avss.n147 1.90702
R5661 avss.n591 avss.n586 1.90702
R5662 avss.n596 avss.n191 1.90702
R5663 avss.n201 avss.n200 1.90702
R5664 avss.n560 avss.n188 1.90702
R5665 avss.n597 avss.n190 1.90702
R5666 avss.n491 avss.n486 1.90702
R5667 avss.n496 avss.n234 1.90702
R5668 avss.n244 avss.n243 1.90702
R5669 avss.n460 avss.n231 1.90702
R5670 avss.n497 avss.n233 1.90702
R5671 avss.n391 avss.n386 1.90702
R5672 avss.n396 avss.n277 1.90702
R5673 avss.n360 avss.n274 1.90702
R5674 avss.n397 avss.n276 1.90702
R5675 avss.n850 avss.n8 1.90702
R5676 2inmux_0.Bit avss.n859 1.54251
R5677 avss.n310 avss.n309 1.3005
R5678 avss.n312 avss.n311 1.3005
R5679 avss.n311 avss.n298 1.3005
R5680 avss.n324 avss.n297 1.3005
R5681 avss.n328 avss.n327 1.3005
R5682 avss.n327 avss.n326 1.3005
R5683 avss.n304 avss.n303 1.3005
R5684 avss.n303 avss.n302 1.3005
R5685 avss.n320 avss.n319 1.3005
R5686 avss.n411 avss.n410 1.3005
R5687 avss.n413 avss.n412 1.3005
R5688 avss.n412 avss.n257 1.3005
R5689 avss.n424 avss.n256 1.3005
R5690 avss.n428 avss.n427 1.3005
R5691 avss.n427 avss.n426 1.3005
R5692 avss.n262 avss.n261 1.3005
R5693 avss.n261 avss.n260 1.3005
R5694 avss.n421 avss.n420 1.3005
R5695 avss.n511 avss.n510 1.3005
R5696 avss.n513 avss.n512 1.3005
R5697 avss.n512 avss.n214 1.3005
R5698 avss.n524 avss.n213 1.3005
R5699 avss.n528 avss.n527 1.3005
R5700 avss.n527 avss.n526 1.3005
R5701 avss.n219 avss.n218 1.3005
R5702 avss.n218 avss.n217 1.3005
R5703 avss.n521 avss.n520 1.3005
R5704 avss.n611 avss.n610 1.3005
R5705 avss.n613 avss.n612 1.3005
R5706 avss.n612 avss.n171 1.3005
R5707 avss.n624 avss.n170 1.3005
R5708 avss.n628 avss.n627 1.3005
R5709 avss.n627 avss.n626 1.3005
R5710 avss.n176 avss.n175 1.3005
R5711 avss.n175 avss.n174 1.3005
R5712 avss.n621 avss.n620 1.3005
R5713 avss.n704 avss.n703 1.3005
R5714 avss.n706 avss.n705 1.3005
R5715 avss.n705 avss.n123 1.3005
R5716 avss.n717 avss.n122 1.3005
R5717 avss.n720 avss.n719 1.3005
R5718 avss.n719 avss.n718 1.3005
R5719 avss.n127 avss.n126 1.3005
R5720 avss.n126 avss.n125 1.3005
R5721 avss.n714 avss.n713 1.3005
R5722 avss.n74 avss.n73 1.3005
R5723 avss.n70 avss.n57 1.3005
R5724 avss.n57 avss.n56 1.3005
R5725 avss.n54 avss.n48 1.3005
R5726 avss.n792 avss.n791 1.3005
R5727 avss.n791 avss.n790 1.3005
R5728 avss.n63 avss.n62 1.3005
R5729 avss.n62 avss.n49 1.3005
R5730 avss.n61 avss.n60 1.3005
R5731 avss.n828 avss.n11 1.3005
R5732 avss.n828 avss.n827 1.3005
R5733 avss.n826 avss.n12 1.3005
R5734 avss.n19 avss.n10 1.3005
R5735 avss.n833 avss.n19 1.3005
R5736 avss.n831 avss.n9 1.3005
R5737 avss.n832 avss.n831 1.3005
R5738 avss.n821 avss.n820 1.3005
R5739 avss.n36 avss.n34 1.3005
R5740 avss.n34 avss.n33 1.3005
R5741 avss.n32 avss.n31 1.3005
R5742 avss.n30 avss.n25 1.3005
R5743 avss.n30 avss.n29 1.3005
R5744 avss.n27 avss.n26 1.3005
R5745 avss.n28 avss.n27 1.3005
R5746 avss.n22 avss.n13 1.3005
R5747 avss.n77 avss.n76 1.3005
R5748 avss.n76 avss.n75 1.3005
R5749 avss.n80 avss.n79 1.3005
R5750 avss.n749 avss.n748 1.3005
R5751 avss.n110 avss.n108 1.3005
R5752 avss.n108 avss.n107 1.3005
R5753 avss.n106 avss.n105 1.3005
R5754 avss.n104 avss.n99 1.3005
R5755 avss.n104 avss.n103 1.3005
R5756 avss.n101 avss.n100 1.3005
R5757 avss.n102 avss.n101 1.3005
R5758 avss.n96 avss.n90 1.3005
R5759 avss.n135 avss.n134 1.3005
R5760 avss.n134 avss.n133 1.3005
R5761 avss.n138 avss.n137 1.3005
R5762 avss.n157 avss.n156 1.3005
R5763 avss.n657 avss.n656 1.3005
R5764 avss.n658 avss.n657 1.3005
R5765 avss.n660 avss.n659 1.3005
R5766 avss.n662 avss.n661 1.3005
R5767 avss.n663 avss.n662 1.3005
R5768 avss.n665 avss.n664 1.3005
R5769 avss.n666 avss.n665 1.3005
R5770 avss.n667 avss.n147 1.3005
R5771 avss.n590 avss.n589 1.3005
R5772 avss.n589 avss.n588 1.3005
R5773 avss.n587 avss.n586 1.3005
R5774 avss.n200 avss.n199 1.3005
R5775 avss.n557 avss.n556 1.3005
R5776 avss.n558 avss.n557 1.3005
R5777 avss.n560 avss.n559 1.3005
R5778 avss.n562 avss.n561 1.3005
R5779 avss.n563 avss.n562 1.3005
R5780 avss.n565 avss.n564 1.3005
R5781 avss.n566 avss.n565 1.3005
R5782 avss.n567 avss.n190 1.3005
R5783 avss.n490 avss.n489 1.3005
R5784 avss.n489 avss.n488 1.3005
R5785 avss.n487 avss.n486 1.3005
R5786 avss.n243 avss.n242 1.3005
R5787 avss.n457 avss.n456 1.3005
R5788 avss.n458 avss.n457 1.3005
R5789 avss.n460 avss.n459 1.3005
R5790 avss.n462 avss.n461 1.3005
R5791 avss.n463 avss.n462 1.3005
R5792 avss.n465 avss.n464 1.3005
R5793 avss.n466 avss.n465 1.3005
R5794 avss.n467 avss.n233 1.3005
R5795 avss.n390 avss.n389 1.3005
R5796 avss.n389 avss.n388 1.3005
R5797 avss.n387 avss.n386 1.3005
R5798 avss.n286 avss.n285 1.3005
R5799 avss.n357 avss.n356 1.3005
R5800 avss.n358 avss.n357 1.3005
R5801 avss.n360 avss.n359 1.3005
R5802 avss.n362 avss.n361 1.3005
R5803 avss.n363 avss.n362 1.3005
R5804 avss.n365 avss.n364 1.3005
R5805 avss.n366 avss.n365 1.3005
R5806 avss.n367 avss.n276 1.3005
R5807 avss.n347 avss.n290 1.3005
R5808 avss.n350 avss.n349 1.3005
R5809 avss.n349 avss.n348 1.3005
R5810 avss.n299 avss.n292 1.3005
R5811 avss.n344 avss.n343 1.3005
R5812 avss.n345 avss.n344 1.3005
R5813 avss.n334 avss.n333 1.3005
R5814 avss.n337 avss.n336 1.3005
R5815 avss.n336 avss.n335 1.3005
R5816 avss.n372 avss.n277 1.3005
R5817 avss.n370 avss.n278 1.3005
R5818 avss.n371 avss.n370 1.3005
R5819 avss.n282 avss.n279 1.3005
R5820 avss.n382 avss.n282 1.3005
R5821 avss.n385 avss.n384 1.3005
R5822 avss.n384 avss.n383 1.3005
R5823 avss.n375 avss.n273 1.3005
R5824 avss.n378 avss.n272 1.3005
R5825 avss.n379 avss.n378 1.3005
R5826 avss.n380 avss.n271 1.3005
R5827 avss.n381 avss.n380 1.3005
R5828 avss.n404 avss.n403 1.3005
R5829 avss.n405 avss.n404 1.3005
R5830 avss.n447 avss.n248 1.3005
R5831 avss.n450 avss.n449 1.3005
R5832 avss.n449 avss.n448 1.3005
R5833 avss.n407 avss.n251 1.3005
R5834 avss.n444 avss.n443 1.3005
R5835 avss.n445 avss.n444 1.3005
R5836 avss.n434 avss.n433 1.3005
R5837 avss.n437 avss.n436 1.3005
R5838 avss.n436 avss.n435 1.3005
R5839 avss.n472 avss.n234 1.3005
R5840 avss.n470 avss.n235 1.3005
R5841 avss.n471 avss.n470 1.3005
R5842 avss.n239 avss.n236 1.3005
R5843 avss.n482 avss.n239 1.3005
R5844 avss.n485 avss.n484 1.3005
R5845 avss.n484 avss.n483 1.3005
R5846 avss.n475 avss.n230 1.3005
R5847 avss.n478 avss.n229 1.3005
R5848 avss.n479 avss.n478 1.3005
R5849 avss.n480 avss.n228 1.3005
R5850 avss.n481 avss.n480 1.3005
R5851 avss.n504 avss.n503 1.3005
R5852 avss.n505 avss.n504 1.3005
R5853 avss.n547 avss.n205 1.3005
R5854 avss.n550 avss.n549 1.3005
R5855 avss.n549 avss.n548 1.3005
R5856 avss.n507 avss.n208 1.3005
R5857 avss.n544 avss.n543 1.3005
R5858 avss.n545 avss.n544 1.3005
R5859 avss.n534 avss.n533 1.3005
R5860 avss.n537 avss.n536 1.3005
R5861 avss.n536 avss.n535 1.3005
R5862 avss.n572 avss.n191 1.3005
R5863 avss.n570 avss.n192 1.3005
R5864 avss.n571 avss.n570 1.3005
R5865 avss.n196 avss.n193 1.3005
R5866 avss.n582 avss.n196 1.3005
R5867 avss.n585 avss.n584 1.3005
R5868 avss.n584 avss.n583 1.3005
R5869 avss.n575 avss.n187 1.3005
R5870 avss.n578 avss.n186 1.3005
R5871 avss.n579 avss.n578 1.3005
R5872 avss.n580 avss.n185 1.3005
R5873 avss.n581 avss.n580 1.3005
R5874 avss.n604 avss.n603 1.3005
R5875 avss.n605 avss.n604 1.3005
R5876 avss.n647 avss.n162 1.3005
R5877 avss.n650 avss.n649 1.3005
R5878 avss.n649 avss.n648 1.3005
R5879 avss.n607 avss.n165 1.3005
R5880 avss.n644 avss.n643 1.3005
R5881 avss.n645 avss.n644 1.3005
R5882 avss.n634 avss.n633 1.3005
R5883 avss.n637 avss.n636 1.3005
R5884 avss.n636 avss.n635 1.3005
R5885 avss.n672 avss.n148 1.3005
R5886 avss.n670 avss.n149 1.3005
R5887 avss.n671 avss.n670 1.3005
R5888 avss.n153 avss.n150 1.3005
R5889 avss.n682 avss.n153 1.3005
R5890 avss.n685 avss.n684 1.3005
R5891 avss.n684 avss.n683 1.3005
R5892 avss.n675 avss.n144 1.3005
R5893 avss.n678 avss.n143 1.3005
R5894 avss.n679 avss.n678 1.3005
R5895 avss.n680 avss.n142 1.3005
R5896 avss.n681 avss.n680 1.3005
R5897 avss.n697 avss.n696 1.3005
R5898 avss.n698 avss.n697 1.3005
R5899 avss.n740 avss.n739 1.3005
R5900 avss.n742 avss.n741 1.3005
R5901 avss.n741 avss.n98 1.3005
R5902 avss.n700 avss.n117 1.3005
R5903 avss.n736 avss.n735 1.3005
R5904 avss.n737 avss.n736 1.3005
R5905 avss.n726 avss.n725 1.3005
R5906 avss.n729 avss.n728 1.3005
R5907 avss.n728 avss.n727 1.3005
R5908 avss.n758 avss.n91 1.3005
R5909 avss.n761 avss.n92 1.3005
R5910 avss.n762 avss.n761 1.3005
R5911 avss.n763 avss.n93 1.3005
R5912 avss.n764 avss.n763 1.3005
R5913 avss.n767 avss.n766 1.3005
R5914 avss.n766 avss.n765 1.3005
R5915 avss.n755 avss.n87 1.3005
R5916 avss.n753 avss.n86 1.3005
R5917 avss.n754 avss.n753 1.3005
R5918 avss.n85 avss.n84 1.3005
R5919 avss.n84 avss.n53 1.3005
R5920 avss.n779 avss.n778 1.3005
R5921 avss.n780 avss.n779 1.3005
R5922 avss.n812 avss.n811 1.3005
R5923 avss.n814 avss.n813 1.3005
R5924 avss.n813 avss.n24 1.3005
R5925 avss.n782 avss.n43 1.3005
R5926 avss.n808 avss.n807 1.3005
R5927 avss.n809 avss.n808 1.3005
R5928 avss.n798 avss.n797 1.3005
R5929 avss.n801 avss.n800 1.3005
R5930 avss.n800 avss.n799 1.3005
R5931 avss.n823 avss.n16 1.3005
R5932 avss.n839 avss.n838 1.3005
R5933 avss.n838 avss.n837 1.3005
R5934 avss.n835 avss.n834 1.3005
R5935 avss.n836 avss.n835 1.3005
R5936 avss.n857 avss.n856 1.3005
R5937 avss.n856 avss.n855 1.3005
R5938 avss.n852 avss.n851 1.3005
R5939 avss.n853 avss.n852 1.3005
R5940 avss.n8 avss.n7 1.3005
R5941 avss.n819 avss.n35 0.990409
R5942 avss.n747 avss.n109 0.990409
R5943 avss.n592 avss.n158 0.990409
R5944 avss.n492 avss.n201 0.990409
R5945 avss.n392 avss.n244 0.990409
R5946 avss.n351 avss.n289 0.92075
R5947 avss.n339 avss.n338 0.92075
R5948 avss.n329 avss.n296 0.92075
R5949 avss.n313 avss.n308 0.92075
R5950 avss.n318 avss.n305 0.92075
R5951 avss.n451 avss.n247 0.92075
R5952 avss.n439 avss.n438 0.92075
R5953 avss.n429 avss.n255 0.92075
R5954 avss.n414 avss.n266 0.92075
R5955 avss.n419 avss.n263 0.92075
R5956 avss.n551 avss.n204 0.92075
R5957 avss.n539 avss.n538 0.92075
R5958 avss.n529 avss.n212 0.92075
R5959 avss.n514 avss.n223 0.92075
R5960 avss.n519 avss.n220 0.92075
R5961 avss.n651 avss.n161 0.92075
R5962 avss.n639 avss.n638 0.92075
R5963 avss.n629 avss.n169 0.92075
R5964 avss.n614 avss.n180 0.92075
R5965 avss.n619 avss.n177 0.92075
R5966 avss.n743 avss.n114 0.92075
R5967 avss.n731 avss.n730 0.92075
R5968 avss.n721 avss.n121 0.92075
R5969 avss.n707 avss.n131 0.92075
R5970 avss.n712 avss.n128 0.92075
R5971 avss.n815 avss.n40 0.92075
R5972 avss.n803 avss.n802 0.92075
R5973 avss.n793 avss.n47 0.92075
R5974 avss.n72 avss.n71 0.92075
R5975 avss.n65 avss.n64 0.92075
R5976 avss.n403 avss.n402 0.771017
R5977 avss.n503 avss.n502 0.771017
R5978 avss.n603 avss.n602 0.771017
R5979 avss.n696 avss.n695 0.771017
R5980 avss.n778 avss.n777 0.771017
R5981 avss.n354 avss.n353 0.709028
R5982 avss.n454 avss.n453 0.709028
R5983 avss.n554 avss.n553 0.709028
R5984 avss.n654 avss.n653 0.709028
R5985 avss.n746 avss.n745 0.709028
R5986 avss.n818 avss.n817 0.709028
R5987 avss.n858 avss.n857 0.471317
R5988 avss.n401 avss.n272 0.463217
R5989 avss.n402 avss.n271 0.463217
R5990 avss.n501 avss.n229 0.463217
R5991 avss.n502 avss.n228 0.463217
R5992 avss.n601 avss.n186 0.463217
R5993 avss.n602 avss.n185 0.463217
R5994 avss.n694 avss.n143 0.463217
R5995 avss.n695 avss.n142 0.463217
R5996 avss.n776 avss.n86 0.463217
R5997 avss.n777 avss.n85 0.463217
R5998 avss.n840 avss.n839 0.463217
R5999 avss.n834 avss.n2 0.463217
R6000 avss.n847 avss.n10 0.463217
R6001 avss.n846 avss.n11 0.463217
R6002 avss.n848 avss.n9 0.463217
R6003 avss.n37 avss.n36 0.463217
R6004 avss.n78 avss.n77 0.463217
R6005 avss.n770 avss.n92 0.463217
R6006 avss.n769 avss.n93 0.463217
R6007 avss.n768 avss.n767 0.463217
R6008 avss.n111 avss.n110 0.463217
R6009 avss.n136 avss.n135 0.463217
R6010 avss.n688 avss.n149 0.463217
R6011 avss.n687 avss.n150 0.463217
R6012 avss.n686 avss.n685 0.463217
R6013 avss.n656 avss.n655 0.463217
R6014 avss.n591 avss.n590 0.463217
R6015 avss.n595 avss.n192 0.463217
R6016 avss.n594 avss.n193 0.463217
R6017 avss.n593 avss.n585 0.463217
R6018 avss.n556 avss.n555 0.463217
R6019 avss.n491 avss.n490 0.463217
R6020 avss.n495 avss.n235 0.463217
R6021 avss.n494 avss.n236 0.463217
R6022 avss.n493 avss.n485 0.463217
R6023 avss.n456 avss.n455 0.463217
R6024 avss.n391 avss.n390 0.463217
R6025 avss.n395 avss.n278 0.463217
R6026 avss.n394 avss.n279 0.463217
R6027 avss.n393 avss.n385 0.463217
R6028 avss.n356 avss.n355 0.463217
R6029 avss.n851 avss.n850 0.463217
R6030 avss.n402 avss.n401 0.3083
R6031 avss.n502 avss.n501 0.3083
R6032 avss.n602 avss.n601 0.3083
R6033 avss.n695 avss.n694 0.3083
R6034 avss.n777 avss.n776 0.3083
R6035 avss.n840 avss.n2 0.3083
R6036 avss.n847 avss.n846 0.3083
R6037 avss.n848 avss.n847 0.3083
R6038 avss.n770 avss.n769 0.3083
R6039 avss.n769 avss.n768 0.3083
R6040 avss.n688 avss.n687 0.3083
R6041 avss.n687 avss.n686 0.3083
R6042 avss.n595 avss.n594 0.3083
R6043 avss.n594 avss.n593 0.3083
R6044 avss.n495 avss.n494 0.3083
R6045 avss.n494 avss.n493 0.3083
R6046 avss.n395 avss.n394 0.3083
R6047 avss.n394 avss.n393 0.3083
R6048 avss.n858 avss.n2 0.3002
R6049 avss.n1 avss.n0 0.252687
R6050 avss.n846 avss.n845 0.2165
R6051 avss.n771 avss.n770 0.2165
R6052 avss.n689 avss.n688 0.2165
R6053 avss.n596 avss.n595 0.2165
R6054 avss.n496 avss.n495 0.2165
R6055 avss.n396 avss.n395 0.2165
R6056 avss.n768 avss.n35 0.1748
R6057 avss.n593 avss.n592 0.1748
R6058 avss.n493 avss.n492 0.1748
R6059 avss.n393 avss.n392 0.1748
R6060 avss.n686 avss.n109 0.17465
R6061 avss.n849 avss.n848 0.1598
R6062 avss.n850 avss.n849 0.152487
R6063 avss.n845 avss.n844 0.148459
R6064 avss.n772 avss.n771 0.148459
R6065 avss.n690 avss.n689 0.148459
R6066 avss.n597 avss.n596 0.148459
R6067 avss.n497 avss.n496 0.148459
R6068 avss.n397 avss.n396 0.148459
R6069 avss.n136 avss.n109 0.13865
R6070 avss.n78 avss.n35 0.1385
R6071 avss.n592 avss.n591 0.1385
R6072 avss.n492 avss.n491 0.1385
R6073 avss.n392 avss.n391 0.1385
R6074 avss.n316 avss.n306 0.122607
R6075 avss.n417 avss.n264 0.122607
R6076 avss.n517 avss.n221 0.122607
R6077 avss.n617 avss.n178 0.122607
R6078 avss.n710 avss.n129 0.122607
R6079 avss.n67 avss.n59 0.122607
R6080 avss.n332 avss.n331 0.10457
R6081 avss.n432 avss.n431 0.10457
R6082 avss.n532 avss.n531 0.10457
R6083 avss.n632 avss.n631 0.10457
R6084 avss.n724 avss.n723 0.10457
R6085 avss.n796 avss.n795 0.10457
R6086 avss.n843 avss.n14 0.073981
R6087 avss.n773 avss.n89 0.073981
R6088 avss.n691 avss.n146 0.073981
R6089 avss.n598 avss.n189 0.073981
R6090 avss.n498 avss.n232 0.073981
R6091 avss.n398 avss.n275 0.073981
R6092 avss.n340 avss.n287 0.0679983
R6093 avss.n440 avss.n245 0.0679983
R6094 avss.n540 avss.n202 0.0679983
R6095 avss.n640 avss.n159 0.0679983
R6096 avss.n732 avss.n112 0.0679983
R6097 avss.n804 avss.n38 0.0679983
R6098 avss.n401 avss.n400 0.0635
R6099 avss.n501 avss.n500 0.0635
R6100 avss.n601 avss.n600 0.0635
R6101 avss.n694 avss.n693 0.0635
R6102 avss.n776 avss.n775 0.0635
R6103 avss.n841 avss.n840 0.0635
R6104 avss.n306 avss.n293 0.0622481
R6105 avss.n264 avss.n252 0.0622481
R6106 avss.n221 avss.n209 0.0622481
R6107 avss.n178 avss.n166 0.0622481
R6108 avss.n129 avss.n118 0.0622481
R6109 avss.n59 avss.n44 0.0622481
R6110 avss.n352 avss.n288 0.0568904
R6111 avss.n452 avss.n246 0.0568904
R6112 avss.n552 avss.n203 0.0568904
R6113 avss.n652 avss.n160 0.0568904
R6114 avss.n744 avss.n113 0.0568904
R6115 avss.n816 avss.n39 0.0568904
R6116 avss.n332 avss.n288 0.054837
R6117 avss.n432 avss.n246 0.054837
R6118 avss.n532 avss.n203 0.054837
R6119 avss.n632 avss.n160 0.054837
R6120 avss.n724 avss.n113 0.054837
R6121 avss.n796 avss.n39 0.054837
R6122 avss.n331 avss.n294 0.0466843
R6123 avss.n431 avss.n253 0.0466843
R6124 avss.n531 avss.n210 0.0466843
R6125 avss.n631 avss.n167 0.0466843
R6126 avss.n723 avss.n119 0.0466843
R6127 avss.n795 avss.n45 0.0466843
R6128 avss.n332 avss.n293 0.0415307
R6129 avss.n432 avss.n252 0.0415307
R6130 avss.n532 avss.n209 0.0415307
R6131 avss.n632 avss.n166 0.0415307
R6132 avss.n724 avss.n118 0.0415307
R6133 avss.n796 avss.n44 0.0415307
R6134 avss.n317 avss.n294 0.0405109
R6135 avss.n314 avss.n307 0.0405109
R6136 avss.n330 avss.n295 0.0405109
R6137 avss.n418 avss.n253 0.0405109
R6138 avss.n415 avss.n265 0.0405109
R6139 avss.n430 avss.n254 0.0405109
R6140 avss.n518 avss.n210 0.0405109
R6141 avss.n515 avss.n222 0.0405109
R6142 avss.n530 avss.n211 0.0405109
R6143 avss.n618 avss.n167 0.0405109
R6144 avss.n615 avss.n179 0.0405109
R6145 avss.n630 avss.n168 0.0405109
R6146 avss.n711 avss.n119 0.0405109
R6147 avss.n708 avss.n130 0.0405109
R6148 avss.n722 avss.n120 0.0405109
R6149 avss.n66 avss.n45 0.0405109
R6150 avss.n69 avss.n58 0.0405109
R6151 avss.n794 avss.n46 0.0405109
R6152 avss.n844 avss.n843 0.0389018
R6153 avss.n773 avss.n772 0.0389018
R6154 avss.n691 avss.n690 0.0389018
R6155 avss.n598 avss.n597 0.0389018
R6156 avss.n498 avss.n497 0.0389018
R6157 avss.n398 avss.n397 0.0389018
R6158 avss.n353 avss.n287 0.035635
R6159 avss.n453 avss.n245 0.035635
R6160 avss.n553 avss.n202 0.035635
R6161 avss.n653 avss.n159 0.035635
R6162 avss.n745 avss.n112 0.035635
R6163 avss.n817 avss.n38 0.035635
R6164 avss.n341 avss.n332 0.0349747
R6165 avss.n441 avss.n432 0.0349747
R6166 avss.n541 avss.n532 0.0349747
R6167 avss.n641 avss.n632 0.0349747
R6168 avss.n733 avss.n724 0.0349747
R6169 avss.n805 avss.n796 0.0349747
R6170 avss.n316 avss.n315 0.0322085
R6171 avss.n315 avss.n293 0.0322085
R6172 avss.n417 avss.n416 0.0322085
R6173 avss.n416 avss.n252 0.0322085
R6174 avss.n517 avss.n516 0.0322085
R6175 avss.n516 avss.n209 0.0322085
R6176 avss.n617 avss.n616 0.0322085
R6177 avss.n616 avss.n166 0.0322085
R6178 avss.n710 avss.n709 0.0322085
R6179 avss.n709 avss.n118 0.0322085
R6180 avss.n68 avss.n67 0.0322085
R6181 avss.n68 avss.n44 0.0322085
R6182 avss.n25 avss.n14 0.0258591
R6183 avss.n26 avss.n14 0.0258591
R6184 avss.n99 avss.n89 0.0258591
R6185 avss.n100 avss.n89 0.0258591
R6186 avss.n661 avss.n146 0.0258591
R6187 avss.n664 avss.n146 0.0258591
R6188 avss.n561 avss.n189 0.0258591
R6189 avss.n564 avss.n189 0.0258591
R6190 avss.n461 avss.n232 0.0258591
R6191 avss.n464 avss.n232 0.0258591
R6192 avss.n361 avss.n275 0.0258591
R6193 avss.n364 avss.n275 0.0258591
R6194 avss.n843 avss.n842 0.023066
R6195 avss.n774 avss.n773 0.023066
R6196 avss.n692 avss.n691 0.023066
R6197 avss.n599 avss.n598 0.023066
R6198 avss.n499 avss.n498 0.023066
R6199 avss.n399 avss.n398 0.023066
R6200 avss.n317 avss.n316 0.0214837
R6201 avss.n315 avss.n295 0.0214837
R6202 avss.n418 avss.n417 0.0214837
R6203 avss.n416 avss.n254 0.0214837
R6204 avss.n518 avss.n517 0.0214837
R6205 avss.n516 avss.n211 0.0214837
R6206 avss.n618 avss.n617 0.0214837
R6207 avss.n616 avss.n168 0.0214837
R6208 avss.n711 avss.n710 0.0214837
R6209 avss.n709 avss.n120 0.0214837
R6210 avss.n67 avss.n66 0.0214837
R6211 avss.n68 avss.n46 0.0214837
R6212 avss.n819 avss.n818 0.0196349
R6213 avss.n747 avss.n746 0.0196349
R6214 avss.n654 avss.n158 0.0196349
R6215 avss.n554 avss.n201 0.0196349
R6216 avss.n454 avss.n244 0.0196349
R6217 avss.n842 avss.n15 0.0163358
R6218 avss.n774 avss.n88 0.0163358
R6219 avss.n692 avss.n145 0.0163358
R6220 avss.n599 avss.n188 0.0163358
R6221 avss.n499 avss.n231 0.0163358
R6222 avss.n399 avss.n274 0.0163358
R6223 avss.n37 avss.n15 0.0139604
R6224 avss.n111 avss.n88 0.0139604
R6225 avss.n655 avss.n145 0.0139604
R6226 avss.n555 avss.n188 0.0139604
R6227 avss.n455 avss.n231 0.0139604
R6228 avss.n355 avss.n274 0.0139604
R6229 avss.n818 avss.n37 0.0130367
R6230 avss.n746 avss.n111 0.0130367
R6231 avss.n655 avss.n654 0.0130367
R6232 avss.n555 avss.n554 0.0130367
R6233 avss.n455 avss.n454 0.0130367
R6234 avss.n355 avss.n354 0.0130367
R6235 avss.n315 avss.n314 0.0121902
R6236 avss.n416 avss.n415 0.0121902
R6237 avss.n516 avss.n515 0.0121902
R6238 avss.n616 avss.n615 0.0121902
R6239 avss.n709 avss.n708 0.0121902
R6240 avss.n69 avss.n68 0.0121902
R6241 avss.n849 avss 0.0118245
R6242 avss.n307 avss.n306 0.00915761
R6243 avss.n265 avss.n264 0.00915761
R6244 avss.n222 avss.n221 0.00915761
R6245 avss.n179 avss.n178 0.00915761
R6246 avss.n130 avss.n129 0.00915761
R6247 avss.n59 avss.n58 0.00915761
R6248 avss.n331 avss.n330 0.00720109
R6249 avss.n431 avss.n430 0.00720109
R6250 avss.n531 avss.n530 0.00720109
R6251 avss.n631 avss.n630 0.00720109
R6252 avss.n723 avss.n722 0.00720109
R6253 avss.n795 avss.n794 0.00720109
R6254 avss.n353 avss.n352 0.00511663
R6255 avss.n453 avss.n452 0.00511663
R6256 avss.n553 avss.n552 0.00511663
R6257 avss.n653 avss.n652 0.00511663
R6258 avss.n745 avss.n744 0.00511663
R6259 avss.n817 avss.n816 0.00511663
R6260 avss.n341 avss.n340 0.000544599
R6261 avss.n441 avss.n440 0.000544599
R6262 avss.n541 avss.n540 0.000544599
R6263 avss.n641 avss.n640 0.000544599
R6264 avss.n733 avss.n732 0.000544599
R6265 avss.n805 avss.n804 0.000544599
R6266 a_48650_3501.n0 a_48650_3501.t4 34.1797
R6267 a_48650_3501.n0 a_48650_3501.t5 19.5798
R6268 a_48650_3501.n1 a_48650_3501.t3 18.7717
R6269 a_48650_3501.n1 a_48650_3501.t1 9.2885
R6270 a_48650_3501.n2 a_48650_3501.n0 4.93379
R6271 a_48650_3501.t0 a_48650_3501.n3 4.23346
R6272 a_48650_3501.n3 a_48650_3501.t2 3.85546
R6273 a_48650_3501.n2 a_48650_3501.n1 0.4055
R6274 a_48650_3501.n3 a_48650_3501.n2 0.352625
R6275 a_6520_1558.n0 a_6520_1558.t5 40.8177
R6276 a_6520_1558.n1 a_6520_1558.t4 40.6313
R6277 a_6520_1558.n1 a_6520_1558.t6 27.3166
R6278 a_6520_1558.n0 a_6520_1558.t7 27.1302
R6279 a_6520_1558.n2 a_6520_1558.n1 19.2576
R6280 a_6520_1558.n3 a_6520_1558.t1 10.0473
R6281 a_6520_1558.t0 a_6520_1558.n5 6.51042
R6282 a_6520_1558.n5 a_6520_1558.n4 6.04952
R6283 a_6520_1558.n2 a_6520_1558.n0 5.91752
R6284 a_6520_1558.n3 a_6520_1558.n2 4.89565
R6285 a_6520_1558.n5 a_6520_1558.n3 0.732092
R6286 a_6520_1558.n4 a_6520_1558.t3 0.7285
R6287 a_6520_1558.n4 a_6520_1558.t2 0.7285
R6288 a_6600_2510.n0 a_6600_2510.t4 41.0041
R6289 a_6600_2510.n1 a_6600_2510.t5 40.8177
R6290 a_6600_2510.n1 a_6600_2510.t7 27.1302
R6291 a_6600_2510.n0 a_6600_2510.t6 26.9438
R6292 a_6600_2510.n2 a_6600_2510.n1 22.5284
R6293 a_6600_2510.n3 a_6600_2510.n2 19.5781
R6294 a_6600_2510.n3 a_6600_2510.t1 10.0473
R6295 a_6600_2510.n4 a_6600_2510.t3 6.51042
R6296 a_6600_2510.n5 a_6600_2510.n4 6.04952
R6297 a_6600_2510.n2 a_6600_2510.n0 5.7305
R6298 a_6600_2510.n4 a_6600_2510.n3 0.732092
R6299 a_6600_2510.t0 a_6600_2510.n5 0.7285
R6300 a_6600_2510.n5 a_6600_2510.t2 0.7285
R6301 a_6520_3763.n1 a_6520_3763.t9 41.0041
R6302 a_6520_3763.n0 a_6520_3763.t5 40.8177
R6303 a_6520_3763.n2 a_6520_3763.t4 40.6313
R6304 a_6520_3763.n2 a_6520_3763.t7 27.3166
R6305 a_6520_3763.n0 a_6520_3763.t8 27.1302
R6306 a_6520_3763.n1 a_6520_3763.t6 26.9438
R6307 a_6520_3763.n3 a_6520_3763.n1 15.6312
R6308 a_6520_3763.n3 a_6520_3763.n2 15.046
R6309 a_6520_3763.n5 a_6520_3763.t3 10.0473
R6310 a_6520_3763.n6 a_6520_3763.t2 6.51042
R6311 a_6520_3763.n7 a_6520_3763.n6 6.04952
R6312 a_6520_3763.n4 a_6520_3763.n0 5.64619
R6313 a_6520_3763.n5 a_6520_3763.n4 5.17851
R6314 a_6520_3763.n4 a_6520_3763.n3 4.5005
R6315 a_6520_3763.n6 a_6520_3763.n5 0.732092
R6316 a_6520_3763.t0 a_6520_3763.n7 0.7285
R6317 a_6520_3763.n7 a_6520_3763.t1 0.7285
R6318 dffrs_1.Q.n3 dffrs_1.Q.t7 40.6313
R6319 dffrs_1.Q.n1 dffrs_1.Q.t4 34.1066
R6320 dffrs_1.Q.n3 dffrs_1.Q.t5 27.3166
R6321 dffrs_1.Q.n0 dffrs_1.Q.t6 19.673
R6322 dffrs_1.Q.n0 dffrs_1.Q.t8 19.4007
R6323 dffrs_1.Q.n7 dffrs_1.Q.n3 14.6967
R6324 dffrs_1.Q.n6 dffrs_1.Q.t2 10.0473
R6325 dffrs_1.Q.n7 dffrs_1.Q.n6 9.39565
R6326 dffrs_1.Q.n2 dffrs_1.Q.n1 6.70486
R6327 dffrs_1.Q.n5 dffrs_1.Q.t1 6.51042
R6328 dffrs_1.Q.n5 dffrs_1.Q.n4 6.04952
R6329 dffrs_1.Q dffrs_1.Q.n2 5.81354
R6330 dffrs_1.Q.n6 dffrs_1.Q.n5 0.732092
R6331 dffrs_1.Q.n4 dffrs_1.Q.t3 0.7285
R6332 dffrs_1.Q.n4 dffrs_1.Q.t0 0.7285
R6333 dffrs_1.Q dffrs_1.Q.n7 0.458082
R6334 dffrs_1.Q.n1 dffrs_1.Q.n0 0.252687
R6335 dffrs_1.Q.n2 2inmux_3.Bit 0.0519286
R6336 a_20234_3501.n0 a_20234_3501.t5 34.1797
R6337 a_20234_3501.n0 a_20234_3501.t4 19.5798
R6338 a_20234_3501.n3 a_20234_3501.t2 18.7717
R6339 a_20234_3501.t0 a_20234_3501.n3 9.2885
R6340 a_20234_3501.n2 a_20234_3501.n0 4.93379
R6341 a_20234_3501.n1 a_20234_3501.t1 4.23346
R6342 a_20234_3501.n1 a_20234_3501.t3 3.85546
R6343 a_20234_3501.n3 a_20234_3501.n2 0.4055
R6344 a_20234_3501.n2 a_20234_3501.n1 0.352625
R6345 2inmux_2.Bit.n3 2inmux_2.Bit.t6 40.6313
R6346 2inmux_2.Bit.n1 2inmux_2.Bit.t5 34.1066
R6347 2inmux_2.Bit.n3 2inmux_2.Bit.t8 27.3166
R6348 2inmux_2.Bit.n0 2inmux_2.Bit.t7 19.673
R6349 2inmux_2.Bit.n0 2inmux_2.Bit.t4 19.4007
R6350 2inmux_2.Bit.n7 2inmux_2.Bit.n3 14.6967
R6351 2inmux_2.Bit.n6 2inmux_2.Bit.t0 10.0473
R6352 2inmux_2.Bit.n7 2inmux_2.Bit.n6 9.39565
R6353 2inmux_2.Bit.n2 2inmux_2.Bit.n1 6.70486
R6354 2inmux_2.Bit.n5 2inmux_2.Bit.t1 6.51042
R6355 2inmux_2.Bit.n5 2inmux_2.Bit.n4 6.04952
R6356 dffrs_0.Q 2inmux_2.Bit.n2 5.81514
R6357 2inmux_2.Bit.n6 2inmux_2.Bit.n5 0.732092
R6358 2inmux_2.Bit.n4 2inmux_2.Bit.t2 0.7285
R6359 2inmux_2.Bit.n4 2inmux_2.Bit.t3 0.7285
R6360 dffrs_0.Q 2inmux_2.Bit.n7 0.458082
R6361 2inmux_2.Bit.n1 2inmux_2.Bit.n0 0.252687
R6362 2inmux_2.Bit.n2 2inmux_2.Bit 0.0519286
R6363 a_1290_3500.n0 a_1290_3500.t4 34.1797
R6364 a_1290_3500.n0 a_1290_3500.t5 19.5798
R6365 a_1290_3500.t0 a_1290_3500.n3 18.7717
R6366 a_1290_3500.n3 a_1290_3500.t1 9.2885
R6367 a_1290_3500.n2 a_1290_3500.n0 4.93379
R6368 a_1290_3500.n1 a_1290_3500.t3 4.23346
R6369 a_1290_3500.n1 a_1290_3500.t2 3.85546
R6370 a_1290_3500.n3 a_1290_3500.n2 0.4055
R6371 a_1290_3500.n2 a_1290_3500.n1 0.352625
R6372 clk.n3 clk.t18 41.0041
R6373 clk.n7 clk.t12 41.0041
R6374 clk.n11 clk.t1 41.0041
R6375 clk.n15 clk.t15 41.0041
R6376 clk.n19 clk.t3 41.0041
R6377 clk.n0 clk.t17 41.0041
R6378 clk.n4 clk.t2 40.8177
R6379 clk.n8 clk.t22 40.8177
R6380 clk.n12 clk.t11 40.8177
R6381 clk.n16 clk.t8 40.8177
R6382 clk.n20 clk.t20 40.8177
R6383 clk.n1 clk.t10 40.8177
R6384 clk.n4 clk.t13 27.1302
R6385 clk.n8 clk.t9 27.1302
R6386 clk.n12 clk.t23 27.1302
R6387 clk.n16 clk.t19 27.1302
R6388 clk.n20 clk.t5 27.1302
R6389 clk.n1 clk.t21 27.1302
R6390 clk.n3 clk.t7 26.9438
R6391 clk.n7 clk.t0 26.9438
R6392 clk.n11 clk.t14 26.9438
R6393 clk.n15 clk.t4 26.9438
R6394 clk.n19 clk.t16 26.9438
R6395 clk.n0 clk.t6 26.9438
R6396 dffrs_5.clk clk.n22 23.2034
R6397 clk.n10 clk.n6 13.9468
R6398 clk.n14 clk.n10 13.9463
R6399 clk.n22 clk.n18 13.9457
R6400 clk.n18 clk.n14 13.9457
R6401 clk.n6 dffrs_0.clk 9.25764
R6402 clk.n10 dffrs_1.clk 9.25764
R6403 clk.n14 dffrs_2.clk 9.25764
R6404 clk.n18 dffrs_3.clk 9.25764
R6405 clk.n22 dffrs_4.clk 9.25764
R6406 clk.n5 clk.n4 7.65746
R6407 clk.n9 clk.n8 7.65746
R6408 clk.n13 clk.n12 7.65746
R6409 clk.n17 clk.n16 7.65746
R6410 clk.n21 clk.n20 7.65746
R6411 clk.n2 clk.n1 7.65746
R6412 clk.n5 clk.n3 7.12229
R6413 clk.n9 clk.n7 7.12229
R6414 clk.n13 clk.n11 7.12229
R6415 clk.n17 clk.n15 7.12229
R6416 clk.n21 clk.n19 7.12229
R6417 clk.n2 clk.n0 7.12229
R6418 clk.n6 clk 3.54742
R6419 dffrs_0.clk clk.n5 0.611214
R6420 dffrs_1.clk clk.n9 0.611214
R6421 dffrs_2.clk clk.n13 0.611214
R6422 dffrs_3.clk clk.n17 0.611214
R6423 dffrs_4.clk clk.n21 0.611214
R6424 dffrs_5.clk clk.n2 0.611214
R6425 a_15992_3763.n1 a_15992_3763.t7 41.0041
R6426 a_15992_3763.n0 a_15992_3763.t5 40.8177
R6427 a_15992_3763.n2 a_15992_3763.t6 40.6313
R6428 a_15992_3763.n2 a_15992_3763.t9 27.3166
R6429 a_15992_3763.n0 a_15992_3763.t8 27.1302
R6430 a_15992_3763.n1 a_15992_3763.t4 26.9438
R6431 a_15992_3763.n3 a_15992_3763.n1 15.6312
R6432 a_15992_3763.n3 a_15992_3763.n2 15.046
R6433 a_15992_3763.n5 a_15992_3763.t1 10.0473
R6434 a_15992_3763.t0 a_15992_3763.n7 6.51042
R6435 a_15992_3763.n7 a_15992_3763.n6 6.04952
R6436 a_15992_3763.n4 a_15992_3763.n0 5.64619
R6437 a_15992_3763.n5 a_15992_3763.n4 5.17851
R6438 a_15992_3763.n4 a_15992_3763.n3 4.5005
R6439 a_15992_3763.n7 a_15992_3763.n5 0.732092
R6440 a_15992_3763.n6 a_15992_3763.t2 0.7285
R6441 a_15992_3763.n6 a_15992_3763.t3 0.7285
R6442 2inmux_1.Bit.n3 2inmux_1.Bit.t8 40.6313
R6443 2inmux_1.Bit.n1 2inmux_1.Bit.t7 34.1066
R6444 2inmux_1.Bit.n3 2inmux_1.Bit.t5 27.3166
R6445 2inmux_1.Bit.n0 2inmux_1.Bit.t4 19.673
R6446 2inmux_1.Bit.n0 2inmux_1.Bit.t6 19.4007
R6447 2inmux_1.Bit.n7 2inmux_1.Bit.n3 14.6967
R6448 2inmux_1.Bit.n6 2inmux_1.Bit.t2 10.0473
R6449 2inmux_1.Bit.n7 2inmux_1.Bit.n6 9.39565
R6450 2inmux_1.Bit.n2 2inmux_1.Bit.n1 6.70486
R6451 2inmux_1.Bit.n5 2inmux_1.Bit.t3 6.51042
R6452 2inmux_1.Bit.n5 2inmux_1.Bit.n4 6.04952
R6453 dffrs_4.Q 2inmux_1.Bit.n2 5.81514
R6454 2inmux_1.Bit.n6 2inmux_1.Bit.n5 0.732092
R6455 2inmux_1.Bit.n4 2inmux_1.Bit.t1 0.7285
R6456 2inmux_1.Bit.n4 2inmux_1.Bit.t0 0.7285
R6457 dffrs_4.Q 2inmux_1.Bit.n7 0.458082
R6458 2inmux_1.Bit.n1 2inmux_1.Bit.n0 0.252687
R6459 2inmux_1.Bit.n2 2inmux_1.Bit 0.0519286
R6460 a_15992_5968.n2 a_15992_5968.t5 40.6313
R6461 a_15992_5968.n2 a_15992_5968.t4 27.3166
R6462 a_15992_5968.n3 a_15992_5968.n2 24.1527
R6463 a_15992_5968.t0 a_15992_5968.n3 10.0473
R6464 a_15992_5968.n1 a_15992_5968.t1 6.51042
R6465 a_15992_5968.n1 a_15992_5968.n0 6.04952
R6466 a_15992_5968.n3 a_15992_5968.n1 0.732092
R6467 a_15992_5968.n0 a_15992_5968.t3 0.7285
R6468 a_15992_5968.n0 a_15992_5968.t2 0.7285
R6469 load.n4 load.t17 34.2529
R6470 load.n10 load.t23 34.2529
R6471 load.n16 load.t28 34.2529
R6472 load.n22 load.t13 34.2529
R6473 load.n28 load.t0 34.2529
R6474 load.n1 load.t9 34.2529
R6475 load.n6 load.t20 34.1797
R6476 load.n12 load.t19 34.1797
R6477 load.n18 load.t14 34.1797
R6478 load.n24 load.t1 34.1797
R6479 load.n30 load.t26 34.1797
R6480 load.n2 load.t3 34.1797
R6481 load.n3 load.t2 19.673
R6482 load.n9 load.t5 19.673
R6483 load.n15 load.t4 19.673
R6484 load.n21 load.t18 19.673
R6485 load.n27 load.t7 19.673
R6486 load.n0 load.t25 19.673
R6487 load.n6 load.t12 19.5798
R6488 load.n12 load.t11 19.5798
R6489 load.n18 load.t6 19.5798
R6490 load.n24 load.t22 19.5798
R6491 load.n30 load.t16 19.5798
R6492 load.n2 load.t24 19.5798
R6493 load.n3 load.t15 19.4007
R6494 load.n9 load.t21 19.4007
R6495 load.n15 load.t27 19.4007
R6496 load.n21 load.t10 19.4007
R6497 load.n27 load.t29 19.4007
R6498 load.n0 load.t8 19.4007
R6499 load.n33 load.n32 15.5531
R6500 load.n8 load.n7 8.46371
R6501 load.n20 load.n19 8.37371
R6502 load.n14 load.n13 8.32871
R6503 load.n26 load.n25 8.32871
R6504 load.n32 load.n31 8.32871
R6505 load.n5 load.n4 7.87164
R6506 load.n11 load.n10 7.87164
R6507 load.n17 load.n16 7.87164
R6508 load.n23 load.n22 7.87164
R6509 load.n29 load.n28 7.87164
R6510 load.n34 load.n1 7.87164
R6511 load.n14 load.n8 7.26762
R6512 load.n32 load.n26 7.22491
R6513 load.n26 load.n20 7.22491
R6514 load.n20 load.n14 7.22491
R6515 load.n7 load.n6 5.00771
R6516 load.n19 load.n18 5.00771
R6517 load.n13 load.n12 4.96432
R6518 load.n25 load.n24 4.96432
R6519 load.n31 load.n30 4.96432
R6520 load.n33 load.n2 4.96432
R6521 load.n13 load.n11 2.11068
R6522 load.n25 load.n23 2.11068
R6523 load.n31 load.n29 2.11068
R6524 load.n34 load.n33 2.11068
R6525 load.n7 load.n5 2.06729
R6526 load.n19 load.n17 2.06729
R6527 load.n5 2inmux_0.Load 0.2255
R6528 load.n11 2inmux_2.Load 0.2255
R6529 load.n17 2inmux_3.Load 0.2255
R6530 load.n23 2inmux_4.Load 0.2255
R6531 load.n29 2inmux_5.Load 0.2255
R6532 2inmux_1.Load load.n34 0.2255
R6533 load.n8 load 0.211008
R6534 load.n4 load.n3 0.106438
R6535 load.n10 load.n9 0.106438
R6536 load.n16 load.n15 0.106438
R6537 load.n22 load.n21 0.106438
R6538 load.n28 load.n27 0.106438
R6539 load.n1 load.n0 0.106438
R6540 a_39178_3501.n0 a_39178_3501.t5 34.1797
R6541 a_39178_3501.n0 a_39178_3501.t4 19.5798
R6542 a_39178_3501.n1 a_39178_3501.t3 18.7717
R6543 a_39178_3501.n1 a_39178_3501.t2 9.2885
R6544 a_39178_3501.n2 a_39178_3501.n0 4.93379
R6545 a_39178_3501.t0 a_39178_3501.n3 4.23346
R6546 a_39178_3501.n3 a_39178_3501.t1 3.85546
R6547 a_39178_3501.n2 a_39178_3501.n1 0.4055
R6548 a_39178_3501.n3 a_39178_3501.n2 0.352625
R6549 dffrs_2.Q.n3 dffrs_2.Q.t8 40.6313
R6550 dffrs_2.Q.n1 dffrs_2.Q.t7 34.1066
R6551 dffrs_2.Q.n3 dffrs_2.Q.t5 27.3166
R6552 dffrs_2.Q.n0 dffrs_2.Q.t4 19.673
R6553 dffrs_2.Q.n0 dffrs_2.Q.t6 19.4007
R6554 dffrs_2.Q.n7 dffrs_2.Q.n3 14.6967
R6555 dffrs_2.Q.n6 dffrs_2.Q.t0 10.0473
R6556 dffrs_2.Q.n7 dffrs_2.Q.n6 9.39565
R6557 dffrs_2.Q.n2 dffrs_2.Q.n1 6.70486
R6558 dffrs_2.Q.n5 dffrs_2.Q.t1 6.51042
R6559 dffrs_2.Q.n5 dffrs_2.Q.n4 6.04952
R6560 dffrs_2.Q dffrs_2.Q.n2 5.81514
R6561 dffrs_2.Q.n6 dffrs_2.Q.n5 0.732092
R6562 dffrs_2.Q.n4 dffrs_2.Q.t3 0.7285
R6563 dffrs_2.Q.n4 dffrs_2.Q.t2 0.7285
R6564 dffrs_2.Q dffrs_2.Q.n7 0.458082
R6565 dffrs_2.Q.n1 dffrs_2.Q.n0 0.252687
R6566 dffrs_2.Q.n2 2inmux_4.Bit 0.0519286
R6567 a_48650_1161.n0 a_48650_1161.t5 34.1797
R6568 a_48650_1161.n0 a_48650_1161.t4 19.5798
R6569 a_48650_1161.t0 a_48650_1161.n3 18.7717
R6570 a_48650_1161.n3 a_48650_1161.t2 9.2885
R6571 a_48650_1161.n2 a_48650_1161.n0 4.93379
R6572 a_48650_1161.n1 a_48650_1161.t3 4.23346
R6573 a_48650_1161.n1 a_48650_1161.t1 3.85546
R6574 a_48650_1161.n3 a_48650_1161.n2 0.4055
R6575 a_48650_1161.n2 a_48650_1161.n1 0.352625
R6576 a_50878_1605.n0 a_50878_1605.t5 34.1797
R6577 a_50878_1605.n0 a_50878_1605.t4 19.5798
R6578 a_50878_1605.t0 a_50878_1605.n3 10.3401
R6579 a_50878_1605.n3 a_50878_1605.t3 9.2885
R6580 a_50878_1605.n2 a_50878_1605.n0 4.93379
R6581 a_50878_1605.n1 a_50878_1605.t2 4.09202
R6582 a_50878_1605.n1 a_50878_1605.t1 3.95079
R6583 a_50878_1605.n3 a_50878_1605.n2 0.599711
R6584 a_50878_1605.n2 a_50878_1605.n1 0.296375
R6585 2inmux_1.OUT.n0 2inmux_1.OUT.t2 41.0041
R6586 2inmux_1.OUT.n0 2inmux_1.OUT.t3 26.9438
R6587 2inmux_1.OUT.n1 2inmux_1.OUT.t1 9.6935
R6588 dffrs_5.d 2inmux_1.OUT.n0 6.55979
R6589 2inmux_1.OUT dffrs_5.d 4.883
R6590 2inmux_1.OUT.n1 2inmux_1.OUT.t0 4.35383
R6591 2inmux_1.OUT 2inmux_1.OUT.n1 0.350857
R6592 a_22462_1605.n0 a_22462_1605.t5 34.1797
R6593 a_22462_1605.n0 a_22462_1605.t4 19.5798
R6594 a_22462_1605.t0 a_22462_1605.n3 10.3401
R6595 a_22462_1605.n3 a_22462_1605.t3 9.2885
R6596 a_22462_1605.n2 a_22462_1605.n0 4.93379
R6597 a_22462_1605.n1 a_22462_1605.t1 4.09202
R6598 a_22462_1605.n1 a_22462_1605.t2 3.95079
R6599 a_22462_1605.n3 a_22462_1605.n2 0.599711
R6600 a_22462_1605.n2 a_22462_1605.n1 0.296375
R6601 a_34936_1559.n0 a_34936_1559.t5 40.8177
R6602 a_34936_1559.n1 a_34936_1559.t6 40.6313
R6603 a_34936_1559.n1 a_34936_1559.t4 27.3166
R6604 a_34936_1559.n0 a_34936_1559.t7 27.1302
R6605 a_34936_1559.n2 a_34936_1559.n1 19.2576
R6606 a_34936_1559.n3 a_34936_1559.t2 10.0473
R6607 a_34936_1559.n4 a_34936_1559.t3 6.51042
R6608 a_34936_1559.n5 a_34936_1559.n4 6.04952
R6609 a_34936_1559.n2 a_34936_1559.n0 5.91752
R6610 a_34936_1559.n3 a_34936_1559.n2 4.89565
R6611 a_34936_1559.n4 a_34936_1559.n3 0.732092
R6612 a_34936_1559.t0 a_34936_1559.n5 0.7285
R6613 a_34936_1559.n5 a_34936_1559.t1 0.7285
R6614 a_34936_3764.n1 a_34936_3764.t8 41.0041
R6615 a_34936_3764.n0 a_34936_3764.t6 40.8177
R6616 a_34936_3764.n2 a_34936_3764.t7 40.6313
R6617 a_34936_3764.n2 a_34936_3764.t4 27.3166
R6618 a_34936_3764.n0 a_34936_3764.t9 27.1302
R6619 a_34936_3764.n1 a_34936_3764.t5 26.9438
R6620 a_34936_3764.n3 a_34936_3764.n1 15.6312
R6621 a_34936_3764.n3 a_34936_3764.n2 15.046
R6622 a_34936_3764.n5 a_34936_3764.t1 10.0473
R6623 a_34936_3764.t0 a_34936_3764.n7 6.51042
R6624 a_34936_3764.n7 a_34936_3764.n6 6.04952
R6625 a_34936_3764.n4 a_34936_3764.n0 5.64619
R6626 a_34936_3764.n5 a_34936_3764.n4 5.17851
R6627 a_34936_3764.n4 a_34936_3764.n3 4.5005
R6628 a_34936_3764.n7 a_34936_3764.n5 0.732092
R6629 a_34936_3764.n6 a_34936_3764.t2 0.7285
R6630 a_34936_3764.n6 a_34936_3764.t3 0.7285
R6631 a_3518_1604.n0 a_3518_1604.t5 34.1797
R6632 a_3518_1604.n0 a_3518_1604.t4 19.5798
R6633 a_3518_1604.n3 a_3518_1604.t3 10.3401
R6634 a_3518_1604.t0 a_3518_1604.n3 9.2885
R6635 a_3518_1604.n2 a_3518_1604.n0 4.93379
R6636 a_3518_1604.n1 a_3518_1604.t2 4.09202
R6637 a_3518_1604.n1 a_3518_1604.t1 3.95079
R6638 a_3518_1604.n3 a_3518_1604.n2 0.599711
R6639 a_3518_1604.n2 a_3518_1604.n1 0.296375
R6640 2inmux_0.OUT.n0 2inmux_0.OUT.t2 41.0041
R6641 2inmux_0.OUT.n0 2inmux_0.OUT.t3 26.9438
R6642 2inmux_0.OUT.n1 2inmux_0.OUT.t1 9.6935
R6643 dffrs_0.d 2inmux_0.OUT.n0 6.55979
R6644 2inmux_0.OUT dffrs_0.d 4.883
R6645 2inmux_0.OUT.n1 2inmux_0.OUT.t0 4.35383
R6646 2inmux_0.OUT 2inmux_0.OUT.n1 0.350857
R6647 a_44408_3764.n1 a_44408_3764.t6 41.0041
R6648 a_44408_3764.n0 a_44408_3764.t5 40.8177
R6649 a_44408_3764.n2 a_44408_3764.t4 40.6313
R6650 a_44408_3764.n2 a_44408_3764.t7 27.3166
R6651 a_44408_3764.n0 a_44408_3764.t9 27.1302
R6652 a_44408_3764.n1 a_44408_3764.t8 26.9438
R6653 a_44408_3764.n3 a_44408_3764.n1 15.6312
R6654 a_44408_3764.n3 a_44408_3764.n2 15.046
R6655 a_44408_3764.n5 a_44408_3764.t1 10.0473
R6656 a_44408_3764.t0 a_44408_3764.n7 6.51042
R6657 a_44408_3764.n7 a_44408_3764.n6 6.04952
R6658 a_44408_3764.n4 a_44408_3764.n0 5.64619
R6659 a_44408_3764.n5 a_44408_3764.n4 5.17851
R6660 a_44408_3764.n4 a_44408_3764.n3 4.5005
R6661 a_44408_3764.n7 a_44408_3764.n5 0.732092
R6662 a_44408_3764.n6 a_44408_3764.t2 0.7285
R6663 a_44408_3764.n6 a_44408_3764.t3 0.7285
R6664 a_20234_1161.n0 a_20234_1161.t4 34.1797
R6665 a_20234_1161.n0 a_20234_1161.t5 19.5798
R6666 a_20234_1161.t0 a_20234_1161.n3 18.7717
R6667 a_20234_1161.n3 a_20234_1161.t3 9.2885
R6668 a_20234_1161.n2 a_20234_1161.n0 4.93379
R6669 a_20234_1161.n1 a_20234_1161.t1 4.23346
R6670 a_20234_1161.n1 a_20234_1161.t2 3.85546
R6671 a_20234_1161.n3 a_20234_1161.n2 0.4055
R6672 a_20234_1161.n2 a_20234_1161.n1 0.352625
R6673 a_29706_1161.n0 a_29706_1161.t4 34.1797
R6674 a_29706_1161.n0 a_29706_1161.t5 19.5798
R6675 a_29706_1161.n1 a_29706_1161.t2 18.7717
R6676 a_29706_1161.n1 a_29706_1161.t1 9.2885
R6677 a_29706_1161.n2 a_29706_1161.n0 4.93379
R6678 a_29706_1161.t0 a_29706_1161.n3 4.23346
R6679 a_29706_1161.n3 a_29706_1161.t3 3.85546
R6680 a_29706_1161.n2 a_29706_1161.n1 0.4055
R6681 a_29706_1161.n3 a_29706_1161.n2 0.352625
R6682 a_25464_3764.n1 a_25464_3764.t5 41.0041
R6683 a_25464_3764.n0 a_25464_3764.t4 40.8177
R6684 a_25464_3764.n2 a_25464_3764.t6 40.6313
R6685 a_25464_3764.n2 a_25464_3764.t9 27.3166
R6686 a_25464_3764.n0 a_25464_3764.t8 27.1302
R6687 a_25464_3764.n1 a_25464_3764.t7 26.9438
R6688 a_25464_3764.n3 a_25464_3764.n1 15.6312
R6689 a_25464_3764.n3 a_25464_3764.n2 15.046
R6690 a_25464_3764.n5 a_25464_3764.t1 10.0473
R6691 a_25464_3764.t0 a_25464_3764.n7 6.51042
R6692 a_25464_3764.n7 a_25464_3764.n6 6.04952
R6693 a_25464_3764.n4 a_25464_3764.n0 5.64619
R6694 a_25464_3764.n5 a_25464_3764.n4 5.17851
R6695 a_25464_3764.n4 a_25464_3764.n3 4.5005
R6696 a_25464_3764.n7 a_25464_3764.n5 0.732092
R6697 a_25464_3764.n6 a_25464_3764.t2 0.7285
R6698 a_25464_3764.n6 a_25464_3764.t3 0.7285
R6699 B6.n1 B6.t1 34.2529
R6700 B6.n0 B6.t0 19.673
R6701 B6.n0 B6.t2 19.4007
R6702 B6.n2 B6.n1 8.05164
R6703 B6.n2 B6 1.87121
R6704 B6.n1 B6.n0 0.106438
R6705 2inmux_0.In B6.n2 0.0455
R6706 a_1290_1160.n0 a_1290_1160.t5 34.1797
R6707 a_1290_1160.n0 a_1290_1160.t4 19.5798
R6708 a_1290_1160.n1 a_1290_1160.t3 18.7717
R6709 a_1290_1160.n1 a_1290_1160.t2 9.2885
R6710 a_1290_1160.n2 a_1290_1160.n0 4.93379
R6711 a_1290_1160.t0 a_1290_1160.n3 4.23346
R6712 a_1290_1160.n3 a_1290_1160.t1 3.85546
R6713 a_1290_1160.n2 a_1290_1160.n1 0.4055
R6714 a_1290_1160.n3 a_1290_1160.n2 0.352625
R6715 a_10762_3500.n0 a_10762_3500.t5 34.1797
R6716 a_10762_3500.n0 a_10762_3500.t4 19.5798
R6717 a_10762_3500.n1 a_10762_3500.t2 18.7717
R6718 a_10762_3500.n1 a_10762_3500.t1 9.2885
R6719 a_10762_3500.n2 a_10762_3500.n0 4.93379
R6720 a_10762_3500.n3 a_10762_3500.t3 4.23346
R6721 a_10762_3500.t0 a_10762_3500.n3 3.85546
R6722 a_10762_3500.n2 a_10762_3500.n1 0.4055
R6723 a_10762_3500.n3 a_10762_3500.n2 0.352625
R6724 a_35016_2511.n0 a_35016_2511.t5 41.0041
R6725 a_35016_2511.n1 a_35016_2511.t6 40.8177
R6726 a_35016_2511.n1 a_35016_2511.t4 27.1302
R6727 a_35016_2511.n0 a_35016_2511.t7 26.9438
R6728 a_35016_2511.n2 a_35016_2511.n1 22.5284
R6729 a_35016_2511.n3 a_35016_2511.n2 19.5781
R6730 a_35016_2511.n3 a_35016_2511.t3 10.0473
R6731 a_35016_2511.n4 a_35016_2511.t2 6.51042
R6732 a_35016_2511.n5 a_35016_2511.n4 6.04952
R6733 a_35016_2511.n2 a_35016_2511.n0 5.7305
R6734 a_35016_2511.n4 a_35016_2511.n3 0.732092
R6735 a_35016_2511.n5 a_35016_2511.t1 0.7285
R6736 a_35016_2511.t0 a_35016_2511.n5 0.7285
R6737 a_41406_1605.n0 a_41406_1605.t5 34.1797
R6738 a_41406_1605.n0 a_41406_1605.t4 19.5798
R6739 a_41406_1605.t0 a_41406_1605.n3 10.3401
R6740 a_41406_1605.n3 a_41406_1605.t3 9.2885
R6741 a_41406_1605.n2 a_41406_1605.n0 4.93379
R6742 a_41406_1605.n1 a_41406_1605.t1 4.09202
R6743 a_41406_1605.n1 a_41406_1605.t2 3.95079
R6744 a_41406_1605.n3 a_41406_1605.n2 0.599711
R6745 a_41406_1605.n2 a_41406_1605.n1 0.296375
R6746 a_44488_2511.n0 a_44488_2511.t7 41.0041
R6747 a_44488_2511.n1 a_44488_2511.t4 40.8177
R6748 a_44488_2511.n1 a_44488_2511.t6 27.1302
R6749 a_44488_2511.n0 a_44488_2511.t5 26.9438
R6750 a_44488_2511.n2 a_44488_2511.n1 22.5284
R6751 a_44488_2511.n3 a_44488_2511.n2 19.5781
R6752 a_44488_2511.n3 a_44488_2511.t1 10.0473
R6753 a_44488_2511.n4 a_44488_2511.t2 6.51042
R6754 a_44488_2511.n5 a_44488_2511.n4 6.04952
R6755 a_44488_2511.n2 a_44488_2511.n0 5.7305
R6756 a_44488_2511.n4 a_44488_2511.n3 0.732092
R6757 a_44488_2511.t0 a_44488_2511.n5 0.7285
R6758 a_44488_2511.n5 a_44488_2511.t3 0.7285
R6759 a_44408_5969.n0 a_44408_5969.t4 40.6313
R6760 a_44408_5969.n0 a_44408_5969.t5 27.3166
R6761 a_44408_5969.n1 a_44408_5969.n0 24.1527
R6762 a_44408_5969.n1 a_44408_5969.t1 10.0473
R6763 a_44408_5969.t0 a_44408_5969.n3 6.51042
R6764 a_44408_5969.n3 a_44408_5969.n2 6.04952
R6765 a_44408_5969.n3 a_44408_5969.n1 0.732092
R6766 a_44408_5969.n2 a_44408_5969.t3 0.7285
R6767 a_44408_5969.n2 a_44408_5969.t2 0.7285
R6768 a_25464_1559.n0 a_25464_1559.t4 40.8177
R6769 a_25464_1559.n1 a_25464_1559.t5 40.6313
R6770 a_25464_1559.n1 a_25464_1559.t7 27.3166
R6771 a_25464_1559.n0 a_25464_1559.t6 27.1302
R6772 a_25464_1559.n2 a_25464_1559.n1 19.2576
R6773 a_25464_1559.n3 a_25464_1559.t1 10.0473
R6774 a_25464_1559.n4 a_25464_1559.t2 6.51042
R6775 a_25464_1559.n5 a_25464_1559.n4 6.04952
R6776 a_25464_1559.n2 a_25464_1559.n0 5.91752
R6777 a_25464_1559.n3 a_25464_1559.n2 4.89565
R6778 a_25464_1559.n4 a_25464_1559.n3 0.732092
R6779 a_25464_1559.t0 a_25464_1559.n5 0.7285
R6780 a_25464_1559.n5 a_25464_1559.t3 0.7285
R6781 a_29706_3501.n0 a_29706_3501.t5 34.1797
R6782 a_29706_3501.n0 a_29706_3501.t4 19.5798
R6783 a_29706_3501.n1 a_29706_3501.t1 18.7717
R6784 a_29706_3501.n1 a_29706_3501.t2 9.2885
R6785 a_29706_3501.n2 a_29706_3501.n0 4.93379
R6786 a_29706_3501.t0 a_29706_3501.n3 4.23346
R6787 a_29706_3501.n3 a_29706_3501.t3 3.85546
R6788 a_29706_3501.n2 a_29706_3501.n1 0.4055
R6789 a_29706_3501.n3 a_29706_3501.n2 0.352625
R6790 dffrs_3.Q.n3 dffrs_3.Q.t6 40.6313
R6791 dffrs_3.Q.n1 dffrs_3.Q.t5 34.1066
R6792 dffrs_3.Q.n3 dffrs_3.Q.t7 27.3166
R6793 dffrs_3.Q.n0 dffrs_3.Q.t8 19.673
R6794 dffrs_3.Q.n0 dffrs_3.Q.t4 19.4007
R6795 dffrs_3.Q.n7 dffrs_3.Q.n3 14.6967
R6796 dffrs_3.Q.n6 dffrs_3.Q.t1 10.0473
R6797 dffrs_3.Q.n7 dffrs_3.Q.n6 9.39565
R6798 dffrs_3.Q.n2 dffrs_3.Q.n1 6.70486
R6799 dffrs_3.Q.n5 dffrs_3.Q.t2 6.51042
R6800 dffrs_3.Q.n5 dffrs_3.Q.n4 6.04952
R6801 dffrs_3.Q dffrs_3.Q.n2 5.81514
R6802 dffrs_3.Q.n6 dffrs_3.Q.n5 0.732092
R6803 dffrs_3.Q.n4 dffrs_3.Q.t0 0.7285
R6804 dffrs_3.Q.n4 dffrs_3.Q.t3 0.7285
R6805 dffrs_3.Q dffrs_3.Q.n7 0.458082
R6806 dffrs_3.Q.n1 dffrs_3.Q.n0 0.252687
R6807 dffrs_3.Q.n2 2inmux_5.Bit 0.0519286
R6808 2inmux_3.OUT.n0 2inmux_3.OUT.t3 41.0041
R6809 2inmux_3.OUT.n0 2inmux_3.OUT.t2 26.9438
R6810 2inmux_3.OUT.n1 2inmux_3.OUT.t1 9.6935
R6811 dffrs_2.d 2inmux_3.OUT.n0 6.55979
R6812 2inmux_3.OUT dffrs_2.d 4.883
R6813 2inmux_3.OUT.n1 2inmux_3.OUT.t0 4.35383
R6814 2inmux_3.OUT 2inmux_3.OUT.n1 0.350857
R6815 a_12990_1604.n0 a_12990_1604.t5 34.1797
R6816 a_12990_1604.n0 a_12990_1604.t4 19.5798
R6817 a_12990_1604.n3 a_12990_1604.t3 10.3401
R6818 a_12990_1604.t0 a_12990_1604.n3 9.2885
R6819 a_12990_1604.n2 a_12990_1604.n0 4.93379
R6820 a_12990_1604.n1 a_12990_1604.t1 4.09202
R6821 a_12990_1604.n1 a_12990_1604.t2 3.95079
R6822 a_12990_1604.n3 a_12990_1604.n2 0.599711
R6823 a_12990_1604.n2 a_12990_1604.n1 0.296375
R6824 a_25464_5969.n0 a_25464_5969.t5 40.6313
R6825 a_25464_5969.n0 a_25464_5969.t4 27.3166
R6826 a_25464_5969.n1 a_25464_5969.n0 24.1527
R6827 a_25464_5969.n1 a_25464_5969.t2 10.0473
R6828 a_25464_5969.n2 a_25464_5969.t3 6.51042
R6829 a_25464_5969.n3 a_25464_5969.n2 6.04952
R6830 a_25464_5969.n2 a_25464_5969.n1 0.732092
R6831 a_25464_5969.n3 a_25464_5969.t1 0.7285
R6832 a_25464_5969.t0 a_25464_5969.n3 0.7285
R6833 a_44408_1559.n0 a_44408_1559.t5 40.8177
R6834 a_44408_1559.n1 a_44408_1559.t4 40.6313
R6835 a_44408_1559.n1 a_44408_1559.t6 27.3166
R6836 a_44408_1559.n0 a_44408_1559.t7 27.1302
R6837 a_44408_1559.n2 a_44408_1559.n1 19.2576
R6838 a_44408_1559.n3 a_44408_1559.t2 10.0473
R6839 a_44408_1559.n4 a_44408_1559.t3 6.51042
R6840 a_44408_1559.n5 a_44408_1559.n4 6.04952
R6841 a_44408_1559.n2 a_44408_1559.n0 5.91752
R6842 a_44408_1559.n3 a_44408_1559.n2 4.89565
R6843 a_44408_1559.n4 a_44408_1559.n3 0.732092
R6844 a_44408_1559.n5 a_44408_1559.t1 0.7285
R6845 a_44408_1559.t0 a_44408_1559.n5 0.7285
R6846 a_53880_1559.n0 a_53880_1559.t6 40.8177
R6847 a_53880_1559.n1 a_53880_1559.t7 40.6313
R6848 a_53880_1559.n1 a_53880_1559.t5 27.3166
R6849 a_53880_1559.n0 a_53880_1559.t4 27.1302
R6850 a_53880_1559.n2 a_53880_1559.n1 19.2576
R6851 a_53880_1559.n3 a_53880_1559.t3 10.0473
R6852 a_53880_1559.n4 a_53880_1559.t2 6.51042
R6853 a_53880_1559.n5 a_53880_1559.n4 6.04952
R6854 a_53880_1559.n2 a_53880_1559.n0 5.91752
R6855 a_53880_1559.n3 a_53880_1559.n2 4.89565
R6856 a_53880_1559.n4 a_53880_1559.n3 0.732092
R6857 a_53880_1559.t0 a_53880_1559.n5 0.7285
R6858 a_53880_1559.n5 a_53880_1559.t1 0.7285
R6859 a_53960_2511.n0 a_53960_2511.t5 41.0041
R6860 a_53960_2511.n1 a_53960_2511.t6 40.8177
R6861 a_53960_2511.n1 a_53960_2511.t4 27.1302
R6862 a_53960_2511.n0 a_53960_2511.t7 26.9438
R6863 a_53960_2511.n2 a_53960_2511.n1 22.5284
R6864 a_53960_2511.n3 a_53960_2511.n2 19.5781
R6865 a_53960_2511.n3 a_53960_2511.t2 10.0473
R6866 a_53960_2511.n4 a_53960_2511.t3 6.51042
R6867 a_53960_2511.n5 a_53960_2511.n4 6.04952
R6868 a_53960_2511.n2 a_53960_2511.n0 5.7305
R6869 a_53960_2511.n4 a_53960_2511.n3 0.732092
R6870 a_53960_2511.n5 a_53960_2511.t1 0.7285
R6871 a_53960_2511.t0 a_53960_2511.n5 0.7285
R6872 a_53880_3764.n3 a_53880_3764.t8 41.0041
R6873 a_53880_3764.n2 a_53880_3764.t7 40.8177
R6874 a_53880_3764.n4 a_53880_3764.t9 40.6313
R6875 a_53880_3764.n4 a_53880_3764.t6 27.3166
R6876 a_53880_3764.n2 a_53880_3764.t4 27.1302
R6877 a_53880_3764.n3 a_53880_3764.t5 26.9438
R6878 a_53880_3764.n5 a_53880_3764.n3 15.6312
R6879 a_53880_3764.n5 a_53880_3764.n4 15.046
R6880 a_53880_3764.t0 a_53880_3764.n7 10.0473
R6881 a_53880_3764.n1 a_53880_3764.t1 6.51042
R6882 a_53880_3764.n1 a_53880_3764.n0 6.04952
R6883 a_53880_3764.n6 a_53880_3764.n2 5.64619
R6884 a_53880_3764.n7 a_53880_3764.n6 5.17851
R6885 a_53880_3764.n6 a_53880_3764.n5 4.5005
R6886 a_53880_3764.n7 a_53880_3764.n1 0.732092
R6887 a_53880_3764.n0 a_53880_3764.t2 0.7285
R6888 a_53880_3764.n0 a_53880_3764.t3 0.7285
R6889 2inmux_2.OUT.n0 2inmux_2.OUT.t2 41.0041
R6890 2inmux_2.OUT.n0 2inmux_2.OUT.t3 26.9438
R6891 2inmux_2.OUT.n1 2inmux_2.OUT.t1 9.6935
R6892 dffrs_1.d 2inmux_2.OUT.n0 6.55979
R6893 2inmux_2.OUT dffrs_1.d 4.883
R6894 2inmux_2.OUT.n1 2inmux_2.OUT.t0 4.35383
R6895 2inmux_2.OUT 2inmux_2.OUT.n1 0.350857
R6896 a_16072_2510.n2 a_16072_2510.t4 41.0041
R6897 a_16072_2510.n3 a_16072_2510.t5 40.8177
R6898 a_16072_2510.n3 a_16072_2510.t7 27.1302
R6899 a_16072_2510.n2 a_16072_2510.t6 26.9438
R6900 a_16072_2510.n4 a_16072_2510.n3 22.5284
R6901 a_16072_2510.n5 a_16072_2510.n4 19.5781
R6902 a_16072_2510.t0 a_16072_2510.n5 10.0473
R6903 a_16072_2510.n1 a_16072_2510.t1 6.51042
R6904 a_16072_2510.n1 a_16072_2510.n0 6.04952
R6905 a_16072_2510.n4 a_16072_2510.n2 5.7305
R6906 a_16072_2510.n5 a_16072_2510.n1 0.732092
R6907 a_16072_2510.n0 a_16072_2510.t2 0.7285
R6908 a_16072_2510.n0 a_16072_2510.t3 0.7285
R6909 a_34936_5969.n0 a_34936_5969.t5 40.6313
R6910 a_34936_5969.n0 a_34936_5969.t4 27.3166
R6911 a_34936_5969.n1 a_34936_5969.n0 24.1527
R6912 a_34936_5969.n1 a_34936_5969.t2 10.0473
R6913 a_34936_5969.n2 a_34936_5969.t1 6.51042
R6914 a_34936_5969.n3 a_34936_5969.n2 6.04952
R6915 a_34936_5969.n2 a_34936_5969.n1 0.732092
R6916 a_34936_5969.t0 a_34936_5969.n3 0.7285
R6917 a_34936_5969.n3 a_34936_5969.t3 0.7285
R6918 a_15992_1558.n2 a_15992_1558.t4 40.8177
R6919 a_15992_1558.n3 a_15992_1558.t5 40.6313
R6920 a_15992_1558.n3 a_15992_1558.t7 27.3166
R6921 a_15992_1558.n2 a_15992_1558.t6 27.1302
R6922 a_15992_1558.n4 a_15992_1558.n3 19.2576
R6923 a_15992_1558.t0 a_15992_1558.n5 10.0473
R6924 a_15992_1558.n1 a_15992_1558.t1 6.51042
R6925 a_15992_1558.n1 a_15992_1558.n0 6.04952
R6926 a_15992_1558.n4 a_15992_1558.n2 5.91752
R6927 a_15992_1558.n5 a_15992_1558.n4 4.89565
R6928 a_15992_1558.n5 a_15992_1558.n1 0.732092
R6929 a_15992_1558.n0 a_15992_1558.t2 0.7285
R6930 a_15992_1558.n0 a_15992_1558.t3 0.7285
R6931 a_53880_5969.n0 a_53880_5969.t4 40.6313
R6932 a_53880_5969.n0 a_53880_5969.t5 27.3166
R6933 a_53880_5969.n1 a_53880_5969.n0 24.1527
R6934 a_53880_5969.n1 a_53880_5969.t2 10.0473
R6935 a_53880_5969.n2 a_53880_5969.t3 6.51042
R6936 a_53880_5969.n3 a_53880_5969.n2 6.04952
R6937 a_53880_5969.n2 a_53880_5969.n1 0.732092
R6938 a_53880_5969.n3 a_53880_5969.t1 0.7285
R6939 a_53880_5969.t0 a_53880_5969.n3 0.7285
R6940 a_31934_1605.n0 a_31934_1605.t5 34.1797
R6941 a_31934_1605.n0 a_31934_1605.t4 19.5798
R6942 a_31934_1605.t0 a_31934_1605.n3 10.3401
R6943 a_31934_1605.n3 a_31934_1605.t3 9.2885
R6944 a_31934_1605.n2 a_31934_1605.n0 4.93379
R6945 a_31934_1605.n1 a_31934_1605.t1 4.09202
R6946 a_31934_1605.n1 a_31934_1605.t2 3.95079
R6947 a_31934_1605.n3 a_31934_1605.n2 0.599711
R6948 a_31934_1605.n2 a_31934_1605.n1 0.296375
R6949 2inmux_4.OUT.n0 2inmux_4.OUT.t2 41.0041
R6950 2inmux_4.OUT.n0 2inmux_4.OUT.t3 26.9438
R6951 2inmux_4.OUT.n1 2inmux_4.OUT.t1 9.6935
R6952 dffrs_3.d 2inmux_4.OUT.n0 6.55979
R6953 2inmux_4.OUT dffrs_3.d 4.883
R6954 2inmux_4.OUT.n1 2inmux_4.OUT.t0 4.35383
R6955 2inmux_4.OUT 2inmux_4.OUT.n1 0.350857
R6956 a_25544_2511.n0 a_25544_2511.t6 41.0041
R6957 a_25544_2511.n1 a_25544_2511.t7 40.8177
R6958 a_25544_2511.n1 a_25544_2511.t5 27.1302
R6959 a_25544_2511.n0 a_25544_2511.t4 26.9438
R6960 a_25544_2511.n2 a_25544_2511.n1 22.5284
R6961 a_25544_2511.n3 a_25544_2511.n2 19.5781
R6962 a_25544_2511.n3 a_25544_2511.t2 10.0473
R6963 a_25544_2511.n4 a_25544_2511.t1 6.51042
R6964 a_25544_2511.n5 a_25544_2511.n4 6.04952
R6965 a_25544_2511.n2 a_25544_2511.n0 5.7305
R6966 a_25544_2511.n4 a_25544_2511.n3 0.732092
R6967 a_25544_2511.n5 a_25544_2511.t3 0.7285
R6968 a_25544_2511.t0 a_25544_2511.n5 0.7285
R6969 B5.n1 B5.t0 34.2529
R6970 B5.n0 B5.t1 19.673
R6971 B5.n0 B5.t2 19.4007
R6972 B5.n2 B5.n1 8.05164
R6973 B5.n2 B5 1.87121
R6974 B5.n1 B5.n0 0.106438
R6975 2inmux_2.In B5.n2 0.0455
R6976 a_10762_1160.n0 a_10762_1160.t5 34.1797
R6977 a_10762_1160.n0 a_10762_1160.t4 19.5798
R6978 a_10762_1160.n1 a_10762_1160.t2 18.7717
R6979 a_10762_1160.n1 a_10762_1160.t1 9.2885
R6980 a_10762_1160.n2 a_10762_1160.n0 4.93379
R6981 a_10762_1160.n3 a_10762_1160.t3 4.23346
R6982 a_10762_1160.t0 a_10762_1160.n3 3.85546
R6983 a_10762_1160.n2 a_10762_1160.n1 0.4055
R6984 a_10762_1160.n3 a_10762_1160.n2 0.352625
R6985 a_6520_5968.n0 a_6520_5968.t4 40.6313
R6986 a_6520_5968.n0 a_6520_5968.t5 27.3166
R6987 a_6520_5968.n1 a_6520_5968.n0 24.1527
R6988 a_6520_5968.n1 a_6520_5968.t2 10.0473
R6989 a_6520_5968.n2 a_6520_5968.t1 6.51042
R6990 a_6520_5968.n3 a_6520_5968.n2 6.04952
R6991 a_6520_5968.n2 a_6520_5968.n1 0.732092
R6992 a_6520_5968.t0 a_6520_5968.n3 0.7285
R6993 a_6520_5968.n3 a_6520_5968.t3 0.7285
R6994 serial_out.n0 serial_out.t4 40.6313
R6995 serial_out.n0 serial_out.t5 27.3166
R6996 serial_out.n4 serial_out.n0 14.6967
R6997 serial_out.n3 serial_out.t3 10.0473
R6998 serial_out.n4 serial_out.n3 9.39565
R6999 serial_out.n2 serial_out.t2 6.51042
R7000 serial_out.n2 serial_out.n1 6.04952
R7001 dffrs_5.Q serial_out 5.90514
R7002 serial_out.n3 serial_out.n2 0.732092
R7003 serial_out.n1 serial_out.t1 0.7285
R7004 serial_out.n1 serial_out.t0 0.7285
R7005 dffrs_5.Q serial_out.n4 0.458082
R7006 B2.n1 B2.t2 34.2529
R7007 B2.n0 B2.t0 19.673
R7008 B2.n0 B2.t1 19.4007
R7009 B2.n2 B2.n1 8.05164
R7010 B2.n2 B2 1.87121
R7011 B2.n1 B2.n0 0.106438
R7012 2inmux_5.In B2.n2 0.0455
R7013 a_39178_1161.n0 a_39178_1161.t5 34.1797
R7014 a_39178_1161.n0 a_39178_1161.t4 19.5798
R7015 a_39178_1161.n1 a_39178_1161.t2 18.7717
R7016 a_39178_1161.n1 a_39178_1161.t1 9.2885
R7017 a_39178_1161.n2 a_39178_1161.n0 4.93379
R7018 a_39178_1161.t0 a_39178_1161.n3 4.23346
R7019 a_39178_1161.n3 a_39178_1161.t3 3.85546
R7020 a_39178_1161.n2 a_39178_1161.n1 0.4055
R7021 a_39178_1161.n3 a_39178_1161.n2 0.352625
R7022 2inmux_5.OUT.n0 2inmux_5.OUT.t3 41.0041
R7023 2inmux_5.OUT.n0 2inmux_5.OUT.t2 26.9438
R7024 2inmux_5.OUT.n1 2inmux_5.OUT.t1 9.6935
R7025 dffrs_4.d 2inmux_5.OUT.n0 6.55979
R7026 2inmux_5.OUT dffrs_4.d 4.883
R7027 2inmux_5.OUT.n1 2inmux_5.OUT.t0 4.35383
R7028 2inmux_5.OUT 2inmux_5.OUT.n1 0.350857
R7029 B4.n1 B4.t1 34.2529
R7030 B4.n0 B4.t0 19.673
R7031 B4.n0 B4.t2 19.4007
R7032 B4.n2 B4.n1 8.05164
R7033 B4.n2 B4 1.87282
R7034 B4.n1 B4.n0 0.106438
R7035 2inmux_3.In B4.n2 0.0455
R7036 B1.n1 B1.t1 34.2529
R7037 B1.n0 B1.t0 19.673
R7038 B1.n0 B1.t2 19.4007
R7039 B1.n2 B1.n1 8.05164
R7040 B1.n2 B1 1.87121
R7041 B1.n1 B1.n0 0.106438
R7042 2inmux_1.In B1.n2 0.0455
R7043 B3.n1 B3.t1 34.2529
R7044 B3.n0 B3.t0 19.673
R7045 B3.n0 B3.t2 19.4007
R7046 B3.n2 B3.n1 8.05164
R7047 B3.n2 B3 1.87121
R7048 B3.n1 B3.n0 0.106438
R7049 2inmux_4.In B3.n2 0.0455
.ends

