magic
tech gf180mcuD
magscale 1 10
timestamp 1757500055
<< nwell >>
rect -1110 -310 1110 310
<< pmos >>
rect -860 -100 -660 100
rect -556 -100 -356 100
rect -252 -100 -52 100
rect 52 -100 252 100
rect 356 -100 556 100
rect 660 -100 860 100
<< pdiff >>
rect -948 87 -860 100
rect -948 -87 -935 87
rect -889 -87 -860 87
rect -948 -100 -860 -87
rect -660 87 -556 100
rect -660 -87 -631 87
rect -585 -87 -556 87
rect -660 -100 -556 -87
rect -356 87 -252 100
rect -356 -87 -327 87
rect -281 -87 -252 87
rect -356 -100 -252 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 252 87 356 100
rect 252 -87 281 87
rect 327 -87 356 87
rect 252 -100 356 -87
rect 556 87 660 100
rect 556 -87 585 87
rect 631 -87 660 87
rect 556 -100 660 -87
rect 860 87 948 100
rect 860 -87 889 87
rect 935 -87 948 87
rect 860 -100 948 -87
<< pdiffc >>
rect -935 -87 -889 87
rect -631 -87 -585 87
rect -327 -87 -281 87
rect -23 -87 23 87
rect 281 -87 327 87
rect 585 -87 631 87
rect 889 -87 935 87
<< nsubdiff >>
rect -1086 214 1086 286
rect -1086 170 -1014 214
rect -1086 -170 -1073 170
rect -1027 -170 -1014 170
rect 1014 170 1086 214
rect -1086 -214 -1014 -170
rect 1014 -170 1027 170
rect 1073 -170 1086 170
rect 1014 -214 1086 -170
rect -1086 -286 1086 -214
<< nsubdiffcont >>
rect -1073 -170 -1027 170
rect 1027 -170 1073 170
<< polysilicon >>
rect -860 179 -660 192
rect -860 133 -847 179
rect -673 133 -660 179
rect -860 100 -660 133
rect -556 179 -356 192
rect -556 133 -543 179
rect -369 133 -356 179
rect -556 100 -356 133
rect -252 179 -52 192
rect -252 133 -239 179
rect -65 133 -52 179
rect -252 100 -52 133
rect 52 179 252 192
rect 52 133 65 179
rect 239 133 252 179
rect 52 100 252 133
rect 356 179 556 192
rect 356 133 369 179
rect 543 133 556 179
rect 356 100 556 133
rect 660 179 860 192
rect 660 133 673 179
rect 847 133 860 179
rect 660 100 860 133
rect -860 -133 -660 -100
rect -860 -179 -847 -133
rect -673 -179 -660 -133
rect -860 -192 -660 -179
rect -556 -133 -356 -100
rect -556 -179 -543 -133
rect -369 -179 -356 -133
rect -556 -192 -356 -179
rect -252 -133 -52 -100
rect -252 -179 -239 -133
rect -65 -179 -52 -133
rect -252 -192 -52 -179
rect 52 -133 252 -100
rect 52 -179 65 -133
rect 239 -179 252 -133
rect 52 -192 252 -179
rect 356 -133 556 -100
rect 356 -179 369 -133
rect 543 -179 556 -133
rect 356 -192 556 -179
rect 660 -133 860 -100
rect 660 -179 673 -133
rect 847 -179 860 -133
rect 660 -192 860 -179
<< polycontact >>
rect -847 133 -673 179
rect -543 133 -369 179
rect -239 133 -65 179
rect 65 133 239 179
rect 369 133 543 179
rect 673 133 847 179
rect -847 -179 -673 -133
rect -543 -179 -369 -133
rect -239 -179 -65 -133
rect 65 -179 239 -133
rect 369 -179 543 -133
rect 673 -179 847 -133
<< metal1 >>
rect -1073 170 -1027 181
rect -858 133 -847 179
rect -673 133 -662 179
rect -554 133 -543 179
rect -369 133 -358 179
rect -250 133 -239 179
rect -65 133 -54 179
rect 54 133 65 179
rect 239 133 250 179
rect 358 133 369 179
rect 543 133 554 179
rect 662 133 673 179
rect 847 133 858 179
rect 1027 170 1073 181
rect -935 87 -889 98
rect -935 -98 -889 -87
rect -631 87 -585 98
rect -631 -98 -585 -87
rect -327 87 -281 98
rect -327 -98 -281 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 281 87 327 98
rect 281 -98 327 -87
rect 585 87 631 98
rect 585 -98 631 -87
rect 889 87 935 98
rect 889 -98 935 -87
rect -1073 -181 -1027 -170
rect -858 -179 -847 -133
rect -673 -179 -662 -133
rect -554 -179 -543 -133
rect -369 -179 -358 -133
rect -250 -179 -239 -133
rect -65 -179 -54 -133
rect 54 -179 65 -133
rect 239 -179 250 -133
rect 358 -179 369 -133
rect 543 -179 554 -133
rect 662 -179 673 -133
rect 847 -179 858 -133
rect 1027 -181 1073 -170
<< properties >>
string FIXED_BBOX -1050 -250 1050 250
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
