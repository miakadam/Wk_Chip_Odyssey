magic
tech gf180mcuD
magscale 1 10
timestamp 1757048890
<< pwell >>
rect -958 -360 958 360
<< nmos >>
rect -708 -150 -508 150
rect -404 -150 -204 150
rect -100 -150 100 150
rect 204 -150 404 150
rect 508 -150 708 150
<< ndiff >>
rect -796 137 -708 150
rect -796 -137 -783 137
rect -737 -137 -708 137
rect -796 -150 -708 -137
rect -508 137 -404 150
rect -508 -137 -479 137
rect -433 -137 -404 137
rect -508 -150 -404 -137
rect -204 137 -100 150
rect -204 -137 -175 137
rect -129 -137 -100 137
rect -204 -150 -100 -137
rect 100 137 204 150
rect 100 -137 129 137
rect 175 -137 204 137
rect 100 -150 204 -137
rect 404 137 508 150
rect 404 -137 433 137
rect 479 -137 508 137
rect 404 -150 508 -137
rect 708 137 796 150
rect 708 -137 737 137
rect 783 -137 796 137
rect 708 -150 796 -137
<< ndiffc >>
rect -783 -137 -737 137
rect -479 -137 -433 137
rect -175 -137 -129 137
rect 129 -137 175 137
rect 433 -137 479 137
rect 737 -137 783 137
<< psubdiff >>
rect -934 264 934 336
rect -934 220 -862 264
rect -934 -220 -921 220
rect -875 -220 -862 220
rect 862 220 934 264
rect -934 -264 -862 -220
rect 862 -220 875 220
rect 921 -220 934 220
rect 862 -264 934 -220
rect -934 -336 934 -264
<< psubdiffcont >>
rect -921 -220 -875 220
rect 875 -220 921 220
<< polysilicon >>
rect -708 229 -508 242
rect -708 183 -695 229
rect -521 183 -508 229
rect -708 150 -508 183
rect -404 229 -204 242
rect -404 183 -391 229
rect -217 183 -204 229
rect -404 150 -204 183
rect -100 229 100 242
rect -100 183 -87 229
rect 87 183 100 229
rect -100 150 100 183
rect 204 229 404 242
rect 204 183 217 229
rect 391 183 404 229
rect 204 150 404 183
rect 508 229 708 242
rect 508 183 521 229
rect 695 183 708 229
rect 508 150 708 183
rect -708 -183 -508 -150
rect -708 -229 -695 -183
rect -521 -229 -508 -183
rect -708 -242 -508 -229
rect -404 -183 -204 -150
rect -404 -229 -391 -183
rect -217 -229 -204 -183
rect -404 -242 -204 -229
rect -100 -183 100 -150
rect -100 -229 -87 -183
rect 87 -229 100 -183
rect -100 -242 100 -229
rect 204 -183 404 -150
rect 204 -229 217 -183
rect 391 -229 404 -183
rect 204 -242 404 -229
rect 508 -183 708 -150
rect 508 -229 521 -183
rect 695 -229 708 -183
rect 508 -242 708 -229
<< polycontact >>
rect -695 183 -521 229
rect -391 183 -217 229
rect -87 183 87 229
rect 217 183 391 229
rect 521 183 695 229
rect -695 -229 -521 -183
rect -391 -229 -217 -183
rect -87 -229 87 -183
rect 217 -229 391 -183
rect 521 -229 695 -183
<< metal1 >>
rect -921 277 921 323
rect -921 220 -875 277
rect -706 183 -695 229
rect -521 183 -510 229
rect -402 183 -391 229
rect -217 183 -206 229
rect -98 183 -87 229
rect 87 183 98 229
rect 206 183 217 229
rect 391 183 402 229
rect 510 183 521 229
rect 695 183 706 229
rect 875 220 921 277
rect -783 137 -737 148
rect -783 -148 -737 -137
rect -479 137 -433 148
rect -479 -148 -433 -137
rect -175 137 -129 148
rect -175 -148 -129 -137
rect 129 137 175 148
rect 129 -148 175 -137
rect 433 137 479 148
rect 433 -148 479 -137
rect 737 137 783 148
rect 737 -148 783 -137
rect -921 -277 -875 -220
rect -706 -229 -695 -183
rect -521 -229 -510 -183
rect -402 -229 -391 -183
rect -217 -229 -206 -183
rect -98 -229 -87 -183
rect 87 -229 98 -183
rect 206 -229 217 -183
rect 391 -229 402 -183
rect 510 -229 521 -183
rect 695 -229 706 -183
rect 875 -277 921 -220
rect -921 -323 921 -277
<< properties >>
string FIXED_BBOX -898 -300 898 300
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.5 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
