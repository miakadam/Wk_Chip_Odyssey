magic
tech gf180mcuD
magscale 1 10
timestamp 1757365333
<< error_p >>
rect -38 -455 -27 -409
<< nwell >>
rect -290 -586 290 586
<< pmos >>
rect -40 -376 40 424
<< pdiff >>
rect -128 411 -40 424
rect -128 -363 -115 411
rect -69 -363 -40 411
rect -128 -376 -40 -363
rect 40 411 128 424
rect 40 -363 69 411
rect 115 -363 128 411
rect 40 -376 128 -363
<< pdiffc >>
rect -115 -363 -69 411
rect 69 -363 115 411
<< nsubdiff >>
rect -266 490 266 562
rect -266 446 -194 490
rect -266 -446 -253 446
rect -207 -446 -194 446
rect 194 446 266 490
rect -266 -490 -194 -446
rect 194 -446 207 446
rect 253 -446 266 446
rect 194 -490 266 -446
rect -266 -562 266 -490
<< nsubdiffcont >>
rect -253 -446 -207 446
rect 207 -446 253 446
<< polysilicon >>
rect -40 424 40 468
rect -40 -409 40 -376
rect -40 -455 -27 -409
rect 27 -455 40 -409
rect -40 -468 40 -455
<< polycontact >>
rect -27 -455 27 -409
<< metal1 >>
rect -253 446 -207 457
rect 207 446 253 457
rect -115 411 -69 422
rect -115 -374 -69 -363
rect 69 411 115 422
rect 69 -374 115 -363
rect -253 -457 -207 -446
rect -38 -455 -27 -409
rect 27 -455 38 -409
rect 207 -457 253 -446
<< properties >>
string FIXED_BBOX -230 -526 230 526
string gencell pfet_03v3
string library gf180mcu
string parameters w 4.0 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
