* NGSPICE file created from dffrs.ext - technology: (null)

.subckt dffrs vdd vss d clk setb resetb Q Qb
X0 a_292_1130 nand3_8.Z a_108_1130 vss.t12 nfet_03v3
**devattr s=10400,304 d=10400,304
X1 a_1778_n3279 nand3_8.C.t4 a_1594_n3279 vss.t21 nfet_03v3
**devattr s=10400,304 d=10400,304
X2 nand3_0.Z setb.t0 vdd.t25 vdd.t24 pfet_03v3
**devattr s=44000,1176 d=26000,604
X3 nand3_0.Z nand3_6.C.t4 vdd.t9 vdd.t8 pfet_03v3
**devattr s=26000,604 d=44000,1176
X4 a_108_n1075 nand3_0.Z vss.t4 vss.t3 nfet_03v3
**devattr s=17600,576 d=10400,304
X5 a_108_n3280 nand3_6.C.t5 vss.t2 vss.t1 nfet_03v3
**devattr s=17600,576 d=10400,304
X6 nand3_6.C.t0 nand3_0.Z vdd.t1 vdd.t0 pfet_03v3
**devattr s=44000,1176 d=26000,604
X7 Q.t2 setb.t1 vdd.t23 vdd.t22 pfet_03v3
**devattr s=44000,1176 d=26000,604
X8 Qb.t0 resetb.t0 vdd.t19 vdd.t18 pfet_03v3
**devattr s=26000,604 d=44000,1176
X9 vdd.t3 resetb.t1 nand3_8.Z vdd.t2 pfet_03v3
**devattr s=26000,604 d=26000,604
X10 nand3_6.C.t2 clk.t0 vdd.t27 vdd.t26 pfet_03v3
**devattr s=26000,604 d=44000,1176
X11 Q.t3 Qb.t4 a_1778_n1075 vss.t20 nfet_03v3
**devattr s=10400,304 d=17600,576
X12 a_1594_n3279 Q.t4 vss.t14 vss.t13 nfet_03v3
**devattr s=17600,576 d=10400,304
X13 nand3_6.C.t1 clk.t1 a_292_n1075 vss.t15 nfet_03v3
**devattr s=10400,304 d=17600,576
X14 vdd.t35 nand3_8.C.t5 Qb.t3 vdd.t34 pfet_03v3
**devattr s=26000,604 d=26000,604
X15 a_108_1130 setb.t2 vss.t19 vss.t18 nfet_03v3
**devattr s=17600,576 d=10400,304
X16 nand3_0.Z nand3_6.C.t6 a_292_1130 vss.t6 nfet_03v3
**devattr s=10400,304 d=17600,576
X17 a_1778_n1075 nand3_6.C.t7 a_1594_n1075 vss.t17 nfet_03v3
**devattr s=10400,304 d=10400,304
X18 nand3_8.C.t1 nand3_8.Z a_292_n3280 vss.t11 nfet_03v3
**devattr s=10400,304 d=17600,576
X19 nand3_8.C.t3 nand3_6.C.t8 vdd.t21 vdd.t20 pfet_03v3
**devattr s=44000,1176 d=26000,604
X20 a_108_n5485 nand3_8.C.t6 vss.t23 vss.t22 nfet_03v3
**devattr s=17600,576 d=10400,304
X21 vdd.t5 nand3_6.C.t9 Q.t0 vdd.t4 pfet_03v3
**devattr s=26000,604 d=26000,604
X22 Qb.t2 Q.t5 vdd.t29 vdd.t28 pfet_03v3
**devattr s=44000,1176 d=26000,604
X23 a_292_n1075 resetb.t2 a_108_n1075 vss.t10 nfet_03v3
**devattr s=10400,304 d=10400,304
X24 a_292_n3280 clk.t2 a_108_n3280 vss.t16 nfet_03v3
**devattr s=10400,304 d=10400,304
X25 a_1594_n1075 setb.t3 vss.t8 vss.t7 nfet_03v3
**devattr s=17600,576 d=10400,304
X26 nand3_8.C.t2 nand3_8.Z vdd.t15 vdd.t14 pfet_03v3
**devattr s=26000,604 d=44000,1176
X27 nand3_8.Z d.t0 a_292_n5485 vss.t0 nfet_03v3
**devattr s=10400,304 d=17600,576
X28 nand3_8.Z nand3_8.C.t7 vdd.t33 vdd.t32 pfet_03v3
**devattr s=44000,1176 d=26000,604
X29 vdd.t13 nand3_8.Z nand3_0.Z vdd.t12 pfet_03v3
**devattr s=26000,604 d=26000,604
X30 vdd.t31 resetb.t3 nand3_6.C.t3 vdd.t30 pfet_03v3
**devattr s=26000,604 d=26000,604
X31 Q.t1 Qb.t5 vdd.t17 vdd.t16 pfet_03v3
**devattr s=26000,604 d=44000,1176
X32 vdd.t7 clk.t3 nand3_8.C.t0 vdd.t6 pfet_03v3
**devattr s=26000,604 d=26000,604
X33 Qb.t1 resetb.t4 a_1778_n3279 vss.t9 nfet_03v3
**devattr s=10400,304 d=17600,576
X34 a_292_n5485 resetb.t5 a_108_n5485 vss.t5 nfet_03v3
**devattr s=10400,304 d=10400,304
X35 nand3_8.Z d.t1 vdd.t11 vdd.t10 pfet_03v3
**devattr s=26000,604 d=44000,1176
R0 vss.n45 vss.n16 25102.2
R1 vss.n15 vss.n14 7590.9
R2 vss.n46 vss.n15 7328.43
R3 vss.n61 vss.n60 5916.76
R4 vss.n47 vss.n46 5557.62
R5 vss.n48 vss.n47 5551.58
R6 vss.n60 vss.n2 4776.36
R7 vss.n16 vss.n2 4776.36
R8 vss.n46 vss.n45 1101.64
R9 vss.n60 vss.n59 943.385
R10 vss.n24 vss.n2 943.385
R11 vss.n17 vss.n16 943.385
R12 vss.n47 vss.n12 832.22
R13 vss.n47 vss.n13 832.101
R14 vss.n10 vss.t0 703.198
R15 vss.n61 vss.t22 703.198
R16 vss.n34 vss.n15 668.225
R17 vss.n34 vss.t20 582.165
R18 vss.t7 vss.n12 582.165
R19 vss.n9 vss.t11 581.712
R20 vss.n59 vss.t1 581.712
R21 vss.t15 vss.n13 581.712
R22 vss.n24 vss.t3 581.712
R23 vss.n44 vss.t6 581.712
R24 vss.n17 vss.t18 581.712
R25 vss.t0 vss.t5 562.559
R26 vss.t5 vss.t22 562.559
R27 vss.t20 vss.t17 465.733
R28 vss.t17 vss.t7 465.733
R29 vss.t11 vss.t16 465.37
R30 vss.t16 vss.t1 465.37
R31 vss.t10 vss.t15 465.37
R32 vss.t3 vss.t10 465.37
R33 vss.t12 vss.t6 465.37
R34 vss.t18 vss.t12 465.37
R35 vss.n49 vss.n48 327.089
R36 vss.n48 vss.n11 267.438
R37 vss.n14 vss.t9 228.663
R38 vss.n49 vss.t13 228.663
R39 vss.n11 vss.n10 183.444
R40 vss.t9 vss.t21 182.931
R41 vss.t21 vss.t13 182.931
R42 vss.n11 vss.n9 151.751
R43 vss.n45 vss.n44 151.751
R44 vss.n43 vss.n18 61.0571
R45 vss.n50 vss.n8 61.0561
R46 vss.n62 vss.n1 61.0561
R47 vss.n58 vss.n3 61.0561
R48 vss.n26 vss.n25 61.0561
R49 vss.n35 vss.n33 61.0561
R50 vss.n64 vss.n0 9.05442
R51 vss.n56 vss.n55 9.0005
R52 vss.n42 vss.n41 9.0005
R53 vss.n40 vss.n20 9.0005
R54 vss.n37 vss.n36 9.0005
R55 vss.n31 vss.n30 9.0005
R56 vss.n28 vss.n27 9.0005
R57 vss.n22 vss.n21 9.0005
R58 vss.n66 vss.n65 9.0005
R59 vss.n7 vss.n4 9.0005
R60 vss.n52 vss.n8 6.9012
R61 vss.n4 vss.n3 6.46296
R62 vss.n27 vss.n26 6.46296
R63 vss.n36 vss.n35 6.46296
R64 vss.n65 vss.n1 6.4618
R65 vss.n43 vss.n42 6.4618
R66 vss.n52 vss.n51 5.47239
R67 vss.n57 vss.n56 5.03414
R68 vss.n64 vss.n63 5.03414
R69 vss.n23 vss.n22 5.03414
R70 vss.n32 vss.n31 5.03414
R71 vss.n20 vss.n19 5.03414
R72 vss.n51 vss.t14 4.7885
R73 vss.n57 vss.t2 4.7885
R74 vss.n63 vss.t23 4.7885
R75 vss.n23 vss.t4 4.7885
R76 vss.n32 vss.t8 4.7885
R77 vss.n19 vss.t19 4.7885
R78 vss.n53 vss.n52 4.28213
R79 vss.n9 vss.n3 1.3005
R80 vss.n58 vss.n57 1.3005
R81 vss.n59 vss.n58 1.3005
R82 vss.n10 vss.n1 1.3005
R83 vss.n63 vss.n62 1.3005
R84 vss.n62 vss.n61 1.3005
R85 vss.n14 vss.n8 1.3005
R86 vss.n51 vss.n50 1.3005
R87 vss.n50 vss.n49 1.3005
R88 vss.n35 vss.n34 1.3005
R89 vss.n33 vss.n32 1.3005
R90 vss.n33 vss.n12 1.3005
R91 vss.n26 vss.n13 1.3005
R92 vss.n25 vss.n23 1.3005
R93 vss.n25 vss.n24 1.3005
R94 vss.n19 vss.n18 1.3005
R95 vss.n18 vss.n17 1.3005
R96 vss.n44 vss.n43 1.3005
R97 vss.n65 vss.n64 0.92075
R98 vss.n56 vss.n4 0.92075
R99 vss.n27 vss.n22 0.92075
R100 vss.n36 vss.n31 0.92075
R101 vss.n42 vss.n20 0.92075
R102 vss.n39 vss.n38 0.122607
R103 vss.n55 vss.n0 0.115241
R104 vss.n54 vss.n5 0.10457
R105 vss.n7 vss.n0 0.0645882
R106 vss.n38 vss.n6 0.0622481
R107 vss.n55 vss.n54 0.054837
R108 vss.n40 vss.n5 0.0466843
R109 vss.n54 vss.n6 0.0415307
R110 vss.n41 vss.n40 0.0405109
R111 vss.n37 vss.n30 0.0405109
R112 vss.n28 vss.n21 0.0405109
R113 vss.n54 vss.n53 0.0349747
R114 vss.n66 vss.n0 0.0347517
R115 vss.n39 vss.n29 0.0322085
R116 vss.n29 vss.n6 0.0322085
R117 vss.n41 vss.n39 0.0214837
R118 vss.n29 vss.n28 0.0214837
R119 vss.n30 vss.n29 0.0121902
R120 vss.n38 vss.n37 0.00915761
R121 vss vss.n66 0.00754658
R122 vss.n21 vss.n5 0.00720109
R123 vss.n53 vss.n7 0.000544599
R124 nand3_8.C.n0 nand3_8.C.t5 40.8177
R125 nand3_8.C.n1 nand3_8.C.t7 40.6313
R126 nand3_8.C.n1 nand3_8.C.t6 27.3166
R127 nand3_8.C.n0 nand3_8.C.t4 27.1302
R128 nand3_8.C.n3 nand3_8.C.n2 14.119
R129 nand3_8.C.n6 nand3_8.C.t1 10.0473
R130 nand3_8.C.n5 nand3_8.C.t2 6.51042
R131 nand3_8.C.n5 nand3_8.C.n4 6.04952
R132 nand3_7.B nand3_8.C.n0 5.47979
R133 nand3_8.C.n2 nand3_8.C.n1 5.13907
R134 nand3_6.Z nand3_8.C.n6 4.72925
R135 nand3_8.C.n6 nand3_8.C.n5 0.732092
R136 nand3_8.C.n4 nand3_8.C.t0 0.7285
R137 nand3_8.C.n4 nand3_8.C.t3 0.7285
R138 nand3_8.C.n3 nand3_7.B 0.438233
R139 nand3_6.Z nand3_8.C.n3 0.166901
R140 nand3_8.C.n2 nand3_8.C 0.0455
R141 setb.n2 setb.t0 40.6313
R142 setb.n0 setb.t1 40.6313
R143 setb.n2 setb.t2 27.3166
R144 setb.n0 setb.t3 27.3166
R145 setb.n3 setb.n1 9.22229
R146 setb.n3 setb.n2 5.14711
R147 setb.n1 setb.n0 5.13907
R148 nand3_0.C setb 0.784786
R149 setb.n1 nand3_2.C 0.0455
R150 nand3_0.C setb.n3 0.0374643
R151 vdd.t8 vdd.n29 250.9
R152 vdd.n30 vdd.t24 250.9
R153 vdd.t26 vdd.n23 250.9
R154 vdd.n24 vdd.t0 250.9
R155 vdd.t16 vdd.n1 250.9
R156 vdd.n2 vdd.t22 250.9
R157 vdd.t14 vdd.n11 250.9
R158 vdd.n12 vdd.t20 250.9
R159 vdd.t18 vdd.n17 250.9
R160 vdd.n18 vdd.t28 250.9
R161 vdd.t10 vdd.n6 250.9
R162 vdd.n7 vdd.t32 250.9
R163 vdd.t12 vdd.t8 200
R164 vdd.t24 vdd.t12 200
R165 vdd.t30 vdd.t26 200
R166 vdd.t0 vdd.t30 200
R167 vdd.t4 vdd.t16 200
R168 vdd.t22 vdd.t4 200
R169 vdd.t6 vdd.t14 200
R170 vdd.t20 vdd.t6 200
R171 vdd.t34 vdd.t18 200
R172 vdd.t28 vdd.t34 200
R173 vdd.t2 vdd.t10 200
R174 vdd.t32 vdd.t2 200
R175 vdd.n30 vdd.n29 68.0765
R176 vdd.n24 vdd.n23 68.0765
R177 vdd.n2 vdd.n1 68.0765
R178 vdd.n12 vdd.n11 68.0765
R179 vdd.n18 vdd.n17 68.0765
R180 vdd.n7 vdd.n6 68.0765
R181 vdd.n15 vdd.n9 13.5406
R182 vdd.n33 vdd.n32 13.5005
R183 vdd.n27 vdd.n26 13.5005
R184 vdd.n27 vdd.n4 13.5005
R185 vdd.n15 vdd.n14 13.5005
R186 vdd.n21 vdd.n20 13.5005
R187 vdd.n32 vdd.n29 6.4802
R188 vdd.n26 vdd.n23 6.4802
R189 vdd.n4 vdd.n1 6.4802
R190 vdd.n14 vdd.n11 6.4802
R191 vdd.n20 vdd.n17 6.4802
R192 vdd.n9 vdd.n6 6.4802
R193 vdd.n32 vdd.n28 6.25878
R194 vdd.n26 vdd.n22 6.25878
R195 vdd.n4 vdd.n0 6.25878
R196 vdd.n14 vdd.n10 6.25878
R197 vdd.n20 vdd.n16 6.25878
R198 vdd.n9 vdd.n5 6.25878
R199 vdd.n32 vdd.n31 5.44497
R200 vdd.n26 vdd.n25 5.44497
R201 vdd.n4 vdd.n3 5.44497
R202 vdd.n14 vdd.n13 5.44497
R203 vdd.n20 vdd.n19 5.44497
R204 vdd.n9 vdd.n8 5.44497
R205 vdd.n31 vdd.t25 1.85637
R206 vdd.n25 vdd.t1 1.85637
R207 vdd.n3 vdd.t23 1.85637
R208 vdd.n13 vdd.t21 1.85637
R209 vdd.n19 vdd.t29 1.85637
R210 vdd.n8 vdd.t33 1.85637
R211 vdd.n31 vdd.n30 1.04105
R212 vdd.n25 vdd.n24 1.04105
R213 vdd.n3 vdd.n2 1.04105
R214 vdd.n13 vdd.n12 1.04105
R215 vdd.n19 vdd.n18 1.04105
R216 vdd.n8 vdd.n7 1.04105
R217 vdd.n28 vdd.t9 0.7285
R218 vdd.n28 vdd.t13 0.7285
R219 vdd.n22 vdd.t27 0.7285
R220 vdd.n22 vdd.t31 0.7285
R221 vdd.n0 vdd.t17 0.7285
R222 vdd.n0 vdd.t5 0.7285
R223 vdd.n10 vdd.t15 0.7285
R224 vdd.n10 vdd.t7 0.7285
R225 vdd.n16 vdd.t19 0.7285
R226 vdd.n16 vdd.t35 0.7285
R227 vdd.n5 vdd.t11 0.7285
R228 vdd.n5 vdd.t3 0.7285
R229 vdd.n33 vdd.n27 0.0405909
R230 vdd.n27 vdd.n21 0.0405727
R231 vdd vdd.n33 0.00297273
R232 vdd.n21 vdd.n15 0.000518182
R233 nand3_6.C.n1 nand3_6.C.t4 41.0041
R234 nand3_6.C.n0 nand3_6.C.t9 40.8177
R235 nand3_6.C.n3 nand3_6.C.t8 40.6313
R236 nand3_6.C.n3 nand3_6.C.t5 27.3166
R237 nand3_6.C.n0 nand3_6.C.t7 27.1302
R238 nand3_6.C.n1 nand3_6.C.t6 26.9438
R239 nand3_6.C.n9 nand3_6.C.t1 10.0473
R240 nand3_6.C.n5 nand3_6.C.n4 9.90747
R241 nand3_6.C.n5 nand3_6.C.n2 9.90116
R242 nand3_6.C.n8 nand3_6.C.t2 6.51042
R243 nand3_6.C.n8 nand3_6.C.n7 6.04952
R244 nand3_6.C.n2 nand3_6.C.n1 5.7305
R245 nand3_2.B nand3_6.C.n0 5.47979
R246 nand3_6.C.n4 nand3_6.C.n3 5.13907
R247 nand3_1.Z nand3_6.C.n9 4.72925
R248 nand3_6.C.n6 nand3_6.C.n5 4.5005
R249 nand3_6.C.n9 nand3_6.C.n8 0.732092
R250 nand3_6.C.n7 nand3_6.C.t3 0.7285
R251 nand3_6.C.n7 nand3_6.C.t0 0.7285
R252 nand3_1.Z nand3_6.C.n6 0.449758
R253 nand3_6.C.n6 nand3_2.B 0.166901
R254 nand3_6.C.n2 nand3_0.A 0.0455
R255 nand3_6.C.n4 nand3_6.C 0.0455
R256 Q.n0 Q.t5 40.6313
R257 Q.n0 Q.t4 27.3166
R258 Q.n3 Q.t3 10.0473
R259 Q.n5 Q.n4 9.55818
R260 Q.n2 Q.t1 6.51042
R261 Q.n2 Q.n1 6.04952
R262 Q.n5 Q.n0 5.13907
R263 nand3_2.Z Q.n3 4.72925
R264 Q.n4 nand3_2.Z 4.6669
R265 Q.n3 Q.n2 0.732092
R266 Q.n1 Q.t0 0.7285
R267 Q.n1 Q.t2 0.7285
R268 Q.n4 Q 0.458082
R269 nand3_7.C Q.n5 0.0455
R270 resetb.n0 resetb.t0 41.0041
R271 resetb.n2 resetb.t1 40.8177
R272 resetb.n1 resetb.t3 40.8177
R273 resetb.n2 resetb.t5 27.1302
R274 resetb.n1 resetb.t2 27.1302
R275 resetb.n0 resetb.t4 26.9438
R276 resetb.n3 nand3_1.B 12.1571
R277 resetb.n5 resetb.n4 7.75389
R278 resetb.n4 resetb.n3 5.93546
R279 resetb.n5 resetb.n0 5.7305
R280 nand3_8.B resetb.n2 5.47979
R281 nand3_1.B resetb.n1 5.47979
R282 resetb.n3 nand3_8.B 5.09593
R283 resetb.n4 resetb 0.136036
R284 nand3_7.A resetb.n5 0.0455
R285 Qb.n0 Qb.t5 41.0041
R286 Qb.n0 Qb.t4 26.9438
R287 Qb.n3 Qb.t1 10.0473
R288 Qb.n5 Qb.n4 9.84255
R289 Qb.n2 Qb.t0 6.51042
R290 Qb.n2 Qb.n1 6.04952
R291 Qb.n5 Qb.n0 5.7305
R292 Qb.n4 nand3_7.Z 4.94976
R293 nand3_7.Z Qb.n3 4.72925
R294 Qb.n3 Qb.n2 0.732092
R295 Qb.n1 Qb.t3 0.7285
R296 Qb.n1 Qb.t2 0.7285
R297 Qb.n4 Qb 0.175225
R298 nand3_2.A Qb.n5 0.0455
R299 clk.n0 clk.t0 41.0041
R300 clk.n1 clk.t3 40.8177
R301 clk.n1 clk.t2 27.1302
R302 clk.n0 clk.t1 26.9438
R303 nand3_1.A clk.n0 5.7755
R304 nand3_6.B clk.n1 5.47979
R305 clk.n2 nand3_6.B 2.17818
R306 nand3_1.A clk.n2 1.34729
R307 clk.n2 clk 0.611214
R308 d.n0 d.t1 41.0041
R309 d.n0 d.t0 26.9438
R310 nand3_8.A d.n0 5.7755
R311 nand3_8.A d 0.784786
.ends

