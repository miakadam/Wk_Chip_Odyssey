magic
tech gf180mcuD
magscale 1 10
timestamp 1757714585
<< metal1 >>
rect 1480 4000 13900 4380
rect 4011 1082 4089 4000
rect 5620 3320 5700 4000
rect 7880 3040 7960 4000
rect 6700 2380 6780 2600
rect 9100 2380 9180 4000
rect 5565 1279 5659 1291
rect 7675 1279 7747 1281
rect 5565 1203 5577 1279
rect 5657 1203 6695 1279
rect 6823 1203 7677 1279
rect 7733 1203 7747 1279
rect 5565 1201 5659 1203
rect 7675 1191 7747 1203
rect 4010 881 4090 1082
rect 3993 864 4106 881
rect 3993 786 4010 864
rect 4090 786 4106 864
rect 3993 775 4106 786
rect 4869 543 7471 546
rect 7891 543 7957 1518
rect 8123 1279 8195 1281
rect 10201 1279 10305 1291
rect 8123 1203 8137 1279
rect 8193 1203 8979 1279
rect 9175 1203 10213 1279
rect 10293 1203 10305 1279
rect 8123 1191 8195 1203
rect 10201 1201 10305 1203
rect 10421 1100 10499 4000
rect 10420 930 10500 1100
rect 10400 750 10520 930
rect 10400 690 10420 750
rect 10500 690 10520 750
rect 11305 552 11463 567
rect 11305 546 11332 552
rect 9182 543 11332 546
rect 3544 483 11332 543
rect 4396 454 4599 483
rect 4869 481 11332 483
rect 4396 365 4454 454
rect 4545 365 4599 454
rect 11305 445 11332 481
rect 11441 546 11463 552
rect 11441 481 11688 546
rect 11441 445 11463 481
rect 11305 434 11463 445
rect 4396 336 4599 365
rect 1470 -3350 6470 -3275
rect 1470 -3675 6470 -3600
rect 9953 -4257 10094 -4241
rect 9953 -4394 9967 -4257
rect 9952 -4467 9967 -4394
rect 10072 -4405 10094 -4257
rect 10072 -4467 10089 -4405
rect 9952 -4485 10089 -4467
rect 1565 -5180 7841 -5100
rect 1039 -5472 13459 -5418
rect 1039 -5473 9964 -5472
rect 1039 -5540 5457 -5473
rect 1039 -5627 4456 -5540
rect 4541 -5560 5457 -5540
rect 5546 -5478 9964 -5473
rect 5546 -5560 6013 -5478
rect 4541 -5627 6013 -5560
rect 1039 -5689 6013 -5627
rect 6368 -5675 9964 -5478
rect 10078 -5526 13459 -5472
rect 10078 -5628 10442 -5526
rect 10546 -5548 13459 -5526
rect 10546 -5628 11332 -5548
rect 10078 -5655 11332 -5628
rect 11441 -5655 13459 -5548
rect 10078 -5675 13459 -5655
rect 6368 -5689 13459 -5675
rect 1039 -5798 13459 -5689
<< via1 >>
rect 5577 1203 5657 1279
rect 7677 1203 7733 1279
rect 4010 786 4090 864
rect 8137 1203 8193 1279
rect 10213 1203 10293 1279
rect 10420 690 10500 750
rect 4454 365 4545 454
rect 11332 445 11441 552
rect 9967 -4467 10072 -4257
rect 4456 -5627 4541 -5540
rect 5457 -5560 5546 -5473
rect 6013 -5689 6368 -5478
rect 9964 -5675 10078 -5472
rect 10442 -5628 10546 -5526
rect 11332 -5655 11441 -5548
<< metal2 >>
rect 1725 2783 5325 2843
rect 5909 2527 7276 2579
rect 5985 2523 7276 2527
rect 7220 2136 7276 2523
rect 5565 1279 5659 1291
rect 7677 1281 7733 1302
rect 8137 1281 8193 1648
rect 5565 1203 5577 1279
rect 5657 1203 5659 1279
rect 5565 1201 5659 1203
rect 7675 1279 7747 1281
rect 7675 1203 7677 1279
rect 7733 1203 7747 1279
rect 3993 864 4106 881
rect 3993 786 4010 864
rect 4090 786 4106 864
rect 3993 775 4106 786
rect 4010 320 4090 775
rect 4446 454 4555 467
rect 4446 365 4454 454
rect 4545 365 4555 454
rect 4446 358 4555 365
rect 4000 300 4100 320
rect 4000 220 4010 300
rect 4090 220 4100 300
rect 4000 210 4100 220
rect 4454 -1018 4545 358
rect 5577 -924 5657 1201
rect 7675 1191 7747 1203
rect 8123 1279 8195 1281
rect 8123 1203 8137 1279
rect 8193 1203 8195 1279
rect 8123 1191 8195 1203
rect 10201 1279 10305 1291
rect 10201 1203 10213 1279
rect 10293 1203 10305 1279
rect 10201 1201 10305 1203
rect 10213 100 10293 1201
rect 10400 790 10520 810
rect 10400 690 10420 790
rect 10500 690 10520 790
rect 10400 670 10520 690
rect 11305 552 11463 567
rect 11305 445 11332 552
rect 11441 445 11463 552
rect 11305 434 11463 445
rect 4456 -5518 4543 -1018
rect 5449 -2466 5894 -2362
rect 9976 -2457 10546 -2353
rect 5457 -5220 5546 -2466
rect 9953 -4257 10094 -4241
rect 9953 -4394 9967 -4257
rect 9952 -4467 9967 -4394
rect 10072 -4405 10094 -4257
rect 10072 -4467 10089 -4405
rect 9952 -4485 10089 -4467
rect 5431 -5473 5583 -5220
rect 6018 -5469 6368 -4778
rect 9970 -5408 10069 -4485
rect 9970 -5453 10087 -5408
rect 9960 -5464 10087 -5453
rect 4432 -5540 4567 -5518
rect 4432 -5627 4456 -5540
rect 4541 -5627 4567 -5540
rect 5431 -5560 5457 -5473
rect 5546 -5560 5583 -5473
rect 5431 -5593 5583 -5560
rect 5999 -5478 6389 -5469
rect 4432 -5642 4567 -5627
rect 5999 -5689 6013 -5478
rect 6368 -5689 6389 -5478
rect 5999 -5710 6389 -5689
rect 9960 -5472 10086 -5464
rect 9960 -5675 9964 -5472
rect 10078 -5675 10086 -5472
rect 10442 -5516 10546 -2457
rect 10431 -5526 10559 -5516
rect 10431 -5628 10442 -5526
rect 10546 -5628 10559 -5526
rect 11332 -5536 11441 434
rect 10431 -5662 10559 -5628
rect 11322 -5548 11450 -5536
rect 11322 -5655 11332 -5548
rect 11441 -5655 11450 -5548
rect 9960 -5694 10086 -5675
rect 11322 -5677 11450 -5655
<< via2 >>
rect 4010 220 4090 300
rect 10420 750 10500 790
rect 10420 710 10500 750
<< metal3 >>
rect 10400 790 10520 810
rect 10400 710 10420 790
rect 10500 710 10520 790
rect 10400 690 10520 710
rect 4000 300 4100 320
rect 4000 220 4010 300
rect 4090 220 4100 300
rect 4000 210 4100 220
rect 4010 26 4090 210
rect 4010 -54 5310 26
rect 10420 -40 10500 690
use lvsclean_SAlatch  x1
timestamp 1757676563
transform 1 0 -9053 0 1 -1780
box 11023 -3410 22953 2129
use rslatch  x2
timestamp 1757675171
transform 1 0 5355 0 1 3480
box 1870 -2178 3290 -420
use inv_mia  x3
timestamp 1757680375
transform 1 0 1295 0 1 2105
box 5150 -1650 5730 322
use osu_sc_buf_4  x4
timestamp 1757675583
transform -1 0 6205 0 1 2073
box 0 -10 1140 1260
use inv_mia  x5
timestamp 1757680375
transform -1 0 14575 0 1 2105
box 5150 -1650 5730 322
<< labels >>
rlabel metal1 1470 -3310 1470 -3310 7 Vin1
port 6 w
rlabel metal1 1470 -3638 1470 -3638 7 Vin2
port 8 w
rlabel space 3494 -2927 3494 -2927 5 off3
port 5 s
rlabel space 1992 -2918 1992 -2918 5 off4
port 7 s
rlabel space 3392 -1380 3392 -1380 1 off2
port 3 n
rlabel space 4035 -1380 4035 -1380 1 off1
port 0 n
rlabel space 11850 -1380 11850 -1380 1 off5
port 9 n
rlabel space 12501 -1380 12501 -1380 1 off6
port 11 n
rlabel space 13866 -2918 13866 -2918 5 off8
port 13 s
rlabel space 12405 -2927 12405 -2927 5 off7
port 12 s
rlabel metal2 5577 172 5577 172 7 out1
rlabel metal2 10293 152 10293 152 3 out2
rlabel metal2 5618 192 5618 192 1 Vout2
port 6 n
rlabel metal1 1565 -5144 1565 -5144 7 CLK
port 4 w
rlabel space 7953 146 7953 146 1 VDD
rlabel space 5790 -4801 5790 -4801 7 VSS
rlabel space 5543 2063 5543 2063 5 VSS
port 2 s
rlabel metal1 7897 1460 7897 1460 5 VSS
rlabel metal1 9203 481 9203 481 5 VSS
rlabel metal1 6775 481 6775 481 5 VSS
rlabel space 9317 2389 9317 2389 1 VDD
rlabel space 6535 2389 6535 2389 1 VDD
rlabel space 7660 3060 7660 3060 1 VDD
rlabel space 5523 3333 5523 3333 1 VDD
port 1 n
rlabel metal2 6801 2579 6801 2579 1 latch
rlabel metal1 8411 1279 8411 1279 1 inv2
rlabel metal1 7231 1279 7231 1279 1 inv1
rlabel metal2 1725 2811 1725 2811 7 Vout
port 10 w
rlabel via1 5645 1229 5645 1229 3 in
port 2 w
rlabel via1 8161 1233 8161 1233 7 out
port 3 w
rlabel metal1 1524 4047 1530 4329 7 VDD
rlabel metal1 1101 -5744 1107 -5462 7 VSS
<< end >>
