* NGSPICE file created from comp_SAR_final.ext - technology: gf180mcuD

.subckt comparator_no_offsetcal VDD VSS CLK Vin1 Vin2 Vout
X0 VDD a_5265_2223# Vout VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 VDD a_6467_n692# a_6379_n600# VDD pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=1u
X2 no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X3 VSS a_7711_n4982# a_7623_n4890# VSS nfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.4u
X4 VDD a_5265_2223# Vout VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VDD no_offsetLatch_0.Vout2 x5.out VDD pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.4u
X6 no_offsetLatch_0.Vp CLK VDD VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X7 a_9403_n600# a_9203_n692# VDD VDD pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=1u
X8 VDD CLK no_offsetLatch_0.Vout2 VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X9 no_offsetLatch_0.Vout2 a_8125_n1848# a_8037_n1756# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X10 no_offsetLatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X11 a_6667_n4104# Vin1 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X12 VDD no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X13 no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X14 no_offsetLatch_0.Vp a_6163_n3233# a_6075_n3141# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X15 no_offsetLatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X16 a_6667_n4104# Vin2 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X17 a_6667_n4104# Vin1 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X18 a_9707_n4104# a_9507_n4196# no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
X19 Vout a_5265_2223# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X20 no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X21 VDD CLK no_offsetLatch_0.Vq VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X22 a_7745_n1756# a_7545_n1848# no_offsetLatch_0.Vout1 VSS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X23 a_5265_2223# x4.A VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X24 no_offsetLatch_0.Vq no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X25 x4.A x2.Vout2 VDD VDD pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X26 x4.A x3.out VSS VSS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X27 no_offsetLatch_0.Vq a_6163_n4196# a_6075_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X28 no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X29 a_6667_n4104# Vin2 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X30 a_6667_n4104# Vin2 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X31 Vout a_5265_2223# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X32 Vout a_5265_2223# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X33 no_offsetLatch_0.Vout1 CLK VDD VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X34 no_offsetLatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X35 no_offsetLatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X36 a_5265_2223# x4.A VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X37 VDD no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X38 no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X39 no_offsetLatch_0.Vp no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X40 a_6667_n4104# Vin1 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X41 Vout a_5265_2223# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X42 no_offsetLatch_0.Vq no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X43 a_9541_n1756# a_9341_n1848# no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X44 no_offsetLatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X45 VDD x4.A x2.Vout2 VDD pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X46 VSS x5.out x2.Vout2 VSS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X47 a_6667_n4104# Vin1 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X48 no_offsetLatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X49 no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X50 no_offsetLatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X51 x3.out no_offsetLatch_0.Vout1 VSS VSS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.4u
X52 no_offsetLatch_0.Vp a_6329_n1848# a_6241_n1756# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X53 a_6667_n4104# CLK VSS VSS nfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.4u
X54 a_8159_n4890# a_8079_n4982# a_6667_n4104# VSS nfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.4u
X55 VSS a_5265_2223# Vout VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X56 VSS no_offsetLatch_0.Vout2 x5.out VSS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.4u
X57 x3.out no_offsetLatch_0.Vout1 VDD VDD pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.4u
X58 VDD no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X59 no_offsetLatch_0.Vout2 no_offsetLatch_0.Vout1 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X60 a_6667_n4104# Vin2 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X61 a_6667_n4104# Vin2 no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X62 VSS a_5265_2223# Vout VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X63 no_offsetLatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X64 no_offsetLatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X65 no_offsetLatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X66 a_6667_n4104# Vin1 no_offsetLatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X67 VDD no_offsetLatch_0.Vout1 no_offsetLatch_0.Vout2 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X68 a_9707_n3141# a_9507_n3233# no_offsetLatch_0.Vq VSS nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
.ends

.subckt inv2 in vdd out vss
X0 out in vdd vdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X1 out in vss vss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
.ends

.subckt adc_PISO load B6 B5 B4 serial_out avdd B3 avss B2 B1 clk
X0 a_44488_8266# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X1 a_50206_2781# a_48650_3501# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X2 a_6600_2510# a_6520_1558# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X3 a_6520_1558# a_6520_3763# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X4 avdd dffrs_1.Q a_20234_3501# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X5 avdd a_6520_3763# 2inmux_2.Bit avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X6 a_2846_2780# a_1290_3500# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X7 dffrs_4.Qb avdd a_46158_3857# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X8 a_15992_3763# clk a_16256_6060# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X9 2inmux_1.Bit dffrs_4.Qb a_46158_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X10 a_10950_2780# 2inmux_2.Bit avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X11 a_15992_5968# a_15992_3763# a_16256_8265# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X12 a_39178_3501# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X13 avss dffrs_2.Q a_29894_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X14 a_50206_441# a_48650_1161# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X15 2inmux_1.OUT a_50878_1605# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X16 avdd a_6520_1558# dffrs_0.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X17 avss a_21790_2781# a_22462_1605# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X18 a_35016_1651# a_34936_1559# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X19 a_35016_3856# a_34936_3764# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X20 2inmux_0.OUT a_3518_1604# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X21 a_22462_1605# a_21790_441# a_22650_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X22 a_29000_1361# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X23 avss a_47944_1361# a_48838_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X24 avdd avdd a_44408_3764# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X25 a_21790_441# a_20234_1161# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X26 a_1478_2780# load a_1290_3500# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X27 avdd a_29000_1361# a_29706_1161# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X28 a_25464_3764# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X29 avdd avdd a_6600_2510# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X30 a_1478_440# B6 a_1290_1160# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X31 avdd a_25464_3764# dffrs_2.Q avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X32 a_35200_6061# avdd a_35016_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X33 avdd 2inmux_2.Bit a_10762_3500# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X34 a_1290_1160# B6 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X35 2inmux_2.Bit dffrs_0.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X36 avdd clk a_6520_1558# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X37 a_35200_8266# a_35016_2511# a_35016_8266# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X38 avss 2inmux_1.Bit a_48838_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X39 avss a_40734_2781# a_41406_1605# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X40 avdd a_44488_2511# a_44408_5969# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X41 avdd a_25464_1559# dffrs_2.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X42 a_31262_2781# a_29706_3501# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X43 a_47944_1361# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X44 a_39366_2781# dffrs_3.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X45 dffrs_0.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X46 avdd a_584_1360# a_1290_1160# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X47 2inmux_3.OUT a_22462_1605# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X48 a_51066_2325# a_50206_441# a_50878_1605# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X49 a_12990_1604# a_12318_440# a_13178_2324# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X50 a_25464_5969# a_25464_3764# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X51 a_44488_2511# a_44408_1559# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X52 avdd avdd a_15992_3763# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X53 a_44408_3764# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X54 a_44408_1559# a_44408_3764# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X55 a_20422_2781# load a_20234_3501# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X56 avdd a_44408_3764# 2inmux_1.Bit avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X57 a_54144_6061# avdd a_53960_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X58 a_55630_3857# a_53880_1559# a_55446_3857# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X59 a_54144_8266# a_53960_2511# a_53960_8266# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X60 avdd a_15992_3763# dffrs_1.Q avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X61 a_25544_6061# a_25464_5969# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X62 a_27030_3857# dffrs_2.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X63 a_25544_8266# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X64 dffrs_2.Q dffrs_2.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X65 a_55630_6061# a_53880_3764# a_55446_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X66 a_3518_1604# a_2846_440# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X67 a_27030_6061# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X68 a_34936_3764# clk a_35200_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X69 a_31262_2781# a_29706_3501# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X70 avdd dffrs_3.Q a_39178_3501# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X71 a_16072_2510# 2inmux_2.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X72 a_34936_5969# a_34936_3764# a_35200_8266# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X73 avdd a_44408_1559# dffrs_4.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X74 a_15992_1558# a_16072_2510# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X75 a_39366_441# a_38472_1361# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X76 a_21790_441# a_20234_1161# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X77 a_1290_1160# B6 a_1478_440# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X78 a_44408_5969# a_44408_3764# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X79 avdd a_15992_1558# dffrs_1.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X80 dffrs_2.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X81 avss a_12318_2780# a_12990_1604# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X82 avdd a_16072_2510# a_15992_5968# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X83 a_53880_3764# a_53880_5969# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X84 a_2846_440# a_1290_1160# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X85 a_44672_1651# avdd a_44488_1651# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X86 2inmux_4.OUT a_31934_1605# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X87 a_44672_3856# clk a_44488_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X88 dffrs_3.Q avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X89 a_45974_3857# 2inmux_1.Bit avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X90 a_10950_2780# load a_10762_3500# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X91 a_25544_2511# 2inmux_3.OUT a_25728_1651# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X92 a_1478_440# a_584_1360# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X93 a_16072_6060# a_15992_5968# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X94 a_25464_1559# a_25544_2511# a_25728_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X95 a_25728_6061# avdd a_25544_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X96 a_45974_6061# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X97 a_53880_3764# clk a_54144_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X98 dffrs_5.Qb avdd a_55630_3857# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X99 a_10762_1160# B5 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X100 a_19528_1361# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X101 a_39366_2781# load a_39178_3501# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X102 avdd avdd a_35016_2511# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X103 a_16072_8265# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X104 a_25728_8266# a_25544_2511# a_25544_8266# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X105 a_53880_5969# a_53880_3764# a_54144_8266# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X106 dffrs_1.Q dffrs_1.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X107 a_6520_3763# clk a_6784_6060# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X108 avdd clk a_34936_1559# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X109 avdd a_12318_2780# a_13178_2324# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X110 a_22462_1605# a_21790_441# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X111 a_53880_5969# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X112 a_6520_5968# a_6520_3763# a_6784_8265# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X113 serial_out dffrs_5.Qb a_55630_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X114 dffrs_3.Qb dffrs_3.Q avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X115 avss a_38472_1361# a_39366_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X116 a_39366_441# B2 a_39178_1161# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X117 dffrs_1.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X118 serial_out avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X119 a_16256_1650# avdd a_16072_1650# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X120 a_44488_2511# 2inmux_5.OUT a_44672_1651# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X121 a_6520_3763# a_6520_5968# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X122 a_16256_3855# clk a_16072_3855# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X123 a_44408_1559# a_44488_2511# a_44672_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X124 avss a_584_1360# a_1478_440# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X125 a_17558_3856# dffrs_1.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X126 avdd avdd a_53960_2511# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X127 a_48650_3501# load a_48838_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X128 a_41406_1605# a_40734_441# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X129 avdd a_34936_3764# dffrs_3.Q avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X130 avdd clk a_53880_1559# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X131 a_25544_2511# a_25464_1559# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X132 a_25464_1559# a_25464_3764# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X133 dffrs_5.Qb serial_out avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X134 a_12990_1604# a_12318_440# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X135 2inmux_1.OUT a_50878_1605# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X136 a_17558_6060# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X137 avss avss a_1478_2780# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X138 a_22650_2325# a_21790_2781# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X139 a_35016_2511# 2inmux_4.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X140 a_34936_1559# a_35016_2511# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X141 2inmux_0.OUT a_3518_1604# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X142 avss a_50206_2781# a_50878_1605# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X143 a_40734_2781# a_39178_3501# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X144 avdd a_34936_1559# dffrs_3.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X145 a_20422_441# B4 a_20234_1161# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X146 a_48838_2781# 2inmux_1.Bit avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X147 a_6520_5968# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X148 a_53960_1651# a_53880_1559# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X149 a_53960_3856# a_53880_3764# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X150 a_12318_440# a_10762_1160# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X151 a_41406_1605# a_40734_441# a_41594_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X152 a_48650_3501# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X153 a_29706_3501# load a_29894_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X154 avdd avdd a_6520_3763# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X155 a_35016_6061# a_34936_5969# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X156 2inmux_2.Bit avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X157 a_16072_2510# a_15992_1558# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X158 a_10056_1360# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X159 a_53960_2511# 2inmux_1.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X160 a_35016_8266# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X161 a_15992_1558# a_15992_3763# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X162 a_40734_2781# a_39178_3501# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X163 avdd avdd a_25544_2511# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X164 a_41594_2325# a_40734_2781# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X165 avdd a_31262_2781# a_32122_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X166 avdd clk a_25464_1559# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X167 a_53880_1559# a_53960_2511# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X168 avdd 2inmux_1.Bit a_48650_3501# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X169 a_6600_2510# 2inmux_0.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X170 a_584_1360# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X171 a_6520_1558# a_6600_2510# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X172 dffrs_3.Qb avdd a_36686_3857# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X173 avss dffrs_1.Q a_20422_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X174 2inmux_3.OUT a_22462_1605# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X175 a_20234_1161# B4 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X176 dffrs_0.Qb 2inmux_2.Bit avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X177 a_20234_1161# B4 a_20422_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X178 dffrs_3.Q dffrs_3.Qb a_36686_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X179 a_12318_2780# a_10762_3500# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X180 avdd a_6600_2510# a_6520_5968# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X181 a_29706_3501# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X182 avss a_2846_2780# a_3518_1604# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X183 2inmux_5.OUT a_41406_1605# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X184 a_44408_3764# a_44408_5969# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X185 a_6600_1650# a_6520_1558# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X186 a_50206_441# a_48650_1161# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X187 a_2846_440# a_1290_1160# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X188 avdd a_19528_1361# a_20234_1161# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X189 a_6600_3855# a_6520_3763# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X190 a_3706_2324# a_2846_440# a_3518_1604# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X191 avss a_10056_1360# a_10950_440# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X192 a_39178_1161# B2 a_39366_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X193 a_20422_441# a_19528_1361# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X194 a_10950_440# B5 a_10762_1160# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X195 a_31934_1605# a_31262_441# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X196 a_15992_3763# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X197 2inmux_1.Bit dffrs_4.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X198 avdd a_2846_2780# a_3706_2324# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X199 a_40734_441# a_39178_1161# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X200 a_39178_1161# B2 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X201 a_8270_3856# a_6520_1558# a_8086_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X202 a_12318_2780# a_10762_3500# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X203 a_13178_2324# a_12318_2780# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X204 a_44408_5969# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X205 a_8270_6060# a_6520_3763# a_8086_6060# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X206 2inmux_4.OUT a_31934_1605# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X207 dffrs_4.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X208 a_21790_2781# a_20234_3501# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X209 a_29894_2781# dffrs_2.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X210 avdd a_10056_1360# a_10762_1160# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X211 2inmux_2.OUT a_12990_1604# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X212 a_31934_1605# a_31262_441# a_32122_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X213 a_15992_5968# a_15992_3763# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X214 a_6784_1650# avdd a_6600_1650# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X215 a_19528_1361# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X216 a_22650_2325# a_21790_441# a_22462_1605# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X217 a_6784_3855# clk a_6600_3855# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X218 a_1290_3500# load a_1478_2780# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X219 a_35016_2511# a_34936_1559# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X220 avdd avdd a_34936_3764# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X221 a_34936_1559# a_34936_3764# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X222 a_44672_6061# avdd a_44488_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X223 a_38472_1361# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X224 a_44672_8266# a_44488_2511# a_44488_8266# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X225 dffrs_0.Qb avdd a_8270_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X226 a_27214_3857# a_25464_1559# a_27030_3857# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X227 a_1478_2780# avss avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X228 avss a_19528_1361# a_20422_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X229 a_25464_3764# clk a_25728_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X230 a_21790_2781# a_20234_3501# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X231 avdd dffrs_2.Q a_29706_3501# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X232 a_25464_5969# a_25464_3764# a_25728_8266# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X233 a_27214_6061# a_25464_3764# a_27030_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X234 a_10762_1160# B5 a_10950_440# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X235 a_10950_440# a_10056_1360# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X236 2inmux_2.Bit dffrs_0.Qb a_8270_6060# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X237 a_50878_1605# a_50206_441# a_51066_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X238 a_44488_1651# a_44408_1559# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X239 avss a_31262_2781# a_31934_1605# avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X240 avdd a_35016_2511# a_34936_5969# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X241 a_1290_3500# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X242 a_44488_3856# a_44408_3764# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X243 a_41594_2325# a_40734_441# a_41406_1605# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X244 avdd avdd a_53880_3764# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X245 a_25464_3764# a_25464_5969# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X246 a_13178_2324# a_12318_440# a_12990_1604# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X247 a_29894_2781# load a_29706_3501# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X248 a_31262_441# a_29706_1161# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X249 avdd a_38472_1361# a_39178_1161# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X250 dffrs_2.Q avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X251 a_34936_3764# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X252 avdd a_53880_3764# serial_out avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X253 a_46158_3857# a_44408_1559# a_45974_3857# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X254 a_16072_2510# 2inmux_2.OUT a_16256_1650# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X255 a_51066_2325# a_50206_2781# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X256 avdd avss a_1290_3500# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X257 a_15992_1558# a_16072_2510# a_16256_3855# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X258 a_29894_441# a_29000_1361# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X259 a_16256_6060# avdd a_16072_6060# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X260 a_44408_3764# clk a_44672_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X261 a_17742_3856# a_15992_1558# a_17558_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X262 a_16256_8265# a_16072_2510# a_16072_8265# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X263 a_44408_5969# a_44408_3764# a_44672_8266# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X264 a_46158_6061# a_44408_3764# a_45974_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X265 dffrs_2.Qb avdd a_27214_3857# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X266 a_17742_6060# a_15992_3763# a_17558_6060# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X267 dffrs_2.Qb dffrs_2.Q avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X268 avdd a_53880_1559# dffrs_5.Qb avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X269 avdd a_53960_2511# a_53880_5969# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X270 dffrs_2.Q dffrs_2.Qb a_27214_6061# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X271 a_25464_5969# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X272 a_10056_1360# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X273 a_34936_5969# a_34936_3764# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X274 a_31262_441# a_29706_1161# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X275 a_15992_3763# a_15992_5968# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X276 avdd avdd a_25464_3764# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X277 2inmux_1.Bit avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X278 a_53880_3764# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X279 a_584_1360# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X280 a_10762_3500# load a_10950_2780# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X281 a_35200_1651# avdd a_35016_1651# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X282 a_6520_3763# clk avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X283 a_53960_6061# a_53880_5969# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X284 a_35200_3856# clk a_35016_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X285 a_53960_8266# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X286 serial_out dffrs_5.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X287 a_36502_3857# dffrs_3.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X288 avdd a_50206_2781# a_51066_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X289 avdd avdd a_44488_2511# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X290 a_29000_1361# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X291 avdd clk a_44408_1559# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X292 a_3706_2324# a_2846_2780# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X293 a_36502_6061# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X294 dffrs_4.Qb 2inmux_1.Bit avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X295 dffrs_1.Qb avdd a_17742_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X296 a_25544_2511# 2inmux_3.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X297 2inmux_5.OUT a_41406_1605# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X298 a_25464_1559# a_25544_2511# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X299 dffrs_5.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X300 a_15992_5968# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X301 a_53880_5969# a_53880_3764# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X302 dffrs_1.Q dffrs_1.Qb a_17742_6060# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X303 avss a_29000_1361# a_29894_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X304 avdd a_25544_2511# a_25464_5969# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X305 a_10762_3500# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X306 a_54144_1651# avdd a_53960_1651# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X307 a_6520_5968# a_6520_3763# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X308 a_25544_1651# a_25464_1559# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X309 a_32122_2325# a_31262_441# a_31934_1605# avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X310 a_25544_3856# a_25464_3764# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X311 a_54144_3856# clk a_53960_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X312 a_55446_3857# serial_out avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X313 a_48838_441# B1 a_48650_1161# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X314 a_47944_1361# load avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X315 a_35016_2511# 2inmux_4.OUT a_35200_1651# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X316 dffrs_1.Q avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X317 a_34936_1559# a_35016_2511# a_35200_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X318 a_50878_1605# a_50206_441# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X319 a_6600_6060# a_6520_5968# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X320 a_55446_6061# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X321 a_36686_3857# a_34936_1559# a_36502_3857# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X322 a_48838_2781# load a_48650_3501# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X323 a_44488_2511# 2inmux_5.OUT avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X324 avdd avdd a_16072_2510# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X325 avdd a_21790_2781# a_22650_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X326 a_6600_8265# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X327 a_36686_6061# a_34936_3764# a_36502_6061# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X328 avdd clk a_15992_1558# avdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X329 a_44408_1559# a_44488_2511# avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X330 dffrs_1.Qb dffrs_1.Q avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X331 avss 2inmux_2.Bit a_10950_2780# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X332 2inmux_2.OUT a_12990_1604# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X333 a_48650_1161# B1 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X334 avss dffrs_3.Q a_39366_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X335 a_16072_1650# a_15992_1558# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X336 a_34936_3764# a_34936_5969# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X337 a_25728_1651# avdd a_25544_1651# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X338 a_29894_441# B3 a_29706_1161# avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X339 a_53960_2511# 2inmux_1.OUT a_54144_1651# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X340 a_40734_441# a_39178_1161# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X341 a_38472_1361# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X342 a_16072_3855# a_15992_3763# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X343 a_53880_1559# a_53960_2511# a_54144_3856# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X344 a_6600_2510# 2inmux_0.OUT a_6784_1650# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X345 avdd a_47944_1361# a_48650_1161# avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X346 a_53960_2511# a_53880_1559# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X347 a_53880_1559# a_53880_3764# avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X348 a_25728_3856# clk a_25544_3856# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X349 a_20234_3501# load a_20422_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X350 a_6520_1558# a_6600_2510# a_6784_3855# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X351 a_8086_3856# 2inmux_2.Bit avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X352 avdd a_40734_2781# a_41594_2325# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X353 dffrs_3.Q dffrs_3.Qb avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X354 a_6784_6060# avdd a_6600_6060# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X355 a_29706_1161# B3 avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X356 a_32122_2325# a_31262_2781# avdd avdd pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X357 a_6784_8265# a_6600_2510# a_6600_8265# avss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X358 a_8086_6060# avdd avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X359 a_48650_1161# B1 a_48838_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X360 a_50206_2781# a_48650_3501# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X361 a_34936_5969# avdd avdd avdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X362 a_20422_2781# dffrs_1.Q avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X363 a_2846_2780# a_1290_3500# avss avss nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.5u
X364 dffrs_3.Qb avdd avdd avdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X365 a_29706_1161# B3 a_29894_441# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X366 a_20234_3501# load avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X367 a_3518_1604# a_2846_440# a_3706_2324# avdd pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X368 a_48838_441# a_47944_1361# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X369 a_39178_3501# load a_39366_2781# avss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X370 a_12318_440# a_10762_1160# avdd avdd pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
X371 a_44488_6061# a_44408_5969# avss avss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
.ends

.subckt SARlogic vdd vss clk reset comp_in d5 d4 d3 d2 d1 d0
X0 dffrs_5.Qb reset a_26858_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X1 a_1150_7058# dffrs_13.nand3_8.Z a_966_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X2 vdd dffrs_12.nand3_8.Z dffrs_12.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X3 dffrs_5.nand3_1.C dffrs_5.nand3_6.C a_25372_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X4 a_14732_12225# dffrs_8.nand3_8.C a_14548_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X5 dffrs_10.nand3_8.C dffrs_10.nand3_8.Z a_21330_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X6 vdd dffrs_12.Q dffrs_11.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X7 a_9020_4853# dffrs_1.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X8 d2 dffrs_2.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X9 a_18774_14429# dffrs_9.nand3_6.C a_18590_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X10 dffrs_10.nand3_6.C d0 a_21330_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X11 a_22632_14429# dffrs_3.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X12 vdd reset dffrs_11.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X13 dffrs_4.nand3_6.C clk a_21330_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X14 a_13246_16634# dffrs_8.nand3_8.Z a_13062_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X15 a_13062_16634# dffrs_1.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X16 dffrs_12.nand3_8.C dffrs_12.nand3_8.Z a_29414_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X17 a_6648_14432# dffrs_14.nand3_6.C a_6464_14432# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X18 dffrs_13.nand3_6.C clk a_1150_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X19 dffrs_12.nand3_6.C vss a_29414_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X20 dffrs_4.Q dffrs_4.Qb a_22816_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X21 a_25188_16634# dffrs_4.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X22 dffrs_11.nand3_8.Z comp_in a_25372_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X23 a_21146_12224# dffrs_10.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X24 dffrs_7.nand3_8.C dffrs_7.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X25 dffrs_0.d dffrs_13.Qb a_2636_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X26 dffrs_9.nand3_8.C dffrs_9.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X27 vdd dffrs_0.nand3_6.C dffrs_0.Q vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X28 dffrs_7.nand3_6.C d3 vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X29 dffrs_9.nand3_6.C dffrs_9.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X30 a_21146_14429# dffrs_10.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X31 dffrs_5.Q vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X32 dffrs_2.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X33 dffrs_1.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X34 a_966_443# dffrs_13.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X35 a_6648_12228# dffrs_14.nand3_8.C a_6464_12228# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X36 dffrs_0.nand3_8.Z dffrs_0.d vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X37 dffrs_2.nand3_1.C dffrs_2.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X38 dffrs_4.Qb reset a_22816_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X39 vdd reset dffrs_3.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X40 dffrs_1.nand3_1.C dffrs_1.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X41 vdd reset dffrs_5.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X42 a_4978_14432# dffrs_14.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X43 a_9020_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X44 dffrs_0.nand3_8.C dffrs_0.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X45 a_17288_10019# reset a_17104_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X46 dffrs_13.Qb vdd a_2636_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X47 vdd clk dffrs_3.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X48 a_4978_4853# dffrs_0.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X49 dffrs_10.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X50 dffrs_12.Q dffrs_12.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X51 vdd clk dffrs_5.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X52 dffrs_4.nand3_1.C dffrs_4.nand3_6.C a_21330_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X53 a_4978_16637# dffrs_13.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X54 vdd dffrs_0.nand3_8.C dffrs_0.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X55 vdd dffrs_12.nand3_6.C dffrs_12.Q vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X56 dffrs_5.nand3_8.Z dffrs_4.Q a_25372_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X57 d0 dffrs_11.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X58 dffrs_5.Qb dffrs_5.Q vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X59 dffrs_13.nand3_1.C dffrs_13.nand3_6.C a_1150_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X60 dffrs_10.nand3_1.C dffrs_10.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X61 a_21330_443# reset a_21146_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X62 vdd dffrs_7.nand3_6.C d4 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X63 d4 dffrs_7.Qb a_10690_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X64 a_9020_443# dffrs_1.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X65 dffrs_1.nand3_8.Z dffrs_0.Q a_9204_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X66 dffrs_12.nand3_1.C dffrs_12.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X67 dffrs_4.nand3_6.C dffrs_4.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X68 dffrs_8.Qb reset a_14732_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X69 dffrs_10.Qb d1 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X70 vdd reset dffrs_8.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X71 dffrs_11.nand3_8.C dffrs_11.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X72 vdd dffrs_9.nand3_8.C dffrs_9.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X73 dffrs_4.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X74 dffrs_8.nand3_8.Z dffrs_8.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X75 d0 dffrs_4.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X76 d2 dffrs_9.Qb a_18774_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X77 a_22816_14429# dffrs_10.nand3_6.C a_22632_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X78 dffrs_11.nand3_6.C dffrs_12.Q vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X79 a_18774_4853# dffrs_3.nand3_6.C a_18590_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X80 a_29230_16634# dffrs_5.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X81 dffrs_4.Q vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X82 dffrs_10.nand3_1.C dffrs_3.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X83 a_25188_443# dffrs_5.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X84 dffrs_11.nand3_8.Z dffrs_11.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X85 a_9204_2648# clk a_9020_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X86 dffrs_2.d dffrs_1.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X87 dffrs_0.d reset vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X88 a_4978_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X89 vdd reset dffrs_4.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X90 vdd dffrs_5.nand3_6.C dffrs_5.Q vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X91 dffrs_13.nand3_6.C dffrs_13.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X92 dffrs_3.nand3_8.C dffrs_3.nand3_8.Z a_17288_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X93 vdd vdd dffrs_13.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X94 a_14548_12225# d3 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X95 vdd d1 dffrs_9.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X96 vdd clk dffrs_4.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X97 a_18774_2649# dffrs_3.nand3_8.C a_18590_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X98 dffrs_13.nand3_1.C reset vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X99 dffrs_5.nand3_8.Z dffrs_4.Q vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X100 vdd reset dffrs_9.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X101 dffrs_4.Qb dffrs_4.Q vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X102 vdd clk dffrs_13.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X103 dffrs_5.nand3_8.C dffrs_5.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X104 dffrs_13.Qb dffrs_0.d vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X105 a_9204_12224# d3 a_9020_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X106 dffrs_1.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X107 a_9020_12224# dffrs_7.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X108 vdd dffrs_5.nand3_8.C dffrs_5.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X109 a_9204_14429# reset a_9020_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X110 a_13246_4853# reset a_13062_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X111 a_9020_14429# dffrs_7.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X112 a_14732_4853# dffrs_2.nand3_6.C a_14548_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X113 dffrs_7.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X114 dffrs_4.d dffrs_3.Qb a_18774_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X115 dffrs_9.nand3_1.C dffrs_9.nand3_6.C a_17288_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X116 a_21330_16634# dffrs_10.nand3_8.Z a_21146_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X117 vdd dffrs_4.nand3_6.C dffrs_4.Q vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X118 vdd reset dffrs_14.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X119 dffrs_2.nand3_8.C dffrs_2.nand3_8.Z a_13246_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X120 vdd dffrs_10.nand3_8.C dffrs_10.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X121 dffrs_9.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X122 dffrs_1.nand3_8.C dffrs_1.nand3_8.Z a_9204_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X123 dffrs_12.nand3_8.Z dffrs_12.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X124 dffrs_1.nand3_8.Z dffrs_1.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X125 vdd dffrs_13.nand3_6.C dffrs_0.d vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X126 a_14732_2649# dffrs_2.nand3_8.C a_14548_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X127 vdd dffrs_11.nand3_6.C d0 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X128 dffrs_12.Q dffrs_5.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X129 dffrs_4.nand3_8.Z dffrs_4.d vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X130 a_29414_16634# dffrs_12.nand3_8.Z a_29230_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X131 dffrs_1.nand3_8.C dffrs_1.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X132 dffrs_4.nand3_8.C dffrs_4.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X133 dffrs_13.nand3_8.Z vss vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X134 a_13246_7058# dffrs_2.nand3_8.Z a_13062_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X135 a_25372_12224# dffrs_12.Q a_25188_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X136 dffrs_3.Qb reset a_18774_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X137 d4 dffrs_0.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X138 a_18590_14429# dffrs_2.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X139 vdd dffrs_4.nand3_8.C dffrs_4.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X140 a_25372_14429# reset a_25188_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X141 dffrs_13.nand3_8.C dffrs_13.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X142 vdd dffrs_7.nand3_8.Z dffrs_7.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X143 dffrs_8.nand3_8.Z comp_in a_13246_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X144 dffrs_7.nand3_1.C dffrs_0.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X145 vdd dffrs_13.nand3_8.C dffrs_13.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X146 a_25188_4853# dffrs_5.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X147 a_10690_4853# dffrs_1.nand3_6.C a_10506_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X148 a_21146_2648# dffrs_4.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X149 a_17104_12224# dffrs_9.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X150 dffrs_7.nand3_8.C dffrs_7.nand3_8.Z a_9204_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X151 vdd d4 dffrs_14.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X152 dffrs_2.nand3_6.C dffrs_2.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X153 dffrs_7.nand3_6.C d3 a_9204_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X154 a_17104_14429# dffrs_9.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X155 dffrs_2.Q dffrs_2.Qb a_14732_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X156 dffrs_0.nand3_8.Z dffrs_0.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X157 dffrs_2.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X158 vdd reset dffrs_0.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X159 dffrs_3.nand3_6.C dffrs_3.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X160 dffrs_0.nand3_8.C dffrs_0.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X161 a_10690_2649# dffrs_1.nand3_8.C a_10506_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X162 vdd dffrs_0.nand3_8.Z dffrs_0.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X163 dffrs_3.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X164 dffrs_10.Qb reset a_22816_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X165 a_966_2648# dffrs_13.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X166 vdd reset dffrs_10.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X167 dffrs_9.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X168 dffrs_4.d vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X169 dffrs_12.Q dffrs_12.Qb a_30900_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X170 d0 dffrs_11.Qb a_26858_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X171 dffrs_2.Qb reset a_14732_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X172 a_25188_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X173 a_30900_14429# dffrs_12.nand3_6.C a_30716_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X174 vdd dffrs_11.nand3_8.Z dffrs_11.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X175 dffrs_10.nand3_1.C dffrs_10.nand3_6.C a_21330_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X176 dffrs_14.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X177 dffrs_8.nand3_8.C dffrs_8.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X178 vdd reset dffrs_12.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X179 a_10690_14429# dffrs_7.nand3_6.C a_10506_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X180 dffrs_8.nand3_6.C d2 vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X181 dffrs_12.nand3_1.C dffrs_12.nand3_6.C a_29414_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X182 dffrs_3.Qb dffrs_4.d vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X183 a_22632_12225# d1 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X184 a_18774_12225# dffrs_9.nand3_8.C a_18590_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X185 dffrs_9.Qb d2 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X186 dffrs_11.nand3_8.C dffrs_11.nand3_8.Z a_25372_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X187 dffrs_11.nand3_6.C dffrs_12.Q a_25372_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X188 a_26674_14429# dffrs_4.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X189 dffrs_7.nand3_1.C dffrs_7.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X190 a_21146_16634# dffrs_3.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X191 dffrs_13.nand3_8.Z vss a_1150_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X192 dffrs_9.nand3_1.C dffrs_2.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X193 dffrs_2.Q vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X194 dffrs_0.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X195 a_17288_12224# d1 a_17104_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X196 dffrs_14.nand3_8.C dffrs_14.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X197 vdd reset dffrs_3.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X198 vdd reset dffrs_5.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X199 vdd reset dffrs_2.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X200 dffrs_0.nand3_1.C dffrs_0.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X201 a_17288_14429# reset a_17104_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X202 vdd dffrs_3.nand3_8.Z dffrs_3.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X203 vdd dffrs_5.nand3_8.Z dffrs_5.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X204 a_13246_10019# reset a_13062_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X205 dffrs_0.Q dffrs_0.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X206 vdd clk dffrs_2.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X207 a_13062_10019# dffrs_8.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X208 dffrs_2.nand3_8.Z dffrs_2.d a_13246_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X209 dffrs_2.Qb dffrs_2.Q vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X210 dffrs_12.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X211 a_25188_10019# dffrs_11.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X212 vdd dffrs_12.nand3_8.C dffrs_12.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X213 dffrs_10.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X214 dffrs_11.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X215 dffrs_11.nand3_1.C dffrs_11.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X216 dffrs_0.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X217 a_6464_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X218 vdd dffrs_7.nand3_8.C dffrs_7.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X219 dffrs_7.Qb reset a_10690_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X220 a_17288_443# reset a_17104_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X221 dffrs_12.nand3_8.Z vss vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X222 a_13062_443# dffrs_2.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X223 a_9204_4853# reset a_9020_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X224 vdd dffrs_8.nand3_6.C d3 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X225 a_13062_2648# dffrs_2.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X226 dffrs_2.d vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X227 a_22816_12225# dffrs_10.nand3_8.C a_22632_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X228 dffrs_9.Qb reset a_18774_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X229 dffrs_11.Qb d0 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X230 dffrs_3.nand3_6.C clk a_17288_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X231 dffrs_10.nand3_8.Z dffrs_10.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X232 a_5162_2648# clk a_4978_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X233 a_25372_443# reset a_25188_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X234 vdd reset dffrs_4.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X235 a_17104_2648# dffrs_3.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X236 a_26858_14429# dffrs_11.nand3_6.C a_26674_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X237 a_30716_14429# dffrs_5.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X238 a_6464_2649# dffrs_0.Q vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X239 vdd vdd dffrs_13.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X240 vdd dffrs_9.nand3_8.Z dffrs_9.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X241 vdd dffrs_4.nand3_8.Z dffrs_4.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X242 dffrs_5.nand3_8.Z dffrs_5.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X243 dffrs_14.nand3_8.Z dffrs_14.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X244 vdd d2 dffrs_8.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X245 dffrs_5.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X246 vdd dffrs_13.nand3_8.Z dffrs_13.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X247 dffrs_8.nand3_8.C dffrs_8.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X248 a_10506_14429# dffrs_0.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X249 dffrs_5.nand3_8.C dffrs_5.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X250 dffrs_1.Qb dffrs_2.d vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X251 vdd reset dffrs_8.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X252 a_9204_443# reset a_9020_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X253 a_9204_16634# dffrs_7.nand3_8.Z a_9020_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X254 dffrs_5.nand3_1.C dffrs_5.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X255 dffrs_8.nand3_6.C dffrs_8.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X256 dffrs_0.nand3_8.Z dffrs_0.d a_5162_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X257 a_9020_16634# dffrs_0.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X258 dffrs_11.nand3_8.C dffrs_11.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X259 dffrs_5.Q dffrs_5.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X260 a_5162_10022# reset a_4978_10022# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X261 dffrs_11.nand3_6.C dffrs_11.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X262 a_9204_7058# dffrs_1.nand3_8.Z a_9020_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X263 a_29230_10019# dffrs_12.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X264 a_5162_12227# d4 a_4978_12227# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X265 a_21146_443# dffrs_4.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X266 dffrs_3.nand3_1.C dffrs_3.nand3_6.C a_17288_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X267 a_6648_4853# dffrs_0.nand3_6.C a_6464_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X268 dffrs_5.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X269 a_4978_443# dffrs_0.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X270 a_26674_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X271 dffrs_2.nand3_6.C clk a_13246_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X272 dffrs_1.nand3_6.C clk a_9204_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X273 dffrs_14.nand3_8.C dffrs_14.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X274 dffrs_1.nand3_6.C dffrs_1.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X275 dffrs_0.nand3_8.C dffrs_0.nand3_8.Z a_5162_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X276 dffrs_4.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X277 a_17288_2648# clk a_17104_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X278 d3 dffrs_8.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X279 a_25372_2648# clk a_25188_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X280 dffrs_1.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X281 a_6648_2649# dffrs_0.nand3_8.C a_6464_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X282 a_25372_16634# dffrs_11.nand3_8.Z a_25188_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X283 dffrs_13.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X284 dffrs_4.nand3_1.C dffrs_4.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X285 a_26674_2649# dffrs_5.Q vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X286 dffrs_8.nand3_8.C dffrs_8.nand3_8.Z a_13246_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X287 dffrs_12.Qb dffrs_12.Q vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X288 vdd dffrs_11.nand3_8.C dffrs_11.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X289 dffrs_4.Q dffrs_4.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X290 dffrs_13.nand3_1.C dffrs_13.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X291 dffrs_8.nand3_6.C d2 a_13246_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X292 dffrs_0.d dffrs_13.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X293 a_18590_12225# d2 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X294 dffrs_7.Qb d4 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X295 vdd reset dffrs_7.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X296 dffrs_12.nand3_8.C dffrs_12.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X297 a_21146_4853# dffrs_4.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X298 vdd reset dffrs_14.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X299 dffrs_7.nand3_8.Z dffrs_7.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X300 d3 dffrs_1.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X301 dffrs_2.nand3_1.C dffrs_2.nand3_6.C a_13246_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X302 dffrs_12.nand3_6.C dffrs_12.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X303 dffrs_1.nand3_1.C dffrs_1.nand3_6.C a_9204_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X304 dffrs_7.nand3_1.C dffrs_7.nand3_6.C a_9204_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X305 a_17104_16634# dffrs_2.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X306 a_21330_10019# reset a_21146_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X307 vdd dffrs_14.nand3_8.Z dffrs_14.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X308 dffrs_9.nand3_8.Z comp_in a_17288_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X309 dffrs_4.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X310 a_22632_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X311 dffrs_13.Qb vdd vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X312 dffrs_0.nand3_6.C dffrs_0.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X313 dffrs_14.nand3_8.Z comp_in a_5162_10022# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X314 a_2452_4853# reset vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X315 dffrs_2.d dffrs_1.Qb a_10690_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X316 a_29414_10019# reset a_29230_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X317 a_26858_4853# dffrs_5.nand3_6.C a_26674_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X318 dffrs_0.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X319 dffrs_14.nand3_8.C dffrs_14.nand3_8.Z a_5162_12227# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X320 a_966_4853# dffrs_13.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X321 a_21330_2648# clk a_21146_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X322 a_22632_2649# dffrs_4.Q vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X323 a_1150_2648# clk a_966_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X324 a_2452_2649# dffrs_0.d vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X325 dffrs_1.Qb reset a_10690_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X326 dffrs_5.nand3_8.C dffrs_5.nand3_8.Z a_25372_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X327 a_21146_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X328 dffrs_12.Qb reset a_30900_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X329 dffrs_8.nand3_1.C dffrs_8.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X330 a_26858_2649# dffrs_5.nand3_8.C a_26674_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X331 a_30900_12225# dffrs_12.nand3_8.C a_30716_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X332 dffrs_11.Qb reset a_26858_12225# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X333 vdd reset dffrs_11.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X334 d5 dffrs_14.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X335 vdd reset dffrs_1.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X336 vdd dffrs_3.nand3_6.C dffrs_4.d vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X337 vdd clk dffrs_1.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X338 dffrs_11.nand3_1.C dffrs_11.nand3_6.C a_25372_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X339 a_10690_12225# dffrs_7.nand3_8.C a_10506_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X340 dffrs_3.nand3_8.Z dffrs_2.Q vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X341 vdd d0 dffrs_10.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X342 dffrs_9.nand3_8.C dffrs_9.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X343 a_14732_14429# dffrs_8.nand3_6.C a_14548_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X344 dffrs_9.nand3_6.C d1 vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X345 vdd reset dffrs_10.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X346 dffrs_3.nand3_8.C dffrs_3.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X347 a_966_7058# reset vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X348 vdd dffrs_3.nand3_8.C dffrs_3.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X349 a_26674_12225# d0 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X350 dffrs_14.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X351 a_22816_4853# dffrs_4.nand3_6.C a_22632_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X352 dffrs_9.nand3_8.Z dffrs_9.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X353 dffrs_7.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X354 vdd vss dffrs_12.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X355 d5 dffrs_13.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X356 dffrs_14.nand3_6.C d4 vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X357 vdd reset dffrs_12.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X358 a_2636_4853# dffrs_13.nand3_6.C a_2452_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X359 dffrs_14.nand3_1.C dffrs_14.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X360 a_17288_16634# dffrs_9.nand3_8.Z a_17104_16634# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X361 dffrs_10.nand3_8.Z comp_in a_21330_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X362 a_13246_12224# d2 a_13062_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X363 a_9020_2648# dffrs_1.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X364 vdd reset dffrs_2.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X365 a_13062_12224# dffrs_8.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X366 a_13246_14429# reset a_13062_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X367 dffrs_4.nand3_8.C dffrs_4.nand3_8.Z a_21330_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X368 vdd dffrs_2.nand3_8.Z dffrs_2.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X369 a_13062_14429# dffrs_8.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X370 dffrs_12.nand3_8.Z vss a_29414_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X371 dffrs_13.nand3_8.C dffrs_13.nand3_8.Z a_1150_2648# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X372 a_22816_2649# dffrs_4.nand3_8.C a_22632_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X373 a_25188_12224# dffrs_11.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X374 dffrs_14.Qb d5 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X375 dffrs_4.nand3_8.Z dffrs_4.d a_21330_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X376 vdd dffrs_2.nand3_6.C dffrs_2.Q vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X377 a_2636_2649# dffrs_13.nand3_8.C a_2452_2649# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X378 a_25188_14429# dffrs_11.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X379 a_1150_443# vdd a_966_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X380 a_21146_10019# dffrs_10.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X381 dffrs_2.nand3_8.Z dffrs_2.d vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X382 dffrs_1.nand3_8.Z dffrs_0.Q vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X383 dffrs_4.d dffrs_3.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X384 d1 dffrs_10.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X385 dffrs_2.nand3_8.C dffrs_2.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X386 dffrs_1.nand3_8.C dffrs_1.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X387 a_13062_4853# dffrs_2.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X388 a_4978_10022# dffrs_14.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X389 vdd dffrs_2.nand3_8.C dffrs_2.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X390 dffrs_11.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X391 a_5162_4853# reset a_4978_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X392 a_4978_12227# dffrs_14.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X393 dffrs_3.nand3_8.Z dffrs_2.Q a_17288_443# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X394 a_17104_4853# dffrs_3.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X395 a_4978_2648# dffrs_0.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X396 dffrs_3.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X397 dffrs_10.nand3_8.C dffrs_10.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X398 vdd dffrs_8.nand3_8.C dffrs_8.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X399 d1 dffrs_3.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X400 d3 dffrs_8.Qb a_14732_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X401 vdd dffrs_9.nand3_6.C d2 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X402 dffrs_10.nand3_6.C d0 vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X403 a_18590_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X404 dffrs_5.nand3_6.C dffrs_5.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X405 vdd dffrs_8.nand3_8.Z dffrs_8.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X406 dffrs_4.nand3_8.Z dffrs_4.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X407 a_30716_12225# dffrs_12.Q vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X408 a_26858_12225# dffrs_11.nand3_8.C a_26674_12225# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X409 dffrs_8.nand3_1.C dffrs_1.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X410 vdd reset dffrs_9.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X411 dffrs_12.nand3_8.C dffrs_12.nand3_8.Z vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X412 vdd dffrs_14.nand3_6.C d5 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X413 vdd dffrs_1.nand3_6.C dffrs_2.d vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X414 dffrs_5.nand3_1.C vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X415 dffrs_12.nand3_6.C vss vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X416 dffrs_4.nand3_8.C dffrs_4.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X417 dffrs_11.nand3_1.C dffrs_4.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X418 a_17104_443# dffrs_3.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X419 a_13062_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X420 a_29230_12224# dffrs_12.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X421 a_10506_12225# d4 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X422 dffrs_10.nand3_8.C dffrs_10.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X423 a_5162_14432# reset a_4978_14432# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X424 dffrs_2.Q dffrs_2.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X425 a_18590_2649# dffrs_4.d vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X426 a_13246_443# reset a_13062_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X427 dffrs_10.nand3_6.C dffrs_10.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X428 a_14548_14429# dffrs_1.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X429 a_29230_14429# dffrs_12.nand3_1.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X430 a_5162_16637# dffrs_14.nand3_8.Z a_4978_16637# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X431 a_5162_7058# dffrs_0.nand3_8.Z a_4978_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X432 a_17104_7058# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X433 dffrs_13.nand3_8.Z dffrs_13.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X434 vdd dffrs_1.nand3_8.C dffrs_1.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X435 vdd dffrs_14.nand3_8.C dffrs_14.Qb vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X436 dffrs_14.nand3_6.C dffrs_14.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X437 dffrs_13.nand3_8.C dffrs_13.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X438 dffrs_2.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X439 a_14548_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X440 dffrs_14.nand3_1.C dffrs_13.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X441 dffrs_0.nand3_6.C clk a_5162_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X442 a_25372_4853# reset a_25188_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X443 a_17288_4853# reset a_17104_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X444 a_5162_443# reset a_4978_443# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X445 a_9204_10019# reset a_9020_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X446 a_9020_10019# dffrs_7.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X447 dffrs_0.Q dffrs_0.Qb a_6648_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X448 d4 dffrs_7.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X449 a_13246_2648# clk a_13062_2648# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X450 dffrs_8.nand3_1.C dffrs_8.nand3_6.C a_13246_16634# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X451 a_14548_2649# dffrs_2.Q vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X452 dffrs_8.Qb reset vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X453 d5 dffrs_14.Qb a_6648_14432# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X454 d2 dffrs_9.Qb vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X455 vdd dffrs_10.nand3_6.C d1 vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X456 dffrs_12.nand3_1.C dffrs_5.Qb vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X457 a_21330_12224# d0 a_21146_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X458 dffrs_9.nand3_8.C dffrs_9.nand3_8.Z a_17288_12224# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X459 dffrs_0.Qb reset a_6648_2649# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X460 a_21330_14429# reset a_21146_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X461 dffrs_9.nand3_6.C d1 a_17288_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X462 dffrs_0.nand3_1.C dffrs_0.nand3_6.C a_5162_7058# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X463 a_17288_7058# dffrs_3.nand3_8.Z a_17104_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X464 a_25372_7058# dffrs_5.nand3_8.Z a_25188_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X465 a_29414_12224# vss a_29230_12224# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X466 dffrs_14.Qb reset a_6648_12228# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X467 dffrs_8.Qb d3 vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X468 a_10506_4853# vdd vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X469 dffrs_14.nand3_6.C d4 a_5162_14432# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X470 a_6464_14432# dffrs_13.Qb vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X471 a_29414_14429# reset a_29230_14429# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X472 dffrs_14.nand3_1.C dffrs_14.nand3_6.C a_5162_16637# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X473 a_21330_4853# reset a_21146_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X474 a_25372_10019# reset a_25188_10019# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X475 vdd d3 dffrs_7.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X476 a_1150_4853# vdd a_966_4853# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X477 dffrs_7.nand3_8.C dffrs_7.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X478 vdd reset dffrs_7.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X479 dffrs_5.nand3_6.C clk a_25372_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X480 dffrs_7.nand3_6.C dffrs_7.nand3_1.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X481 a_25188_2648# dffrs_5.nand3_6.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X482 a_10506_2649# dffrs_2.d vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X483 a_6464_12228# d5 vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X484 dffrs_0.Q vdd vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X485 dffrs_2.nand3_8.Z dffrs_2.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X486 dffrs_5.Q dffrs_5.Qb a_26858_4853# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X487 vdd reset dffrs_1.nand3_6.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X488 a_17104_10019# dffrs_9.nand3_8.C vss vss nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X489 dffrs_7.nand3_8.Z comp_in a_9204_10019# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X490 dffrs_8.nand3_8.Z comp_in vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X491 dffrs_2.nand3_8.C dffrs_2.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X492 vdd reset dffrs_0.nand3_8.Z vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X493 d1 dffrs_10.Qb a_22816_14429# vss nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X494 dffrs_3.nand3_8.Z dffrs_3.nand3_8.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X495 vdd dffrs_1.nand3_8.Z dffrs_1.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X496 dffrs_9.nand3_1.C dffrs_9.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X497 vdd dffrs_10.nand3_8.Z dffrs_10.nand3_1.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X498 dffrs_3.nand3_6.C clk vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
X499 vdd clk dffrs_0.nand3_8.C vdd pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X500 dffrs_3.nand3_8.C dffrs_3.nand3_6.C vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X501 a_21330_7058# dffrs_4.nand3_8.Z a_21146_7058# vss nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
X502 dffrs_0.Qb dffrs_0.Q vdd vdd pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X503 dffrs_3.nand3_1.C dffrs_3.nand3_6.C vdd vdd pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
.ends

.subckt comp_SAR_final Vdd Vss Clk Vin1 Vin2 Comp_out Reset SAR_in Load Clk_piso Piso_out
Xcomparator_no_offsetcal_0 Vdd Vss Clk Vin1 Vin2 Comp_out comparator_no_offsetcal
Xinv2_0 Load Vdd inv2_0/out Vss inv2
Xadc_PISO_0 inv2_0/out adc_PISO_0/B6 adc_PISO_0/B5 adc_PISO_0/B4 Piso_out Vdd adc_PISO_0/B3
+ Vss adc_PISO_0/B2 adc_PISO_0/B1 Clk_piso adc_PISO
XSARlogic_0 Vdd Vss Clk Reset SAR_in adc_PISO_0/B6 adc_PISO_0/B5 adc_PISO_0/B4 adc_PISO_0/B3
+ adc_PISO_0/B2 adc_PISO_0/B1 SARlogic
.ends

