magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -2718 -23370 2718 23370
<< nmos >>
rect -2468 19160 -2068 23160
rect -1964 19160 -1564 23160
rect -1460 19160 -1060 23160
rect -956 19160 -556 23160
rect -452 19160 -52 23160
rect 52 19160 452 23160
rect 556 19160 956 23160
rect 1060 19160 1460 23160
rect 1564 19160 1964 23160
rect 2068 19160 2468 23160
rect -2468 14928 -2068 18928
rect -1964 14928 -1564 18928
rect -1460 14928 -1060 18928
rect -956 14928 -556 18928
rect -452 14928 -52 18928
rect 52 14928 452 18928
rect 556 14928 956 18928
rect 1060 14928 1460 18928
rect 1564 14928 1964 18928
rect 2068 14928 2468 18928
rect -2468 10696 -2068 14696
rect -1964 10696 -1564 14696
rect -1460 10696 -1060 14696
rect -956 10696 -556 14696
rect -452 10696 -52 14696
rect 52 10696 452 14696
rect 556 10696 956 14696
rect 1060 10696 1460 14696
rect 1564 10696 1964 14696
rect 2068 10696 2468 14696
rect -2468 6464 -2068 10464
rect -1964 6464 -1564 10464
rect -1460 6464 -1060 10464
rect -956 6464 -556 10464
rect -452 6464 -52 10464
rect 52 6464 452 10464
rect 556 6464 956 10464
rect 1060 6464 1460 10464
rect 1564 6464 1964 10464
rect 2068 6464 2468 10464
rect -2468 2232 -2068 6232
rect -1964 2232 -1564 6232
rect -1460 2232 -1060 6232
rect -956 2232 -556 6232
rect -452 2232 -52 6232
rect 52 2232 452 6232
rect 556 2232 956 6232
rect 1060 2232 1460 6232
rect 1564 2232 1964 6232
rect 2068 2232 2468 6232
rect -2468 -2000 -2068 2000
rect -1964 -2000 -1564 2000
rect -1460 -2000 -1060 2000
rect -956 -2000 -556 2000
rect -452 -2000 -52 2000
rect 52 -2000 452 2000
rect 556 -2000 956 2000
rect 1060 -2000 1460 2000
rect 1564 -2000 1964 2000
rect 2068 -2000 2468 2000
rect -2468 -6232 -2068 -2232
rect -1964 -6232 -1564 -2232
rect -1460 -6232 -1060 -2232
rect -956 -6232 -556 -2232
rect -452 -6232 -52 -2232
rect 52 -6232 452 -2232
rect 556 -6232 956 -2232
rect 1060 -6232 1460 -2232
rect 1564 -6232 1964 -2232
rect 2068 -6232 2468 -2232
rect -2468 -10464 -2068 -6464
rect -1964 -10464 -1564 -6464
rect -1460 -10464 -1060 -6464
rect -956 -10464 -556 -6464
rect -452 -10464 -52 -6464
rect 52 -10464 452 -6464
rect 556 -10464 956 -6464
rect 1060 -10464 1460 -6464
rect 1564 -10464 1964 -6464
rect 2068 -10464 2468 -6464
rect -2468 -14696 -2068 -10696
rect -1964 -14696 -1564 -10696
rect -1460 -14696 -1060 -10696
rect -956 -14696 -556 -10696
rect -452 -14696 -52 -10696
rect 52 -14696 452 -10696
rect 556 -14696 956 -10696
rect 1060 -14696 1460 -10696
rect 1564 -14696 1964 -10696
rect 2068 -14696 2468 -10696
rect -2468 -18928 -2068 -14928
rect -1964 -18928 -1564 -14928
rect -1460 -18928 -1060 -14928
rect -956 -18928 -556 -14928
rect -452 -18928 -52 -14928
rect 52 -18928 452 -14928
rect 556 -18928 956 -14928
rect 1060 -18928 1460 -14928
rect 1564 -18928 1964 -14928
rect 2068 -18928 2468 -14928
rect -2468 -23160 -2068 -19160
rect -1964 -23160 -1564 -19160
rect -1460 -23160 -1060 -19160
rect -956 -23160 -556 -19160
rect -452 -23160 -52 -19160
rect 52 -23160 452 -19160
rect 556 -23160 956 -19160
rect 1060 -23160 1460 -19160
rect 1564 -23160 1964 -19160
rect 2068 -23160 2468 -19160
<< ndiff >>
rect -2556 23147 -2468 23160
rect -2556 19173 -2543 23147
rect -2497 19173 -2468 23147
rect -2556 19160 -2468 19173
rect -2068 23147 -1964 23160
rect -2068 19173 -2039 23147
rect -1993 19173 -1964 23147
rect -2068 19160 -1964 19173
rect -1564 23147 -1460 23160
rect -1564 19173 -1535 23147
rect -1489 19173 -1460 23147
rect -1564 19160 -1460 19173
rect -1060 23147 -956 23160
rect -1060 19173 -1031 23147
rect -985 19173 -956 23147
rect -1060 19160 -956 19173
rect -556 23147 -452 23160
rect -556 19173 -527 23147
rect -481 19173 -452 23147
rect -556 19160 -452 19173
rect -52 23147 52 23160
rect -52 19173 -23 23147
rect 23 19173 52 23147
rect -52 19160 52 19173
rect 452 23147 556 23160
rect 452 19173 481 23147
rect 527 19173 556 23147
rect 452 19160 556 19173
rect 956 23147 1060 23160
rect 956 19173 985 23147
rect 1031 19173 1060 23147
rect 956 19160 1060 19173
rect 1460 23147 1564 23160
rect 1460 19173 1489 23147
rect 1535 19173 1564 23147
rect 1460 19160 1564 19173
rect 1964 23147 2068 23160
rect 1964 19173 1993 23147
rect 2039 19173 2068 23147
rect 1964 19160 2068 19173
rect 2468 23147 2556 23160
rect 2468 19173 2497 23147
rect 2543 19173 2556 23147
rect 2468 19160 2556 19173
rect -2556 18915 -2468 18928
rect -2556 14941 -2543 18915
rect -2497 14941 -2468 18915
rect -2556 14928 -2468 14941
rect -2068 18915 -1964 18928
rect -2068 14941 -2039 18915
rect -1993 14941 -1964 18915
rect -2068 14928 -1964 14941
rect -1564 18915 -1460 18928
rect -1564 14941 -1535 18915
rect -1489 14941 -1460 18915
rect -1564 14928 -1460 14941
rect -1060 18915 -956 18928
rect -1060 14941 -1031 18915
rect -985 14941 -956 18915
rect -1060 14928 -956 14941
rect -556 18915 -452 18928
rect -556 14941 -527 18915
rect -481 14941 -452 18915
rect -556 14928 -452 14941
rect -52 18915 52 18928
rect -52 14941 -23 18915
rect 23 14941 52 18915
rect -52 14928 52 14941
rect 452 18915 556 18928
rect 452 14941 481 18915
rect 527 14941 556 18915
rect 452 14928 556 14941
rect 956 18915 1060 18928
rect 956 14941 985 18915
rect 1031 14941 1060 18915
rect 956 14928 1060 14941
rect 1460 18915 1564 18928
rect 1460 14941 1489 18915
rect 1535 14941 1564 18915
rect 1460 14928 1564 14941
rect 1964 18915 2068 18928
rect 1964 14941 1993 18915
rect 2039 14941 2068 18915
rect 1964 14928 2068 14941
rect 2468 18915 2556 18928
rect 2468 14941 2497 18915
rect 2543 14941 2556 18915
rect 2468 14928 2556 14941
rect -2556 14683 -2468 14696
rect -2556 10709 -2543 14683
rect -2497 10709 -2468 14683
rect -2556 10696 -2468 10709
rect -2068 14683 -1964 14696
rect -2068 10709 -2039 14683
rect -1993 10709 -1964 14683
rect -2068 10696 -1964 10709
rect -1564 14683 -1460 14696
rect -1564 10709 -1535 14683
rect -1489 10709 -1460 14683
rect -1564 10696 -1460 10709
rect -1060 14683 -956 14696
rect -1060 10709 -1031 14683
rect -985 10709 -956 14683
rect -1060 10696 -956 10709
rect -556 14683 -452 14696
rect -556 10709 -527 14683
rect -481 10709 -452 14683
rect -556 10696 -452 10709
rect -52 14683 52 14696
rect -52 10709 -23 14683
rect 23 10709 52 14683
rect -52 10696 52 10709
rect 452 14683 556 14696
rect 452 10709 481 14683
rect 527 10709 556 14683
rect 452 10696 556 10709
rect 956 14683 1060 14696
rect 956 10709 985 14683
rect 1031 10709 1060 14683
rect 956 10696 1060 10709
rect 1460 14683 1564 14696
rect 1460 10709 1489 14683
rect 1535 10709 1564 14683
rect 1460 10696 1564 10709
rect 1964 14683 2068 14696
rect 1964 10709 1993 14683
rect 2039 10709 2068 14683
rect 1964 10696 2068 10709
rect 2468 14683 2556 14696
rect 2468 10709 2497 14683
rect 2543 10709 2556 14683
rect 2468 10696 2556 10709
rect -2556 10451 -2468 10464
rect -2556 6477 -2543 10451
rect -2497 6477 -2468 10451
rect -2556 6464 -2468 6477
rect -2068 10451 -1964 10464
rect -2068 6477 -2039 10451
rect -1993 6477 -1964 10451
rect -2068 6464 -1964 6477
rect -1564 10451 -1460 10464
rect -1564 6477 -1535 10451
rect -1489 6477 -1460 10451
rect -1564 6464 -1460 6477
rect -1060 10451 -956 10464
rect -1060 6477 -1031 10451
rect -985 6477 -956 10451
rect -1060 6464 -956 6477
rect -556 10451 -452 10464
rect -556 6477 -527 10451
rect -481 6477 -452 10451
rect -556 6464 -452 6477
rect -52 10451 52 10464
rect -52 6477 -23 10451
rect 23 6477 52 10451
rect -52 6464 52 6477
rect 452 10451 556 10464
rect 452 6477 481 10451
rect 527 6477 556 10451
rect 452 6464 556 6477
rect 956 10451 1060 10464
rect 956 6477 985 10451
rect 1031 6477 1060 10451
rect 956 6464 1060 6477
rect 1460 10451 1564 10464
rect 1460 6477 1489 10451
rect 1535 6477 1564 10451
rect 1460 6464 1564 6477
rect 1964 10451 2068 10464
rect 1964 6477 1993 10451
rect 2039 6477 2068 10451
rect 1964 6464 2068 6477
rect 2468 10451 2556 10464
rect 2468 6477 2497 10451
rect 2543 6477 2556 10451
rect 2468 6464 2556 6477
rect -2556 6219 -2468 6232
rect -2556 2245 -2543 6219
rect -2497 2245 -2468 6219
rect -2556 2232 -2468 2245
rect -2068 6219 -1964 6232
rect -2068 2245 -2039 6219
rect -1993 2245 -1964 6219
rect -2068 2232 -1964 2245
rect -1564 6219 -1460 6232
rect -1564 2245 -1535 6219
rect -1489 2245 -1460 6219
rect -1564 2232 -1460 2245
rect -1060 6219 -956 6232
rect -1060 2245 -1031 6219
rect -985 2245 -956 6219
rect -1060 2232 -956 2245
rect -556 6219 -452 6232
rect -556 2245 -527 6219
rect -481 2245 -452 6219
rect -556 2232 -452 2245
rect -52 6219 52 6232
rect -52 2245 -23 6219
rect 23 2245 52 6219
rect -52 2232 52 2245
rect 452 6219 556 6232
rect 452 2245 481 6219
rect 527 2245 556 6219
rect 452 2232 556 2245
rect 956 6219 1060 6232
rect 956 2245 985 6219
rect 1031 2245 1060 6219
rect 956 2232 1060 2245
rect 1460 6219 1564 6232
rect 1460 2245 1489 6219
rect 1535 2245 1564 6219
rect 1460 2232 1564 2245
rect 1964 6219 2068 6232
rect 1964 2245 1993 6219
rect 2039 2245 2068 6219
rect 1964 2232 2068 2245
rect 2468 6219 2556 6232
rect 2468 2245 2497 6219
rect 2543 2245 2556 6219
rect 2468 2232 2556 2245
rect -2556 1987 -2468 2000
rect -2556 -1987 -2543 1987
rect -2497 -1987 -2468 1987
rect -2556 -2000 -2468 -1987
rect -2068 1987 -1964 2000
rect -2068 -1987 -2039 1987
rect -1993 -1987 -1964 1987
rect -2068 -2000 -1964 -1987
rect -1564 1987 -1460 2000
rect -1564 -1987 -1535 1987
rect -1489 -1987 -1460 1987
rect -1564 -2000 -1460 -1987
rect -1060 1987 -956 2000
rect -1060 -1987 -1031 1987
rect -985 -1987 -956 1987
rect -1060 -2000 -956 -1987
rect -556 1987 -452 2000
rect -556 -1987 -527 1987
rect -481 -1987 -452 1987
rect -556 -2000 -452 -1987
rect -52 1987 52 2000
rect -52 -1987 -23 1987
rect 23 -1987 52 1987
rect -52 -2000 52 -1987
rect 452 1987 556 2000
rect 452 -1987 481 1987
rect 527 -1987 556 1987
rect 452 -2000 556 -1987
rect 956 1987 1060 2000
rect 956 -1987 985 1987
rect 1031 -1987 1060 1987
rect 956 -2000 1060 -1987
rect 1460 1987 1564 2000
rect 1460 -1987 1489 1987
rect 1535 -1987 1564 1987
rect 1460 -2000 1564 -1987
rect 1964 1987 2068 2000
rect 1964 -1987 1993 1987
rect 2039 -1987 2068 1987
rect 1964 -2000 2068 -1987
rect 2468 1987 2556 2000
rect 2468 -1987 2497 1987
rect 2543 -1987 2556 1987
rect 2468 -2000 2556 -1987
rect -2556 -2245 -2468 -2232
rect -2556 -6219 -2543 -2245
rect -2497 -6219 -2468 -2245
rect -2556 -6232 -2468 -6219
rect -2068 -2245 -1964 -2232
rect -2068 -6219 -2039 -2245
rect -1993 -6219 -1964 -2245
rect -2068 -6232 -1964 -6219
rect -1564 -2245 -1460 -2232
rect -1564 -6219 -1535 -2245
rect -1489 -6219 -1460 -2245
rect -1564 -6232 -1460 -6219
rect -1060 -2245 -956 -2232
rect -1060 -6219 -1031 -2245
rect -985 -6219 -956 -2245
rect -1060 -6232 -956 -6219
rect -556 -2245 -452 -2232
rect -556 -6219 -527 -2245
rect -481 -6219 -452 -2245
rect -556 -6232 -452 -6219
rect -52 -2245 52 -2232
rect -52 -6219 -23 -2245
rect 23 -6219 52 -2245
rect -52 -6232 52 -6219
rect 452 -2245 556 -2232
rect 452 -6219 481 -2245
rect 527 -6219 556 -2245
rect 452 -6232 556 -6219
rect 956 -2245 1060 -2232
rect 956 -6219 985 -2245
rect 1031 -6219 1060 -2245
rect 956 -6232 1060 -6219
rect 1460 -2245 1564 -2232
rect 1460 -6219 1489 -2245
rect 1535 -6219 1564 -2245
rect 1460 -6232 1564 -6219
rect 1964 -2245 2068 -2232
rect 1964 -6219 1993 -2245
rect 2039 -6219 2068 -2245
rect 1964 -6232 2068 -6219
rect 2468 -2245 2556 -2232
rect 2468 -6219 2497 -2245
rect 2543 -6219 2556 -2245
rect 2468 -6232 2556 -6219
rect -2556 -6477 -2468 -6464
rect -2556 -10451 -2543 -6477
rect -2497 -10451 -2468 -6477
rect -2556 -10464 -2468 -10451
rect -2068 -6477 -1964 -6464
rect -2068 -10451 -2039 -6477
rect -1993 -10451 -1964 -6477
rect -2068 -10464 -1964 -10451
rect -1564 -6477 -1460 -6464
rect -1564 -10451 -1535 -6477
rect -1489 -10451 -1460 -6477
rect -1564 -10464 -1460 -10451
rect -1060 -6477 -956 -6464
rect -1060 -10451 -1031 -6477
rect -985 -10451 -956 -6477
rect -1060 -10464 -956 -10451
rect -556 -6477 -452 -6464
rect -556 -10451 -527 -6477
rect -481 -10451 -452 -6477
rect -556 -10464 -452 -10451
rect -52 -6477 52 -6464
rect -52 -10451 -23 -6477
rect 23 -10451 52 -6477
rect -52 -10464 52 -10451
rect 452 -6477 556 -6464
rect 452 -10451 481 -6477
rect 527 -10451 556 -6477
rect 452 -10464 556 -10451
rect 956 -6477 1060 -6464
rect 956 -10451 985 -6477
rect 1031 -10451 1060 -6477
rect 956 -10464 1060 -10451
rect 1460 -6477 1564 -6464
rect 1460 -10451 1489 -6477
rect 1535 -10451 1564 -6477
rect 1460 -10464 1564 -10451
rect 1964 -6477 2068 -6464
rect 1964 -10451 1993 -6477
rect 2039 -10451 2068 -6477
rect 1964 -10464 2068 -10451
rect 2468 -6477 2556 -6464
rect 2468 -10451 2497 -6477
rect 2543 -10451 2556 -6477
rect 2468 -10464 2556 -10451
rect -2556 -10709 -2468 -10696
rect -2556 -14683 -2543 -10709
rect -2497 -14683 -2468 -10709
rect -2556 -14696 -2468 -14683
rect -2068 -10709 -1964 -10696
rect -2068 -14683 -2039 -10709
rect -1993 -14683 -1964 -10709
rect -2068 -14696 -1964 -14683
rect -1564 -10709 -1460 -10696
rect -1564 -14683 -1535 -10709
rect -1489 -14683 -1460 -10709
rect -1564 -14696 -1460 -14683
rect -1060 -10709 -956 -10696
rect -1060 -14683 -1031 -10709
rect -985 -14683 -956 -10709
rect -1060 -14696 -956 -14683
rect -556 -10709 -452 -10696
rect -556 -14683 -527 -10709
rect -481 -14683 -452 -10709
rect -556 -14696 -452 -14683
rect -52 -10709 52 -10696
rect -52 -14683 -23 -10709
rect 23 -14683 52 -10709
rect -52 -14696 52 -14683
rect 452 -10709 556 -10696
rect 452 -14683 481 -10709
rect 527 -14683 556 -10709
rect 452 -14696 556 -14683
rect 956 -10709 1060 -10696
rect 956 -14683 985 -10709
rect 1031 -14683 1060 -10709
rect 956 -14696 1060 -14683
rect 1460 -10709 1564 -10696
rect 1460 -14683 1489 -10709
rect 1535 -14683 1564 -10709
rect 1460 -14696 1564 -14683
rect 1964 -10709 2068 -10696
rect 1964 -14683 1993 -10709
rect 2039 -14683 2068 -10709
rect 1964 -14696 2068 -14683
rect 2468 -10709 2556 -10696
rect 2468 -14683 2497 -10709
rect 2543 -14683 2556 -10709
rect 2468 -14696 2556 -14683
rect -2556 -14941 -2468 -14928
rect -2556 -18915 -2543 -14941
rect -2497 -18915 -2468 -14941
rect -2556 -18928 -2468 -18915
rect -2068 -14941 -1964 -14928
rect -2068 -18915 -2039 -14941
rect -1993 -18915 -1964 -14941
rect -2068 -18928 -1964 -18915
rect -1564 -14941 -1460 -14928
rect -1564 -18915 -1535 -14941
rect -1489 -18915 -1460 -14941
rect -1564 -18928 -1460 -18915
rect -1060 -14941 -956 -14928
rect -1060 -18915 -1031 -14941
rect -985 -18915 -956 -14941
rect -1060 -18928 -956 -18915
rect -556 -14941 -452 -14928
rect -556 -18915 -527 -14941
rect -481 -18915 -452 -14941
rect -556 -18928 -452 -18915
rect -52 -14941 52 -14928
rect -52 -18915 -23 -14941
rect 23 -18915 52 -14941
rect -52 -18928 52 -18915
rect 452 -14941 556 -14928
rect 452 -18915 481 -14941
rect 527 -18915 556 -14941
rect 452 -18928 556 -18915
rect 956 -14941 1060 -14928
rect 956 -18915 985 -14941
rect 1031 -18915 1060 -14941
rect 956 -18928 1060 -18915
rect 1460 -14941 1564 -14928
rect 1460 -18915 1489 -14941
rect 1535 -18915 1564 -14941
rect 1460 -18928 1564 -18915
rect 1964 -14941 2068 -14928
rect 1964 -18915 1993 -14941
rect 2039 -18915 2068 -14941
rect 1964 -18928 2068 -18915
rect 2468 -14941 2556 -14928
rect 2468 -18915 2497 -14941
rect 2543 -18915 2556 -14941
rect 2468 -18928 2556 -18915
rect -2556 -19173 -2468 -19160
rect -2556 -23147 -2543 -19173
rect -2497 -23147 -2468 -19173
rect -2556 -23160 -2468 -23147
rect -2068 -19173 -1964 -19160
rect -2068 -23147 -2039 -19173
rect -1993 -23147 -1964 -19173
rect -2068 -23160 -1964 -23147
rect -1564 -19173 -1460 -19160
rect -1564 -23147 -1535 -19173
rect -1489 -23147 -1460 -19173
rect -1564 -23160 -1460 -23147
rect -1060 -19173 -956 -19160
rect -1060 -23147 -1031 -19173
rect -985 -23147 -956 -19173
rect -1060 -23160 -956 -23147
rect -556 -19173 -452 -19160
rect -556 -23147 -527 -19173
rect -481 -23147 -452 -19173
rect -556 -23160 -452 -23147
rect -52 -19173 52 -19160
rect -52 -23147 -23 -19173
rect 23 -23147 52 -19173
rect -52 -23160 52 -23147
rect 452 -19173 556 -19160
rect 452 -23147 481 -19173
rect 527 -23147 556 -19173
rect 452 -23160 556 -23147
rect 956 -19173 1060 -19160
rect 956 -23147 985 -19173
rect 1031 -23147 1060 -19173
rect 956 -23160 1060 -23147
rect 1460 -19173 1564 -19160
rect 1460 -23147 1489 -19173
rect 1535 -23147 1564 -19173
rect 1460 -23160 1564 -23147
rect 1964 -19173 2068 -19160
rect 1964 -23147 1993 -19173
rect 2039 -23147 2068 -19173
rect 1964 -23160 2068 -23147
rect 2468 -19173 2556 -19160
rect 2468 -23147 2497 -19173
rect 2543 -23147 2556 -19173
rect 2468 -23160 2556 -23147
<< ndiffc >>
rect -2543 19173 -2497 23147
rect -2039 19173 -1993 23147
rect -1535 19173 -1489 23147
rect -1031 19173 -985 23147
rect -527 19173 -481 23147
rect -23 19173 23 23147
rect 481 19173 527 23147
rect 985 19173 1031 23147
rect 1489 19173 1535 23147
rect 1993 19173 2039 23147
rect 2497 19173 2543 23147
rect -2543 14941 -2497 18915
rect -2039 14941 -1993 18915
rect -1535 14941 -1489 18915
rect -1031 14941 -985 18915
rect -527 14941 -481 18915
rect -23 14941 23 18915
rect 481 14941 527 18915
rect 985 14941 1031 18915
rect 1489 14941 1535 18915
rect 1993 14941 2039 18915
rect 2497 14941 2543 18915
rect -2543 10709 -2497 14683
rect -2039 10709 -1993 14683
rect -1535 10709 -1489 14683
rect -1031 10709 -985 14683
rect -527 10709 -481 14683
rect -23 10709 23 14683
rect 481 10709 527 14683
rect 985 10709 1031 14683
rect 1489 10709 1535 14683
rect 1993 10709 2039 14683
rect 2497 10709 2543 14683
rect -2543 6477 -2497 10451
rect -2039 6477 -1993 10451
rect -1535 6477 -1489 10451
rect -1031 6477 -985 10451
rect -527 6477 -481 10451
rect -23 6477 23 10451
rect 481 6477 527 10451
rect 985 6477 1031 10451
rect 1489 6477 1535 10451
rect 1993 6477 2039 10451
rect 2497 6477 2543 10451
rect -2543 2245 -2497 6219
rect -2039 2245 -1993 6219
rect -1535 2245 -1489 6219
rect -1031 2245 -985 6219
rect -527 2245 -481 6219
rect -23 2245 23 6219
rect 481 2245 527 6219
rect 985 2245 1031 6219
rect 1489 2245 1535 6219
rect 1993 2245 2039 6219
rect 2497 2245 2543 6219
rect -2543 -1987 -2497 1987
rect -2039 -1987 -1993 1987
rect -1535 -1987 -1489 1987
rect -1031 -1987 -985 1987
rect -527 -1987 -481 1987
rect -23 -1987 23 1987
rect 481 -1987 527 1987
rect 985 -1987 1031 1987
rect 1489 -1987 1535 1987
rect 1993 -1987 2039 1987
rect 2497 -1987 2543 1987
rect -2543 -6219 -2497 -2245
rect -2039 -6219 -1993 -2245
rect -1535 -6219 -1489 -2245
rect -1031 -6219 -985 -2245
rect -527 -6219 -481 -2245
rect -23 -6219 23 -2245
rect 481 -6219 527 -2245
rect 985 -6219 1031 -2245
rect 1489 -6219 1535 -2245
rect 1993 -6219 2039 -2245
rect 2497 -6219 2543 -2245
rect -2543 -10451 -2497 -6477
rect -2039 -10451 -1993 -6477
rect -1535 -10451 -1489 -6477
rect -1031 -10451 -985 -6477
rect -527 -10451 -481 -6477
rect -23 -10451 23 -6477
rect 481 -10451 527 -6477
rect 985 -10451 1031 -6477
rect 1489 -10451 1535 -6477
rect 1993 -10451 2039 -6477
rect 2497 -10451 2543 -6477
rect -2543 -14683 -2497 -10709
rect -2039 -14683 -1993 -10709
rect -1535 -14683 -1489 -10709
rect -1031 -14683 -985 -10709
rect -527 -14683 -481 -10709
rect -23 -14683 23 -10709
rect 481 -14683 527 -10709
rect 985 -14683 1031 -10709
rect 1489 -14683 1535 -10709
rect 1993 -14683 2039 -10709
rect 2497 -14683 2543 -10709
rect -2543 -18915 -2497 -14941
rect -2039 -18915 -1993 -14941
rect -1535 -18915 -1489 -14941
rect -1031 -18915 -985 -14941
rect -527 -18915 -481 -14941
rect -23 -18915 23 -14941
rect 481 -18915 527 -14941
rect 985 -18915 1031 -14941
rect 1489 -18915 1535 -14941
rect 1993 -18915 2039 -14941
rect 2497 -18915 2543 -14941
rect -2543 -23147 -2497 -19173
rect -2039 -23147 -1993 -19173
rect -1535 -23147 -1489 -19173
rect -1031 -23147 -985 -19173
rect -527 -23147 -481 -19173
rect -23 -23147 23 -19173
rect 481 -23147 527 -19173
rect 985 -23147 1031 -19173
rect 1489 -23147 1535 -19173
rect 1993 -23147 2039 -19173
rect 2497 -23147 2543 -19173
<< psubdiff >>
rect -2694 23274 2694 23346
rect -2694 23230 -2622 23274
rect -2694 -23230 -2681 23230
rect -2635 -23230 -2622 23230
rect 2622 23230 2694 23274
rect -2694 -23274 -2622 -23230
rect 2622 -23230 2635 23230
rect 2681 -23230 2694 23230
rect 2622 -23274 2694 -23230
rect -2694 -23346 2694 -23274
<< psubdiffcont >>
rect -2681 -23230 -2635 23230
rect 2635 -23230 2681 23230
<< polysilicon >>
rect -2468 23239 -2068 23252
rect -2468 23193 -2455 23239
rect -2081 23193 -2068 23239
rect -2468 23160 -2068 23193
rect -1964 23239 -1564 23252
rect -1964 23193 -1951 23239
rect -1577 23193 -1564 23239
rect -1964 23160 -1564 23193
rect -1460 23239 -1060 23252
rect -1460 23193 -1447 23239
rect -1073 23193 -1060 23239
rect -1460 23160 -1060 23193
rect -956 23239 -556 23252
rect -956 23193 -943 23239
rect -569 23193 -556 23239
rect -956 23160 -556 23193
rect -452 23239 -52 23252
rect -452 23193 -439 23239
rect -65 23193 -52 23239
rect -452 23160 -52 23193
rect 52 23239 452 23252
rect 52 23193 65 23239
rect 439 23193 452 23239
rect 52 23160 452 23193
rect 556 23239 956 23252
rect 556 23193 569 23239
rect 943 23193 956 23239
rect 556 23160 956 23193
rect 1060 23239 1460 23252
rect 1060 23193 1073 23239
rect 1447 23193 1460 23239
rect 1060 23160 1460 23193
rect 1564 23239 1964 23252
rect 1564 23193 1577 23239
rect 1951 23193 1964 23239
rect 1564 23160 1964 23193
rect 2068 23239 2468 23252
rect 2068 23193 2081 23239
rect 2455 23193 2468 23239
rect 2068 23160 2468 23193
rect -2468 19127 -2068 19160
rect -2468 19081 -2455 19127
rect -2081 19081 -2068 19127
rect -2468 19068 -2068 19081
rect -1964 19127 -1564 19160
rect -1964 19081 -1951 19127
rect -1577 19081 -1564 19127
rect -1964 19068 -1564 19081
rect -1460 19127 -1060 19160
rect -1460 19081 -1447 19127
rect -1073 19081 -1060 19127
rect -1460 19068 -1060 19081
rect -956 19127 -556 19160
rect -956 19081 -943 19127
rect -569 19081 -556 19127
rect -956 19068 -556 19081
rect -452 19127 -52 19160
rect -452 19081 -439 19127
rect -65 19081 -52 19127
rect -452 19068 -52 19081
rect 52 19127 452 19160
rect 52 19081 65 19127
rect 439 19081 452 19127
rect 52 19068 452 19081
rect 556 19127 956 19160
rect 556 19081 569 19127
rect 943 19081 956 19127
rect 556 19068 956 19081
rect 1060 19127 1460 19160
rect 1060 19081 1073 19127
rect 1447 19081 1460 19127
rect 1060 19068 1460 19081
rect 1564 19127 1964 19160
rect 1564 19081 1577 19127
rect 1951 19081 1964 19127
rect 1564 19068 1964 19081
rect 2068 19127 2468 19160
rect 2068 19081 2081 19127
rect 2455 19081 2468 19127
rect 2068 19068 2468 19081
rect -2468 19007 -2068 19020
rect -2468 18961 -2455 19007
rect -2081 18961 -2068 19007
rect -2468 18928 -2068 18961
rect -1964 19007 -1564 19020
rect -1964 18961 -1951 19007
rect -1577 18961 -1564 19007
rect -1964 18928 -1564 18961
rect -1460 19007 -1060 19020
rect -1460 18961 -1447 19007
rect -1073 18961 -1060 19007
rect -1460 18928 -1060 18961
rect -956 19007 -556 19020
rect -956 18961 -943 19007
rect -569 18961 -556 19007
rect -956 18928 -556 18961
rect -452 19007 -52 19020
rect -452 18961 -439 19007
rect -65 18961 -52 19007
rect -452 18928 -52 18961
rect 52 19007 452 19020
rect 52 18961 65 19007
rect 439 18961 452 19007
rect 52 18928 452 18961
rect 556 19007 956 19020
rect 556 18961 569 19007
rect 943 18961 956 19007
rect 556 18928 956 18961
rect 1060 19007 1460 19020
rect 1060 18961 1073 19007
rect 1447 18961 1460 19007
rect 1060 18928 1460 18961
rect 1564 19007 1964 19020
rect 1564 18961 1577 19007
rect 1951 18961 1964 19007
rect 1564 18928 1964 18961
rect 2068 19007 2468 19020
rect 2068 18961 2081 19007
rect 2455 18961 2468 19007
rect 2068 18928 2468 18961
rect -2468 14895 -2068 14928
rect -2468 14849 -2455 14895
rect -2081 14849 -2068 14895
rect -2468 14836 -2068 14849
rect -1964 14895 -1564 14928
rect -1964 14849 -1951 14895
rect -1577 14849 -1564 14895
rect -1964 14836 -1564 14849
rect -1460 14895 -1060 14928
rect -1460 14849 -1447 14895
rect -1073 14849 -1060 14895
rect -1460 14836 -1060 14849
rect -956 14895 -556 14928
rect -956 14849 -943 14895
rect -569 14849 -556 14895
rect -956 14836 -556 14849
rect -452 14895 -52 14928
rect -452 14849 -439 14895
rect -65 14849 -52 14895
rect -452 14836 -52 14849
rect 52 14895 452 14928
rect 52 14849 65 14895
rect 439 14849 452 14895
rect 52 14836 452 14849
rect 556 14895 956 14928
rect 556 14849 569 14895
rect 943 14849 956 14895
rect 556 14836 956 14849
rect 1060 14895 1460 14928
rect 1060 14849 1073 14895
rect 1447 14849 1460 14895
rect 1060 14836 1460 14849
rect 1564 14895 1964 14928
rect 1564 14849 1577 14895
rect 1951 14849 1964 14895
rect 1564 14836 1964 14849
rect 2068 14895 2468 14928
rect 2068 14849 2081 14895
rect 2455 14849 2468 14895
rect 2068 14836 2468 14849
rect -2468 14775 -2068 14788
rect -2468 14729 -2455 14775
rect -2081 14729 -2068 14775
rect -2468 14696 -2068 14729
rect -1964 14775 -1564 14788
rect -1964 14729 -1951 14775
rect -1577 14729 -1564 14775
rect -1964 14696 -1564 14729
rect -1460 14775 -1060 14788
rect -1460 14729 -1447 14775
rect -1073 14729 -1060 14775
rect -1460 14696 -1060 14729
rect -956 14775 -556 14788
rect -956 14729 -943 14775
rect -569 14729 -556 14775
rect -956 14696 -556 14729
rect -452 14775 -52 14788
rect -452 14729 -439 14775
rect -65 14729 -52 14775
rect -452 14696 -52 14729
rect 52 14775 452 14788
rect 52 14729 65 14775
rect 439 14729 452 14775
rect 52 14696 452 14729
rect 556 14775 956 14788
rect 556 14729 569 14775
rect 943 14729 956 14775
rect 556 14696 956 14729
rect 1060 14775 1460 14788
rect 1060 14729 1073 14775
rect 1447 14729 1460 14775
rect 1060 14696 1460 14729
rect 1564 14775 1964 14788
rect 1564 14729 1577 14775
rect 1951 14729 1964 14775
rect 1564 14696 1964 14729
rect 2068 14775 2468 14788
rect 2068 14729 2081 14775
rect 2455 14729 2468 14775
rect 2068 14696 2468 14729
rect -2468 10663 -2068 10696
rect -2468 10617 -2455 10663
rect -2081 10617 -2068 10663
rect -2468 10604 -2068 10617
rect -1964 10663 -1564 10696
rect -1964 10617 -1951 10663
rect -1577 10617 -1564 10663
rect -1964 10604 -1564 10617
rect -1460 10663 -1060 10696
rect -1460 10617 -1447 10663
rect -1073 10617 -1060 10663
rect -1460 10604 -1060 10617
rect -956 10663 -556 10696
rect -956 10617 -943 10663
rect -569 10617 -556 10663
rect -956 10604 -556 10617
rect -452 10663 -52 10696
rect -452 10617 -439 10663
rect -65 10617 -52 10663
rect -452 10604 -52 10617
rect 52 10663 452 10696
rect 52 10617 65 10663
rect 439 10617 452 10663
rect 52 10604 452 10617
rect 556 10663 956 10696
rect 556 10617 569 10663
rect 943 10617 956 10663
rect 556 10604 956 10617
rect 1060 10663 1460 10696
rect 1060 10617 1073 10663
rect 1447 10617 1460 10663
rect 1060 10604 1460 10617
rect 1564 10663 1964 10696
rect 1564 10617 1577 10663
rect 1951 10617 1964 10663
rect 1564 10604 1964 10617
rect 2068 10663 2468 10696
rect 2068 10617 2081 10663
rect 2455 10617 2468 10663
rect 2068 10604 2468 10617
rect -2468 10543 -2068 10556
rect -2468 10497 -2455 10543
rect -2081 10497 -2068 10543
rect -2468 10464 -2068 10497
rect -1964 10543 -1564 10556
rect -1964 10497 -1951 10543
rect -1577 10497 -1564 10543
rect -1964 10464 -1564 10497
rect -1460 10543 -1060 10556
rect -1460 10497 -1447 10543
rect -1073 10497 -1060 10543
rect -1460 10464 -1060 10497
rect -956 10543 -556 10556
rect -956 10497 -943 10543
rect -569 10497 -556 10543
rect -956 10464 -556 10497
rect -452 10543 -52 10556
rect -452 10497 -439 10543
rect -65 10497 -52 10543
rect -452 10464 -52 10497
rect 52 10543 452 10556
rect 52 10497 65 10543
rect 439 10497 452 10543
rect 52 10464 452 10497
rect 556 10543 956 10556
rect 556 10497 569 10543
rect 943 10497 956 10543
rect 556 10464 956 10497
rect 1060 10543 1460 10556
rect 1060 10497 1073 10543
rect 1447 10497 1460 10543
rect 1060 10464 1460 10497
rect 1564 10543 1964 10556
rect 1564 10497 1577 10543
rect 1951 10497 1964 10543
rect 1564 10464 1964 10497
rect 2068 10543 2468 10556
rect 2068 10497 2081 10543
rect 2455 10497 2468 10543
rect 2068 10464 2468 10497
rect -2468 6431 -2068 6464
rect -2468 6385 -2455 6431
rect -2081 6385 -2068 6431
rect -2468 6372 -2068 6385
rect -1964 6431 -1564 6464
rect -1964 6385 -1951 6431
rect -1577 6385 -1564 6431
rect -1964 6372 -1564 6385
rect -1460 6431 -1060 6464
rect -1460 6385 -1447 6431
rect -1073 6385 -1060 6431
rect -1460 6372 -1060 6385
rect -956 6431 -556 6464
rect -956 6385 -943 6431
rect -569 6385 -556 6431
rect -956 6372 -556 6385
rect -452 6431 -52 6464
rect -452 6385 -439 6431
rect -65 6385 -52 6431
rect -452 6372 -52 6385
rect 52 6431 452 6464
rect 52 6385 65 6431
rect 439 6385 452 6431
rect 52 6372 452 6385
rect 556 6431 956 6464
rect 556 6385 569 6431
rect 943 6385 956 6431
rect 556 6372 956 6385
rect 1060 6431 1460 6464
rect 1060 6385 1073 6431
rect 1447 6385 1460 6431
rect 1060 6372 1460 6385
rect 1564 6431 1964 6464
rect 1564 6385 1577 6431
rect 1951 6385 1964 6431
rect 1564 6372 1964 6385
rect 2068 6431 2468 6464
rect 2068 6385 2081 6431
rect 2455 6385 2468 6431
rect 2068 6372 2468 6385
rect -2468 6311 -2068 6324
rect -2468 6265 -2455 6311
rect -2081 6265 -2068 6311
rect -2468 6232 -2068 6265
rect -1964 6311 -1564 6324
rect -1964 6265 -1951 6311
rect -1577 6265 -1564 6311
rect -1964 6232 -1564 6265
rect -1460 6311 -1060 6324
rect -1460 6265 -1447 6311
rect -1073 6265 -1060 6311
rect -1460 6232 -1060 6265
rect -956 6311 -556 6324
rect -956 6265 -943 6311
rect -569 6265 -556 6311
rect -956 6232 -556 6265
rect -452 6311 -52 6324
rect -452 6265 -439 6311
rect -65 6265 -52 6311
rect -452 6232 -52 6265
rect 52 6311 452 6324
rect 52 6265 65 6311
rect 439 6265 452 6311
rect 52 6232 452 6265
rect 556 6311 956 6324
rect 556 6265 569 6311
rect 943 6265 956 6311
rect 556 6232 956 6265
rect 1060 6311 1460 6324
rect 1060 6265 1073 6311
rect 1447 6265 1460 6311
rect 1060 6232 1460 6265
rect 1564 6311 1964 6324
rect 1564 6265 1577 6311
rect 1951 6265 1964 6311
rect 1564 6232 1964 6265
rect 2068 6311 2468 6324
rect 2068 6265 2081 6311
rect 2455 6265 2468 6311
rect 2068 6232 2468 6265
rect -2468 2199 -2068 2232
rect -2468 2153 -2455 2199
rect -2081 2153 -2068 2199
rect -2468 2140 -2068 2153
rect -1964 2199 -1564 2232
rect -1964 2153 -1951 2199
rect -1577 2153 -1564 2199
rect -1964 2140 -1564 2153
rect -1460 2199 -1060 2232
rect -1460 2153 -1447 2199
rect -1073 2153 -1060 2199
rect -1460 2140 -1060 2153
rect -956 2199 -556 2232
rect -956 2153 -943 2199
rect -569 2153 -556 2199
rect -956 2140 -556 2153
rect -452 2199 -52 2232
rect -452 2153 -439 2199
rect -65 2153 -52 2199
rect -452 2140 -52 2153
rect 52 2199 452 2232
rect 52 2153 65 2199
rect 439 2153 452 2199
rect 52 2140 452 2153
rect 556 2199 956 2232
rect 556 2153 569 2199
rect 943 2153 956 2199
rect 556 2140 956 2153
rect 1060 2199 1460 2232
rect 1060 2153 1073 2199
rect 1447 2153 1460 2199
rect 1060 2140 1460 2153
rect 1564 2199 1964 2232
rect 1564 2153 1577 2199
rect 1951 2153 1964 2199
rect 1564 2140 1964 2153
rect 2068 2199 2468 2232
rect 2068 2153 2081 2199
rect 2455 2153 2468 2199
rect 2068 2140 2468 2153
rect -2468 2079 -2068 2092
rect -2468 2033 -2455 2079
rect -2081 2033 -2068 2079
rect -2468 2000 -2068 2033
rect -1964 2079 -1564 2092
rect -1964 2033 -1951 2079
rect -1577 2033 -1564 2079
rect -1964 2000 -1564 2033
rect -1460 2079 -1060 2092
rect -1460 2033 -1447 2079
rect -1073 2033 -1060 2079
rect -1460 2000 -1060 2033
rect -956 2079 -556 2092
rect -956 2033 -943 2079
rect -569 2033 -556 2079
rect -956 2000 -556 2033
rect -452 2079 -52 2092
rect -452 2033 -439 2079
rect -65 2033 -52 2079
rect -452 2000 -52 2033
rect 52 2079 452 2092
rect 52 2033 65 2079
rect 439 2033 452 2079
rect 52 2000 452 2033
rect 556 2079 956 2092
rect 556 2033 569 2079
rect 943 2033 956 2079
rect 556 2000 956 2033
rect 1060 2079 1460 2092
rect 1060 2033 1073 2079
rect 1447 2033 1460 2079
rect 1060 2000 1460 2033
rect 1564 2079 1964 2092
rect 1564 2033 1577 2079
rect 1951 2033 1964 2079
rect 1564 2000 1964 2033
rect 2068 2079 2468 2092
rect 2068 2033 2081 2079
rect 2455 2033 2468 2079
rect 2068 2000 2468 2033
rect -2468 -2033 -2068 -2000
rect -2468 -2079 -2455 -2033
rect -2081 -2079 -2068 -2033
rect -2468 -2092 -2068 -2079
rect -1964 -2033 -1564 -2000
rect -1964 -2079 -1951 -2033
rect -1577 -2079 -1564 -2033
rect -1964 -2092 -1564 -2079
rect -1460 -2033 -1060 -2000
rect -1460 -2079 -1447 -2033
rect -1073 -2079 -1060 -2033
rect -1460 -2092 -1060 -2079
rect -956 -2033 -556 -2000
rect -956 -2079 -943 -2033
rect -569 -2079 -556 -2033
rect -956 -2092 -556 -2079
rect -452 -2033 -52 -2000
rect -452 -2079 -439 -2033
rect -65 -2079 -52 -2033
rect -452 -2092 -52 -2079
rect 52 -2033 452 -2000
rect 52 -2079 65 -2033
rect 439 -2079 452 -2033
rect 52 -2092 452 -2079
rect 556 -2033 956 -2000
rect 556 -2079 569 -2033
rect 943 -2079 956 -2033
rect 556 -2092 956 -2079
rect 1060 -2033 1460 -2000
rect 1060 -2079 1073 -2033
rect 1447 -2079 1460 -2033
rect 1060 -2092 1460 -2079
rect 1564 -2033 1964 -2000
rect 1564 -2079 1577 -2033
rect 1951 -2079 1964 -2033
rect 1564 -2092 1964 -2079
rect 2068 -2033 2468 -2000
rect 2068 -2079 2081 -2033
rect 2455 -2079 2468 -2033
rect 2068 -2092 2468 -2079
rect -2468 -2153 -2068 -2140
rect -2468 -2199 -2455 -2153
rect -2081 -2199 -2068 -2153
rect -2468 -2232 -2068 -2199
rect -1964 -2153 -1564 -2140
rect -1964 -2199 -1951 -2153
rect -1577 -2199 -1564 -2153
rect -1964 -2232 -1564 -2199
rect -1460 -2153 -1060 -2140
rect -1460 -2199 -1447 -2153
rect -1073 -2199 -1060 -2153
rect -1460 -2232 -1060 -2199
rect -956 -2153 -556 -2140
rect -956 -2199 -943 -2153
rect -569 -2199 -556 -2153
rect -956 -2232 -556 -2199
rect -452 -2153 -52 -2140
rect -452 -2199 -439 -2153
rect -65 -2199 -52 -2153
rect -452 -2232 -52 -2199
rect 52 -2153 452 -2140
rect 52 -2199 65 -2153
rect 439 -2199 452 -2153
rect 52 -2232 452 -2199
rect 556 -2153 956 -2140
rect 556 -2199 569 -2153
rect 943 -2199 956 -2153
rect 556 -2232 956 -2199
rect 1060 -2153 1460 -2140
rect 1060 -2199 1073 -2153
rect 1447 -2199 1460 -2153
rect 1060 -2232 1460 -2199
rect 1564 -2153 1964 -2140
rect 1564 -2199 1577 -2153
rect 1951 -2199 1964 -2153
rect 1564 -2232 1964 -2199
rect 2068 -2153 2468 -2140
rect 2068 -2199 2081 -2153
rect 2455 -2199 2468 -2153
rect 2068 -2232 2468 -2199
rect -2468 -6265 -2068 -6232
rect -2468 -6311 -2455 -6265
rect -2081 -6311 -2068 -6265
rect -2468 -6324 -2068 -6311
rect -1964 -6265 -1564 -6232
rect -1964 -6311 -1951 -6265
rect -1577 -6311 -1564 -6265
rect -1964 -6324 -1564 -6311
rect -1460 -6265 -1060 -6232
rect -1460 -6311 -1447 -6265
rect -1073 -6311 -1060 -6265
rect -1460 -6324 -1060 -6311
rect -956 -6265 -556 -6232
rect -956 -6311 -943 -6265
rect -569 -6311 -556 -6265
rect -956 -6324 -556 -6311
rect -452 -6265 -52 -6232
rect -452 -6311 -439 -6265
rect -65 -6311 -52 -6265
rect -452 -6324 -52 -6311
rect 52 -6265 452 -6232
rect 52 -6311 65 -6265
rect 439 -6311 452 -6265
rect 52 -6324 452 -6311
rect 556 -6265 956 -6232
rect 556 -6311 569 -6265
rect 943 -6311 956 -6265
rect 556 -6324 956 -6311
rect 1060 -6265 1460 -6232
rect 1060 -6311 1073 -6265
rect 1447 -6311 1460 -6265
rect 1060 -6324 1460 -6311
rect 1564 -6265 1964 -6232
rect 1564 -6311 1577 -6265
rect 1951 -6311 1964 -6265
rect 1564 -6324 1964 -6311
rect 2068 -6265 2468 -6232
rect 2068 -6311 2081 -6265
rect 2455 -6311 2468 -6265
rect 2068 -6324 2468 -6311
rect -2468 -6385 -2068 -6372
rect -2468 -6431 -2455 -6385
rect -2081 -6431 -2068 -6385
rect -2468 -6464 -2068 -6431
rect -1964 -6385 -1564 -6372
rect -1964 -6431 -1951 -6385
rect -1577 -6431 -1564 -6385
rect -1964 -6464 -1564 -6431
rect -1460 -6385 -1060 -6372
rect -1460 -6431 -1447 -6385
rect -1073 -6431 -1060 -6385
rect -1460 -6464 -1060 -6431
rect -956 -6385 -556 -6372
rect -956 -6431 -943 -6385
rect -569 -6431 -556 -6385
rect -956 -6464 -556 -6431
rect -452 -6385 -52 -6372
rect -452 -6431 -439 -6385
rect -65 -6431 -52 -6385
rect -452 -6464 -52 -6431
rect 52 -6385 452 -6372
rect 52 -6431 65 -6385
rect 439 -6431 452 -6385
rect 52 -6464 452 -6431
rect 556 -6385 956 -6372
rect 556 -6431 569 -6385
rect 943 -6431 956 -6385
rect 556 -6464 956 -6431
rect 1060 -6385 1460 -6372
rect 1060 -6431 1073 -6385
rect 1447 -6431 1460 -6385
rect 1060 -6464 1460 -6431
rect 1564 -6385 1964 -6372
rect 1564 -6431 1577 -6385
rect 1951 -6431 1964 -6385
rect 1564 -6464 1964 -6431
rect 2068 -6385 2468 -6372
rect 2068 -6431 2081 -6385
rect 2455 -6431 2468 -6385
rect 2068 -6464 2468 -6431
rect -2468 -10497 -2068 -10464
rect -2468 -10543 -2455 -10497
rect -2081 -10543 -2068 -10497
rect -2468 -10556 -2068 -10543
rect -1964 -10497 -1564 -10464
rect -1964 -10543 -1951 -10497
rect -1577 -10543 -1564 -10497
rect -1964 -10556 -1564 -10543
rect -1460 -10497 -1060 -10464
rect -1460 -10543 -1447 -10497
rect -1073 -10543 -1060 -10497
rect -1460 -10556 -1060 -10543
rect -956 -10497 -556 -10464
rect -956 -10543 -943 -10497
rect -569 -10543 -556 -10497
rect -956 -10556 -556 -10543
rect -452 -10497 -52 -10464
rect -452 -10543 -439 -10497
rect -65 -10543 -52 -10497
rect -452 -10556 -52 -10543
rect 52 -10497 452 -10464
rect 52 -10543 65 -10497
rect 439 -10543 452 -10497
rect 52 -10556 452 -10543
rect 556 -10497 956 -10464
rect 556 -10543 569 -10497
rect 943 -10543 956 -10497
rect 556 -10556 956 -10543
rect 1060 -10497 1460 -10464
rect 1060 -10543 1073 -10497
rect 1447 -10543 1460 -10497
rect 1060 -10556 1460 -10543
rect 1564 -10497 1964 -10464
rect 1564 -10543 1577 -10497
rect 1951 -10543 1964 -10497
rect 1564 -10556 1964 -10543
rect 2068 -10497 2468 -10464
rect 2068 -10543 2081 -10497
rect 2455 -10543 2468 -10497
rect 2068 -10556 2468 -10543
rect -2468 -10617 -2068 -10604
rect -2468 -10663 -2455 -10617
rect -2081 -10663 -2068 -10617
rect -2468 -10696 -2068 -10663
rect -1964 -10617 -1564 -10604
rect -1964 -10663 -1951 -10617
rect -1577 -10663 -1564 -10617
rect -1964 -10696 -1564 -10663
rect -1460 -10617 -1060 -10604
rect -1460 -10663 -1447 -10617
rect -1073 -10663 -1060 -10617
rect -1460 -10696 -1060 -10663
rect -956 -10617 -556 -10604
rect -956 -10663 -943 -10617
rect -569 -10663 -556 -10617
rect -956 -10696 -556 -10663
rect -452 -10617 -52 -10604
rect -452 -10663 -439 -10617
rect -65 -10663 -52 -10617
rect -452 -10696 -52 -10663
rect 52 -10617 452 -10604
rect 52 -10663 65 -10617
rect 439 -10663 452 -10617
rect 52 -10696 452 -10663
rect 556 -10617 956 -10604
rect 556 -10663 569 -10617
rect 943 -10663 956 -10617
rect 556 -10696 956 -10663
rect 1060 -10617 1460 -10604
rect 1060 -10663 1073 -10617
rect 1447 -10663 1460 -10617
rect 1060 -10696 1460 -10663
rect 1564 -10617 1964 -10604
rect 1564 -10663 1577 -10617
rect 1951 -10663 1964 -10617
rect 1564 -10696 1964 -10663
rect 2068 -10617 2468 -10604
rect 2068 -10663 2081 -10617
rect 2455 -10663 2468 -10617
rect 2068 -10696 2468 -10663
rect -2468 -14729 -2068 -14696
rect -2468 -14775 -2455 -14729
rect -2081 -14775 -2068 -14729
rect -2468 -14788 -2068 -14775
rect -1964 -14729 -1564 -14696
rect -1964 -14775 -1951 -14729
rect -1577 -14775 -1564 -14729
rect -1964 -14788 -1564 -14775
rect -1460 -14729 -1060 -14696
rect -1460 -14775 -1447 -14729
rect -1073 -14775 -1060 -14729
rect -1460 -14788 -1060 -14775
rect -956 -14729 -556 -14696
rect -956 -14775 -943 -14729
rect -569 -14775 -556 -14729
rect -956 -14788 -556 -14775
rect -452 -14729 -52 -14696
rect -452 -14775 -439 -14729
rect -65 -14775 -52 -14729
rect -452 -14788 -52 -14775
rect 52 -14729 452 -14696
rect 52 -14775 65 -14729
rect 439 -14775 452 -14729
rect 52 -14788 452 -14775
rect 556 -14729 956 -14696
rect 556 -14775 569 -14729
rect 943 -14775 956 -14729
rect 556 -14788 956 -14775
rect 1060 -14729 1460 -14696
rect 1060 -14775 1073 -14729
rect 1447 -14775 1460 -14729
rect 1060 -14788 1460 -14775
rect 1564 -14729 1964 -14696
rect 1564 -14775 1577 -14729
rect 1951 -14775 1964 -14729
rect 1564 -14788 1964 -14775
rect 2068 -14729 2468 -14696
rect 2068 -14775 2081 -14729
rect 2455 -14775 2468 -14729
rect 2068 -14788 2468 -14775
rect -2468 -14849 -2068 -14836
rect -2468 -14895 -2455 -14849
rect -2081 -14895 -2068 -14849
rect -2468 -14928 -2068 -14895
rect -1964 -14849 -1564 -14836
rect -1964 -14895 -1951 -14849
rect -1577 -14895 -1564 -14849
rect -1964 -14928 -1564 -14895
rect -1460 -14849 -1060 -14836
rect -1460 -14895 -1447 -14849
rect -1073 -14895 -1060 -14849
rect -1460 -14928 -1060 -14895
rect -956 -14849 -556 -14836
rect -956 -14895 -943 -14849
rect -569 -14895 -556 -14849
rect -956 -14928 -556 -14895
rect -452 -14849 -52 -14836
rect -452 -14895 -439 -14849
rect -65 -14895 -52 -14849
rect -452 -14928 -52 -14895
rect 52 -14849 452 -14836
rect 52 -14895 65 -14849
rect 439 -14895 452 -14849
rect 52 -14928 452 -14895
rect 556 -14849 956 -14836
rect 556 -14895 569 -14849
rect 943 -14895 956 -14849
rect 556 -14928 956 -14895
rect 1060 -14849 1460 -14836
rect 1060 -14895 1073 -14849
rect 1447 -14895 1460 -14849
rect 1060 -14928 1460 -14895
rect 1564 -14849 1964 -14836
rect 1564 -14895 1577 -14849
rect 1951 -14895 1964 -14849
rect 1564 -14928 1964 -14895
rect 2068 -14849 2468 -14836
rect 2068 -14895 2081 -14849
rect 2455 -14895 2468 -14849
rect 2068 -14928 2468 -14895
rect -2468 -18961 -2068 -18928
rect -2468 -19007 -2455 -18961
rect -2081 -19007 -2068 -18961
rect -2468 -19020 -2068 -19007
rect -1964 -18961 -1564 -18928
rect -1964 -19007 -1951 -18961
rect -1577 -19007 -1564 -18961
rect -1964 -19020 -1564 -19007
rect -1460 -18961 -1060 -18928
rect -1460 -19007 -1447 -18961
rect -1073 -19007 -1060 -18961
rect -1460 -19020 -1060 -19007
rect -956 -18961 -556 -18928
rect -956 -19007 -943 -18961
rect -569 -19007 -556 -18961
rect -956 -19020 -556 -19007
rect -452 -18961 -52 -18928
rect -452 -19007 -439 -18961
rect -65 -19007 -52 -18961
rect -452 -19020 -52 -19007
rect 52 -18961 452 -18928
rect 52 -19007 65 -18961
rect 439 -19007 452 -18961
rect 52 -19020 452 -19007
rect 556 -18961 956 -18928
rect 556 -19007 569 -18961
rect 943 -19007 956 -18961
rect 556 -19020 956 -19007
rect 1060 -18961 1460 -18928
rect 1060 -19007 1073 -18961
rect 1447 -19007 1460 -18961
rect 1060 -19020 1460 -19007
rect 1564 -18961 1964 -18928
rect 1564 -19007 1577 -18961
rect 1951 -19007 1964 -18961
rect 1564 -19020 1964 -19007
rect 2068 -18961 2468 -18928
rect 2068 -19007 2081 -18961
rect 2455 -19007 2468 -18961
rect 2068 -19020 2468 -19007
rect -2468 -19081 -2068 -19068
rect -2468 -19127 -2455 -19081
rect -2081 -19127 -2068 -19081
rect -2468 -19160 -2068 -19127
rect -1964 -19081 -1564 -19068
rect -1964 -19127 -1951 -19081
rect -1577 -19127 -1564 -19081
rect -1964 -19160 -1564 -19127
rect -1460 -19081 -1060 -19068
rect -1460 -19127 -1447 -19081
rect -1073 -19127 -1060 -19081
rect -1460 -19160 -1060 -19127
rect -956 -19081 -556 -19068
rect -956 -19127 -943 -19081
rect -569 -19127 -556 -19081
rect -956 -19160 -556 -19127
rect -452 -19081 -52 -19068
rect -452 -19127 -439 -19081
rect -65 -19127 -52 -19081
rect -452 -19160 -52 -19127
rect 52 -19081 452 -19068
rect 52 -19127 65 -19081
rect 439 -19127 452 -19081
rect 52 -19160 452 -19127
rect 556 -19081 956 -19068
rect 556 -19127 569 -19081
rect 943 -19127 956 -19081
rect 556 -19160 956 -19127
rect 1060 -19081 1460 -19068
rect 1060 -19127 1073 -19081
rect 1447 -19127 1460 -19081
rect 1060 -19160 1460 -19127
rect 1564 -19081 1964 -19068
rect 1564 -19127 1577 -19081
rect 1951 -19127 1964 -19081
rect 1564 -19160 1964 -19127
rect 2068 -19081 2468 -19068
rect 2068 -19127 2081 -19081
rect 2455 -19127 2468 -19081
rect 2068 -19160 2468 -19127
rect -2468 -23193 -2068 -23160
rect -2468 -23239 -2455 -23193
rect -2081 -23239 -2068 -23193
rect -2468 -23252 -2068 -23239
rect -1964 -23193 -1564 -23160
rect -1964 -23239 -1951 -23193
rect -1577 -23239 -1564 -23193
rect -1964 -23252 -1564 -23239
rect -1460 -23193 -1060 -23160
rect -1460 -23239 -1447 -23193
rect -1073 -23239 -1060 -23193
rect -1460 -23252 -1060 -23239
rect -956 -23193 -556 -23160
rect -956 -23239 -943 -23193
rect -569 -23239 -556 -23193
rect -956 -23252 -556 -23239
rect -452 -23193 -52 -23160
rect -452 -23239 -439 -23193
rect -65 -23239 -52 -23193
rect -452 -23252 -52 -23239
rect 52 -23193 452 -23160
rect 52 -23239 65 -23193
rect 439 -23239 452 -23193
rect 52 -23252 452 -23239
rect 556 -23193 956 -23160
rect 556 -23239 569 -23193
rect 943 -23239 956 -23193
rect 556 -23252 956 -23239
rect 1060 -23193 1460 -23160
rect 1060 -23239 1073 -23193
rect 1447 -23239 1460 -23193
rect 1060 -23252 1460 -23239
rect 1564 -23193 1964 -23160
rect 1564 -23239 1577 -23193
rect 1951 -23239 1964 -23193
rect 1564 -23252 1964 -23239
rect 2068 -23193 2468 -23160
rect 2068 -23239 2081 -23193
rect 2455 -23239 2468 -23193
rect 2068 -23252 2468 -23239
<< polycontact >>
rect -2455 23193 -2081 23239
rect -1951 23193 -1577 23239
rect -1447 23193 -1073 23239
rect -943 23193 -569 23239
rect -439 23193 -65 23239
rect 65 23193 439 23239
rect 569 23193 943 23239
rect 1073 23193 1447 23239
rect 1577 23193 1951 23239
rect 2081 23193 2455 23239
rect -2455 19081 -2081 19127
rect -1951 19081 -1577 19127
rect -1447 19081 -1073 19127
rect -943 19081 -569 19127
rect -439 19081 -65 19127
rect 65 19081 439 19127
rect 569 19081 943 19127
rect 1073 19081 1447 19127
rect 1577 19081 1951 19127
rect 2081 19081 2455 19127
rect -2455 18961 -2081 19007
rect -1951 18961 -1577 19007
rect -1447 18961 -1073 19007
rect -943 18961 -569 19007
rect -439 18961 -65 19007
rect 65 18961 439 19007
rect 569 18961 943 19007
rect 1073 18961 1447 19007
rect 1577 18961 1951 19007
rect 2081 18961 2455 19007
rect -2455 14849 -2081 14895
rect -1951 14849 -1577 14895
rect -1447 14849 -1073 14895
rect -943 14849 -569 14895
rect -439 14849 -65 14895
rect 65 14849 439 14895
rect 569 14849 943 14895
rect 1073 14849 1447 14895
rect 1577 14849 1951 14895
rect 2081 14849 2455 14895
rect -2455 14729 -2081 14775
rect -1951 14729 -1577 14775
rect -1447 14729 -1073 14775
rect -943 14729 -569 14775
rect -439 14729 -65 14775
rect 65 14729 439 14775
rect 569 14729 943 14775
rect 1073 14729 1447 14775
rect 1577 14729 1951 14775
rect 2081 14729 2455 14775
rect -2455 10617 -2081 10663
rect -1951 10617 -1577 10663
rect -1447 10617 -1073 10663
rect -943 10617 -569 10663
rect -439 10617 -65 10663
rect 65 10617 439 10663
rect 569 10617 943 10663
rect 1073 10617 1447 10663
rect 1577 10617 1951 10663
rect 2081 10617 2455 10663
rect -2455 10497 -2081 10543
rect -1951 10497 -1577 10543
rect -1447 10497 -1073 10543
rect -943 10497 -569 10543
rect -439 10497 -65 10543
rect 65 10497 439 10543
rect 569 10497 943 10543
rect 1073 10497 1447 10543
rect 1577 10497 1951 10543
rect 2081 10497 2455 10543
rect -2455 6385 -2081 6431
rect -1951 6385 -1577 6431
rect -1447 6385 -1073 6431
rect -943 6385 -569 6431
rect -439 6385 -65 6431
rect 65 6385 439 6431
rect 569 6385 943 6431
rect 1073 6385 1447 6431
rect 1577 6385 1951 6431
rect 2081 6385 2455 6431
rect -2455 6265 -2081 6311
rect -1951 6265 -1577 6311
rect -1447 6265 -1073 6311
rect -943 6265 -569 6311
rect -439 6265 -65 6311
rect 65 6265 439 6311
rect 569 6265 943 6311
rect 1073 6265 1447 6311
rect 1577 6265 1951 6311
rect 2081 6265 2455 6311
rect -2455 2153 -2081 2199
rect -1951 2153 -1577 2199
rect -1447 2153 -1073 2199
rect -943 2153 -569 2199
rect -439 2153 -65 2199
rect 65 2153 439 2199
rect 569 2153 943 2199
rect 1073 2153 1447 2199
rect 1577 2153 1951 2199
rect 2081 2153 2455 2199
rect -2455 2033 -2081 2079
rect -1951 2033 -1577 2079
rect -1447 2033 -1073 2079
rect -943 2033 -569 2079
rect -439 2033 -65 2079
rect 65 2033 439 2079
rect 569 2033 943 2079
rect 1073 2033 1447 2079
rect 1577 2033 1951 2079
rect 2081 2033 2455 2079
rect -2455 -2079 -2081 -2033
rect -1951 -2079 -1577 -2033
rect -1447 -2079 -1073 -2033
rect -943 -2079 -569 -2033
rect -439 -2079 -65 -2033
rect 65 -2079 439 -2033
rect 569 -2079 943 -2033
rect 1073 -2079 1447 -2033
rect 1577 -2079 1951 -2033
rect 2081 -2079 2455 -2033
rect -2455 -2199 -2081 -2153
rect -1951 -2199 -1577 -2153
rect -1447 -2199 -1073 -2153
rect -943 -2199 -569 -2153
rect -439 -2199 -65 -2153
rect 65 -2199 439 -2153
rect 569 -2199 943 -2153
rect 1073 -2199 1447 -2153
rect 1577 -2199 1951 -2153
rect 2081 -2199 2455 -2153
rect -2455 -6311 -2081 -6265
rect -1951 -6311 -1577 -6265
rect -1447 -6311 -1073 -6265
rect -943 -6311 -569 -6265
rect -439 -6311 -65 -6265
rect 65 -6311 439 -6265
rect 569 -6311 943 -6265
rect 1073 -6311 1447 -6265
rect 1577 -6311 1951 -6265
rect 2081 -6311 2455 -6265
rect -2455 -6431 -2081 -6385
rect -1951 -6431 -1577 -6385
rect -1447 -6431 -1073 -6385
rect -943 -6431 -569 -6385
rect -439 -6431 -65 -6385
rect 65 -6431 439 -6385
rect 569 -6431 943 -6385
rect 1073 -6431 1447 -6385
rect 1577 -6431 1951 -6385
rect 2081 -6431 2455 -6385
rect -2455 -10543 -2081 -10497
rect -1951 -10543 -1577 -10497
rect -1447 -10543 -1073 -10497
rect -943 -10543 -569 -10497
rect -439 -10543 -65 -10497
rect 65 -10543 439 -10497
rect 569 -10543 943 -10497
rect 1073 -10543 1447 -10497
rect 1577 -10543 1951 -10497
rect 2081 -10543 2455 -10497
rect -2455 -10663 -2081 -10617
rect -1951 -10663 -1577 -10617
rect -1447 -10663 -1073 -10617
rect -943 -10663 -569 -10617
rect -439 -10663 -65 -10617
rect 65 -10663 439 -10617
rect 569 -10663 943 -10617
rect 1073 -10663 1447 -10617
rect 1577 -10663 1951 -10617
rect 2081 -10663 2455 -10617
rect -2455 -14775 -2081 -14729
rect -1951 -14775 -1577 -14729
rect -1447 -14775 -1073 -14729
rect -943 -14775 -569 -14729
rect -439 -14775 -65 -14729
rect 65 -14775 439 -14729
rect 569 -14775 943 -14729
rect 1073 -14775 1447 -14729
rect 1577 -14775 1951 -14729
rect 2081 -14775 2455 -14729
rect -2455 -14895 -2081 -14849
rect -1951 -14895 -1577 -14849
rect -1447 -14895 -1073 -14849
rect -943 -14895 -569 -14849
rect -439 -14895 -65 -14849
rect 65 -14895 439 -14849
rect 569 -14895 943 -14849
rect 1073 -14895 1447 -14849
rect 1577 -14895 1951 -14849
rect 2081 -14895 2455 -14849
rect -2455 -19007 -2081 -18961
rect -1951 -19007 -1577 -18961
rect -1447 -19007 -1073 -18961
rect -943 -19007 -569 -18961
rect -439 -19007 -65 -18961
rect 65 -19007 439 -18961
rect 569 -19007 943 -18961
rect 1073 -19007 1447 -18961
rect 1577 -19007 1951 -18961
rect 2081 -19007 2455 -18961
rect -2455 -19127 -2081 -19081
rect -1951 -19127 -1577 -19081
rect -1447 -19127 -1073 -19081
rect -943 -19127 -569 -19081
rect -439 -19127 -65 -19081
rect 65 -19127 439 -19081
rect 569 -19127 943 -19081
rect 1073 -19127 1447 -19081
rect 1577 -19127 1951 -19081
rect 2081 -19127 2455 -19081
rect -2455 -23239 -2081 -23193
rect -1951 -23239 -1577 -23193
rect -1447 -23239 -1073 -23193
rect -943 -23239 -569 -23193
rect -439 -23239 -65 -23193
rect 65 -23239 439 -23193
rect 569 -23239 943 -23193
rect 1073 -23239 1447 -23193
rect 1577 -23239 1951 -23193
rect 2081 -23239 2455 -23193
<< metal1 >>
rect -2681 23287 2681 23333
rect -2681 23230 -2635 23287
rect -2466 23193 -2455 23239
rect -2081 23193 -2070 23239
rect -1962 23193 -1951 23239
rect -1577 23193 -1566 23239
rect -1458 23193 -1447 23239
rect -1073 23193 -1062 23239
rect -954 23193 -943 23239
rect -569 23193 -558 23239
rect -450 23193 -439 23239
rect -65 23193 -54 23239
rect 54 23193 65 23239
rect 439 23193 450 23239
rect 558 23193 569 23239
rect 943 23193 954 23239
rect 1062 23193 1073 23239
rect 1447 23193 1458 23239
rect 1566 23193 1577 23239
rect 1951 23193 1962 23239
rect 2070 23193 2081 23239
rect 2455 23193 2466 23239
rect 2635 23230 2681 23287
rect -2543 23147 -2497 23158
rect -2543 19162 -2497 19173
rect -2039 23147 -1993 23158
rect -2039 19162 -1993 19173
rect -1535 23147 -1489 23158
rect -1535 19162 -1489 19173
rect -1031 23147 -985 23158
rect -1031 19162 -985 19173
rect -527 23147 -481 23158
rect -527 19162 -481 19173
rect -23 23147 23 23158
rect -23 19162 23 19173
rect 481 23147 527 23158
rect 481 19162 527 19173
rect 985 23147 1031 23158
rect 985 19162 1031 19173
rect 1489 23147 1535 23158
rect 1489 19162 1535 19173
rect 1993 23147 2039 23158
rect 1993 19162 2039 19173
rect 2497 23147 2543 23158
rect 2497 19162 2543 19173
rect -2466 19081 -2455 19127
rect -2081 19081 -2070 19127
rect -1962 19081 -1951 19127
rect -1577 19081 -1566 19127
rect -1458 19081 -1447 19127
rect -1073 19081 -1062 19127
rect -954 19081 -943 19127
rect -569 19081 -558 19127
rect -450 19081 -439 19127
rect -65 19081 -54 19127
rect 54 19081 65 19127
rect 439 19081 450 19127
rect 558 19081 569 19127
rect 943 19081 954 19127
rect 1062 19081 1073 19127
rect 1447 19081 1458 19127
rect 1566 19081 1577 19127
rect 1951 19081 1962 19127
rect 2070 19081 2081 19127
rect 2455 19081 2466 19127
rect -2466 18961 -2455 19007
rect -2081 18961 -2070 19007
rect -1962 18961 -1951 19007
rect -1577 18961 -1566 19007
rect -1458 18961 -1447 19007
rect -1073 18961 -1062 19007
rect -954 18961 -943 19007
rect -569 18961 -558 19007
rect -450 18961 -439 19007
rect -65 18961 -54 19007
rect 54 18961 65 19007
rect 439 18961 450 19007
rect 558 18961 569 19007
rect 943 18961 954 19007
rect 1062 18961 1073 19007
rect 1447 18961 1458 19007
rect 1566 18961 1577 19007
rect 1951 18961 1962 19007
rect 2070 18961 2081 19007
rect 2455 18961 2466 19007
rect -2543 18915 -2497 18926
rect -2543 14930 -2497 14941
rect -2039 18915 -1993 18926
rect -2039 14930 -1993 14941
rect -1535 18915 -1489 18926
rect -1535 14930 -1489 14941
rect -1031 18915 -985 18926
rect -1031 14930 -985 14941
rect -527 18915 -481 18926
rect -527 14930 -481 14941
rect -23 18915 23 18926
rect -23 14930 23 14941
rect 481 18915 527 18926
rect 481 14930 527 14941
rect 985 18915 1031 18926
rect 985 14930 1031 14941
rect 1489 18915 1535 18926
rect 1489 14930 1535 14941
rect 1993 18915 2039 18926
rect 1993 14930 2039 14941
rect 2497 18915 2543 18926
rect 2497 14930 2543 14941
rect -2466 14849 -2455 14895
rect -2081 14849 -2070 14895
rect -1962 14849 -1951 14895
rect -1577 14849 -1566 14895
rect -1458 14849 -1447 14895
rect -1073 14849 -1062 14895
rect -954 14849 -943 14895
rect -569 14849 -558 14895
rect -450 14849 -439 14895
rect -65 14849 -54 14895
rect 54 14849 65 14895
rect 439 14849 450 14895
rect 558 14849 569 14895
rect 943 14849 954 14895
rect 1062 14849 1073 14895
rect 1447 14849 1458 14895
rect 1566 14849 1577 14895
rect 1951 14849 1962 14895
rect 2070 14849 2081 14895
rect 2455 14849 2466 14895
rect -2466 14729 -2455 14775
rect -2081 14729 -2070 14775
rect -1962 14729 -1951 14775
rect -1577 14729 -1566 14775
rect -1458 14729 -1447 14775
rect -1073 14729 -1062 14775
rect -954 14729 -943 14775
rect -569 14729 -558 14775
rect -450 14729 -439 14775
rect -65 14729 -54 14775
rect 54 14729 65 14775
rect 439 14729 450 14775
rect 558 14729 569 14775
rect 943 14729 954 14775
rect 1062 14729 1073 14775
rect 1447 14729 1458 14775
rect 1566 14729 1577 14775
rect 1951 14729 1962 14775
rect 2070 14729 2081 14775
rect 2455 14729 2466 14775
rect -2543 14683 -2497 14694
rect -2543 10698 -2497 10709
rect -2039 14683 -1993 14694
rect -2039 10698 -1993 10709
rect -1535 14683 -1489 14694
rect -1535 10698 -1489 10709
rect -1031 14683 -985 14694
rect -1031 10698 -985 10709
rect -527 14683 -481 14694
rect -527 10698 -481 10709
rect -23 14683 23 14694
rect -23 10698 23 10709
rect 481 14683 527 14694
rect 481 10698 527 10709
rect 985 14683 1031 14694
rect 985 10698 1031 10709
rect 1489 14683 1535 14694
rect 1489 10698 1535 10709
rect 1993 14683 2039 14694
rect 1993 10698 2039 10709
rect 2497 14683 2543 14694
rect 2497 10698 2543 10709
rect -2466 10617 -2455 10663
rect -2081 10617 -2070 10663
rect -1962 10617 -1951 10663
rect -1577 10617 -1566 10663
rect -1458 10617 -1447 10663
rect -1073 10617 -1062 10663
rect -954 10617 -943 10663
rect -569 10617 -558 10663
rect -450 10617 -439 10663
rect -65 10617 -54 10663
rect 54 10617 65 10663
rect 439 10617 450 10663
rect 558 10617 569 10663
rect 943 10617 954 10663
rect 1062 10617 1073 10663
rect 1447 10617 1458 10663
rect 1566 10617 1577 10663
rect 1951 10617 1962 10663
rect 2070 10617 2081 10663
rect 2455 10617 2466 10663
rect -2466 10497 -2455 10543
rect -2081 10497 -2070 10543
rect -1962 10497 -1951 10543
rect -1577 10497 -1566 10543
rect -1458 10497 -1447 10543
rect -1073 10497 -1062 10543
rect -954 10497 -943 10543
rect -569 10497 -558 10543
rect -450 10497 -439 10543
rect -65 10497 -54 10543
rect 54 10497 65 10543
rect 439 10497 450 10543
rect 558 10497 569 10543
rect 943 10497 954 10543
rect 1062 10497 1073 10543
rect 1447 10497 1458 10543
rect 1566 10497 1577 10543
rect 1951 10497 1962 10543
rect 2070 10497 2081 10543
rect 2455 10497 2466 10543
rect -2543 10451 -2497 10462
rect -2543 6466 -2497 6477
rect -2039 10451 -1993 10462
rect -2039 6466 -1993 6477
rect -1535 10451 -1489 10462
rect -1535 6466 -1489 6477
rect -1031 10451 -985 10462
rect -1031 6466 -985 6477
rect -527 10451 -481 10462
rect -527 6466 -481 6477
rect -23 10451 23 10462
rect -23 6466 23 6477
rect 481 10451 527 10462
rect 481 6466 527 6477
rect 985 10451 1031 10462
rect 985 6466 1031 6477
rect 1489 10451 1535 10462
rect 1489 6466 1535 6477
rect 1993 10451 2039 10462
rect 1993 6466 2039 6477
rect 2497 10451 2543 10462
rect 2497 6466 2543 6477
rect -2466 6385 -2455 6431
rect -2081 6385 -2070 6431
rect -1962 6385 -1951 6431
rect -1577 6385 -1566 6431
rect -1458 6385 -1447 6431
rect -1073 6385 -1062 6431
rect -954 6385 -943 6431
rect -569 6385 -558 6431
rect -450 6385 -439 6431
rect -65 6385 -54 6431
rect 54 6385 65 6431
rect 439 6385 450 6431
rect 558 6385 569 6431
rect 943 6385 954 6431
rect 1062 6385 1073 6431
rect 1447 6385 1458 6431
rect 1566 6385 1577 6431
rect 1951 6385 1962 6431
rect 2070 6385 2081 6431
rect 2455 6385 2466 6431
rect -2466 6265 -2455 6311
rect -2081 6265 -2070 6311
rect -1962 6265 -1951 6311
rect -1577 6265 -1566 6311
rect -1458 6265 -1447 6311
rect -1073 6265 -1062 6311
rect -954 6265 -943 6311
rect -569 6265 -558 6311
rect -450 6265 -439 6311
rect -65 6265 -54 6311
rect 54 6265 65 6311
rect 439 6265 450 6311
rect 558 6265 569 6311
rect 943 6265 954 6311
rect 1062 6265 1073 6311
rect 1447 6265 1458 6311
rect 1566 6265 1577 6311
rect 1951 6265 1962 6311
rect 2070 6265 2081 6311
rect 2455 6265 2466 6311
rect -2543 6219 -2497 6230
rect -2543 2234 -2497 2245
rect -2039 6219 -1993 6230
rect -2039 2234 -1993 2245
rect -1535 6219 -1489 6230
rect -1535 2234 -1489 2245
rect -1031 6219 -985 6230
rect -1031 2234 -985 2245
rect -527 6219 -481 6230
rect -527 2234 -481 2245
rect -23 6219 23 6230
rect -23 2234 23 2245
rect 481 6219 527 6230
rect 481 2234 527 2245
rect 985 6219 1031 6230
rect 985 2234 1031 2245
rect 1489 6219 1535 6230
rect 1489 2234 1535 2245
rect 1993 6219 2039 6230
rect 1993 2234 2039 2245
rect 2497 6219 2543 6230
rect 2497 2234 2543 2245
rect -2466 2153 -2455 2199
rect -2081 2153 -2070 2199
rect -1962 2153 -1951 2199
rect -1577 2153 -1566 2199
rect -1458 2153 -1447 2199
rect -1073 2153 -1062 2199
rect -954 2153 -943 2199
rect -569 2153 -558 2199
rect -450 2153 -439 2199
rect -65 2153 -54 2199
rect 54 2153 65 2199
rect 439 2153 450 2199
rect 558 2153 569 2199
rect 943 2153 954 2199
rect 1062 2153 1073 2199
rect 1447 2153 1458 2199
rect 1566 2153 1577 2199
rect 1951 2153 1962 2199
rect 2070 2153 2081 2199
rect 2455 2153 2466 2199
rect -2466 2033 -2455 2079
rect -2081 2033 -2070 2079
rect -1962 2033 -1951 2079
rect -1577 2033 -1566 2079
rect -1458 2033 -1447 2079
rect -1073 2033 -1062 2079
rect -954 2033 -943 2079
rect -569 2033 -558 2079
rect -450 2033 -439 2079
rect -65 2033 -54 2079
rect 54 2033 65 2079
rect 439 2033 450 2079
rect 558 2033 569 2079
rect 943 2033 954 2079
rect 1062 2033 1073 2079
rect 1447 2033 1458 2079
rect 1566 2033 1577 2079
rect 1951 2033 1962 2079
rect 2070 2033 2081 2079
rect 2455 2033 2466 2079
rect -2543 1987 -2497 1998
rect -2543 -1998 -2497 -1987
rect -2039 1987 -1993 1998
rect -2039 -1998 -1993 -1987
rect -1535 1987 -1489 1998
rect -1535 -1998 -1489 -1987
rect -1031 1987 -985 1998
rect -1031 -1998 -985 -1987
rect -527 1987 -481 1998
rect -527 -1998 -481 -1987
rect -23 1987 23 1998
rect -23 -1998 23 -1987
rect 481 1987 527 1998
rect 481 -1998 527 -1987
rect 985 1987 1031 1998
rect 985 -1998 1031 -1987
rect 1489 1987 1535 1998
rect 1489 -1998 1535 -1987
rect 1993 1987 2039 1998
rect 1993 -1998 2039 -1987
rect 2497 1987 2543 1998
rect 2497 -1998 2543 -1987
rect -2466 -2079 -2455 -2033
rect -2081 -2079 -2070 -2033
rect -1962 -2079 -1951 -2033
rect -1577 -2079 -1566 -2033
rect -1458 -2079 -1447 -2033
rect -1073 -2079 -1062 -2033
rect -954 -2079 -943 -2033
rect -569 -2079 -558 -2033
rect -450 -2079 -439 -2033
rect -65 -2079 -54 -2033
rect 54 -2079 65 -2033
rect 439 -2079 450 -2033
rect 558 -2079 569 -2033
rect 943 -2079 954 -2033
rect 1062 -2079 1073 -2033
rect 1447 -2079 1458 -2033
rect 1566 -2079 1577 -2033
rect 1951 -2079 1962 -2033
rect 2070 -2079 2081 -2033
rect 2455 -2079 2466 -2033
rect -2466 -2199 -2455 -2153
rect -2081 -2199 -2070 -2153
rect -1962 -2199 -1951 -2153
rect -1577 -2199 -1566 -2153
rect -1458 -2199 -1447 -2153
rect -1073 -2199 -1062 -2153
rect -954 -2199 -943 -2153
rect -569 -2199 -558 -2153
rect -450 -2199 -439 -2153
rect -65 -2199 -54 -2153
rect 54 -2199 65 -2153
rect 439 -2199 450 -2153
rect 558 -2199 569 -2153
rect 943 -2199 954 -2153
rect 1062 -2199 1073 -2153
rect 1447 -2199 1458 -2153
rect 1566 -2199 1577 -2153
rect 1951 -2199 1962 -2153
rect 2070 -2199 2081 -2153
rect 2455 -2199 2466 -2153
rect -2543 -2245 -2497 -2234
rect -2543 -6230 -2497 -6219
rect -2039 -2245 -1993 -2234
rect -2039 -6230 -1993 -6219
rect -1535 -2245 -1489 -2234
rect -1535 -6230 -1489 -6219
rect -1031 -2245 -985 -2234
rect -1031 -6230 -985 -6219
rect -527 -2245 -481 -2234
rect -527 -6230 -481 -6219
rect -23 -2245 23 -2234
rect -23 -6230 23 -6219
rect 481 -2245 527 -2234
rect 481 -6230 527 -6219
rect 985 -2245 1031 -2234
rect 985 -6230 1031 -6219
rect 1489 -2245 1535 -2234
rect 1489 -6230 1535 -6219
rect 1993 -2245 2039 -2234
rect 1993 -6230 2039 -6219
rect 2497 -2245 2543 -2234
rect 2497 -6230 2543 -6219
rect -2466 -6311 -2455 -6265
rect -2081 -6311 -2070 -6265
rect -1962 -6311 -1951 -6265
rect -1577 -6311 -1566 -6265
rect -1458 -6311 -1447 -6265
rect -1073 -6311 -1062 -6265
rect -954 -6311 -943 -6265
rect -569 -6311 -558 -6265
rect -450 -6311 -439 -6265
rect -65 -6311 -54 -6265
rect 54 -6311 65 -6265
rect 439 -6311 450 -6265
rect 558 -6311 569 -6265
rect 943 -6311 954 -6265
rect 1062 -6311 1073 -6265
rect 1447 -6311 1458 -6265
rect 1566 -6311 1577 -6265
rect 1951 -6311 1962 -6265
rect 2070 -6311 2081 -6265
rect 2455 -6311 2466 -6265
rect -2466 -6431 -2455 -6385
rect -2081 -6431 -2070 -6385
rect -1962 -6431 -1951 -6385
rect -1577 -6431 -1566 -6385
rect -1458 -6431 -1447 -6385
rect -1073 -6431 -1062 -6385
rect -954 -6431 -943 -6385
rect -569 -6431 -558 -6385
rect -450 -6431 -439 -6385
rect -65 -6431 -54 -6385
rect 54 -6431 65 -6385
rect 439 -6431 450 -6385
rect 558 -6431 569 -6385
rect 943 -6431 954 -6385
rect 1062 -6431 1073 -6385
rect 1447 -6431 1458 -6385
rect 1566 -6431 1577 -6385
rect 1951 -6431 1962 -6385
rect 2070 -6431 2081 -6385
rect 2455 -6431 2466 -6385
rect -2543 -6477 -2497 -6466
rect -2543 -10462 -2497 -10451
rect -2039 -6477 -1993 -6466
rect -2039 -10462 -1993 -10451
rect -1535 -6477 -1489 -6466
rect -1535 -10462 -1489 -10451
rect -1031 -6477 -985 -6466
rect -1031 -10462 -985 -10451
rect -527 -6477 -481 -6466
rect -527 -10462 -481 -10451
rect -23 -6477 23 -6466
rect -23 -10462 23 -10451
rect 481 -6477 527 -6466
rect 481 -10462 527 -10451
rect 985 -6477 1031 -6466
rect 985 -10462 1031 -10451
rect 1489 -6477 1535 -6466
rect 1489 -10462 1535 -10451
rect 1993 -6477 2039 -6466
rect 1993 -10462 2039 -10451
rect 2497 -6477 2543 -6466
rect 2497 -10462 2543 -10451
rect -2466 -10543 -2455 -10497
rect -2081 -10543 -2070 -10497
rect -1962 -10543 -1951 -10497
rect -1577 -10543 -1566 -10497
rect -1458 -10543 -1447 -10497
rect -1073 -10543 -1062 -10497
rect -954 -10543 -943 -10497
rect -569 -10543 -558 -10497
rect -450 -10543 -439 -10497
rect -65 -10543 -54 -10497
rect 54 -10543 65 -10497
rect 439 -10543 450 -10497
rect 558 -10543 569 -10497
rect 943 -10543 954 -10497
rect 1062 -10543 1073 -10497
rect 1447 -10543 1458 -10497
rect 1566 -10543 1577 -10497
rect 1951 -10543 1962 -10497
rect 2070 -10543 2081 -10497
rect 2455 -10543 2466 -10497
rect -2466 -10663 -2455 -10617
rect -2081 -10663 -2070 -10617
rect -1962 -10663 -1951 -10617
rect -1577 -10663 -1566 -10617
rect -1458 -10663 -1447 -10617
rect -1073 -10663 -1062 -10617
rect -954 -10663 -943 -10617
rect -569 -10663 -558 -10617
rect -450 -10663 -439 -10617
rect -65 -10663 -54 -10617
rect 54 -10663 65 -10617
rect 439 -10663 450 -10617
rect 558 -10663 569 -10617
rect 943 -10663 954 -10617
rect 1062 -10663 1073 -10617
rect 1447 -10663 1458 -10617
rect 1566 -10663 1577 -10617
rect 1951 -10663 1962 -10617
rect 2070 -10663 2081 -10617
rect 2455 -10663 2466 -10617
rect -2543 -10709 -2497 -10698
rect -2543 -14694 -2497 -14683
rect -2039 -10709 -1993 -10698
rect -2039 -14694 -1993 -14683
rect -1535 -10709 -1489 -10698
rect -1535 -14694 -1489 -14683
rect -1031 -10709 -985 -10698
rect -1031 -14694 -985 -14683
rect -527 -10709 -481 -10698
rect -527 -14694 -481 -14683
rect -23 -10709 23 -10698
rect -23 -14694 23 -14683
rect 481 -10709 527 -10698
rect 481 -14694 527 -14683
rect 985 -10709 1031 -10698
rect 985 -14694 1031 -14683
rect 1489 -10709 1535 -10698
rect 1489 -14694 1535 -14683
rect 1993 -10709 2039 -10698
rect 1993 -14694 2039 -14683
rect 2497 -10709 2543 -10698
rect 2497 -14694 2543 -14683
rect -2466 -14775 -2455 -14729
rect -2081 -14775 -2070 -14729
rect -1962 -14775 -1951 -14729
rect -1577 -14775 -1566 -14729
rect -1458 -14775 -1447 -14729
rect -1073 -14775 -1062 -14729
rect -954 -14775 -943 -14729
rect -569 -14775 -558 -14729
rect -450 -14775 -439 -14729
rect -65 -14775 -54 -14729
rect 54 -14775 65 -14729
rect 439 -14775 450 -14729
rect 558 -14775 569 -14729
rect 943 -14775 954 -14729
rect 1062 -14775 1073 -14729
rect 1447 -14775 1458 -14729
rect 1566 -14775 1577 -14729
rect 1951 -14775 1962 -14729
rect 2070 -14775 2081 -14729
rect 2455 -14775 2466 -14729
rect -2466 -14895 -2455 -14849
rect -2081 -14895 -2070 -14849
rect -1962 -14895 -1951 -14849
rect -1577 -14895 -1566 -14849
rect -1458 -14895 -1447 -14849
rect -1073 -14895 -1062 -14849
rect -954 -14895 -943 -14849
rect -569 -14895 -558 -14849
rect -450 -14895 -439 -14849
rect -65 -14895 -54 -14849
rect 54 -14895 65 -14849
rect 439 -14895 450 -14849
rect 558 -14895 569 -14849
rect 943 -14895 954 -14849
rect 1062 -14895 1073 -14849
rect 1447 -14895 1458 -14849
rect 1566 -14895 1577 -14849
rect 1951 -14895 1962 -14849
rect 2070 -14895 2081 -14849
rect 2455 -14895 2466 -14849
rect -2543 -14941 -2497 -14930
rect -2543 -18926 -2497 -18915
rect -2039 -14941 -1993 -14930
rect -2039 -18926 -1993 -18915
rect -1535 -14941 -1489 -14930
rect -1535 -18926 -1489 -18915
rect -1031 -14941 -985 -14930
rect -1031 -18926 -985 -18915
rect -527 -14941 -481 -14930
rect -527 -18926 -481 -18915
rect -23 -14941 23 -14930
rect -23 -18926 23 -18915
rect 481 -14941 527 -14930
rect 481 -18926 527 -18915
rect 985 -14941 1031 -14930
rect 985 -18926 1031 -18915
rect 1489 -14941 1535 -14930
rect 1489 -18926 1535 -18915
rect 1993 -14941 2039 -14930
rect 1993 -18926 2039 -18915
rect 2497 -14941 2543 -14930
rect 2497 -18926 2543 -18915
rect -2466 -19007 -2455 -18961
rect -2081 -19007 -2070 -18961
rect -1962 -19007 -1951 -18961
rect -1577 -19007 -1566 -18961
rect -1458 -19007 -1447 -18961
rect -1073 -19007 -1062 -18961
rect -954 -19007 -943 -18961
rect -569 -19007 -558 -18961
rect -450 -19007 -439 -18961
rect -65 -19007 -54 -18961
rect 54 -19007 65 -18961
rect 439 -19007 450 -18961
rect 558 -19007 569 -18961
rect 943 -19007 954 -18961
rect 1062 -19007 1073 -18961
rect 1447 -19007 1458 -18961
rect 1566 -19007 1577 -18961
rect 1951 -19007 1962 -18961
rect 2070 -19007 2081 -18961
rect 2455 -19007 2466 -18961
rect -2466 -19127 -2455 -19081
rect -2081 -19127 -2070 -19081
rect -1962 -19127 -1951 -19081
rect -1577 -19127 -1566 -19081
rect -1458 -19127 -1447 -19081
rect -1073 -19127 -1062 -19081
rect -954 -19127 -943 -19081
rect -569 -19127 -558 -19081
rect -450 -19127 -439 -19081
rect -65 -19127 -54 -19081
rect 54 -19127 65 -19081
rect 439 -19127 450 -19081
rect 558 -19127 569 -19081
rect 943 -19127 954 -19081
rect 1062 -19127 1073 -19081
rect 1447 -19127 1458 -19081
rect 1566 -19127 1577 -19081
rect 1951 -19127 1962 -19081
rect 2070 -19127 2081 -19081
rect 2455 -19127 2466 -19081
rect -2543 -19173 -2497 -19162
rect -2543 -23158 -2497 -23147
rect -2039 -19173 -1993 -19162
rect -2039 -23158 -1993 -23147
rect -1535 -19173 -1489 -19162
rect -1535 -23158 -1489 -23147
rect -1031 -19173 -985 -19162
rect -1031 -23158 -985 -23147
rect -527 -19173 -481 -19162
rect -527 -23158 -481 -23147
rect -23 -19173 23 -19162
rect -23 -23158 23 -23147
rect 481 -19173 527 -19162
rect 481 -23158 527 -23147
rect 985 -19173 1031 -19162
rect 985 -23158 1031 -23147
rect 1489 -19173 1535 -19162
rect 1489 -23158 1535 -23147
rect 1993 -19173 2039 -19162
rect 1993 -23158 2039 -23147
rect 2497 -19173 2543 -19162
rect 2497 -23158 2543 -23147
rect -2681 -23287 -2635 -23230
rect -2466 -23239 -2455 -23193
rect -2081 -23239 -2070 -23193
rect -1962 -23239 -1951 -23193
rect -1577 -23239 -1566 -23193
rect -1458 -23239 -1447 -23193
rect -1073 -23239 -1062 -23193
rect -954 -23239 -943 -23193
rect -569 -23239 -558 -23193
rect -450 -23239 -439 -23193
rect -65 -23239 -54 -23193
rect 54 -23239 65 -23193
rect 439 -23239 450 -23193
rect 558 -23239 569 -23193
rect 943 -23239 954 -23193
rect 1062 -23239 1073 -23193
rect 1447 -23239 1458 -23193
rect 1566 -23239 1577 -23193
rect 1951 -23239 1962 -23193
rect 2070 -23239 2081 -23193
rect 2455 -23239 2466 -23193
rect 2635 -23287 2681 -23230
rect -2681 -23333 2681 -23287
<< properties >>
string FIXED_BBOX -2658 -23310 2658 23310
string gencell nfet_03v3
string library gf180mcu
string parameters w 20.0 l 2.0 m 11 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
