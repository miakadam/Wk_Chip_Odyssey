magic
tech gf180mcuD
magscale 1 10
timestamp 1755256602
<< error_p >>
rect -34 133 -23 179
rect 23 133 34 144
rect -80 -98 -57 -87
rect 57 -98 80 -87
rect -34 -179 -23 -133
<< pwell >>
rect -278 -310 278 310
<< nmos >>
rect -28 -100 28 100
<< ndiff >>
rect -116 87 -28 100
rect -116 -87 -103 87
rect -57 -87 -28 87
rect -116 -100 -28 -87
rect 28 87 116 100
rect 28 -87 57 87
rect 103 -87 116 87
rect 28 -100 116 -87
<< ndiffc >>
rect -103 -87 -57 87
rect 57 -87 103 87
<< psubdiff >>
rect -254 214 254 286
rect -254 170 -182 214
rect -254 -170 -241 170
rect -195 -170 -182 170
rect 182 170 254 214
rect -254 -214 -182 -170
rect 182 -170 195 170
rect 241 -170 254 170
rect 182 -214 254 -170
rect -254 -286 254 -214
<< psubdiffcont >>
rect -241 -170 -195 170
rect 195 -170 241 170
<< polysilicon >>
rect -36 179 36 192
rect -36 133 -23 179
rect 23 133 36 179
rect -36 120 36 133
rect -28 100 28 120
rect -28 -120 28 -100
rect -36 -133 36 -120
rect -36 -179 -23 -133
rect 23 -179 36 -133
rect -36 -192 36 -179
<< polycontact >>
rect -23 133 23 179
rect -23 -179 23 -133
<< metal1 >>
rect -241 227 241 273
rect -241 170 -195 227
rect -34 133 -23 179
rect 23 133 34 179
rect 195 170 241 227
rect -103 87 -57 98
rect -103 -98 -57 -87
rect 57 87 103 98
rect 57 -98 103 -87
rect -241 -227 -195 -170
rect -34 -179 -23 -133
rect 23 -179 34 -133
rect 195 -227 241 -170
rect -241 -273 241 -227
<< properties >>
string FIXED_BBOX -218 -250 218 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
