magic
tech gf180mcuD
magscale 1 10
timestamp 1757925391
<< nwell >>
rect 1290 -140 1890 880
rect 2178 -140 2778 880
<< pwell >>
rect 1290 -860 2778 -240
<< nmos >>
rect 1540 -650 1640 -450
rect 1744 -650 1844 -450
rect 2224 -650 2324 -450
rect 2428 -650 2528 -450
<< pmos >>
rect 1540 70 1640 670
rect 2428 70 2528 670
<< ndiff >>
rect 1452 -463 1540 -450
rect 1452 -637 1465 -463
rect 1511 -637 1540 -463
rect 1452 -650 1540 -637
rect 1640 -463 1744 -450
rect 1640 -637 1669 -463
rect 1715 -637 1744 -463
rect 1640 -650 1744 -637
rect 1844 -463 1932 -450
rect 1844 -637 1873 -463
rect 1919 -637 1932 -463
rect 1844 -650 1932 -637
rect 2136 -463 2224 -450
rect 2136 -637 2149 -463
rect 2195 -637 2224 -463
rect 2136 -650 2224 -637
rect 2324 -463 2428 -450
rect 2324 -637 2353 -463
rect 2399 -637 2428 -463
rect 2324 -650 2428 -637
rect 2528 -463 2616 -450
rect 2528 -637 2557 -463
rect 2603 -637 2616 -463
rect 2528 -650 2616 -637
<< pdiff >>
rect 1452 657 1540 670
rect 1452 83 1465 657
rect 1511 83 1540 657
rect 1452 70 1540 83
rect 1640 657 1728 670
rect 1640 83 1669 657
rect 1715 83 1728 657
rect 1640 70 1728 83
rect 2340 657 2428 670
rect 2340 83 2353 657
rect 2399 83 2428 657
rect 2340 70 2428 83
rect 2528 657 2616 670
rect 2528 83 2557 657
rect 2603 83 2616 657
rect 2528 70 2616 83
<< ndiffc >>
rect 1465 -637 1511 -463
rect 1669 -637 1715 -463
rect 1873 -637 1919 -463
rect 2149 -637 2195 -463
rect 2353 -637 2399 -463
rect 2557 -637 2603 -463
<< pdiffc >>
rect 1465 83 1511 657
rect 1669 83 1715 657
rect 2353 83 2399 657
rect 2557 83 2603 657
<< psubdiff >>
rect 1314 -336 2754 -264
rect 1314 -380 1386 -336
rect 1314 -720 1327 -380
rect 1373 -720 1386 -380
rect 1998 -380 2070 -336
rect 1314 -764 1386 -720
rect 1998 -720 2011 -380
rect 2057 -720 2070 -380
rect 2682 -380 2754 -336
rect 1998 -764 2070 -720
rect 2682 -720 2695 -380
rect 2741 -720 2754 -380
rect 2682 -764 2754 -720
rect 1314 -836 2754 -764
<< nsubdiff >>
rect 1314 784 1866 856
rect 1314 740 1386 784
rect 1314 0 1327 740
rect 1373 0 1386 740
rect 1794 740 1866 784
rect 1314 -44 1386 0
rect 1794 0 1807 740
rect 1853 0 1866 740
rect 1794 -44 1866 0
rect 1314 -116 1866 -44
rect 2202 784 2754 856
rect 2202 740 2274 784
rect 2202 0 2215 740
rect 2261 0 2274 740
rect 2682 740 2754 784
rect 2202 -44 2274 0
rect 2682 0 2695 740
rect 2741 0 2754 740
rect 2682 -44 2754 0
rect 2202 -116 2754 -44
<< psubdiffcont >>
rect 1327 -720 1373 -380
rect 2011 -720 2057 -380
rect 2695 -720 2741 -380
<< nsubdiffcont >>
rect 1327 0 1373 740
rect 1807 0 1853 740
rect 2215 0 2261 740
rect 2695 0 2741 740
<< polysilicon >>
rect 1540 749 1640 762
rect 1540 703 1553 749
rect 1627 703 1640 749
rect 1540 670 1640 703
rect 1540 37 1640 70
rect 1540 -9 1553 37
rect 1627 -9 1640 37
rect 1540 -22 1640 -9
rect 2428 749 2528 762
rect 2428 703 2441 749
rect 2515 703 2528 749
rect 2428 670 2528 703
rect 2428 37 2528 70
rect 2428 -9 2441 37
rect 2515 -9 2528 37
rect 2428 -22 2528 -9
rect 1540 -371 1640 -358
rect 1540 -417 1553 -371
rect 1627 -417 1640 -371
rect 1540 -450 1640 -417
rect 1744 -371 1844 -358
rect 1744 -417 1757 -371
rect 1831 -417 1844 -371
rect 1744 -450 1844 -417
rect 1540 -683 1640 -650
rect 1540 -729 1553 -683
rect 1627 -729 1640 -683
rect 1540 -742 1640 -729
rect 1744 -683 1844 -650
rect 1744 -729 1757 -683
rect 1831 -729 1844 -683
rect 1744 -742 1844 -729
rect 2224 -371 2324 -358
rect 2224 -417 2237 -371
rect 2311 -417 2324 -371
rect 2224 -450 2324 -417
rect 2428 -371 2528 -358
rect 2428 -417 2441 -371
rect 2515 -417 2528 -371
rect 2428 -450 2528 -417
rect 2224 -683 2324 -650
rect 2224 -729 2237 -683
rect 2311 -729 2324 -683
rect 2224 -742 2324 -729
rect 2428 -683 2528 -650
rect 2428 -729 2441 -683
rect 2515 -729 2528 -683
rect 2428 -742 2528 -729
<< polycontact >>
rect 1553 703 1627 749
rect 1553 -9 1627 37
rect 2441 703 2515 749
rect 2441 -9 2515 37
rect 1553 -417 1627 -371
rect 1757 -417 1831 -371
rect 1553 -729 1627 -683
rect 1757 -729 1831 -683
rect 2237 -417 2311 -371
rect 2441 -417 2515 -371
rect 2237 -729 2311 -683
rect 2441 -729 2515 -683
<< metal1 >>
rect 1290 880 2778 1080
rect 1327 740 1373 751
rect 1542 749 1638 780
rect 1542 703 1553 749
rect 1627 703 1638 749
rect 1807 740 2261 880
rect 1465 657 1511 668
rect 1448 373 1465 383
rect 1669 657 1807 668
rect 1511 373 1528 383
rect 1448 133 1460 373
rect 1516 133 1528 373
rect 1448 123 1465 133
rect 1511 123 1528 133
rect 1465 72 1511 83
rect 1715 83 1807 657
rect 1669 72 1807 83
rect 1327 -11 1373 0
rect 1542 -9 1553 37
rect 1627 -9 1638 37
rect 1542 -84 1638 -9
rect 1853 72 2215 740
rect 1807 -11 1853 0
rect 2430 749 2526 780
rect 2430 703 2441 749
rect 2515 703 2526 749
rect 2695 740 2741 751
rect 2261 657 2399 668
rect 2261 83 2353 657
rect 2557 657 2603 668
rect 2540 373 2557 383
rect 2603 373 2620 383
rect 2540 133 2552 373
rect 2608 133 2620 373
rect 2540 123 2557 133
rect 2261 72 2399 83
rect 2603 123 2620 133
rect 2557 72 2603 83
rect 2215 -11 2261 0
rect 2430 -9 2441 37
rect 2515 -9 2526 37
rect 1542 -140 1562 -84
rect 1618 -140 1638 -84
rect 1542 -358 1638 -140
rect 2430 -228 2526 -9
rect 2695 -11 2741 0
rect 2362 -240 2526 -228
rect 2362 -296 2374 -240
rect 2430 -296 2526 -240
rect 2362 -308 2526 -296
rect 2430 -358 2526 -308
rect 1327 -380 1373 -369
rect 1542 -371 1842 -358
rect 1542 -417 1553 -371
rect 1627 -404 1757 -371
rect 1627 -417 1638 -404
rect 1746 -417 1757 -404
rect 1831 -417 1842 -371
rect 2011 -380 2057 -369
rect 1373 -463 1511 -452
rect 1373 -637 1465 -463
rect 1669 -463 1715 -452
rect 1652 -522 1669 -512
rect 1873 -463 2011 -452
rect 1715 -522 1732 -512
rect 1652 -578 1664 -522
rect 1720 -578 1732 -522
rect 1652 -588 1669 -578
rect 1373 -648 1511 -637
rect 1715 -588 1732 -578
rect 1669 -648 1715 -637
rect 1919 -637 2011 -463
rect 1873 -648 2011 -637
rect 1327 -860 1373 -720
rect 1542 -729 1553 -683
rect 1627 -729 1638 -683
rect 1542 -760 1638 -729
rect 1746 -729 1757 -683
rect 1831 -729 1842 -683
rect 1746 -760 1842 -729
rect 2226 -371 2526 -358
rect 2226 -417 2237 -371
rect 2311 -404 2441 -371
rect 2311 -417 2322 -404
rect 2430 -417 2441 -404
rect 2515 -417 2526 -371
rect 2695 -380 2741 -369
rect 2149 -463 2195 -452
rect 2132 -522 2149 -512
rect 2353 -463 2399 -452
rect 2195 -522 2212 -512
rect 2132 -578 2144 -522
rect 2200 -578 2212 -522
rect 2132 -588 2149 -578
rect 2195 -588 2212 -578
rect 2336 -522 2353 -512
rect 2557 -463 2603 -452
rect 2399 -522 2416 -512
rect 2336 -578 2348 -522
rect 2404 -578 2416 -522
rect 2336 -588 2353 -578
rect 2149 -648 2195 -637
rect 2399 -588 2416 -578
rect 2540 -522 2557 -512
rect 2603 -522 2620 -512
rect 2540 -578 2552 -522
rect 2608 -578 2620 -522
rect 2540 -588 2557 -578
rect 2353 -648 2399 -637
rect 2603 -588 2620 -578
rect 2557 -648 2603 -637
rect 2011 -860 2057 -720
rect 2226 -729 2237 -683
rect 2311 -729 2322 -683
rect 2226 -760 2322 -729
rect 2430 -729 2441 -683
rect 2515 -729 2526 -683
rect 2430 -760 2526 -729
rect 2695 -860 2741 -720
rect 1290 -1060 2778 -860
<< via1 >>
rect 1460 133 1465 373
rect 1465 133 1511 373
rect 1511 133 1516 373
rect 2552 133 2557 373
rect 2557 133 2603 373
rect 2603 133 2608 373
rect 1562 -140 1618 -84
rect 2374 -296 2430 -240
rect 1664 -578 1669 -522
rect 1669 -578 1715 -522
rect 1715 -578 1720 -522
rect 2144 -578 2149 -522
rect 2149 -578 2195 -522
rect 2195 -578 2200 -522
rect 2348 -578 2353 -522
rect 2353 -578 2399 -522
rect 2399 -578 2404 -522
rect 2552 -578 2557 -522
rect 2557 -578 2603 -522
rect 2603 -578 2608 -522
<< metal2 >>
rect 1448 373 2620 383
rect 1448 133 1460 373
rect 1516 133 2552 373
rect 2608 133 2620 373
rect 1448 123 2620 133
rect 1542 -84 1620 -72
rect 1203 -140 1562 -84
rect 1618 -140 1620 -84
rect 1542 -152 1620 -140
rect 2540 -162 2620 123
rect 2540 -218 2778 -162
rect 2362 -240 2432 -228
rect 1203 -296 2374 -240
rect 2430 -296 2432 -240
rect 2362 -308 2432 -296
rect 1652 -522 1732 -512
rect 1652 -578 1664 -522
rect 1720 -578 1732 -522
rect 1652 -764 1732 -578
rect 2132 -522 2212 -512
rect 2132 -578 2144 -522
rect 2200 -578 2212 -522
rect 2132 -588 2212 -578
rect 2336 -522 2416 -512
rect 2336 -578 2348 -522
rect 2404 -578 2416 -522
rect 2336 -764 2416 -578
rect 2540 -522 2620 -218
rect 2540 -578 2552 -522
rect 2608 -578 2620 -522
rect 2540 -588 2620 -578
rect 1652 -836 2416 -764
<< via2 >>
rect 2144 -578 2200 -522
rect 2552 -578 2608 -522
<< metal3 >>
rect 2132 -522 2620 -512
rect 2132 -578 2144 -522
rect 2200 -578 2552 -522
rect 2608 -578 2620 -522
rect 2132 -588 2620 -578
<< labels >>
rlabel metal1 2026 1080 2026 1080 1 VDD
port 0 n
rlabel metal2 2778 -190 2778 -190 3 OUT
port 1 e
rlabel metal2 1203 -271 1203 -271 7 A
port 2 w
rlabel metal2 1203 -113 1203 -113 7 B
port 3 w
rlabel metal1 2035 -1060 2035 -1060 5 VSS
port 4 s
<< end >>
