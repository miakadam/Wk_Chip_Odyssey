* NGSPICE file created from nand3_1.ext - technology: gf180mcuD

.subckt nand3_1 A B Y VDD VSS C
X0 a_390_210# B a_280_210# VSS nfet_03v3 ad=0.10625p pd=1.1u as=0.10625p ps=1.1u w=0.85u l=0.3u
X1 Y A VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 VDD B Y VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X3 VSS C a_390_210# VSS nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X4 Y C VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 a_280_210# A Y VSS nfet_03v3 ad=0.10625p pd=1.1u as=0.425p ps=2.7u w=0.85u l=0.3u
.ends

