* NGSPICE file created from SARlogic.ext - technology: (null)

.subckt SARlogic vdd vss clk reset comp_in d5 d4 d3 d2 d1 d0
X0 dffrs_5.Qb.t1 reset.t0 a_26858_2649 vss.t304 nfet_03v3
**devattr s=10400,304 d=17600,576
X1 a_1150_7058 dffrs_13.nand3_8.Z.t4 a_966_7058 vss.t45 nfet_03v3
**devattr s=10400,304 d=10400,304
X2 vdd.t67 dffrs_12.nand3_8.Z dffrs_12.nand3_1.C vdd.t66 pfet_03v3
**devattr s=26000,604 d=26000,604
X3 dffrs_5.nand3_1.C.t1 dffrs_5.nand3_6.C.t4 a_25372_7058 vss.t216 nfet_03v3
**devattr s=10400,304 d=17600,576
X4 a_14732_12225 dffrs_8.nand3_8.C.t4 a_14548_12225 vss.t48 nfet_03v3
**devattr s=10400,304 d=10400,304
X5 dffrs_10.nand3_8.C.t1 dffrs_10.nand3_8.Z a_21330_12224 vss.t192 nfet_03v3
**devattr s=10400,304 d=17600,576
X6 vdd.t158 dffrs_12.Q.t4 dffrs_11.nand3_8.C.t0 vdd.t157 pfet_03v3
**devattr s=26000,604 d=26000,604
X7 a_9020_4853 dffrs_1.nand3_1.C.t4 vss.t115 vss.t114 nfet_03v3
**devattr s=17600,576 d=10400,304
X8 d2.t2 dffrs_2.Qb.t4 vdd.t178 vdd.t177 pfet_03v3
**devattr s=44000,1176 d=26000,604
X9 a_18774_14429 dffrs_9.nand3_6.C.t4 a_18590_14429 vss.t218 nfet_03v3
**devattr s=10400,304 d=10400,304
X10 dffrs_10.nand3_6.C.t1 d0.t4 a_21330_14429 vss.t226 nfet_03v3
**devattr s=10400,304 d=17600,576
X11 a_22632_14429 dffrs_3.Qb.t4 vss.t308 vss.t307 nfet_03v3
**devattr s=17600,576 d=10400,304
X12 vdd.t454 reset.t1 dffrs_11.nand3_6.C.t3 vdd.t453 pfet_03v3
**devattr s=26000,604 d=26000,604
X13 dffrs_4.nand3_6.C.t1 clk.t0 a_21330_4853 vss.t92 nfet_03v3
**devattr s=10400,304 d=17600,576
X14 a_13246_16634 dffrs_8.nand3_8.Z a_13062_16634 vss.t178 nfet_03v3
**devattr s=10400,304 d=10400,304
X15 a_13062_16634 dffrs_1.Qb.t4 vss.t117 vss.t116 nfet_03v3
**devattr s=17600,576 d=10400,304
X16 dffrs_12.nand3_8.C.t0 dffrs_12.nand3_8.Z a_29414_12224 vss.t54 nfet_03v3
**devattr s=10400,304 d=17600,576
X17 a_6648_14432 dffrs_14.nand3_6.C.t4 a_6464_14432 vss.t134 nfet_03v3
**devattr s=10400,304 d=10400,304
X18 dffrs_13.nand3_6.C.t1 clk.t1 a_1150_4853 vss.t93 nfet_03v3
**devattr s=10400,304 d=17600,576
X19 dffrs_12.nand3_6.C.t1 vss.t214 a_29414_14429 vss.t215 nfet_03v3
**devattr s=10400,304 d=17600,576
X20 dffrs_4.Q.t3 dffrs_4.Qb.t4 a_22816_4853 vss.t11 nfet_03v3
**devattr s=10400,304 d=17600,576
X21 a_25188_16634 dffrs_4.Qb.t5 vss.t13 vss.t12 nfet_03v3
**devattr s=17600,576 d=10400,304
X22 dffrs_11.nand3_8.Z comp_in.t0 a_25372_10019 vss.t231 nfet_03v3
**devattr s=10400,304 d=17600,576
X23 a_21146_12224 dffrs_10.nand3_6.C.t4 vss.t322 vss.t321 nfet_03v3
**devattr s=17600,576 d=10400,304
X24 dffrs_7.nand3_8.C.t0 dffrs_7.nand3_8.Z vdd.t49 vdd.t48 pfet_03v3
**devattr s=26000,604 d=44000,1176
X25 dffrs_0.d.t0 dffrs_13.Qb.t4 a_2636_4853 vss.t242 nfet_03v3
**devattr s=10400,304 d=17600,576
X26 dffrs_9.nand3_8.C.t3 dffrs_9.nand3_6.C.t5 vdd.t320 vdd.t319 pfet_03v3
**devattr s=44000,1176 d=26000,604
X27 vdd.t138 dffrs_0.nand3_6.C.t4 dffrs_0.Q.t2 vdd.t137 pfet_03v3
**devattr s=26000,604 d=26000,604
X28 dffrs_7.nand3_6.C.t0 d3.t4 vdd.t350 vdd.t349 pfet_03v3
**devattr s=26000,604 d=44000,1176
X29 dffrs_9.nand3_6.C.t0 dffrs_9.nand3_1.C vdd.t63 vdd.t62 pfet_03v3
**devattr s=44000,1176 d=26000,604
X30 a_21146_14429 dffrs_10.nand3_1.C vss.t32 vss.t31 nfet_03v3
**devattr s=17600,576 d=10400,304
X31 dffrs_5.Q.t1 vdd.t126 vdd.t128 vdd.t127 pfet_03v3
**devattr s=44000,1176 d=26000,604
X32 dffrs_2.nand3_6.C.t0 clk.t2 vdd.t166 vdd.t165 pfet_03v3
**devattr s=26000,604 d=44000,1176
X33 dffrs_1.nand3_6.C.t0 clk.t3 vdd.t482 vdd.t481 pfet_03v3
**devattr s=26000,604 d=44000,1176
X34 a_966_443 dffrs_13.nand3_8.C.t4 vss.t1 vss.t0 nfet_03v3
**devattr s=17600,576 d=10400,304
X35 a_6648_12228 dffrs_14.nand3_8.C.t4 a_6464_12228 vss.t207 nfet_03v3
**devattr s=10400,304 d=10400,304
X36 dffrs_0.nand3_8.Z.t1 dffrs_0.d.t4 vdd.t152 vdd.t151 pfet_03v3
**devattr s=26000,604 d=44000,1176
X37 dffrs_2.nand3_1.C.t2 dffrs_2.nand3_6.C.t4 vdd.t9 vdd.t8 pfet_03v3
**devattr s=26000,604 d=44000,1176
X38 dffrs_4.Qb.t1 reset.t2 a_22816_2649 vss.t303 nfet_03v3
**devattr s=10400,304 d=17600,576
X39 vdd.t452 reset.t3 dffrs_3.nand3_8.Z.t3 vdd.t451 pfet_03v3
**devattr s=26000,604 d=26000,604
X40 dffrs_1.nand3_1.C.t3 dffrs_1.nand3_6.C.t4 vdd.t458 vdd.t457 pfet_03v3
**devattr s=26000,604 d=44000,1176
X41 vdd.t450 reset.t4 dffrs_5.nand3_8.Z.t3 vdd.t449 pfet_03v3
**devattr s=26000,604 d=26000,604
X42 a_4978_14432 dffrs_14.nand3_1.C vss.t66 vss.t65 nfet_03v3
**devattr s=17600,576 d=10400,304
X43 a_9020_7058 vdd.t519 vss.t183 vss.t182 nfet_03v3
**devattr s=17600,576 d=10400,304
X44 dffrs_0.nand3_8.C.t1 dffrs_0.nand3_8.Z.t4 vdd.t366 vdd.t365 pfet_03v3
**devattr s=26000,604 d=44000,1176
X45 a_17288_10019 reset.t5 a_17104_10019 vss.t302 nfet_03v3
**devattr s=10400,304 d=10400,304
X46 dffrs_13.Qb.t2 vdd.t520 a_2636_2649 vss.t184 nfet_03v3
**devattr s=10400,304 d=17600,576
X47 vdd.t484 clk.t4 dffrs_3.nand3_8.C.t3 vdd.t483 pfet_03v3
**devattr s=26000,604 d=26000,604
X48 a_4978_4853 dffrs_0.nand3_1.C.t4 vss.t237 vss.t236 nfet_03v3
**devattr s=17600,576 d=10400,304
X49 dffrs_10.Qb reset.t6 vdd.t448 vdd.t447 pfet_03v3
**devattr s=26000,604 d=44000,1176
X50 dffrs_12.Q.t1 dffrs_12.Qb vdd.t270 vdd.t269 pfet_03v3
**devattr s=26000,604 d=44000,1176
X51 vdd.t486 clk.t5 dffrs_5.nand3_8.C.t1 vdd.t485 pfet_03v3
**devattr s=26000,604 d=26000,604
X52 dffrs_4.nand3_1.C.t0 dffrs_4.nand3_6.C.t4 a_21330_7058 vss.t133 nfet_03v3
**devattr s=10400,304 d=17600,576
X53 a_4978_16637 dffrs_13.Qb.t5 vss.t77 vss.t76 nfet_03v3
**devattr s=17600,576 d=10400,304
X54 vdd.t188 dffrs_0.nand3_8.C.t4 dffrs_0.Qb.t0 vdd.t187 pfet_03v3
**devattr s=26000,604 d=26000,604
X55 vdd.t170 dffrs_12.nand3_6.C.t4 dffrs_12.Q.t0 vdd.t169 pfet_03v3
**devattr s=26000,604 d=26000,604
X56 dffrs_5.nand3_8.Z.t1 dffrs_4.Q.t4 a_25372_443 vss.t71 nfet_03v3
**devattr s=10400,304 d=17600,576
X57 d0.t0 dffrs_11.Qb vdd.t3 vdd.t2 pfet_03v3
**devattr s=26000,604 d=44000,1176
X58 dffrs_5.Qb.t0 dffrs_5.Q.t4 vdd.t21 vdd.t20 pfet_03v3
**devattr s=44000,1176 d=26000,604
X59 dffrs_13.nand3_1.C.t0 dffrs_13.nand3_6.C.t4 a_1150_7058 vss.t7 nfet_03v3
**devattr s=10400,304 d=17600,576
X60 dffrs_10.nand3_1.C dffrs_10.nand3_6.C.t5 vdd.t468 vdd.t467 pfet_03v3
**devattr s=26000,604 d=44000,1176
X61 a_21330_443 reset.t7 a_21146_443 vss.t301 nfet_03v3
**devattr s=10400,304 d=10400,304
X62 vdd.t456 dffrs_7.nand3_6.C.t4 d4.t3 vdd.t455 pfet_03v3
**devattr s=26000,604 d=26000,604
X63 d4.t1 dffrs_7.Qb a_10690_14429 vss.t36 nfet_03v3
**devattr s=10400,304 d=17600,576
X64 a_9020_443 dffrs_1.nand3_8.C.t4 vss.t82 vss.t81 nfet_03v3
**devattr s=17600,576 d=10400,304
X65 dffrs_1.nand3_8.Z.t3 dffrs_0.Q.t4 a_9204_443 vss.t199 nfet_03v3
**devattr s=10400,304 d=17600,576
X66 dffrs_12.nand3_1.C dffrs_12.nand3_6.C.t5 vdd.t504 vdd.t503 pfet_03v3
**devattr s=26000,604 d=44000,1176
X67 dffrs_4.nand3_6.C.t2 dffrs_4.nand3_1.C.t4 vdd.t244 vdd.t243 pfet_03v3
**devattr s=44000,1176 d=26000,604
X68 dffrs_8.Qb reset.t8 a_14732_12225 vss.t300 nfet_03v3
**devattr s=10400,304 d=17600,576
X69 dffrs_10.Qb d1.t4 vdd.t246 vdd.t245 pfet_03v3
**devattr s=44000,1176 d=26000,604
X70 vdd.t446 reset.t9 dffrs_8.nand3_8.Z vdd.t445 pfet_03v3
**devattr s=26000,604 d=26000,604
X71 dffrs_11.nand3_8.C.t3 dffrs_11.nand3_8.Z vdd.t274 vdd.t273 pfet_03v3
**devattr s=26000,604 d=44000,1176
X72 vdd.t73 dffrs_9.nand3_8.C.t4 dffrs_9.Qb vdd.t72 pfet_03v3
**devattr s=26000,604 d=26000,604
X73 dffrs_4.nand3_1.C.t2 vdd.t123 vdd.t125 vdd.t124 pfet_03v3
**devattr s=44000,1176 d=26000,604
X74 dffrs_8.nand3_8.Z dffrs_8.nand3_8.C.t5 vdd.t61 vdd.t60 pfet_03v3
**devattr s=44000,1176 d=26000,604
X75 d0.t2 dffrs_4.Qb.t6 vdd.t13 vdd.t12 pfet_03v3
**devattr s=44000,1176 d=26000,604
X76 d2.t0 dffrs_9.Qb a_18774_14429 vss.t30 nfet_03v3
**devattr s=10400,304 d=17600,576
X77 a_22816_14429 dffrs_10.nand3_6.C.t6 a_22632_14429 vss.t314 nfet_03v3
**devattr s=10400,304 d=10400,304
X78 dffrs_11.nand3_6.C.t1 dffrs_12.Q.t5 vdd.t77 vdd.t76 pfet_03v3
**devattr s=26000,604 d=44000,1176
X79 a_18774_4853 dffrs_3.nand3_6.C.t4 a_18590_4853 vss.t8 nfet_03v3
**devattr s=10400,304 d=10400,304
X80 a_29230_16634 dffrs_5.Qb.t4 vss.t250 vss.t249 nfet_03v3
**devattr s=17600,576 d=10400,304
X81 dffrs_4.Q.t1 vdd.t120 vdd.t122 vdd.t121 pfet_03v3
**devattr s=44000,1176 d=26000,604
X82 dffrs_10.nand3_1.C dffrs_3.Qb.t5 vdd.t464 vdd.t463 pfet_03v3
**devattr s=44000,1176 d=26000,604
X83 a_25188_443 dffrs_5.nand3_8.C.t4 vss.t339 vss.t338 nfet_03v3
**devattr s=17600,576 d=10400,304
X84 dffrs_11.nand3_8.Z dffrs_11.nand3_8.C.t4 vdd.t474 vdd.t473 pfet_03v3
**devattr s=44000,1176 d=26000,604
X85 a_9204_2648 clk.t6 a_9020_2648 vss.t323 nfet_03v3
**devattr s=10400,304 d=10400,304
X86 dffrs_2.d.t2 dffrs_1.Qb.t5 vdd.t204 vdd.t203 pfet_03v3
**devattr s=26000,604 d=44000,1176
X87 dffrs_0.d.t3 reset.t10 vdd.t444 vdd.t443 pfet_03v3
**devattr s=44000,1176 d=26000,604
X88 a_4978_7058 vdd.t521 vss.t186 vss.t185 nfet_03v3
**devattr s=17600,576 d=10400,304
X89 vdd.t442 reset.t11 dffrs_4.nand3_8.Z.t3 vdd.t441 pfet_03v3
**devattr s=26000,604 d=26000,604
X90 vdd.t314 dffrs_5.nand3_6.C.t5 dffrs_5.Q.t0 vdd.t313 pfet_03v3
**devattr s=26000,604 d=26000,604
X91 dffrs_13.nand3_6.C.t3 dffrs_13.nand3_1.C.t4 vdd.t264 vdd.t263 pfet_03v3
**devattr s=44000,1176 d=26000,604
X92 dffrs_3.nand3_8.C.t2 dffrs_3.nand3_8.Z.t4 a_17288_2648 vss.t197 nfet_03v3
**devattr s=10400,304 d=17600,576
X93 vdd.t119 vdd.t117 dffrs_13.nand3_8.Z.t1 vdd.t118 pfet_03v3
**devattr s=26000,604 d=26000,604
X94 a_14548_12225 d3.t5 vss.t244 vss.t243 nfet_03v3
**devattr s=17600,576 d=10400,304
X95 vdd.t254 d1.t5 dffrs_9.nand3_8.C.t2 vdd.t253 pfet_03v3
**devattr s=26000,604 d=26000,604
X96 vdd.t488 clk.t7 dffrs_4.nand3_8.C.t1 vdd.t487 pfet_03v3
**devattr s=26000,604 d=26000,604
X97 a_18774_2649 dffrs_3.nand3_8.C.t4 a_18590_2649 vss.t161 nfet_03v3
**devattr s=10400,304 d=10400,304
X98 dffrs_13.nand3_1.C.t3 reset.t12 vdd.t440 vdd.t439 pfet_03v3
**devattr s=44000,1176 d=26000,604
X99 dffrs_5.nand3_8.Z.t2 dffrs_4.Q.t5 vdd.t136 vdd.t135 pfet_03v3
**devattr s=26000,604 d=44000,1176
X100 vdd.t438 reset.t13 dffrs_9.nand3_6.C.t3 vdd.t437 pfet_03v3
**devattr s=26000,604 d=26000,604
X101 dffrs_4.Qb.t0 dffrs_4.Q.t6 vdd.t134 vdd.t133 pfet_03v3
**devattr s=44000,1176 d=26000,604
X102 vdd.t490 clk.t8 dffrs_13.nand3_8.C.t0 vdd.t489 pfet_03v3
**devattr s=26000,604 d=26000,604
X103 dffrs_5.nand3_8.C.t2 dffrs_5.nand3_8.Z.t4 vdd.t284 vdd.t283 pfet_03v3
**devattr s=26000,604 d=44000,1176
X104 dffrs_13.Qb.t3 dffrs_0.d.t5 vdd.t498 vdd.t497 pfet_03v3
**devattr s=44000,1176 d=26000,604
X105 a_9204_12224 d3.t6 a_9020_12224 vss.t245 nfet_03v3
**devattr s=10400,304 d=10400,304
X106 dffrs_1.Qb.t1 reset.t14 vdd.t436 vdd.t435 pfet_03v3
**devattr s=26000,604 d=44000,1176
X107 a_9020_12224 dffrs_7.nand3_6.C.t5 vss.t4 vss.t3 nfet_03v3
**devattr s=17600,576 d=10400,304
X108 vdd.t518 dffrs_5.nand3_8.C.t5 dffrs_5.Qb.t3 vdd.t517 pfet_03v3
**devattr s=26000,604 d=26000,604
X109 a_9204_14429 reset.t15 a_9020_14429 vss.t299 nfet_03v3
**devattr s=10400,304 d=10400,304
X110 a_13246_4853 reset.t16 a_13062_4853 vss.t298 nfet_03v3
**devattr s=10400,304 d=10400,304
X111 a_9020_14429 dffrs_7.nand3_1.C vss.t254 vss.t253 nfet_03v3
**devattr s=17600,576 d=10400,304
X112 a_14732_4853 dffrs_2.nand3_6.C.t5 a_14548_4853 vss.t6 nfet_03v3
**devattr s=10400,304 d=10400,304
X113 dffrs_7.Qb reset.t17 vdd.t434 vdd.t433 pfet_03v3
**devattr s=26000,604 d=44000,1176
X114 dffrs_4.d.t0 dffrs_3.Qb.t6 a_18774_4853 vss.t309 nfet_03v3
**devattr s=10400,304 d=17600,576
X115 dffrs_9.nand3_1.C dffrs_9.nand3_6.C.t6 a_17288_16634 vss.t219 nfet_03v3
**devattr s=10400,304 d=17600,576
X116 a_21330_16634 dffrs_10.nand3_8.Z a_21146_16634 vss.t191 nfet_03v3
**devattr s=10400,304 d=10400,304
X117 vdd.t216 dffrs_4.nand3_6.C.t5 dffrs_4.Q.t0 vdd.t215 pfet_03v3
**devattr s=26000,604 d=26000,604
X118 vdd.t432 reset.t18 dffrs_14.nand3_8.Z vdd.t431 pfet_03v3
**devattr s=26000,604 d=26000,604
X119 dffrs_2.nand3_8.C.t3 dffrs_2.nand3_8.Z.t4 a_13246_2648 vss.t312 nfet_03v3
**devattr s=10400,304 d=17600,576
X120 dffrs_9.Qb reset.t19 vdd.t430 vdd.t429 pfet_03v3
**devattr s=26000,604 d=44000,1176
X121 vdd.t154 dffrs_10.nand3_8.C.t4 dffrs_10.Qb vdd.t153 pfet_03v3
**devattr s=26000,604 d=26000,604
X122 dffrs_12.nand3_8.Z dffrs_12.nand3_8.C.t4 vdd.t212 vdd.t211 pfet_03v3
**devattr s=44000,1176 d=26000,604
X123 dffrs_1.nand3_8.C.t1 dffrs_1.nand3_8.Z.t4 a_9204_2648 vss.t166 nfet_03v3
**devattr s=10400,304 d=17600,576
X124 vdd.t11 dffrs_13.nand3_6.C.t5 dffrs_0.d.t2 vdd.t10 pfet_03v3
**devattr s=26000,604 d=26000,604
X125 dffrs_1.nand3_8.Z.t0 dffrs_1.nand3_8.C.t5 vdd.t184 vdd.t183 pfet_03v3
**devattr s=44000,1176 d=26000,604
X126 a_14732_2649 dffrs_2.nand3_8.C.t4 a_14548_2649 vss.t85 nfet_03v3
**devattr s=10400,304 d=10400,304
X127 dffrs_4.nand3_8.Z.t1 dffrs_4.d.t4 vdd.t230 vdd.t229 pfet_03v3
**devattr s=26000,604 d=44000,1176
X128 dffrs_12.Q.t3 dffrs_5.Qb.t5 vdd.t356 vdd.t355 pfet_03v3
**devattr s=44000,1176 d=26000,604
X129 vdd.t196 dffrs_11.nand3_6.C.t4 d0.t3 vdd.t195 pfet_03v3
**devattr s=26000,604 d=26000,604
X130 dffrs_1.nand3_8.C.t3 dffrs_1.nand3_6.C.t5 vdd.t460 vdd.t459 pfet_03v3
**devattr s=44000,1176 d=26000,604
X131 a_29414_16634 dffrs_12.nand3_8.Z a_29230_16634 vss.t53 nfet_03v3
**devattr s=10400,304 d=10400,304
X132 a_25372_12224 dffrs_12.Q.t6 a_25188_12224 vss.t58 nfet_03v3
**devattr s=10400,304 d=10400,304
X133 a_13246_7058 dffrs_2.nand3_8.Z.t5 a_13062_7058 vss.t313 nfet_03v3
**devattr s=10400,304 d=10400,304
X134 dffrs_13.nand3_8.Z.t2 vss.t340 vdd.t312 vdd.t311 pfet_03v3
**devattr s=26000,604 d=44000,1176
X135 dffrs_4.nand3_8.C.t2 dffrs_4.nand3_8.Z.t4 vdd.t358 vdd.t357 pfet_03v3
**devattr s=26000,604 d=44000,1176
X136 dffrs_3.Qb.t3 reset.t20 a_18774_2649 vss.t297 nfet_03v3
**devattr s=10400,304 d=17600,576
X137 vdd.t480 dffrs_4.nand3_8.C.t4 dffrs_4.Qb.t3 vdd.t479 pfet_03v3
**devattr s=26000,604 d=26000,604
X138 a_18590_14429 dffrs_2.Qb.t5 vss.t104 vss.t103 nfet_03v3
**devattr s=17600,576 d=10400,304
X139 d4.t2 dffrs_0.Qb.t4 vdd.t69 vdd.t68 pfet_03v3
**devattr s=44000,1176 d=26000,604
X140 dffrs_13.nand3_8.C.t2 dffrs_13.nand3_8.Z.t5 vdd.t258 vdd.t257 pfet_03v3
**devattr s=26000,604 d=44000,1176
X141 a_25372_14429 reset.t21 a_25188_14429 vss.t296 nfet_03v3
**devattr s=10400,304 d=10400,304
X142 dffrs_8.nand3_8.Z comp_in.t1 a_13246_10019 vss.t232 nfet_03v3
**devattr s=10400,304 d=17600,576
X143 vdd.t47 dffrs_7.nand3_8.Z dffrs_7.nand3_1.C vdd.t46 pfet_03v3
**devattr s=26000,604 d=26000,604
X144 vdd.t1 dffrs_13.nand3_8.C.t5 dffrs_13.Qb.t0 vdd.t0 pfet_03v3
**devattr s=26000,604 d=26000,604
X145 dffrs_7.nand3_1.C dffrs_0.Qb.t5 vdd.t71 vdd.t70 pfet_03v3
**devattr s=44000,1176 d=26000,604
X146 a_25188_4853 dffrs_5.nand3_1.C.t4 vss.t44 vss.t43 nfet_03v3
**devattr s=17600,576 d=10400,304
X147 a_10690_4853 dffrs_1.nand3_6.C.t6 a_10506_4853 vss.t305 nfet_03v3
**devattr s=10400,304 d=10400,304
X148 vdd.t160 d4.t4 dffrs_14.nand3_8.C.t1 vdd.t159 pfet_03v3
**devattr s=26000,604 d=26000,604
X149 dffrs_7.nand3_8.C.t1 dffrs_7.nand3_8.Z a_9204_12224 vss.t42 nfet_03v3
**devattr s=10400,304 d=17600,576
X150 a_17104_12224 dffrs_9.nand3_6.C.t7 vss.t221 vss.t220 nfet_03v3
**devattr s=17600,576 d=10400,304
X151 a_21146_2648 dffrs_4.nand3_6.C.t6 vss.t128 vss.t127 nfet_03v3
**devattr s=17600,576 d=10400,304
X152 dffrs_2.nand3_6.C.t2 dffrs_2.nand3_1.C.t4 vdd.t288 vdd.t287 pfet_03v3
**devattr s=44000,1176 d=26000,604
X153 dffrs_2.Q.t2 dffrs_2.Qb.t6 a_14732_4853 vss.t105 nfet_03v3
**devattr s=10400,304 d=17600,576
X154 a_17104_14429 dffrs_9.nand3_1.C vss.t50 vss.t49 nfet_03v3
**devattr s=17600,576 d=10400,304
X155 dffrs_7.nand3_6.C.t1 d3.t7 a_9204_14429 vss.t141 nfet_03v3
**devattr s=10400,304 d=17600,576
X156 dffrs_2.nand3_1.C.t0 vdd.t114 vdd.t116 vdd.t115 pfet_03v3
**devattr s=44000,1176 d=26000,604
X157 dffrs_0.nand3_8.Z.t0 dffrs_0.nand3_8.C.t5 vdd.t190 vdd.t189 pfet_03v3
**devattr s=44000,1176 d=26000,604
X158 vdd.t428 reset.t22 dffrs_0.nand3_6.C.t3 vdd.t427 pfet_03v3
**devattr s=26000,604 d=26000,604
X159 dffrs_3.nand3_6.C.t2 dffrs_3.nand3_1.C.t4 vdd.t228 vdd.t227 pfet_03v3
**devattr s=44000,1176 d=26000,604
X160 dffrs_0.nand3_8.C.t3 dffrs_0.nand3_6.C.t5 vdd.t140 vdd.t139 pfet_03v3
**devattr s=44000,1176 d=26000,604
X161 a_10690_2649 dffrs_1.nand3_8.C.t6 a_10506_2649 vss.t108 nfet_03v3
**devattr s=10400,304 d=10400,304
X162 vdd.t368 dffrs_0.nand3_8.Z.t5 dffrs_0.nand3_1.C.t1 vdd.t367 pfet_03v3
**devattr s=26000,604 d=26000,604
X163 dffrs_3.nand3_1.C.t3 vdd.t111 vdd.t113 vdd.t112 pfet_03v3
**devattr s=44000,1176 d=26000,604
X164 dffrs_10.Qb reset.t23 a_22816_12225 vss.t295 nfet_03v3
**devattr s=10400,304 d=17600,576
X165 dffrs_9.nand3_8.Z comp_in.t2 vdd.t336 vdd.t335 pfet_03v3
**devattr s=26000,604 d=44000,1176
X166 vdd.t426 reset.t24 dffrs_10.nand3_8.Z vdd.t425 pfet_03v3
**devattr s=26000,604 d=26000,604
X167 a_966_2648 dffrs_13.nand3_6.C.t6 vss.t326 vss.t325 nfet_03v3
**devattr s=17600,576 d=10400,304
X168 dffrs_12.Q.t2 dffrs_12.Qb a_30900_14429 vss.t179 nfet_03v3
**devattr s=10400,304 d=17600,576
X169 dffrs_4.d.t3 vdd.t108 vdd.t110 vdd.t109 pfet_03v3
**devattr s=44000,1176 d=26000,604
X170 a_30900_14429 dffrs_12.nand3_6.C.t6 a_30716_14429 vss.t331 nfet_03v3
**devattr s=10400,304 d=10400,304
X171 a_25188_7058 vdd.t522 vss.t188 vss.t187 nfet_03v3
**devattr s=17600,576 d=10400,304
X172 dffrs_2.Qb.t2 reset.t25 a_14732_2649 vss.t294 nfet_03v3
**devattr s=10400,304 d=17600,576
X173 d0.t1 dffrs_11.Qb a_26858_14429 vss.t2 nfet_03v3
**devattr s=10400,304 d=17600,576
X174 dffrs_14.nand3_8.Z comp_in.t3 vdd.t338 vdd.t337 pfet_03v3
**devattr s=26000,604 d=44000,1176
X175 dffrs_10.nand3_1.C dffrs_10.nand3_6.C.t7 a_21330_16634 vss.t315 nfet_03v3
**devattr s=10400,304 d=17600,576
X176 vdd.t272 dffrs_11.nand3_8.Z dffrs_11.nand3_1.C vdd.t271 pfet_03v3
**devattr s=26000,604 d=26000,604
X177 dffrs_8.nand3_8.C.t2 dffrs_8.nand3_8.Z vdd.t268 vdd.t267 pfet_03v3
**devattr s=26000,604 d=44000,1176
X178 vdd.t424 reset.t26 dffrs_12.nand3_8.Z vdd.t423 pfet_03v3
**devattr s=26000,604 d=26000,604
X179 a_10690_14429 dffrs_7.nand3_6.C.t6 a_10506_14429 vss.t5 nfet_03v3
**devattr s=10400,304 d=10400,304
X180 dffrs_8.nand3_6.C.t1 d2.t4 vdd.t514 vdd.t513 pfet_03v3
**devattr s=26000,604 d=44000,1176
X181 dffrs_12.nand3_1.C dffrs_12.nand3_6.C.t7 a_29414_16634 vss.t332 nfet_03v3
**devattr s=10400,304 d=17600,576
X182 dffrs_3.Qb.t0 dffrs_4.d.t5 vdd.t39 vdd.t38 pfet_03v3
**devattr s=44000,1176 d=26000,604
X183 dffrs_9.Qb d2.t5 vdd.t516 vdd.t515 pfet_03v3
**devattr s=44000,1176 d=26000,604
X184 a_18774_12225 dffrs_9.nand3_8.C.t5 a_18590_12225 vss.t55 nfet_03v3
**devattr s=10400,304 d=10400,304
X185 a_22632_12225 d1.t6 vss.t169 vss.t168 nfet_03v3
**devattr s=17600,576 d=10400,304
X186 dffrs_11.nand3_8.C.t2 dffrs_11.nand3_8.Z a_25372_12224 vss.t181 nfet_03v3
**devattr s=10400,304 d=17600,576
X187 a_26674_14429 dffrs_4.Qb.t7 vss.t15 vss.t14 nfet_03v3
**devattr s=17600,576 d=10400,304
X188 dffrs_11.nand3_6.C.t0 dffrs_12.Q.t7 a_25372_14429 vss.t59 nfet_03v3
**devattr s=10400,304 d=17600,576
X189 dffrs_13.nand3_8.Z.t3 vss.t212 a_1150_443 vss.t213 nfet_03v3
**devattr s=10400,304 d=17600,576
X190 a_21146_16634 dffrs_3.Qb.t7 vss.t311 vss.t310 nfet_03v3
**devattr s=17600,576 d=10400,304
X191 dffrs_7.nand3_1.C dffrs_7.nand3_6.C.t7 vdd.t7 vdd.t6 pfet_03v3
**devattr s=26000,604 d=44000,1176
X192 dffrs_9.nand3_1.C dffrs_2.Qb.t7 vdd.t180 vdd.t179 pfet_03v3
**devattr s=44000,1176 d=26000,604
X193 dffrs_2.Q.t0 vdd.t105 vdd.t107 vdd.t106 pfet_03v3
**devattr s=44000,1176 d=26000,604
X194 dffrs_0.nand3_6.C.t0 clk.t9 vdd.t172 vdd.t171 pfet_03v3
**devattr s=26000,604 d=44000,1176
X195 dffrs_14.nand3_8.C.t3 dffrs_14.nand3_8.Z vdd.t328 vdd.t327 pfet_03v3
**devattr s=26000,604 d=44000,1176
X196 a_17288_12224 d1.t7 a_17104_12224 vss.t170 nfet_03v3
**devattr s=10400,304 d=10400,304
X197 vdd.t422 reset.t27 dffrs_3.nand3_6.C.t3 vdd.t421 pfet_03v3
**devattr s=26000,604 d=26000,604
X198 vdd.t420 reset.t28 dffrs_5.nand3_6.C.t3 vdd.t419 pfet_03v3
**devattr s=26000,604 d=26000,604
X199 dffrs_0.nand3_1.C.t2 dffrs_0.nand3_6.C.t6 vdd.t142 vdd.t141 pfet_03v3
**devattr s=26000,604 d=44000,1176
X200 vdd.t418 reset.t29 dffrs_2.nand3_8.Z.t3 vdd.t417 pfet_03v3
**devattr s=26000,604 d=26000,604
X201 a_17288_14429 reset.t30 a_17104_14429 vss.t293 nfet_03v3
**devattr s=10400,304 d=10400,304
X202 vdd.t292 dffrs_3.nand3_8.Z.t5 dffrs_3.nand3_1.C.t2 vdd.t291 pfet_03v3
**devattr s=26000,604 d=26000,604
X203 a_13246_10019 reset.t31 a_13062_10019 vss.t292 nfet_03v3
**devattr s=10400,304 d=10400,304
X204 vdd.t286 dffrs_5.nand3_8.Z.t5 dffrs_5.nand3_1.C.t3 vdd.t285 pfet_03v3
**devattr s=26000,604 d=26000,604
X205 dffrs_0.Q.t1 dffrs_0.Qb.t6 vdd.t348 vdd.t347 pfet_03v3
**devattr s=26000,604 d=44000,1176
X206 vdd.t174 clk.t10 dffrs_2.nand3_8.C.t0 vdd.t173 pfet_03v3
**devattr s=26000,604 d=26000,604
X207 a_13062_10019 dffrs_8.nand3_8.C.t6 vss.t47 vss.t46 nfet_03v3
**devattr s=17600,576 d=10400,304
X208 dffrs_2.nand3_8.Z.t1 dffrs_2.d.t4 a_13246_443 vss.t316 nfet_03v3
**devattr s=10400,304 d=17600,576
X209 dffrs_2.Qb.t1 dffrs_2.Q.t4 vdd.t298 vdd.t297 pfet_03v3
**devattr s=44000,1176 d=26000,604
X210 dffrs_12.Qb reset.t32 vdd.t416 vdd.t415 pfet_03v3
**devattr s=26000,604 d=44000,1176
X211 vdd.t214 dffrs_12.nand3_8.C.t5 dffrs_12.Qb vdd.t213 pfet_03v3
**devattr s=26000,604 d=26000,604
X212 a_25188_10019 dffrs_11.nand3_8.C.t5 vss.t63 vss.t62 nfet_03v3
**devattr s=17600,576 d=10400,304
X213 dffrs_11.Qb reset.t33 vdd.t414 vdd.t413 pfet_03v3
**devattr s=26000,604 d=44000,1176
X214 dffrs_10.nand3_8.Z comp_in.t4 vdd.t340 vdd.t339 pfet_03v3
**devattr s=26000,604 d=44000,1176
X215 dffrs_0.Qb.t2 reset.t34 vdd.t412 vdd.t411 pfet_03v3
**devattr s=26000,604 d=44000,1176
X216 dffrs_11.nand3_1.C dffrs_11.nand3_6.C.t5 vdd.t198 vdd.t197 pfet_03v3
**devattr s=26000,604 d=44000,1176
X217 vdd.t500 dffrs_7.nand3_8.C.t4 dffrs_7.Qb vdd.t499 pfet_03v3
**devattr s=26000,604 d=26000,604
X218 a_6464_4853 vdd.t523 vss.t190 vss.t189 nfet_03v3
**devattr s=17600,576 d=10400,304
X219 dffrs_7.Qb reset.t35 a_10690_12225 vss.t291 nfet_03v3
**devattr s=10400,304 d=17600,576
X220 dffrs_12.nand3_8.Z vss.t341 vdd.t310 vdd.t309 pfet_03v3
**devattr s=26000,604 d=44000,1176
X221 a_17288_443 reset.t36 a_17104_443 vss.t290 nfet_03v3
**devattr s=10400,304 d=10400,304
X222 a_9204_4853 reset.t37 a_9020_4853 vss.t289 nfet_03v3
**devattr s=10400,304 d=10400,304
X223 a_13062_443 dffrs_2.nand3_8.C.t5 vss.t87 vss.t86 nfet_03v3
**devattr s=17600,576 d=10400,304
X224 vdd.t238 dffrs_8.nand3_6.C.t4 d3.t2 vdd.t237 pfet_03v3
**devattr s=26000,604 d=26000,604
X225 a_13062_2648 dffrs_2.nand3_6.C.t6 vss.t20 vss.t19 nfet_03v3
**devattr s=17600,576 d=10400,304
X226 dffrs_2.d.t0 vdd.t102 vdd.t104 vdd.t103 pfet_03v3
**devattr s=44000,1176 d=26000,604
X227 dffrs_11.Qb d0.t5 vdd.t508 vdd.t507 pfet_03v3
**devattr s=44000,1176 d=26000,604
X228 dffrs_9.Qb reset.t38 a_18774_12225 vss.t288 nfet_03v3
**devattr s=10400,304 d=17600,576
X229 a_22816_12225 dffrs_10.nand3_8.C.t5 a_22632_12225 vss.t80 nfet_03v3
**devattr s=10400,304 d=10400,304
X230 dffrs_10.nand3_8.Z dffrs_10.nand3_8.C.t6 vdd.t156 vdd.t155 pfet_03v3
**devattr s=44000,1176 d=26000,604
X231 dffrs_3.nand3_6.C.t1 clk.t11 a_17288_4853 vss.t100 nfet_03v3
**devattr s=10400,304 d=17600,576
X232 a_5162_2648 clk.t12 a_4978_2648 vss.t101 nfet_03v3
**devattr s=10400,304 d=10400,304
X233 vdd.t410 reset.t40 dffrs_4.nand3_6.C.t3 vdd.t409 pfet_03v3
**devattr s=26000,604 d=26000,604
X234 a_25372_443 reset.t39 a_25188_443 vss.t287 nfet_03v3
**devattr s=10400,304 d=10400,304
X235 a_17104_2648 dffrs_3.nand3_6.C.t5 vss.t10 vss.t9 nfet_03v3
**devattr s=17600,576 d=10400,304
X236 a_30716_14429 dffrs_5.Qb.t6 vss.t248 vss.t247 nfet_03v3
**devattr s=17600,576 d=10400,304
X237 a_26858_14429 dffrs_11.nand3_6.C.t6 a_26674_14429 vss.t113 nfet_03v3
**devattr s=10400,304 d=10400,304
X238 a_6464_2649 dffrs_0.Q.t5 vss.t140 vss.t139 nfet_03v3
**devattr s=17600,576 d=10400,304
X239 vdd.t101 vdd.t99 dffrs_13.nand3_6.C.t2 vdd.t100 pfet_03v3
**devattr s=26000,604 d=26000,604
X240 vdd.t360 dffrs_4.nand3_8.Z.t5 dffrs_4.nand3_1.C.t3 vdd.t359 pfet_03v3
**devattr s=26000,604 d=26000,604
X241 vdd.t132 dffrs_9.nand3_8.Z dffrs_9.nand3_1.C vdd.t131 pfet_03v3
**devattr s=26000,604 d=26000,604
X242 dffrs_5.nand3_8.Z.t0 dffrs_5.nand3_8.C.t6 vdd.t144 vdd.t143 pfet_03v3
**devattr s=44000,1176 d=26000,604
X243 vdd.t210 d2.t6 dffrs_8.nand3_8.C.t0 vdd.t209 pfet_03v3
**devattr s=26000,604 d=26000,604
X244 dffrs_14.nand3_8.Z dffrs_14.nand3_8.C.t5 vdd.t302 vdd.t301 pfet_03v3
**devattr s=44000,1176 d=26000,604
X245 dffrs_5.nand3_6.C.t2 clk.t13 vdd.t176 vdd.t175 pfet_03v3
**devattr s=26000,604 d=44000,1176
X246 vdd.t256 dffrs_13.nand3_8.Z.t6 dffrs_13.nand3_1.C.t2 vdd.t255 pfet_03v3
**devattr s=26000,604 d=26000,604
X247 dffrs_8.nand3_8.C.t1 dffrs_8.nand3_6.C.t5 vdd.t260 vdd.t259 pfet_03v3
**devattr s=44000,1176 d=26000,604
X248 dffrs_1.Qb.t3 dffrs_2.d.t5 vdd.t476 vdd.t475 pfet_03v3
**devattr s=44000,1176 d=26000,604
X249 dffrs_5.nand3_8.C.t0 dffrs_5.nand3_6.C.t6 vdd.t316 vdd.t315 pfet_03v3
**devattr s=44000,1176 d=26000,604
X250 a_10506_14429 dffrs_0.Qb.t7 vss.t239 vss.t238 nfet_03v3
**devattr s=17600,576 d=10400,304
X251 a_9204_443 reset.t42 a_9020_443 vss.t286 nfet_03v3
**devattr s=10400,304 d=10400,304
X252 vdd.t408 reset.t41 dffrs_8.nand3_6.C.t3 vdd.t407 pfet_03v3
**devattr s=26000,604 d=26000,604
X253 dffrs_5.nand3_1.C.t0 dffrs_5.nand3_6.C.t7 vdd.t318 vdd.t317 pfet_03v3
**devattr s=26000,604 d=44000,1176
X254 a_9204_16634 dffrs_7.nand3_8.Z a_9020_16634 vss.t41 nfet_03v3
**devattr s=10400,304 d=10400,304
X255 dffrs_8.nand3_6.C.t0 dffrs_8.nand3_1.C vdd.t45 vdd.t44 pfet_03v3
**devattr s=44000,1176 d=26000,604
X256 dffrs_0.nand3_8.Z.t2 dffrs_0.d.t6 a_5162_443 vss.t328 nfet_03v3
**devattr s=10400,304 d=17600,576
X257 dffrs_11.nand3_8.C.t1 dffrs_11.nand3_6.C.t7 vdd.t200 vdd.t199 pfet_03v3
**devattr s=44000,1176 d=26000,604
X258 a_9020_16634 dffrs_0.Qb.t8 vss.t241 vss.t240 nfet_03v3
**devattr s=17600,576 d=10400,304
X259 dffrs_5.Q.t2 dffrs_5.Qb.t7 vdd.t354 vdd.t353 pfet_03v3
**devattr s=26000,604 d=44000,1176
X260 a_5162_10022 reset.t43 a_4978_10022 vss.t285 nfet_03v3
**devattr s=10400,304 d=10400,304
X261 a_9204_7058 dffrs_1.nand3_8.Z.t5 a_9020_7058 vss.t167 nfet_03v3
**devattr s=10400,304 d=10400,304
X262 dffrs_11.nand3_6.C.t2 dffrs_11.nand3_1.C vdd.t344 vdd.t343 pfet_03v3
**devattr s=44000,1176 d=26000,604
X263 a_29230_10019 dffrs_12.nand3_8.C.t6 vss.t125 vss.t124 nfet_03v3
**devattr s=17600,576 d=10400,304
X264 a_5162_12227 d4.t5 a_4978_12227 vss.t260 nfet_03v3
**devattr s=10400,304 d=10400,304
X265 a_21146_443 dffrs_4.nand3_8.C.t5 vss.t320 vss.t319 nfet_03v3
**devattr s=17600,576 d=10400,304
X266 dffrs_3.nand3_1.C.t1 dffrs_3.nand3_6.C.t6 a_17288_7058 vss.t24 nfet_03v3
**devattr s=10400,304 d=17600,576
X267 a_6648_4853 dffrs_0.nand3_6.C.t7 a_6464_4853 vss.t72 nfet_03v3
**devattr s=10400,304 d=10400,304
X268 a_4978_443 dffrs_0.nand3_8.C.t6 vss.t201 vss.t200 nfet_03v3
**devattr s=17600,576 d=10400,304
X269 dffrs_5.Qb.t2 reset.t44 vdd.t406 vdd.t405 pfet_03v3
**devattr s=26000,604 d=44000,1176
X270 dffrs_2.nand3_6.C.t1 clk.t14 a_13246_4853 vss.t102 nfet_03v3
**devattr s=10400,304 d=17600,576
X271 a_26674_4853 vdd.t524 vss.t143 vss.t142 nfet_03v3
**devattr s=17600,576 d=10400,304
X272 dffrs_1.nand3_6.C.t1 clk.t15 a_9204_4853 vss.t109 nfet_03v3
**devattr s=10400,304 d=17600,576
X273 dffrs_14.nand3_8.C.t0 dffrs_14.nand3_6.C.t5 vdd.t224 vdd.t223 pfet_03v3
**devattr s=44000,1176 d=26000,604
X274 dffrs_1.nand3_6.C.t2 dffrs_1.nand3_1.C.t5 vdd.t202 vdd.t201 pfet_03v3
**devattr s=44000,1176 d=26000,604
X275 dffrs_4.nand3_6.C.t0 clk.t16 vdd.t192 vdd.t191 pfet_03v3
**devattr s=26000,604 d=44000,1176
X276 dffrs_0.nand3_8.C.t2 dffrs_0.nand3_8.Z.t6 a_5162_2648 vss.t259 nfet_03v3
**devattr s=10400,304 d=17600,576
X277 a_17288_2648 clk.t17 a_17104_2648 vss.t110 nfet_03v3
**devattr s=10400,304 d=10400,304
X278 dffrs_1.nand3_1.C.t1 vdd.t96 vdd.t98 vdd.t97 pfet_03v3
**devattr s=44000,1176 d=26000,604
X279 a_25372_2648 clk.t18 a_25188_2648 vss.t111 nfet_03v3
**devattr s=10400,304 d=10400,304
X280 d3.t0 dffrs_8.Qb vdd.t33 vdd.t32 pfet_03v3
**devattr s=26000,604 d=44000,1176
X281 a_6648_2649 dffrs_0.nand3_8.C.t7 a_6464_2649 vss.t202 nfet_03v3
**devattr s=10400,304 d=10400,304
X282 dffrs_4.nand3_1.C.t1 dffrs_4.nand3_6.C.t7 vdd.t218 vdd.t217 pfet_03v3
**devattr s=26000,604 d=44000,1176
X283 dffrs_13.nand3_6.C.t0 clk.t19 vdd.t194 vdd.t193 pfet_03v3
**devattr s=26000,604 d=44000,1176
X284 a_25372_16634 dffrs_11.nand3_8.Z a_25188_16634 vss.t180 nfet_03v3
**devattr s=10400,304 d=10400,304
X285 a_26674_2649 dffrs_5.Q.t5 vss.t23 vss.t22 nfet_03v3
**devattr s=17600,576 d=10400,304
X286 vdd.t81 dffrs_11.nand3_8.C.t6 dffrs_11.Qb vdd.t80 pfet_03v3
**devattr s=26000,604 d=26000,604
X287 dffrs_12.Qb dffrs_12.Q.t8 vdd.t79 vdd.t78 pfet_03v3
**devattr s=44000,1176 d=26000,604
X288 dffrs_8.nand3_8.C.t3 dffrs_8.nand3_8.Z a_13246_12224 vss.t177 nfet_03v3
**devattr s=10400,304 d=17600,576
X289 dffrs_4.Q.t2 dffrs_4.Qb.t8 vdd.t15 vdd.t14 pfet_03v3
**devattr s=26000,604 d=44000,1176
X290 dffrs_13.nand3_1.C.t1 dffrs_13.nand3_6.C.t7 vdd.t492 vdd.t491 pfet_03v3
**devattr s=26000,604 d=44000,1176
X291 dffrs_8.nand3_6.C.t2 d2.t7 a_13246_14429 vss.t120 nfet_03v3
**devattr s=10400,304 d=17600,576
X292 dffrs_0.d.t1 dffrs_13.Qb.t6 vdd.t146 vdd.t145 pfet_03v3
**devattr s=26000,604 d=44000,1176
X293 dffrs_7.Qb d4.t6 vdd.t370 vdd.t369 pfet_03v3
**devattr s=44000,1176 d=26000,604
X294 a_18590_12225 d2.t8 vss.t122 vss.t121 nfet_03v3
**devattr s=17600,576 d=10400,304
X295 dffrs_12.nand3_8.C.t3 dffrs_12.nand3_6.C.t8 vdd.t506 vdd.t505 pfet_03v3
**devattr s=44000,1176 d=26000,604
X296 vdd.t404 reset.t45 dffrs_7.nand3_8.Z vdd.t403 pfet_03v3
**devattr s=26000,604 d=26000,604
X297 a_21146_4853 dffrs_4.nand3_1.C.t5 vss.t163 vss.t162 nfet_03v3
**devattr s=17600,576 d=10400,304
X298 dffrs_7.nand3_8.Z dffrs_7.nand3_8.C.t5 vdd.t332 vdd.t331 pfet_03v3
**devattr s=44000,1176 d=26000,604
X299 vdd.t402 reset.t46 dffrs_14.nand3_6.C.t3 vdd.t401 pfet_03v3
**devattr s=26000,604 d=26000,604
X300 dffrs_2.nand3_1.C.t1 dffrs_2.nand3_6.C.t7 a_13246_7058 vss.t21 nfet_03v3
**devattr s=10400,304 d=17600,576
X301 d3.t3 dffrs_1.Qb.t6 vdd.t206 vdd.t205 pfet_03v3
**devattr s=44000,1176 d=26000,604
X302 dffrs_1.nand3_1.C.t0 dffrs_1.nand3_6.C.t7 a_9204_7058 vss.t16 nfet_03v3
**devattr s=10400,304 d=17600,576
X303 dffrs_12.nand3_6.C.t0 dffrs_12.nand3_1.C vdd.t232 vdd.t231 pfet_03v3
**devattr s=44000,1176 d=26000,604
X304 a_21330_10019 reset.t47 a_21146_10019 vss.t284 nfet_03v3
**devattr s=10400,304 d=10400,304
X305 a_17104_16634 dffrs_2.Qb.t8 vss.t107 vss.t106 nfet_03v3
**devattr s=17600,576 d=10400,304
X306 dffrs_7.nand3_1.C dffrs_7.nand3_6.C.t8 a_9204_16634 vss.t306 nfet_03v3
**devattr s=10400,304 d=17600,576
X307 dffrs_9.nand3_8.Z comp_in.t5 a_17288_10019 vss.t25 nfet_03v3
**devattr s=10400,304 d=17600,576
X308 vdd.t326 dffrs_14.nand3_8.Z dffrs_14.nand3_1.C vdd.t325 pfet_03v3
**devattr s=26000,604 d=26000,604
X309 dffrs_4.Qb.t2 reset.t48 vdd.t400 vdd.t399 pfet_03v3
**devattr s=26000,604 d=44000,1176
X310 a_22632_4853 vdd.t525 vss.t145 vss.t144 nfet_03v3
**devattr s=17600,576 d=10400,304
X311 dffrs_14.nand3_8.Z comp_in.t6 a_5162_10022 vss.t26 nfet_03v3
**devattr s=10400,304 d=17600,576
X312 dffrs_0.nand3_6.C.t2 dffrs_0.nand3_1.C.t5 vdd.t346 vdd.t345 pfet_03v3
**devattr s=44000,1176 d=26000,604
X313 dffrs_13.Qb.t1 vdd.t93 vdd.t95 vdd.t94 pfet_03v3
**devattr s=26000,604 d=44000,1176
X314 a_2452_4853 reset.t49 vss.t283 vss.t282 nfet_03v3
**devattr s=17600,576 d=10400,304
X315 dffrs_2.d.t3 dffrs_1.Qb.t7 a_10690_4853 vss.t118 nfet_03v3
**devattr s=10400,304 d=17600,576
X316 a_29414_10019 reset.t50 a_29230_10019 vss.t281 nfet_03v3
**devattr s=10400,304 d=10400,304
X317 dffrs_14.nand3_8.C.t2 dffrs_14.nand3_8.Z a_5162_12227 vss.t225 nfet_03v3
**devattr s=10400,304 d=17600,576
X318 dffrs_0.nand3_1.C.t0 vdd.t90 vdd.t92 vdd.t91 pfet_03v3
**devattr s=44000,1176 d=26000,604
X319 a_26858_4853 dffrs_5.nand3_6.C.t8 a_26674_4853 vss.t217 nfet_03v3
**devattr s=10400,304 d=10400,304
X320 a_966_4853 dffrs_13.nand3_1.C.t5 vss.t173 vss.t172 nfet_03v3
**devattr s=17600,576 d=10400,304
X321 a_21330_2648 clk.t20 a_21146_2648 vss.t112 nfet_03v3
**devattr s=10400,304 d=10400,304
X322 a_22632_2649 dffrs_4.Q.t7 vss.t70 vss.t69 nfet_03v3
**devattr s=17600,576 d=10400,304
X323 a_1150_2648 clk.t21 a_966_2648 vss.t88 nfet_03v3
**devattr s=10400,304 d=10400,304
X324 dffrs_5.nand3_8.C.t3 dffrs_5.nand3_8.Z.t6 a_25372_2648 vss.t193 nfet_03v3
**devattr s=10400,304 d=17600,576
X325 dffrs_1.Qb.t2 reset.t51 a_10690_2649 vss.t280 nfet_03v3
**devattr s=10400,304 d=17600,576
X326 a_2452_2649 dffrs_0.d.t7 vss.t330 vss.t329 nfet_03v3
**devattr s=17600,576 d=10400,304
X327 dffrs_12.Qb reset.t52 a_30900_12225 vss.t279 nfet_03v3
**devattr s=10400,304 d=17600,576
X328 a_21146_7058 vdd.t526 vss.t147 vss.t146 nfet_03v3
**devattr s=17600,576 d=10400,304
X329 dffrs_8.nand3_1.C dffrs_8.nand3_6.C.t6 vdd.t262 vdd.t261 pfet_03v3
**devattr s=26000,604 d=44000,1176
X330 dffrs_11.Qb reset.t53 a_26858_12225 vss.t278 nfet_03v3
**devattr s=10400,304 d=17600,576
X331 a_30900_12225 dffrs_12.nand3_8.C.t7 a_30716_12225 vss.t126 nfet_03v3
**devattr s=10400,304 d=10400,304
X332 a_26858_2649 dffrs_5.nand3_8.C.t7 a_26674_2649 vss.t75 nfet_03v3
**devattr s=10400,304 d=10400,304
X333 vdd.t398 reset.t54 dffrs_11.nand3_8.Z vdd.t397 pfet_03v3
**devattr s=26000,604 d=26000,604
X334 vdd.t23 dffrs_3.nand3_6.C.t7 dffrs_4.d.t2 vdd.t22 pfet_03v3
**devattr s=26000,604 d=26000,604
X335 vdd.t396 reset.t55 dffrs_1.nand3_8.Z.t1 vdd.t395 pfet_03v3
**devattr s=26000,604 d=26000,604
X336 d5.t2 dffrs_14.Qb vdd.t208 vdd.t207 pfet_03v3
**devattr s=26000,604 d=44000,1176
X337 vdd.t162 clk.t22 dffrs_1.nand3_8.C.t0 vdd.t161 pfet_03v3
**devattr s=26000,604 d=26000,604
X338 dffrs_11.nand3_1.C dffrs_11.nand3_6.C.t8 a_25372_16634 vss.t96 nfet_03v3
**devattr s=10400,304 d=17600,576
X339 a_10690_12225 dffrs_7.nand3_8.C.t6 a_10506_12225 vss.t227 nfet_03v3
**devattr s=10400,304 d=10400,304
X340 dffrs_9.nand3_8.C.t0 dffrs_9.nand3_8.Z vdd.t130 vdd.t129 pfet_03v3
**devattr s=26000,604 d=44000,1176
X341 vdd.t510 d0.t6 dffrs_10.nand3_8.C.t3 vdd.t509 pfet_03v3
**devattr s=26000,604 d=26000,604
X342 dffrs_3.nand3_8.Z.t1 dffrs_2.Q.t5 vdd.t300 vdd.t299 pfet_03v3
**devattr s=26000,604 d=44000,1176
X343 a_14732_14429 dffrs_8.nand3_6.C.t7 a_14548_14429 vss.t171 nfet_03v3
**devattr s=10400,304 d=10400,304
X344 a_966_7058 reset.t57 vss.t277 vss.t276 nfet_03v3
**devattr s=17600,576 d=10400,304
X345 dffrs_3.nand3_8.C.t1 dffrs_3.nand3_8.Z.t6 vdd.t290 vdd.t289 pfet_03v3
**devattr s=26000,604 d=44000,1176
X346 vdd.t394 reset.t56 dffrs_10.nand3_6.C.t3 vdd.t393 pfet_03v3
**devattr s=26000,604 d=26000,604
X347 dffrs_9.nand3_6.C.t1 d1.t8 vdd.t296 vdd.t295 pfet_03v3
**devattr s=26000,604 d=44000,1176
X348 dffrs_14.Qb reset.t58 vdd.t392 vdd.t391 pfet_03v3
**devattr s=26000,604 d=44000,1176
X349 a_26674_12225 d0.t7 vss.t336 vss.t335 nfet_03v3
**devattr s=17600,576 d=10400,304
X350 vdd.t248 dffrs_3.nand3_8.C.t5 dffrs_3.Qb.t1 vdd.t247 pfet_03v3
**devattr s=26000,604 d=26000,604
X351 vdd.t308 vss.t342 dffrs_12.nand3_8.C.t2 vdd.t307 pfet_03v3
**devattr s=26000,604 d=26000,604
X352 dffrs_7.nand3_8.Z comp_in.t7 vdd.t27 vdd.t26 pfet_03v3
**devattr s=26000,604 d=44000,1176
X353 dffrs_9.nand3_8.Z dffrs_9.nand3_8.C.t6 vdd.t75 vdd.t74 pfet_03v3
**devattr s=44000,1176 d=26000,604
X354 a_22816_4853 dffrs_4.nand3_6.C.t8 a_22632_4853 vss.t129 nfet_03v3
**devattr s=10400,304 d=10400,304
X355 d5.t0 dffrs_13.Qb.t7 vdd.t148 vdd.t147 pfet_03v3
**devattr s=44000,1176 d=26000,604
X356 dffrs_14.nand3_6.C.t2 d4.t7 vdd.t372 vdd.t371 pfet_03v3
**devattr s=26000,604 d=44000,1176
X357 vdd.t390 reset.t59 dffrs_12.nand3_6.C.t3 vdd.t389 pfet_03v3
**devattr s=26000,604 d=26000,604
X358 a_2636_4853 dffrs_13.nand3_6.C.t8 a_2452_4853 vss.t327 nfet_03v3
**devattr s=10400,304 d=10400,304
X359 dffrs_10.nand3_8.Z comp_in.t8 a_21330_10019 vss.t27 nfet_03v3
**devattr s=10400,304 d=17600,576
X360 a_17288_16634 dffrs_9.nand3_8.Z a_17104_16634 vss.t68 nfet_03v3
**devattr s=10400,304 d=10400,304
X361 dffrs_14.nand3_1.C dffrs_14.nand3_6.C.t6 vdd.t226 vdd.t225 pfet_03v3
**devattr s=26000,604 d=44000,1176
X362 a_13246_12224 d2.t9 a_13062_12224 vss.t123 nfet_03v3
**devattr s=10400,304 d=10400,304
X363 vdd.t388 reset.t60 dffrs_2.nand3_6.C.t3 vdd.t387 pfet_03v3
**devattr s=26000,604 d=26000,604
X364 a_9020_2648 dffrs_1.nand3_6.C.t8 vss.t18 vss.t17 nfet_03v3
**devattr s=17600,576 d=10400,304
X365 a_13062_12224 dffrs_8.nand3_6.C.t8 vss.t257 vss.t256 nfet_03v3
**devattr s=17600,576 d=10400,304
X366 dffrs_4.nand3_8.C.t3 dffrs_4.nand3_8.Z.t6 a_21330_2648 vss.t252 nfet_03v3
**devattr s=10400,304 d=17600,576
X367 a_13246_14429 reset.t61 a_13062_14429 vss.t275 nfet_03v3
**devattr s=10400,304 d=10400,304
X368 vdd.t276 dffrs_2.nand3_8.Z.t6 dffrs_2.nand3_1.C.t3 vdd.t275 pfet_03v3
**devattr s=26000,604 d=26000,604
X369 dffrs_12.nand3_8.Z vss.t210 a_29414_10019 vss.t211 nfet_03v3
**devattr s=10400,304 d=17600,576
X370 a_13062_14429 dffrs_8.nand3_1.C vss.t40 vss.t39 nfet_03v3
**devattr s=17600,576 d=10400,304
X371 a_22816_2649 dffrs_4.nand3_8.C.t6 a_22632_2649 vss.t255 nfet_03v3
**devattr s=10400,304 d=10400,304
X372 dffrs_13.nand3_8.C.t3 dffrs_13.nand3_8.Z.t7 a_1150_2648 vss.t99 nfet_03v3
**devattr s=10400,304 d=17600,576
X373 dffrs_14.Qb d5.t4 vdd.t43 vdd.t42 pfet_03v3
**devattr s=44000,1176 d=26000,604
X374 a_25188_12224 dffrs_11.nand3_6.C.t9 vss.t98 vss.t97 nfet_03v3
**devattr s=17600,576 d=10400,304
X375 vdd.t19 dffrs_2.nand3_6.C.t8 dffrs_2.Q.t3 vdd.t18 pfet_03v3
**devattr s=26000,604 d=26000,604
X376 dffrs_4.nand3_8.Z.t0 dffrs_4.d.t6 a_21330_443 vss.t33 nfet_03v3
**devattr s=10400,304 d=17600,576
X377 a_2636_2649 dffrs_13.nand3_8.C.t6 a_2452_2649 vss.t28 nfet_03v3
**devattr s=10400,304 d=10400,304
X378 a_1150_443 vdd.t527 a_966_443 vss.t148 nfet_03v3
**devattr s=10400,304 d=10400,304
X379 a_25188_14429 dffrs_11.nand3_1.C vss.t235 vss.t234 nfet_03v3
**devattr s=17600,576 d=10400,304
X380 a_21146_10019 dffrs_10.nand3_8.C.t7 vss.t57 vss.t56 nfet_03v3
**devattr s=17600,576 d=10400,304
X381 dffrs_2.nand3_8.Z.t2 dffrs_2.d.t6 vdd.t478 vdd.t477 pfet_03v3
**devattr s=26000,604 d=44000,1176
X382 dffrs_4.d.t1 dffrs_3.Qb.t8 vdd.t466 vdd.t465 pfet_03v3
**devattr s=26000,604 d=44000,1176
X383 dffrs_1.nand3_8.Z.t2 dffrs_0.Q.t6 vdd.t234 vdd.t233 pfet_03v3
**devattr s=26000,604 d=44000,1176
X384 d1.t3 dffrs_10.Qb vdd.t342 vdd.t341 pfet_03v3
**devattr s=26000,604 d=44000,1176
X385 dffrs_2.nand3_8.C.t2 dffrs_2.nand3_8.Z.t7 vdd.t278 vdd.t277 pfet_03v3
**devattr s=26000,604 d=44000,1176
X386 a_13062_4853 dffrs_2.nand3_1.C.t5 vss.t195 vss.t194 nfet_03v3
**devattr s=17600,576 d=10400,304
X387 dffrs_1.nand3_8.C.t2 dffrs_1.nand3_8.Z.t6 vdd.t252 vdd.t251 pfet_03v3
**devattr s=26000,604 d=44000,1176
X388 a_4978_10022 dffrs_14.nand3_8.C.t6 vss.t206 vss.t205 nfet_03v3
**devattr s=17600,576 d=10400,304
X389 dffrs_11.nand3_8.Z comp_in.t9 vdd.t29 vdd.t28 pfet_03v3
**devattr s=26000,604 d=44000,1176
X390 vdd.t53 dffrs_2.nand3_8.C.t6 dffrs_2.Qb.t0 vdd.t52 pfet_03v3
**devattr s=26000,604 d=26000,604
X391 a_4978_12227 dffrs_14.nand3_6.C.t7 vss.t131 vss.t130 nfet_03v3
**devattr s=17600,576 d=10400,304
X392 a_5162_4853 reset.t62 a_4978_4853 vss.t274 nfet_03v3
**devattr s=10400,304 d=10400,304
X393 dffrs_3.nand3_8.Z.t2 dffrs_2.Q.t6 a_17288_443 vss.t204 nfet_03v3
**devattr s=10400,304 d=17600,576
X394 a_17104_4853 dffrs_3.nand3_1.C.t5 vss.t136 vss.t135 nfet_03v3
**devattr s=17600,576 d=10400,304
X395 a_4978_2648 dffrs_0.nand3_6.C.t8 vss.t74 vss.t73 nfet_03v3
**devattr s=17600,576 d=10400,304
X396 dffrs_3.Qb.t2 reset.t63 vdd.t386 vdd.t385 pfet_03v3
**devattr s=26000,604 d=44000,1176
X397 vdd.t59 dffrs_8.nand3_8.C.t7 dffrs_8.Qb vdd.t58 pfet_03v3
**devattr s=26000,604 d=26000,604
X398 dffrs_10.nand3_8.C.t0 dffrs_10.nand3_8.Z vdd.t282 vdd.t281 pfet_03v3
**devattr s=26000,604 d=44000,1176
X399 d3.t1 dffrs_8.Qb a_14732_14429 vss.t29 nfet_03v3
**devattr s=10400,304 d=17600,576
X400 d1.t0 dffrs_3.Qb.t9 vdd.t330 vdd.t329 pfet_03v3
**devattr s=44000,1176 d=26000,604
X401 a_18590_4853 vdd.t528 vss.t150 vss.t149 nfet_03v3
**devattr s=17600,576 d=10400,304
X402 dffrs_10.nand3_6.C.t2 d0.t8 vdd.t512 vdd.t511 pfet_03v3
**devattr s=26000,604 d=44000,1176
X403 vdd.t322 dffrs_9.nand3_6.C.t8 d2.t3 vdd.t321 pfet_03v3
**devattr s=26000,604 d=26000,604
X404 dffrs_5.nand3_6.C.t0 dffrs_5.nand3_1.C.t5 vdd.t57 vdd.t56 pfet_03v3
**devattr s=44000,1176 d=26000,604
X405 vdd.t266 dffrs_8.nand3_8.Z dffrs_8.nand3_1.C vdd.t265 pfet_03v3
**devattr s=26000,604 d=26000,604
X406 a_26858_12225 dffrs_11.nand3_8.C.t7 a_26674_12225 vss.t64 nfet_03v3
**devattr s=10400,304 d=10400,304
X407 a_30716_12225 dffrs_12.Q.t9 vss.t61 vss.t60 nfet_03v3
**devattr s=17600,576 d=10400,304
X408 dffrs_4.nand3_8.Z.t2 dffrs_4.nand3_8.C.t7 vdd.t364 vdd.t363 pfet_03v3
**devattr s=44000,1176 d=26000,604
X409 dffrs_8.nand3_1.C dffrs_1.Qb.t8 vdd.t168 vdd.t167 pfet_03v3
**devattr s=44000,1176 d=26000,604
X410 vdd.t384 reset.t64 dffrs_9.nand3_8.Z vdd.t383 pfet_03v3
**devattr s=26000,604 d=26000,604
X411 dffrs_12.nand3_8.C.t1 dffrs_12.nand3_8.Z vdd.t65 vdd.t64 pfet_03v3
**devattr s=26000,604 d=44000,1176
X412 vdd.t222 dffrs_14.nand3_6.C.t8 d5.t1 vdd.t221 pfet_03v3
**devattr s=26000,604 d=26000,604
X413 vdd.t17 dffrs_1.nand3_6.C.t9 dffrs_2.d.t1 vdd.t16 pfet_03v3
**devattr s=26000,604 d=26000,604
X414 dffrs_5.nand3_1.C.t2 vdd.t87 vdd.t89 vdd.t88 pfet_03v3
**devattr s=44000,1176 d=26000,604
X415 dffrs_12.nand3_6.C.t2 vss.t343 vdd.t306 vdd.t305 pfet_03v3
**devattr s=26000,604 d=44000,1176
X416 dffrs_4.nand3_8.C.t0 dffrs_4.nand3_6.C.t9 vdd.t220 vdd.t219 pfet_03v3
**devattr s=44000,1176 d=26000,604
X417 dffrs_11.nand3_1.C dffrs_4.Qb.t9 vdd.t502 vdd.t501 pfet_03v3
**devattr s=44000,1176 d=26000,604
X418 a_17104_443 dffrs_3.nand3_8.C.t6 vss.t165 vss.t164 nfet_03v3
**devattr s=17600,576 d=10400,304
X419 a_13062_7058 vdd.t529 vss.t152 vss.t151 nfet_03v3
**devattr s=17600,576 d=10400,304
X420 a_29230_12224 dffrs_12.nand3_6.C.t9 vss.t334 vss.t333 nfet_03v3
**devattr s=17600,576 d=10400,304
X421 a_10506_12225 d4.t8 vss.t175 vss.t174 nfet_03v3
**devattr s=17600,576 d=10400,304
X422 dffrs_10.nand3_8.C.t2 dffrs_10.nand3_6.C.t8 vdd.t470 vdd.t469 pfet_03v3
**devattr s=44000,1176 d=26000,604
X423 a_5162_14432 reset.t65 a_4978_14432 vss.t273 nfet_03v3
**devattr s=10400,304 d=10400,304
X424 dffrs_2.Q.t1 dffrs_2.Qb.t9 vdd.t182 vdd.t181 pfet_03v3
**devattr s=26000,604 d=44000,1176
X425 a_18590_2649 dffrs_4.d.t7 vss.t35 vss.t34 nfet_03v3
**devattr s=17600,576 d=10400,304
X426 a_13246_443 reset.t66 a_13062_443 vss.t272 nfet_03v3
**devattr s=10400,304 d=10400,304
X427 dffrs_10.nand3_6.C.t0 dffrs_10.nand3_1.C vdd.t37 vdd.t36 pfet_03v3
**devattr s=44000,1176 d=26000,604
X428 a_14548_14429 dffrs_1.Qb.t9 vss.t95 vss.t94 nfet_03v3
**devattr s=17600,576 d=10400,304
X429 a_29230_14429 dffrs_12.nand3_1.C vss.t138 vss.t137 nfet_03v3
**devattr s=17600,576 d=10400,304
X430 a_5162_16637 dffrs_14.nand3_8.Z a_4978_16637 vss.t224 nfet_03v3
**devattr s=10400,304 d=10400,304
X431 a_5162_7058 dffrs_0.nand3_8.Z.t7 a_4978_7058 vss.t160 nfet_03v3
**devattr s=10400,304 d=10400,304
X432 a_17104_7058 vdd.t530 vss.t154 vss.t153 nfet_03v3
**devattr s=17600,576 d=10400,304
X433 dffrs_13.nand3_8.Z.t0 dffrs_13.nand3_8.C.t7 vdd.t31 vdd.t30 pfet_03v3
**devattr s=44000,1176 d=26000,604
X434 vdd.t186 dffrs_1.nand3_8.C.t7 dffrs_1.Qb.t0 vdd.t185 pfet_03v3
**devattr s=26000,604 d=26000,604
X435 vdd.t304 dffrs_14.nand3_8.C.t7 dffrs_14.Qb vdd.t303 pfet_03v3
**devattr s=26000,604 d=26000,604
X436 dffrs_14.nand3_6.C.t0 dffrs_14.nand3_1.C vdd.t83 vdd.t82 pfet_03v3
**devattr s=44000,1176 d=26000,604
X437 dffrs_13.nand3_8.C.t1 dffrs_13.nand3_6.C.t9 vdd.t494 vdd.t493 pfet_03v3
**devattr s=44000,1176 d=26000,604
X438 dffrs_2.Qb.t3 reset.t67 vdd.t382 vdd.t381 pfet_03v3
**devattr s=26000,604 d=44000,1176
X439 a_14548_4853 vdd.t531 vss.t156 vss.t155 nfet_03v3
**devattr s=17600,576 d=10400,304
X440 dffrs_14.nand3_1.C dffrs_13.Qb.t8 vdd.t150 vdd.t149 pfet_03v3
**devattr s=44000,1176 d=26000,604
X441 dffrs_0.nand3_6.C.t1 clk.t23 a_5162_4853 vss.t89 nfet_03v3
**devattr s=10400,304 d=17600,576
X442 a_25372_4853 reset.t68 a_25188_4853 vss.t271 nfet_03v3
**devattr s=10400,304 d=10400,304
X443 a_17288_4853 reset.t69 a_17104_4853 vss.t270 nfet_03v3
**devattr s=10400,304 d=10400,304
X444 a_5162_443 reset.t70 a_4978_443 vss.t269 nfet_03v3
**devattr s=10400,304 d=10400,304
X445 a_9204_10019 reset.t71 a_9020_10019 vss.t268 nfet_03v3
**devattr s=10400,304 d=10400,304
X446 a_9020_10019 dffrs_7.nand3_8.C.t7 vss.t229 vss.t228 nfet_03v3
**devattr s=17600,576 d=10400,304
X447 dffrs_0.Q.t3 dffrs_0.Qb.t9 a_6648_4853 vss.t324 nfet_03v3
**devattr s=10400,304 d=17600,576
X448 d4.t0 dffrs_7.Qb vdd.t41 vdd.t40 pfet_03v3
**devattr s=26000,604 d=44000,1176
X449 a_13246_2648 clk.t24 a_13062_2648 vss.t90 nfet_03v3
**devattr s=10400,304 d=10400,304
X450 dffrs_8.nand3_1.C dffrs_8.nand3_6.C.t9 a_13246_16634 vss.t258 nfet_03v3
**devattr s=10400,304 d=17600,576
X451 a_14548_2649 dffrs_2.Q.t7 vss.t84 vss.t83 nfet_03v3
**devattr s=17600,576 d=10400,304
X452 dffrs_8.Qb reset.t72 vdd.t380 vdd.t379 pfet_03v3
**devattr s=26000,604 d=44000,1176
X453 d5.t3 dffrs_14.Qb a_6648_14432 vss.t119 nfet_03v3
**devattr s=10400,304 d=17600,576
X454 d2.t1 dffrs_9.Qb vdd.t35 vdd.t34 pfet_03v3
**devattr s=26000,604 d=44000,1176
X455 vdd.t472 dffrs_10.nand3_6.C.t9 d1.t1 vdd.t471 pfet_03v3
**devattr s=26000,604 d=26000,604
X456 dffrs_12.nand3_1.C dffrs_5.Qb.t8 vdd.t352 vdd.t351 pfet_03v3
**devattr s=44000,1176 d=26000,604
X457 a_21330_12224 d0.t9 a_21146_12224 vss.t337 nfet_03v3
**devattr s=10400,304 d=10400,304
X458 dffrs_9.nand3_8.C.t1 dffrs_9.nand3_8.Z a_17288_12224 vss.t67 nfet_03v3
**devattr s=10400,304 d=17600,576
X459 dffrs_0.Qb.t1 reset.t73 a_6648_2649 vss.t267 nfet_03v3
**devattr s=10400,304 d=17600,576
X460 a_21330_14429 reset.t74 a_21146_14429 vss.t266 nfet_03v3
**devattr s=10400,304 d=10400,304
X461 dffrs_9.nand3_6.C.t2 d1.t9 a_17288_14429 vss.t203 nfet_03v3
**devattr s=10400,304 d=17600,576
X462 dffrs_0.nand3_1.C.t3 dffrs_0.nand3_6.C.t9 a_5162_7058 vss.t251 nfet_03v3
**devattr s=10400,304 d=17600,576
X463 a_17288_7058 dffrs_3.nand3_8.Z.t7 a_17104_7058 vss.t196 nfet_03v3
**devattr s=10400,304 d=10400,304
X464 a_25372_7058 dffrs_5.nand3_8.Z.t7 a_25188_7058 vss.t198 nfet_03v3
**devattr s=10400,304 d=10400,304
X465 a_29414_12224 vss.t208 a_29230_12224 vss.t209 nfet_03v3
**devattr s=10400,304 d=10400,304
X466 dffrs_14.Qb reset.t75 a_6648_12228 vss.t265 nfet_03v3
**devattr s=10400,304 d=17600,576
X467 dffrs_8.Qb d3.t8 vdd.t240 vdd.t239 pfet_03v3
**devattr s=44000,1176 d=26000,604
X468 a_10506_4853 vdd.t532 vss.t158 vss.t157 nfet_03v3
**devattr s=17600,576 d=10400,304
X469 dffrs_14.nand3_6.C.t1 d4.t9 a_5162_14432 vss.t176 nfet_03v3
**devattr s=10400,304 d=17600,576
X470 a_6464_14432 dffrs_13.Qb.t9 vss.t79 vss.t78 nfet_03v3
**devattr s=17600,576 d=10400,304
X471 a_29414_14429 reset.t76 a_29230_14429 vss.t264 nfet_03v3
**devattr s=10400,304 d=10400,304
X472 dffrs_14.nand3_1.C dffrs_14.nand3_6.C.t9 a_5162_16637 vss.t132 nfet_03v3
**devattr s=10400,304 d=17600,576
X473 a_21330_4853 reset.t77 a_21146_4853 vss.t263 nfet_03v3
**devattr s=10400,304 d=10400,304
X474 a_25372_10019 reset.t78 a_25188_10019 vss.t262 nfet_03v3
**devattr s=10400,304 d=10400,304
X475 vdd.t242 d3.t9 dffrs_7.nand3_8.C.t2 vdd.t241 pfet_03v3
**devattr s=26000,604 d=26000,604
X476 a_1150_4853 vdd.t533 a_966_4853 vss.t159 nfet_03v3
**devattr s=10400,304 d=10400,304
X477 dffrs_7.nand3_8.C.t3 dffrs_7.nand3_6.C.t9 vdd.t462 vdd.t461 pfet_03v3
**devattr s=44000,1176 d=26000,604
X478 vdd.t378 reset.t79 dffrs_7.nand3_6.C.t3 vdd.t377 pfet_03v3
**devattr s=26000,604 d=26000,604
X479 dffrs_5.nand3_6.C.t1 clk.t25 a_25372_4853 vss.t91 nfet_03v3
**devattr s=10400,304 d=17600,576
X480 dffrs_7.nand3_6.C.t2 dffrs_7.nand3_1.C vdd.t362 vdd.t361 pfet_03v3
**devattr s=44000,1176 d=26000,604
X481 a_25188_2648 dffrs_5.nand3_6.C.t9 vss.t223 vss.t222 nfet_03v3
**devattr s=17600,576 d=10400,304
X482 a_10506_2649 dffrs_2.d.t7 vss.t318 vss.t317 nfet_03v3
**devattr s=17600,576 d=10400,304
X483 a_6464_12228 d5.t5 vss.t38 vss.t37 nfet_03v3
**devattr s=17600,576 d=10400,304
X484 dffrs_0.Q.t0 vdd.t84 vdd.t86 vdd.t85 pfet_03v3
**devattr s=44000,1176 d=26000,604
X485 dffrs_2.nand3_8.Z.t0 dffrs_2.nand3_8.C.t7 vdd.t55 vdd.t54 pfet_03v3
**devattr s=44000,1176 d=26000,604
X486 dffrs_5.Q.t3 dffrs_5.Qb.t9 a_26858_4853 vss.t246 nfet_03v3
**devattr s=10400,304 d=17600,576
X487 vdd.t376 reset.t80 dffrs_1.nand3_6.C.t3 vdd.t375 pfet_03v3
**devattr s=26000,604 d=26000,604
X488 a_17104_10019 dffrs_9.nand3_8.C.t7 vss.t52 vss.t51 nfet_03v3
**devattr s=17600,576 d=10400,304
X489 dffrs_7.nand3_8.Z comp_in.t10 a_9204_10019 vss.t230 nfet_03v3
**devattr s=10400,304 d=17600,576
X490 dffrs_8.nand3_8.Z comp_in.t11 vdd.t334 vdd.t333 pfet_03v3
**devattr s=26000,604 d=44000,1176
X491 dffrs_2.nand3_8.C.t1 dffrs_2.nand3_6.C.t9 vdd.t5 vdd.t4 pfet_03v3
**devattr s=44000,1176 d=26000,604
X492 vdd.t374 reset.t81 dffrs_0.nand3_8.Z.t3 vdd.t373 pfet_03v3
**devattr s=26000,604 d=26000,604
X493 d1.t2 dffrs_10.Qb a_22816_14429 vss.t233 nfet_03v3
**devattr s=10400,304 d=17600,576
X494 dffrs_3.nand3_8.Z.t0 dffrs_3.nand3_8.C.t7 vdd.t250 vdd.t249 pfet_03v3
**devattr s=44000,1176 d=26000,604
X495 vdd.t294 dffrs_1.nand3_8.Z.t7 dffrs_1.nand3_1.C.t2 vdd.t293 pfet_03v3
**devattr s=26000,604 d=26000,604
X496 dffrs_9.nand3_1.C dffrs_9.nand3_6.C.t9 vdd.t324 vdd.t323 pfet_03v3
**devattr s=26000,604 d=44000,1176
X497 vdd.t280 dffrs_10.nand3_8.Z dffrs_10.nand3_1.C vdd.t279 pfet_03v3
**devattr s=26000,604 d=26000,604
X498 dffrs_3.nand3_6.C.t0 clk.t26 vdd.t164 vdd.t163 pfet_03v3
**devattr s=26000,604 d=44000,1176
X499 vdd.t496 clk.t27 dffrs_0.nand3_8.C.t0 vdd.t495 pfet_03v3
**devattr s=26000,604 d=26000,604
X500 dffrs_3.nand3_8.C.t0 dffrs_3.nand3_6.C.t8 vdd.t25 vdd.t24 pfet_03v3
**devattr s=44000,1176 d=26000,604
X501 a_21330_7058 dffrs_4.nand3_8.Z.t7 a_21146_7058 vss.t261 nfet_03v3
**devattr s=10400,304 d=10400,304
X502 dffrs_0.Qb.t3 dffrs_0.Q.t7 vdd.t236 vdd.t235 pfet_03v3
**devattr s=44000,1176 d=26000,604
X503 dffrs_3.nand3_1.C.t0 dffrs_3.nand3_6.C.t9 vdd.t51 vdd.t50 pfet_03v3
**devattr s=26000,604 d=44000,1176
R0 reset.n11 reset.t58 41.0041
R1 reset.n17 reset.t34 41.0041
R2 reset.n25 reset.t17 41.0041
R3 reset.n31 reset.t14 41.0041
R4 reset.n39 reset.t72 41.0041
R5 reset.n45 reset.t67 41.0041
R6 reset.n53 reset.t19 41.0041
R7 reset.n59 reset.t63 41.0041
R8 reset.n67 reset.t6 41.0041
R9 reset.n73 reset.t48 41.0041
R10 reset.n81 reset.t33 41.0041
R11 reset.n87 reset.t44 41.0041
R12 reset.n0 reset.t32 41.0041
R13 reset.n14 reset.t18 40.8177
R14 reset.n13 reset.t46 40.8177
R15 reset.n20 reset.t81 40.8177
R16 reset.n19 reset.t22 40.8177
R17 reset.n28 reset.t45 40.8177
R18 reset.n27 reset.t79 40.8177
R19 reset.n34 reset.t55 40.8177
R20 reset.n33 reset.t80 40.8177
R21 reset.n42 reset.t9 40.8177
R22 reset.n41 reset.t41 40.8177
R23 reset.n48 reset.t29 40.8177
R24 reset.n47 reset.t60 40.8177
R25 reset.n56 reset.t64 40.8177
R26 reset.n55 reset.t13 40.8177
R27 reset.n62 reset.t3 40.8177
R28 reset.n61 reset.t27 40.8177
R29 reset.n70 reset.t24 40.8177
R30 reset.n69 reset.t56 40.8177
R31 reset.n76 reset.t11 40.8177
R32 reset.n75 reset.t40 40.8177
R33 reset.n84 reset.t54 40.8177
R34 reset.n83 reset.t1 40.8177
R35 reset.n90 reset.t4 40.8177
R36 reset.n89 reset.t28 40.8177
R37 reset.n3 reset.t26 40.8177
R38 reset.n2 reset.t59 40.8177
R39 reset.n8 reset.t12 40.6313
R40 reset.n6 reset.t10 40.6313
R41 reset.n8 reset.t57 27.3166
R42 reset.n6 reset.t49 27.3166
R43 reset.n14 reset.t43 27.1302
R44 reset.n13 reset.t65 27.1302
R45 reset.n20 reset.t70 27.1302
R46 reset.n19 reset.t62 27.1302
R47 reset.n28 reset.t71 27.1302
R48 reset.n27 reset.t15 27.1302
R49 reset.n34 reset.t42 27.1302
R50 reset.n33 reset.t37 27.1302
R51 reset.n42 reset.t31 27.1302
R52 reset.n41 reset.t61 27.1302
R53 reset.n48 reset.t66 27.1302
R54 reset.n47 reset.t16 27.1302
R55 reset.n56 reset.t5 27.1302
R56 reset.n55 reset.t30 27.1302
R57 reset.n62 reset.t36 27.1302
R58 reset.n61 reset.t69 27.1302
R59 reset.n70 reset.t47 27.1302
R60 reset.n69 reset.t74 27.1302
R61 reset.n76 reset.t7 27.1302
R62 reset.n75 reset.t77 27.1302
R63 reset.n84 reset.t78 27.1302
R64 reset.n83 reset.t21 27.1302
R65 reset.n90 reset.t39 27.1302
R66 reset.n89 reset.t68 27.1302
R67 reset.n3 reset.t50 27.1302
R68 reset.n2 reset.t76 27.1302
R69 reset.n11 reset.t75 26.9438
R70 reset.n17 reset.t73 26.9438
R71 reset.n25 reset.t35 26.9438
R72 reset.n31 reset.t51 26.9438
R73 reset.n39 reset.t8 26.9438
R74 reset.n45 reset.t25 26.9438
R75 reset.n53 reset.t38 26.9438
R76 reset.n59 reset.t20 26.9438
R77 reset.n67 reset.t23 26.9438
R78 reset.n73 reset.t2 26.9438
R79 reset.n81 reset.t53 26.9438
R80 reset.n87 reset.t0 26.9438
R81 reset.n0 reset.t52 26.9438
R82 reset.n37 dffrs_1.resetb 19.0901
R83 reset.n51 dffrs_2.resetb 19.0901
R84 reset.n65 dffrs_3.resetb 19.0901
R85 reset.n79 dffrs_4.resetb 19.0901
R86 reset.n93 dffrs_5.resetb 19.0901
R87 reset.n23 dffrs_0.resetb 19.0467
R88 dffrs_12.resetb reset.n94 14.0622
R89 reset.n15 dffrs_14.nand3_1.B 12.1571
R90 reset.n21 dffrs_0.nand3_1.B 12.1571
R91 reset.n29 dffrs_7.nand3_1.B 12.1571
R92 reset.n35 dffrs_1.nand3_1.B 12.1571
R93 reset.n43 dffrs_8.nand3_1.B 12.1571
R94 reset.n49 dffrs_2.nand3_1.B 12.1571
R95 reset.n57 dffrs_9.nand3_1.B 12.1571
R96 reset.n63 dffrs_3.nand3_1.B 12.1571
R97 reset.n71 dffrs_10.nand3_1.B 12.1571
R98 reset.n77 dffrs_4.nand3_1.B 12.1571
R99 reset.n85 dffrs_11.nand3_1.B 12.1571
R100 reset.n91 dffrs_5.nand3_1.B 12.1571
R101 reset.n4 dffrs_12.nand3_1.B 12.1571
R102 reset.n9 reset.n7 9.22229
R103 reset.n24 reset.n10 7.9889
R104 reset.n16 reset.n12 7.75389
R105 reset.n22 reset.n18 7.75389
R106 reset.n30 reset.n26 7.75389
R107 reset.n36 reset.n32 7.75389
R108 reset.n44 reset.n40 7.75389
R109 reset.n50 reset.n46 7.75389
R110 reset.n58 reset.n54 7.75389
R111 reset.n64 reset.n60 7.75389
R112 reset.n72 reset.n68 7.75389
R113 reset.n78 reset.n74 7.75389
R114 reset.n86 reset.n82 7.75389
R115 reset.n92 reset.n88 7.75389
R116 reset.n5 reset.n1 7.75389
R117 reset.n10 dffrs_13.setb 6.43164
R118 reset.n16 reset.n15 5.93546
R119 reset.n22 reset.n21 5.93546
R120 reset.n30 reset.n29 5.93546
R121 reset.n36 reset.n35 5.93546
R122 reset.n44 reset.n43 5.93546
R123 reset.n50 reset.n49 5.93546
R124 reset.n58 reset.n57 5.93546
R125 reset.n64 reset.n63 5.93546
R126 reset.n72 reset.n71 5.93546
R127 reset.n78 reset.n77 5.93546
R128 reset.n86 reset.n85 5.93546
R129 reset.n92 reset.n91 5.93546
R130 reset.n5 reset.n4 5.93546
R131 reset.n37 dffrs_7.resetb 5.93246
R132 reset.n51 dffrs_8.resetb 5.93246
R133 reset.n65 dffrs_9.resetb 5.93246
R134 reset.n79 dffrs_10.resetb 5.93246
R135 reset.n93 dffrs_11.resetb 5.93246
R136 reset.n23 dffrs_14.resetb 5.88425
R137 reset.n12 reset.n11 5.7305
R138 reset.n18 reset.n17 5.7305
R139 reset.n26 reset.n25 5.7305
R140 reset.n32 reset.n31 5.7305
R141 reset.n40 reset.n39 5.7305
R142 reset.n46 reset.n45 5.7305
R143 reset.n54 reset.n53 5.7305
R144 reset.n60 reset.n59 5.7305
R145 reset.n68 reset.n67 5.7305
R146 reset.n74 reset.n73 5.7305
R147 reset.n82 reset.n81 5.7305
R148 reset.n88 reset.n87 5.7305
R149 reset.n1 reset.n0 5.7305
R150 dffrs_14.nand3_8.B reset.n14 5.47979
R151 dffrs_14.nand3_1.B reset.n13 5.47979
R152 dffrs_0.nand3_8.B reset.n20 5.47979
R153 dffrs_0.nand3_1.B reset.n19 5.47979
R154 dffrs_7.nand3_8.B reset.n28 5.47979
R155 dffrs_7.nand3_1.B reset.n27 5.47979
R156 dffrs_1.nand3_8.B reset.n34 5.47979
R157 dffrs_1.nand3_1.B reset.n33 5.47979
R158 dffrs_8.nand3_8.B reset.n42 5.47979
R159 dffrs_8.nand3_1.B reset.n41 5.47979
R160 dffrs_2.nand3_8.B reset.n48 5.47979
R161 dffrs_2.nand3_1.B reset.n47 5.47979
R162 dffrs_9.nand3_8.B reset.n56 5.47979
R163 dffrs_9.nand3_1.B reset.n55 5.47979
R164 dffrs_3.nand3_8.B reset.n62 5.47979
R165 dffrs_3.nand3_1.B reset.n61 5.47979
R166 dffrs_10.nand3_8.B reset.n70 5.47979
R167 dffrs_10.nand3_1.B reset.n69 5.47979
R168 dffrs_4.nand3_8.B reset.n76 5.47979
R169 dffrs_4.nand3_1.B reset.n75 5.47979
R170 dffrs_11.nand3_8.B reset.n84 5.47979
R171 dffrs_11.nand3_1.B reset.n83 5.47979
R172 dffrs_5.nand3_8.B reset.n90 5.47979
R173 dffrs_5.nand3_1.B reset.n89 5.47979
R174 dffrs_12.nand3_8.B reset.n3 5.47979
R175 dffrs_12.nand3_1.B reset.n2 5.47979
R176 reset.n9 reset.n8 5.14711
R177 reset.n7 reset.n6 5.13907
R178 reset.n15 dffrs_14.nand3_8.B 5.09593
R179 reset.n21 dffrs_0.nand3_8.B 5.09593
R180 reset.n29 dffrs_7.nand3_8.B 5.09593
R181 reset.n35 dffrs_1.nand3_8.B 5.09593
R182 reset.n43 dffrs_8.nand3_8.B 5.09593
R183 reset.n49 dffrs_2.nand3_8.B 5.09593
R184 reset.n57 dffrs_9.nand3_8.B 5.09593
R185 reset.n63 dffrs_3.nand3_8.B 5.09593
R186 reset.n71 dffrs_10.nand3_8.B 5.09593
R187 reset.n77 dffrs_4.nand3_8.B 5.09593
R188 reset.n85 dffrs_11.nand3_8.B 5.09593
R189 reset.n91 dffrs_5.nand3_8.B 5.09593
R190 reset.n4 dffrs_12.nand3_8.B 5.09593
R191 reset.n94 reset.n93 4.5005
R192 reset.n80 reset.n79 4.5005
R193 reset.n66 reset.n65 4.5005
R194 reset.n52 reset.n51 4.5005
R195 reset.n38 reset.n37 4.5005
R196 reset.n24 reset.n23 4.5005
R197 reset.n94 reset.n80 3.6383
R198 reset.n80 reset.n66 3.6383
R199 reset.n66 reset.n52 3.6383
R200 reset.n52 reset.n38 3.6383
R201 reset.n38 reset.n24 3.6113
R202 dffrs_13.setb dffrs_13.nand3_0.C 0.783821
R203 reset.n10 reset 0.13775
R204 dffrs_14.resetb reset.n16 0.136036
R205 dffrs_0.resetb reset.n22 0.136036
R206 dffrs_7.resetb reset.n30 0.136036
R207 dffrs_1.resetb reset.n36 0.136036
R208 dffrs_8.resetb reset.n44 0.136036
R209 dffrs_2.resetb reset.n50 0.136036
R210 dffrs_9.resetb reset.n58 0.136036
R211 dffrs_3.resetb reset.n64 0.136036
R212 dffrs_10.resetb reset.n72 0.136036
R213 dffrs_4.resetb reset.n78 0.136036
R214 dffrs_11.resetb reset.n86 0.136036
R215 dffrs_5.resetb reset.n92 0.136036
R216 dffrs_12.resetb reset.n5 0.136036
R217 reset.n7 dffrs_13.nand3_2.C 0.0455
R218 reset.n12 dffrs_14.nand3_7.A 0.0455
R219 reset.n18 dffrs_0.nand3_7.A 0.0455
R220 reset.n26 dffrs_7.nand3_7.A 0.0455
R221 reset.n32 dffrs_1.nand3_7.A 0.0455
R222 reset.n40 dffrs_8.nand3_7.A 0.0455
R223 reset.n46 dffrs_2.nand3_7.A 0.0455
R224 reset.n54 dffrs_9.nand3_7.A 0.0455
R225 reset.n60 dffrs_3.nand3_7.A 0.0455
R226 reset.n68 dffrs_10.nand3_7.A 0.0455
R227 reset.n74 dffrs_4.nand3_7.A 0.0455
R228 reset.n82 dffrs_11.nand3_7.A 0.0455
R229 reset.n88 dffrs_5.nand3_7.A 0.0455
R230 reset.n1 dffrs_12.nand3_7.A 0.0455
R231 dffrs_13.nand3_0.C reset.n9 0.0374643
R232 dffrs_5.Qb.n0 dffrs_5.Qb.t7 41.0041
R233 dffrs_5.Qb.n4 dffrs_5.Qb.t8 40.6313
R234 dffrs_5.Qb.n2 dffrs_5.Qb.t5 40.6313
R235 dffrs_5.Qb dffrs_12.setb 28.013
R236 dffrs_5.Qb.n4 dffrs_5.Qb.t4 27.3166
R237 dffrs_5.Qb.n2 dffrs_5.Qb.t6 27.3166
R238 dffrs_5.Qb.n0 dffrs_5.Qb.t9 26.9438
R239 dffrs_5.Qb.n9 dffrs_5.Qb.t1 10.0473
R240 dffrs_5.Qb.n6 dffrs_5.Qb.n1 9.84255
R241 dffrs_5.Qb.n5 dffrs_5.Qb.n3 9.22229
R242 dffrs_5.Qb.n8 dffrs_5.Qb.t2 6.51042
R243 dffrs_5.Qb.n8 dffrs_5.Qb.n7 6.04952
R244 dffrs_5.Qb.n1 dffrs_5.Qb.n0 5.7305
R245 dffrs_5.Qb.n5 dffrs_5.Qb.n4 5.14711
R246 dffrs_5.Qb.n3 dffrs_5.Qb.n2 5.13907
R247 dffrs_5.nand3_7.Z dffrs_5.Qb.n6 4.94976
R248 dffrs_5.nand3_7.Z dffrs_5.Qb.n9 4.72925
R249 dffrs_12.setb dffrs_12.nand3_0.C 0.784786
R250 dffrs_5.Qb.n9 dffrs_5.Qb.n8 0.732092
R251 dffrs_5.Qb.n7 dffrs_5.Qb.t3 0.7285
R252 dffrs_5.Qb.n7 dffrs_5.Qb.t0 0.7285
R253 dffrs_5.Qb.n6 dffrs_5.Qb 0.175225
R254 dffrs_5.Qb.n1 dffrs_5.nand3_2.A 0.0455
R255 dffrs_5.Qb.n3 dffrs_12.nand3_2.C 0.0455
R256 dffrs_12.nand3_0.C dffrs_5.Qb.n5 0.0374643
R257 vss.n754 vss.n134 6961.73
R258 vss.n764 vss.n132 6188.84
R259 vss.n320 vss.n319 5575.1
R260 vss.n140 vss.n91 5557.62
R261 vss.n915 vss.n24 5557.62
R262 vss.n366 vss.n263 5557.62
R263 vss.n529 vss.n201 5557.62
R264 vss.n576 vss.n182 5557.62
R265 vss.n162 vss.n27 5557.62
R266 vss.n617 vss.n164 5557.62
R267 vss.n673 vss.n672 5557.62
R268 vss.n753 vss.n733 5557.62
R269 vss.n882 vss.n58 5557.62
R270 vss.n317 vss.n237 5557.62
R271 vss.n378 vss.n253 5557.62
R272 vss.n463 vss.n434 5557.62
R273 vss.n418 vss.n237 5551.58
R274 vss.n366 vss.n201 5551.58
R275 vss.n182 vss.n24 5551.58
R276 vss.n617 vss.n162 5551.58
R277 vss.n672 vss.n140 5551.58
R278 vss.n754 vss.n753 5551.58
R279 vss.n848 vss.n58 5551.58
R280 vss.n733 vss.n732 5551.58
R281 vss.n812 vss.n91 5551.58
R282 vss.n561 vss.n164 5551.58
R283 vss.n576 vss.n575 5551.58
R284 vss.n529 vss.n528 5551.58
R285 vss.n384 vss.n378 5551.58
R286 vss.n463 vss.n462 5551.58
R287 vss.n674 vss.n132 4595.28
R288 vss.n316 vss.n307 4591.35
R289 vss.n678 vss.n677 4448.54
R290 vss.n869 vss.n868 4272.42
R291 vss.n317 vss.n316 3944.59
R292 vss.n79 vss.n57 3217.05
R293 vss.n856 vss.n839 3214.99
R294 vss.n335 vss.n334 3157.03
R295 vss.n917 vss.n916 3157.03
R296 vss.n912 vss.n911 3157.03
R297 vss.n150 vss.n139 3157.03
R298 vss.n780 vss.n122 3157.03
R299 vss.n651 vss.n99 3157.03
R300 vss.n610 vss.n609 3157.03
R301 vss.n919 vss.n19 3157.03
R302 vss.n931 vss.n8 3157.03
R303 vss.n396 vss.n245 3157.03
R304 vss.n931 vss.n7 3155.01
R305 vss.n919 vss.n918 3155.01
R306 vss.n610 vss.n28 3155.01
R307 vss.n652 vss.n651 3155.01
R308 vss.n718 vss.n717 3155.01
R309 vss.n798 vss.n797 3155.01
R310 vss.n608 vss.n167 3155.01
R311 vss.n536 vss.n535 3155.01
R312 vss.n515 vss.n514 3155.01
R313 vss.n397 vss.n228 3155.01
R314 vss.n780 vss.n121 3148.94
R315 vss.n883 vss.n56 2696.12
R316 vss.n870 vss.n56 2696.12
R317 vss.n870 vss.n869 2696.12
R318 vss.n134 vss.n132 2425.47
R319 vss.n281 vss.n280 2370
R320 vss.n347 vss.n23 2370
R321 vss.n336 vss.n332 2370
R322 vss.n914 vss.n913 2370
R323 vss.n440 vss.n227 2289.83
R324 vss.n678 vss.n132 2247.51
R325 vss.n335 vss.n263 1873.97
R326 vss.n916 vss.n915 1873.97
R327 vss.n912 vss.n27 1873.97
R328 vss.n673 vss.n139 1873.97
R329 vss.n253 vss.n245 1873.97
R330 vss.n883 vss.n882 1861.56
R331 vss.n884 vss.n55 1639.91
R332 vss.n59 vss.n56 1555.45
R333 vss.n871 vss.n870 1555.45
R334 vss.n869 vss.n69 1555.45
R335 vss.n764 vss.n763 1399.38
R336 vss.n763 vss.n55 1399.38
R337 vss.n420 vss.n228 1336.25
R338 vss.n742 vss.n57 1314.68
R339 vss.n433 vss.n432 1230.04
R340 vss.n316 vss.n315 1111.18
R341 vss.n883 vss.n57 1095.12
R342 vss.n433 vss.n228 1094.63
R343 vss.n304 vss.n227 1057.6
R344 vss.n434 vss.n433 978.216
R345 vss.n319 vss.n317 929.813
R346 vss.n306 vss.n305 904.735
R347 vss.n367 vss.n366 832.22
R348 vss.n672 vss.n664 832.22
R349 vss.n356 vss.n24 832.22
R350 vss.n162 vss.n160 832.22
R351 vss.n754 vss.n691 832.22
R352 vss.n830 vss.n58 832.22
R353 vss.n733 vss.n698 832.22
R354 vss.n105 vss.n91 832.22
R355 vss.n599 vss.n164 832.22
R356 vss.n577 vss.n576 832.22
R357 vss.n529 vss.n202 832.22
R358 vss.n308 vss.n237 832.22
R359 vss.n378 vss.n254 832.22
R360 vss.n464 vss.n463 832.22
R361 vss.n366 vss.n365 832.101
R362 vss.n272 vss.n24 832.101
R363 vss.n162 vss.n161 832.101
R364 vss.n672 vss.n671 832.101
R365 vss.n755 vss.n754 832.101
R366 vss.n68 vss.n58 832.101
R367 vss.n733 vss.n699 832.101
R368 vss.n710 vss.n91 832.101
R369 vss.n164 vss.n163 832.101
R370 vss.n576 vss.n183 832.101
R371 vss.n530 vss.n529 832.101
R372 vss.n244 vss.n237 832.101
R373 vss.n378 vss.n377 832.101
R374 vss.n463 vss.n435 832.101
R375 vss.n718 vss.n709 808.29
R376 vss.n798 vss.n98 808.29
R377 vss.n555 vss.n167 808.29
R378 vss.n536 vss.n198 808.29
R379 vss.n515 vss.n210 808.29
R380 vss.n856 vss.n855 794.258
R381 vss.n719 vss.n718 752.159
R382 vss.n799 vss.n798 752.159
R383 vss.n546 vss.n167 752.159
R384 vss.n537 vss.n536 752.159
R385 vss.n516 vss.n515 752.159
R386 vss.n336 vss.n335 745.506
R387 vss.n916 vss.n23 745.506
R388 vss.n913 vss.n912 745.506
R389 vss.n281 vss.n139 745.506
R390 vss.n320 vss.n245 745.506
R391 vss.n857 vss.n856 738.126
R392 vss.n884 vss.n883 648.605
R393 vss.n526 vss.t33 589.511
R394 vss.t319 vss.n193 589.511
R395 vss.n573 vss.t204 589.511
R396 vss.n545 vss.t164 589.511
R397 vss.n554 vss.t316 589.511
R398 vss.n800 vss.t86 589.511
R399 vss.n810 vss.t199 589.511
R400 vss.n704 vss.t81 589.511
R401 vss.n730 vss.t328 589.511
R402 vss.n858 vss.t200 589.511
R403 vss.n840 vss.t213 589.511
R404 vss.n868 vss.t0 589.511
R405 vss.n460 vss.t71 589.511
R406 vss.n517 vss.t338 589.511
R407 vss.n333 vss.t233 582.165
R408 vss.n367 vss.t307 582.165
R409 vss.n149 vss.t36 582.165
R410 vss.n664 vss.t238 582.165
R411 vss.t30 vss.n22 582.165
R412 vss.n356 vss.t103 582.165
R413 vss.n910 vss.t29 582.165
R414 vss.n160 vss.t94 582.165
R415 vss.n676 vss.t119 582.165
R416 vss.n691 vss.t78 582.165
R417 vss.n831 vss.t242 582.165
R418 vss.t282 vss.n830 582.165
R419 vss.n692 vss.t324 582.165
R420 vss.n698 vss.t189 582.165
R421 vss.t118 vss.n104 582.165
R422 vss.n105 vss.t157 582.165
R423 vss.t105 vss.n166 582.165
R424 vss.n599 vss.t155 582.165
R425 vss.n578 vss.t309 582.165
R426 vss.t149 vss.n577 582.165
R427 vss.n215 vss.t11 582.165
R428 vss.t144 vss.n202 582.165
R429 vss.n315 vss.t179 582.165
R430 vss.n308 vss.t247 582.165
R431 vss.n395 vss.t2 582.165
R432 vss.n254 vss.t14 582.165
R433 vss.n465 vss.t246 582.165
R434 vss.t142 vss.n464 582.165
R435 vss.t54 vss.n419 581.712
R436 vss.n420 vss.t333 581.712
R437 vss.n459 vss.t193 581.712
R438 vss.t222 vss.n209 581.712
R439 vss.n204 vss.t252 581.712
R440 vss.n538 vss.t127 581.712
R441 vss.t197 vss.n185 581.712
R442 vss.n547 vss.t9 581.712
R443 vss.n563 vss.t312 581.712
R444 vss.t19 vss.n97 581.712
R445 vss.t166 vss.n92 581.712
R446 vss.n720 vss.t17 581.712
R447 vss.n729 vss.t259 581.712
R448 vss.t73 vss.n78 581.712
R449 vss.n783 vss.t16 581.712
R450 vss.t182 vss.n782 581.712
R451 vss.n490 vss.t24 581.712
R452 vss.n484 vss.t153 581.712
R453 vss.n584 vss.t133 581.712
R454 vss.t146 vss.n17 581.712
R455 vss.n922 vss.t192 581.712
R456 vss.t321 vss.n921 581.712
R457 vss.n383 vss.t181 581.712
R458 vss.t97 vss.n5 581.712
R459 vss.n474 vss.t216 581.712
R460 vss.t187 vss.n6 581.712
R461 vss.t315 vss.n348 581.712
R462 vss.n349 vss.t310 581.712
R463 vss.n338 vss.t96 581.712
R464 vss.t12 vss.n337 581.712
R465 vss.n365 vss.t226 581.712
R466 vss.t31 vss.n21 581.712
R467 vss.n493 vss.t67 581.712
R468 vss.t220 vss.n492 581.712
R469 vss.n279 vss.t258 581.712
R470 vss.n282 vss.t116 581.712
R471 vss.t42 vss.n117 581.712
R472 vss.n119 vss.t3 581.712
R473 vss.t306 vss.n675 581.712
R474 vss.n679 vss.t240 581.712
R475 vss.n133 vss.t132 581.712
R476 vss.n765 vss.t76 581.712
R477 vss.n741 vss.t225 581.712
R478 vss.n735 vss.t130 581.712
R479 vss.n750 vss.t251 581.712
R480 vss.n742 vss.t185 581.712
R481 vss.n272 vss.t203 581.712
R482 vss.t49 vss.n271 581.712
R483 vss.t219 vss.n25 581.712
R484 vss.n26 vss.t106 581.712
R485 vss.n161 vss.t120 581.712
R486 vss.n653 vss.t39 581.712
R487 vss.n619 vss.t177 581.712
R488 vss.t256 vss.n152 581.712
R489 vss.n621 vss.t21 581.712
R490 vss.t151 vss.n153 581.712
R491 vss.n671 vss.t141 581.712
R492 vss.n665 vss.t253 581.712
R493 vss.n755 vss.t176 581.712
R494 vss.n762 vss.t65 581.712
R495 vss.n881 vss.t7 581.712
R496 vss.n59 vss.t276 581.712
R497 vss.t93 vss.n68 581.712
R498 vss.n871 vss.t172 581.712
R499 vss.n846 vss.t99 581.712
R500 vss.t325 vss.n69 581.712
R501 vss.n699 vss.t89 581.712
R502 vss.n838 vss.t236 581.712
R503 vss.n710 vss.t109 581.712
R504 vss.n716 vss.t114 581.712
R505 vss.n163 vss.t102 581.712
R506 vss.n796 vss.t194 581.712
R507 vss.n183 vss.t100 581.712
R508 vss.n607 vss.t135 581.712
R509 vss.n530 vss.t92 581.712
R510 vss.n534 vss.t162 581.712
R511 vss.t215 vss.n244 581.712
R512 vss.n398 vss.t137 581.712
R513 vss.n318 vss.t332 581.712
R514 vss.n321 vss.t249 581.712
R515 vss.n377 vss.t59 581.712
R516 vss.n255 vss.t234 581.712
R517 vss.n435 vss.t91 581.712
R518 vss.n513 vss.t43 581.712
R519 vss.n882 vss.n881 548.236
R520 vss.n419 vss.n418 548.058
R521 vss.n384 vss.n383 548.058
R522 vss.n418 vss.n417 484.702
R523 vss.n385 vss.n384 484.702
R524 vss.t33 vss.t301 471.61
R525 vss.t301 vss.t319 471.61
R526 vss.t290 vss.t204 471.61
R527 vss.t164 vss.t290 471.61
R528 vss.t316 vss.t272 471.61
R529 vss.t272 vss.t86 471.61
R530 vss.t286 vss.t199 471.61
R531 vss.t81 vss.t286 471.61
R532 vss.t328 vss.t269 471.61
R533 vss.t269 vss.t200 471.61
R534 vss.t213 vss.t148 471.61
R535 vss.t148 vss.t0 471.61
R536 vss.t71 vss.t287 471.61
R537 vss.t287 vss.t338 471.61
R538 vss.t233 vss.t314 465.733
R539 vss.t314 vss.t307 465.733
R540 vss.t36 vss.t5 465.733
R541 vss.t5 vss.t238 465.733
R542 vss.t218 vss.t30 465.733
R543 vss.t103 vss.t218 465.733
R544 vss.t171 vss.t29 465.733
R545 vss.t94 vss.t171 465.733
R546 vss.t119 vss.t134 465.733
R547 vss.t134 vss.t78 465.733
R548 vss.t242 vss.t327 465.733
R549 vss.t327 vss.t282 465.733
R550 vss.t324 vss.t72 465.733
R551 vss.t72 vss.t189 465.733
R552 vss.t305 vss.t118 465.733
R553 vss.t157 vss.t305 465.733
R554 vss.t6 vss.t105 465.733
R555 vss.t155 vss.t6 465.733
R556 vss.t309 vss.t8 465.733
R557 vss.t8 vss.t149 465.733
R558 vss.t11 vss.t129 465.733
R559 vss.t129 vss.t144 465.733
R560 vss.t331 vss.t179 465.733
R561 vss.t247 vss.t331 465.733
R562 vss.t113 vss.t2 465.733
R563 vss.t14 vss.t113 465.733
R564 vss.t246 vss.t217 465.733
R565 vss.t217 vss.t142 465.733
R566 vss.t209 vss.t54 465.37
R567 vss.t333 vss.t209 465.37
R568 vss.t193 vss.t111 465.37
R569 vss.t111 vss.t222 465.37
R570 vss.t252 vss.t112 465.37
R571 vss.t112 vss.t127 465.37
R572 vss.t110 vss.t197 465.37
R573 vss.t9 vss.t110 465.37
R574 vss.t312 vss.t90 465.37
R575 vss.t90 vss.t19 465.37
R576 vss.t323 vss.t166 465.37
R577 vss.t17 vss.t323 465.37
R578 vss.t259 vss.t101 465.37
R579 vss.t101 vss.t73 465.37
R580 vss.t16 vss.t167 465.37
R581 vss.t167 vss.t182 465.37
R582 vss.t196 vss.t24 465.37
R583 vss.t153 vss.t196 465.37
R584 vss.t133 vss.t261 465.37
R585 vss.t261 vss.t146 465.37
R586 vss.t192 vss.t337 465.37
R587 vss.t337 vss.t321 465.37
R588 vss.t181 vss.t58 465.37
R589 vss.t58 vss.t97 465.37
R590 vss.t216 vss.t198 465.37
R591 vss.t198 vss.t187 465.37
R592 vss.t191 vss.t315 465.37
R593 vss.t310 vss.t191 465.37
R594 vss.t96 vss.t180 465.37
R595 vss.t180 vss.t12 465.37
R596 vss.t226 vss.t266 465.37
R597 vss.t266 vss.t31 465.37
R598 vss.t67 vss.t170 465.37
R599 vss.t170 vss.t220 465.37
R600 vss.t258 vss.t178 465.37
R601 vss.t178 vss.t116 465.37
R602 vss.t245 vss.t42 465.37
R603 vss.t3 vss.t245 465.37
R604 vss.t41 vss.t306 465.37
R605 vss.t240 vss.t41 465.37
R606 vss.t132 vss.t224 465.37
R607 vss.t224 vss.t76 465.37
R608 vss.t260 vss.t225 465.37
R609 vss.t130 vss.t260 465.37
R610 vss.t160 vss.t251 465.37
R611 vss.t185 vss.t160 465.37
R612 vss.t203 vss.t293 465.37
R613 vss.t293 vss.t49 465.37
R614 vss.t68 vss.t219 465.37
R615 vss.t106 vss.t68 465.37
R616 vss.t120 vss.t275 465.37
R617 vss.t275 vss.t39 465.37
R618 vss.t177 vss.t123 465.37
R619 vss.t123 vss.t256 465.37
R620 vss.t21 vss.t313 465.37
R621 vss.t313 vss.t151 465.37
R622 vss.t299 vss.t141 465.37
R623 vss.t253 vss.t299 465.37
R624 vss.t176 vss.t273 465.37
R625 vss.t273 vss.t65 465.37
R626 vss.t45 vss.t7 465.37
R627 vss.t276 vss.t45 465.37
R628 vss.t159 vss.t93 465.37
R629 vss.t172 vss.t159 465.37
R630 vss.t99 vss.t88 465.37
R631 vss.t88 vss.t325 465.37
R632 vss.t89 vss.t274 465.37
R633 vss.t274 vss.t236 465.37
R634 vss.t109 vss.t289 465.37
R635 vss.t289 vss.t114 465.37
R636 vss.t102 vss.t298 465.37
R637 vss.t298 vss.t194 465.37
R638 vss.t100 vss.t270 465.37
R639 vss.t270 vss.t135 465.37
R640 vss.t92 vss.t263 465.37
R641 vss.t263 vss.t162 465.37
R642 vss.t264 vss.t215 465.37
R643 vss.t137 vss.t264 465.37
R644 vss.t332 vss.t53 465.37
R645 vss.t53 vss.t249 465.37
R646 vss.t296 vss.t59 465.37
R647 vss.t234 vss.t296 465.37
R648 vss.t91 vss.t271 465.37
R649 vss.t271 vss.t43 465.37
R650 vss.n931 vss.n930 435.214
R651 vss.n919 vss.n20 435.214
R652 vss.n611 vss.n610 435.214
R653 vss.n651 vss.n650 435.214
R654 vss.n780 vss.n779 435.012
R655 vss.n932 vss.n931 404.991
R656 vss.n920 vss.n919 404.991
R657 vss.n610 vss.n165 404.991
R658 vss.n651 vss.n644 404.991
R659 vss.n781 vss.n780 404.803
R660 vss.n934 vss.t231 366.243
R661 vss.t62 vss.n933 366.243
R662 vss.n478 vss.t27 366.243
R663 vss.t56 vss.n18 366.243
R664 vss.n496 vss.t25 366.243
R665 vss.t51 vss.n495 366.243
R666 vss.n633 vss.t230 366.243
R667 vss.t228 vss.n120 366.243
R668 vss.n618 vss.t232 366.243
R669 vss.n643 vss.t46 366.243
R670 vss.n751 vss.t26 365.705
R671 vss.n885 vss.t205 365.705
R672 vss.n307 vss.t279 338.849
R673 vss.n417 vss.t60 338.849
R674 vss.t278 vss.n229 338.849
R675 vss.n385 vss.t335 338.849
R676 vss.n849 vss.n848 307.786
R677 vss.n732 vss.n700 307.786
R678 vss.n813 vss.n812 307.786
R679 vss.n561 vss.n560 307.786
R680 vss.n575 vss.n184 307.786
R681 vss.n528 vss.n203 307.786
R682 vss.n462 vss.n436 307.786
R683 vss.t231 vss.t262 292.995
R684 vss.t262 vss.t62 292.995
R685 vss.t27 vss.t284 292.995
R686 vss.t284 vss.t56 292.995
R687 vss.t25 vss.t302 292.995
R688 vss.t302 vss.t51 292.995
R689 vss.t230 vss.t268 292.995
R690 vss.t268 vss.t228 292.995
R691 vss.t232 vss.t292 292.995
R692 vss.t292 vss.t46 292.995
R693 vss.t26 vss.t285 292.565
R694 vss.t285 vss.t205 292.565
R695 vss.t126 vss.t60 271.079
R696 vss.t64 vss.t278 271.079
R697 vss.t335 vss.t64 271.079
R698 vss.n848 vss.n847 251.655
R699 vss.n732 vss.n731 251.655
R700 vss.n812 vss.n811 251.655
R701 vss.n562 vss.n561 251.655
R702 vss.n575 vss.n574 251.655
R703 vss.n528 vss.n527 251.655
R704 vss.n462 vss.n461 251.655
R705 vss.n347 vss.n263 249.429
R706 vss.n915 vss.n914 249.429
R707 vss.n280 vss.n27 249.429
R708 vss.n674 vss.n673 249.429
R709 vss.n332 vss.n253 249.429
R710 vss.n855 vss.t184 215.171
R711 vss.n849 vss.t329 215.171
R712 vss.n709 vss.t267 215.171
R713 vss.t139 vss.n700 215.171
R714 vss.n98 vss.t280 215.171
R715 vss.n813 vss.t317 215.171
R716 vss.n555 vss.t294 215.171
R717 vss.n560 vss.t83 215.171
R718 vss.n198 vss.t297 215.171
R719 vss.t34 vss.n184 215.171
R720 vss.n210 vss.t303 215.171
R721 vss.t69 vss.n203 215.171
R722 vss.n440 vss.t304 215.171
R723 vss.t22 vss.n436 215.171
R724 vss.n434 vss.n4 205.9
R725 vss.n433 vss.n229 178.264
R726 vss.n432 vss.t124 176.048
R727 vss.t28 vss.t184 172.137
R728 vss.t329 vss.t28 172.137
R729 vss.t267 vss.t202 172.137
R730 vss.t202 vss.t139 172.137
R731 vss.t280 vss.t108 172.137
R732 vss.t108 vss.t317 172.137
R733 vss.t294 vss.t85 172.137
R734 vss.t85 vss.t83 172.137
R735 vss.t297 vss.t161 172.137
R736 vss.t161 vss.t34 172.137
R737 vss.t303 vss.t255 172.137
R738 vss.t255 vss.t69 172.137
R739 vss.t304 vss.t75 172.137
R740 vss.t75 vss.t22 172.137
R741 vss.n201 vss.n200 165.725
R742 vss.n182 vss.n181 165.725
R743 vss.n617 vss.n616 165.725
R744 vss.n645 vss.n140 165.725
R745 vss.n753 vss.n734 165.648
R746 vss.n306 vss.t126 162.059
R747 vss.n527 vss.n526 153.786
R748 vss.n537 vss.n193 153.786
R749 vss.n574 vss.n573 153.786
R750 vss.n546 vss.n545 153.786
R751 vss.n562 vss.n554 153.786
R752 vss.n800 vss.n799 153.786
R753 vss.n811 vss.n810 153.786
R754 vss.n719 vss.n704 153.786
R755 vss.n731 vss.n730 153.786
R756 vss.n858 vss.n857 153.786
R757 vss.n847 vss.n840 153.786
R758 vss.n461 vss.n460 153.786
R759 vss.n517 vss.n516 153.786
R760 vss.n334 vss.n333 151.869
R761 vss.n150 vss.n149 151.869
R762 vss.n917 vss.n22 151.869
R763 vss.n911 vss.n910 151.869
R764 vss.n677 vss.n676 151.869
R765 vss.n831 vss.n79 151.869
R766 vss.n692 vss.n122 151.869
R767 vss.n104 vss.n99 151.869
R768 vss.n609 vss.n166 151.869
R769 vss.n578 vss.n19 151.869
R770 vss.n215 vss.n8 151.869
R771 vss.n396 vss.n395 151.869
R772 vss.n465 vss.n227 151.869
R773 vss.n461 vss.n459 151.751
R774 vss.n516 vss.n209 151.751
R775 vss.n527 vss.n204 151.751
R776 vss.n538 vss.n537 151.751
R777 vss.n574 vss.n185 151.751
R778 vss.n547 vss.n546 151.751
R779 vss.n563 vss.n562 151.751
R780 vss.n799 vss.n97 151.751
R781 vss.n811 vss.n92 151.751
R782 vss.n720 vss.n719 151.751
R783 vss.n731 vss.n729 151.751
R784 vss.n857 vss.n78 151.751
R785 vss.n783 vss.n116 151.751
R786 vss.n782 vss.n781 151.751
R787 vss.n494 vss.n490 151.751
R788 vss.n484 vss.n165 151.751
R789 vss.n584 vss.n16 151.751
R790 vss.n920 vss.n17 151.751
R791 vss.n922 vss.n16 151.751
R792 vss.n921 vss.n920 151.751
R793 vss.n932 vss.n5 151.751
R794 vss.n474 vss.n4 151.751
R795 vss.n932 vss.n6 151.751
R796 vss.n348 vss.n347 151.751
R797 vss.n349 vss.n23 151.751
R798 vss.n338 vss.n332 151.751
R799 vss.n337 vss.n336 151.751
R800 vss.n918 vss.n21 151.751
R801 vss.n494 vss.n493 151.751
R802 vss.n492 vss.n165 151.751
R803 vss.n280 vss.n279 151.751
R804 vss.n282 vss.n281 151.751
R805 vss.n117 vss.n116 151.751
R806 vss.n781 vss.n119 151.751
R807 vss.n675 vss.n674 151.751
R808 vss.n679 vss.n678 151.751
R809 vss.n134 vss.n133 151.751
R810 vss.n765 vss.n764 151.751
R811 vss.n752 vss.n741 151.751
R812 vss.n735 vss.n55 151.751
R813 vss.n752 vss.n750 151.751
R814 vss.n271 vss.n28 151.751
R815 vss.n914 vss.n25 151.751
R816 vss.n913 vss.n26 151.751
R817 vss.n653 vss.n652 151.751
R818 vss.n620 vss.n619 151.751
R819 vss.n644 vss.n152 151.751
R820 vss.n621 vss.n620 151.751
R821 vss.n644 vss.n153 151.751
R822 vss.n665 vss.n121 151.751
R823 vss.n763 vss.n762 151.751
R824 vss.n847 vss.n846 151.751
R825 vss.n839 vss.n838 151.751
R826 vss.n717 vss.n716 151.751
R827 vss.n797 vss.n796 151.751
R828 vss.n608 vss.n607 151.751
R829 vss.n535 vss.n534 151.751
R830 vss.n398 vss.n397 151.751
R831 vss.n319 vss.n318 151.751
R832 vss.n321 vss.n320 151.751
R833 vss.n255 vss.n7 151.751
R834 vss.n514 vss.n513 151.751
R835 vss.t211 vss.t281 140.839
R836 vss.t281 vss.t124 140.839
R837 vss.n201 vss.n16 135.501
R838 vss.n494 vss.n182 135.501
R839 vss.n620 vss.n617 135.501
R840 vss.n140 vss.n116 135.501
R841 vss.n753 vss.n752 135.439
R842 vss.n930 vss.t295 115.856
R843 vss.n200 vss.t168 115.856
R844 vss.t288 vss.n20 115.856
R845 vss.n181 vss.t121 115.856
R846 vss.n611 vss.t300 115.856
R847 vss.n616 vss.t243 115.856
R848 vss.n650 vss.t291 115.856
R849 vss.n645 vss.t174 115.856
R850 vss.n779 vss.t265 115.802
R851 vss.n734 vss.t37 115.802
R852 vss.t279 vss.n306 109.022
R853 vss.n304 vss.t211 102.567
R854 vss.n934 vss.n4 95.5419
R855 vss.n933 vss.n932 95.5419
R856 vss.n478 vss.n16 95.5419
R857 vss.n920 vss.n18 95.5419
R858 vss.n496 vss.n494 95.5419
R859 vss.n495 vss.n165 95.5419
R860 vss.n633 vss.n116 95.5419
R861 vss.n781 vss.n120 95.5419
R862 vss.n620 vss.n618 95.5419
R863 vss.n644 vss.n643 95.5419
R864 vss.n752 vss.n751 95.4017
R865 vss.n885 vss.n884 95.4017
R866 vss.t80 vss.t295 92.6849
R867 vss.t168 vss.t80 92.6849
R868 vss.t55 vss.t288 92.6849
R869 vss.t121 vss.t55 92.6849
R870 vss.t300 vss.t48 92.6849
R871 vss.t48 vss.t243 92.6849
R872 vss.t227 vss.t291 92.6849
R873 vss.t174 vss.t227 92.6849
R874 vss.t207 vss.t265 92.6419
R875 vss.t37 vss.t207 92.6419
R876 vss.n305 vss.n304 73.4814
R877 vss.n416 vss.n238 61.0571
R878 vss.n350 vss.n346 61.0571
R879 vss.n480 vss.n479 61.0571
R880 vss.n491 vss.n41 61.0571
R881 vss.n497 vss.n483 61.0571
R882 vss.n283 vss.n278 61.0571
R883 vss.n118 vss.n48 61.0571
R884 vss.n635 vss.n634 61.0571
R885 vss.n663 vss.n141 61.0571
R886 vss.n680 vss.n138 61.0571
R887 vss.n766 vss.n131 61.0571
R888 vss.n740 vss.n736 61.0571
R889 vss.n749 vss.n743 61.0571
R890 vss.n867 vss.n70 61.0571
R891 vss.n106 vss.n103 61.0571
R892 vss.n217 vss.n216 61.0571
R893 vss.n518 vss.n208 61.0571
R894 vss.n442 vss.n441 61.0561
R895 vss.n512 vss.n211 61.0561
R896 vss.n466 vss.n226 61.0561
R897 vss.n431 vss.n230 61.0561
R898 vss.n387 vss.n386 61.0561
R899 vss.n376 vss.n256 61.0561
R900 vss.n394 vss.n246 61.0561
R901 vss.n322 vss.n303 61.0561
R902 vss.n399 vss.n243 61.0561
R903 vss.n314 vss.n309 61.0561
R904 vss.n421 vss.n236 61.0561
R905 vss.n450 vss.n449 61.0561
R906 vss.n458 vss.n437 61.0561
R907 vss.n533 vss.n531 61.0561
R908 vss.n197 vss.n194 61.0561
R909 vss.n525 vss.n205 61.0561
R910 vss.n539 vss.n192 61.0561
R911 vss.n606 vss.n168 61.0561
R912 vss.n559 vss.n556 61.0561
R913 vss.n572 vss.n186 61.0561
R914 vss.n548 vss.n544 61.0561
R915 vss.n795 vss.n100 61.0561
R916 vss.n601 vss.n600 61.0561
R917 vss.n814 vss.n90 61.0561
R918 vss.n801 vss.n96 61.0561
R919 vss.n564 vss.n553 61.0561
R920 vss.n715 vss.n711 61.0561
R921 vss.n708 vss.n705 61.0561
R922 vss.n809 vss.n93 61.0561
R923 vss.n721 vss.n703 61.0561
R924 vss.n837 vss.n80 61.0561
R925 vss.n697 vss.n693 61.0561
R926 vss.n845 vss.n841 61.0561
R927 vss.n854 vss.n850 61.0561
R928 vss.n859 vss.n77 61.0561
R929 vss.n728 vss.n701 61.0561
R930 vss.n872 vss.n67 61.0561
R931 vss.n880 vss.n60 61.0561
R932 vss.n886 vss.n54 61.0561
R933 vss.n778 vss.n123 61.0561
R934 vss.n761 vss.n756 61.0561
R935 vss.n690 vss.n135 61.0561
R936 vss.n670 vss.n666 61.0561
R937 vss.n649 vss.n646 61.0561
R938 vss.n784 vss.n115 61.0561
R939 vss.n642 vss.n154 61.0561
R940 vss.n624 vss.n622 61.0561
R941 vss.n151 vss.n44 61.0561
R942 vss.n615 vss.n612 61.0561
R943 vss.n654 vss.n148 61.0561
R944 vss.n909 vss.n29 61.0561
R945 vss.n293 vss.n291 61.0561
R946 vss.n180 vss.n178 61.0561
R947 vss.n489 vss.n485 61.0561
R948 vss.n273 vss.n270 61.0561
R949 vss.n358 vss.n357 61.0561
R950 vss.n923 vss.n15 61.0561
R951 vss.n586 vss.n585 61.0561
R952 vss.n929 vss.n9 61.0561
R953 vss.n935 vss.n3 61.0561
R954 vss.n475 vss.n473 61.0561
R955 vss.n382 vss.n380 61.0561
R956 vss.n364 vss.n264 61.0561
R957 vss.n368 vss.n262 61.0561
R958 vss.n339 vss.n331 61.0561
R959 vss.n832 vss.n829 61.0561
R960 vss.n579 vss.n177 61.0561
R961 vss.n401 vss.t343 41.0041
R962 vss.n427 vss.t341 41.0041
R963 vss.n72 vss.t340 41.0041
R964 vss.n402 vss.t342 40.8177
R965 vss.n402 vss.t208 27.1302
R966 vss.n401 vss.t214 26.9438
R967 vss.n427 vss.t210 26.9438
R968 vss.n72 vss.t212 26.9438
R969 vss.n864 dffrs_13.d 13.7563
R970 vss.n404 dffrs_12.clk 13.599
R971 vss.n428 dffrs_12.d 13.599
R972 vss.n865 vss.n864 9.04466
R973 vss.n429 vss.n428 9.04027
R974 vss.n232 vss.n231 9.03475
R975 vss.n438 vss.n207 9.03475
R976 vss.n325 vss.n324 9.0005
R977 vss.n406 vss.n405 9.0005
R978 vss.n412 vss.n235 9.0005
R979 vss.n793 vss.n792 9.0005
R980 vss.n835 vss.n834 9.0005
R981 vss.n250 vss.n248 9.0005
R982 vss.n363 vss.n362 9.0005
R983 vss.n345 vss.n344 9.0005
R984 vss.n370 vss.n259 9.0005
R985 vss.n372 vss.n371 9.0005
R986 vss.n372 vss.n258 9.0005
R987 vss.n375 vss.n374 9.0005
R988 vss.n341 vss.n340 9.0005
R989 vss.n329 vss.n260 9.0005
R990 vss.n500 vss.n499 9.0005
R991 vss.n900 vss.n899 9.0005
R992 vss.n631 vss.n155 9.0005
R993 vss.n297 vss.n296 9.0005
R994 vss.n275 vss.n274 9.0005
R995 vss.n34 vss.n31 9.0005
R996 vss.n286 vss.n285 9.0005
R997 vss.n657 vss.n656 9.0005
R998 vss.n897 vss.n896 9.0005
R999 vss.n640 vss.n639 9.0005
R1000 vss.n894 vss.n893 9.0005
R1001 vss.n637 vss.n53 9.0005
R1002 vss.n669 vss.n136 9.0005
R1003 vss.n661 vss.n660 9.0005
R1004 vss.n144 vss.n137 9.0005
R1005 vss.n770 vss.n769 9.0005
R1006 vss.n757 vss.n128 9.0005
R1007 vss.n688 vss.n127 9.0005
R1008 vss.n738 vss.n51 9.0005
R1009 vss.n888 vss.n52 9.0005
R1010 vss.n759 vss.n758 9.0005
R1011 vss.n768 vss.n130 9.0005
R1012 vss.n668 vss.n126 9.0005
R1013 vss.n687 vss.n686 9.0005
R1014 vss.n683 vss.n682 9.0005
R1015 vss.n748 vss.n747 9.0005
R1016 vss.n890 vss.n889 9.0005
R1017 vss.n739 vss.n50 9.0005
R1018 vss.n639 vss.n638 9.0005
R1019 vss.n896 vss.n895 9.0005
R1020 vss.n657 vss.n142 9.0005
R1021 vss.n147 vss.n146 9.0005
R1022 vss.n288 vss.n287 9.0005
R1023 vss.n907 vss.n33 9.0005
R1024 vss.n908 vss.n907 9.0005
R1025 vss.n295 vss.n292 9.0005
R1026 vss.n628 vss.n627 9.0005
R1027 vss.n632 vss.n631 9.0005
R1028 vss.n899 vss.n898 9.0005
R1029 vss.n499 vss.n498 9.0005
R1030 vss.n902 vss.n13 9.0005
R1031 vss.n902 vss.n901 9.0005
R1032 vss.n360 vss.n266 9.0005
R1033 vss.n353 vss.n352 9.0005
R1034 vss.n360 vss.n359 9.0005
R1035 vss.n354 vss.n268 9.0005
R1036 vss.n66 vss.n65 9.0005
R1037 vss.n879 vss.n878 9.0005
R1038 vss.n877 vss.n62 9.0005
R1039 vss.n875 vss.n874 9.0005
R1040 vss.n827 vss.n826 9.0005
R1041 vss.n843 vss.n74 9.0005
R1042 vss.n862 vss.n861 9.0005
R1043 vss.n862 vss.n71 9.0005
R1044 vss.n726 vss.n75 9.0005
R1045 vss.n844 vss.n75 9.0005
R1046 vss.n834 vss.n833 9.0005
R1047 vss.n745 vss.n82 9.0005
R1048 vss.n822 vss.n81 9.0005
R1049 vss.n695 vss.n84 9.0005
R1050 vss.n790 vss.n789 9.0005
R1051 vss.n712 vss.n108 9.0005
R1052 vss.n786 vss.n785 9.0005
R1053 vss.n713 vss.n85 9.0005
R1054 vss.n694 vss.n85 9.0005
R1055 vss.n113 vss.n112 9.0005
R1056 vss.n807 vss.n805 9.0005
R1057 vss.n805 vss.n76 9.0005
R1058 vss.n724 vss.n723 9.0005
R1059 vss.n727 vss.n724 9.0005
R1060 vss.n804 vss.n803 9.0005
R1061 vss.n808 vss.n804 9.0005
R1062 vss.n551 vss.n89 9.0005
R1063 vss.n702 vss.n89 9.0005
R1064 vss.n792 vss.n791 9.0005
R1065 vss.n626 vss.n623 9.0005
R1066 vss.n158 vss.n101 9.0005
R1067 vss.n597 vss.n596 9.0005
R1068 vss.n507 vss.n506 9.0005
R1069 vss.n199 vss.n173 9.0005
R1070 vss.n583 vss.n172 9.0005
R1071 vss.n502 vss.n1 9.0005
R1072 vss.n502 vss.n501 9.0005
R1073 vss.n925 vss.n11 9.0005
R1074 vss.n925 vss.n924 9.0005
R1075 vss.n937 vss.n936 9.0005
R1076 vss.n381 vss.n233 9.0005
R1077 vss.n393 vss.n392 9.0005
R1078 vss.n424 vss.n423 9.0005
R1079 vss.n302 vss.n301 9.0005
R1080 vss.n408 vss.n407 9.0005
R1081 vss.n313 vss.n310 9.0005
R1082 vss.n312 vss.n241 9.0005
R1083 vss.n457 vss.n439 9.0005
R1084 vss.n468 vss.n467 9.0005
R1085 vss.n224 vss.n223 9.0005
R1086 vss.n220 vss.n212 9.0005
R1087 vss.n477 vss.n476 9.0005
R1088 vss.n510 vss.n509 9.0005
R1089 vss.n509 vss.n508 9.0005
R1090 vss.n471 vss.n219 9.0005
R1091 vss.n521 vss.n520 9.0005
R1092 vss.n524 vss.n521 9.0005
R1093 vss.n456 vss.n454 9.0005
R1094 vss.n454 vss.n191 9.0005
R1095 vss.n523 vss.n187 9.0005
R1096 vss.n571 vss.n187 9.0005
R1097 vss.n542 vss.n541 9.0005
R1098 vss.n543 vss.n542 9.0005
R1099 vss.n581 vss.n174 9.0005
R1100 vss.n581 vss.n580 9.0005
R1101 vss.n589 vss.n588 9.0005
R1102 vss.n175 vss.n171 9.0005
R1103 vss.n593 vss.n169 9.0005
R1104 vss.n488 vss.n157 9.0005
R1105 vss.n604 vss.n603 9.0005
R1106 vss.n603 vss.n602 9.0005
R1107 vss.n487 vss.n156 9.0005
R1108 vss.n570 vss.n568 9.0005
R1109 vss.n568 vss.n95 9.0005
R1110 vss.n566 vss.n550 9.0005
R1111 vss.n566 vss.n565 9.0005
R1112 vss.n677 vss.n121 8.08508
R1113 vss.n444 vss.n441 6.9012
R1114 vss.n414 vss.n238 6.9012
R1115 vss.n388 vss.n387 6.9012
R1116 vss.n452 vss.n449 6.9012
R1117 vss.n197 vss.n196 6.9012
R1118 vss.n557 vss.n556 6.9012
R1119 vss.n816 vss.n90 6.9012
R1120 vss.n708 vss.n707 6.9012
R1121 vss.n854 vss.n853 6.9012
R1122 vss.n178 vss.n39 6.9012
R1123 vss.n929 vss.n928 6.9012
R1124 vss.n613 vss.n612 6.9012
R1125 vss.n649 vss.n648 6.9012
R1126 vss.n778 vss.n777 6.9012
R1127 vss.n212 vss.n211 6.46296
R1128 vss.n467 vss.n466 6.46296
R1129 vss.n407 vss.n243 6.46296
R1130 vss.n236 vss.n235 6.46296
R1131 vss.n458 vss.n457 6.46296
R1132 vss.n531 vss.n199 6.46296
R1133 vss.n192 vss.n191 6.46296
R1134 vss.n169 vss.n168 6.46296
R1135 vss.n544 vss.n543 6.46296
R1136 vss.n101 vss.n100 6.46296
R1137 vss.n565 vss.n564 6.46296
R1138 vss.n712 vss.n711 6.46296
R1139 vss.n703 vss.n702 6.46296
R1140 vss.n81 vss.n80 6.46296
R1141 vss.n845 vss.n844 6.46296
R1142 vss.n728 vss.n727 6.46296
R1143 vss.n924 vss.n923 6.46296
R1144 vss.n382 vss.n381 6.46296
R1145 vss.n394 vss.n393 6.46296
R1146 vss.n364 vss.n363 6.46296
R1147 vss.n371 vss.n262 6.46296
R1148 vss.n376 vss.n375 6.46296
R1149 vss.n901 vss.n41 6.46296
R1150 vss.n274 vss.n273 6.46296
R1151 vss.n909 vss.n908 6.46296
R1152 vss.n148 vss.n147 6.46296
R1153 vss.n898 vss.n44 6.46296
R1154 vss.n895 vss.n48 6.46296
R1155 vss.n670 vss.n669 6.46296
R1156 vss.n142 vss.n141 6.46296
R1157 vss.n757 vss.n756 6.46296
R1158 vss.n687 vss.n135 6.46296
R1159 vss.n740 vss.n739 6.46296
R1160 vss.n359 vss.n358 6.46296
R1161 vss.n67 vss.n66 6.46296
R1162 vss.n833 vss.n832 6.46296
R1163 vss.n694 vss.n693 6.46296
R1164 vss.n791 vss.n103 6.46296
R1165 vss.n602 vss.n601 6.46296
R1166 vss.n580 vss.n579 6.46296
R1167 vss.n508 vss.n216 6.46296
R1168 vss.n314 vss.n313 6.46296
R1169 vss.n303 vss.n302 6.4618
R1170 vss.n231 vss.n230 6.4618
R1171 vss.n525 vss.n524 6.4618
R1172 vss.n572 vss.n571 6.4618
R1173 vss.n96 vss.n95 6.4618
R1174 vss.n809 vss.n808 6.4618
R1175 vss.n77 vss.n76 6.4618
R1176 vss.n785 vss.n784 6.4618
R1177 vss.n489 vss.n488 6.4618
R1178 vss.n585 vss.n583 6.4618
R1179 vss.n936 vss.n935 6.4618
R1180 vss.n476 vss.n475 6.4618
R1181 vss.n346 vss.n345 6.4618
R1182 vss.n340 vss.n339 6.4618
R1183 vss.n501 vss.n479 6.4618
R1184 vss.n498 vss.n497 6.4618
R1185 vss.n296 vss.n291 6.4618
R1186 vss.n287 vss.n278 6.4618
R1187 vss.n632 vss.n154 6.4618
R1188 vss.n638 vss.n634 6.4618
R1189 vss.n138 vss.n137 6.4618
R1190 vss.n769 vss.n131 6.4618
R1191 vss.n889 vss.n54 6.4618
R1192 vss.n749 vss.n748 6.4618
R1193 vss.n627 vss.n622 6.4618
R1194 vss.n880 vss.n879 6.4618
R1195 vss.n71 vss.n70 6.4618
R1196 vss.n208 vss.n207 6.4618
R1197 dffrs_12.nand3_1.A vss.n401 5.7755
R1198 dffrs_12.nand3_8.A vss.n427 5.7755
R1199 dffrs_13.nand3_8.A vss.n72 5.7755
R1200 dffrs_12.nand3_6.B vss.n402 5.47979
R1201 vss.n444 vss.n443 5.47239
R1202 vss.n415 vss.n414 5.47239
R1203 vss.n452 vss.n451 5.47239
R1204 vss.n196 vss.n195 5.47239
R1205 vss.n558 vss.n557 5.47239
R1206 vss.n816 vss.n815 5.47239
R1207 vss.n707 vss.n706 5.47239
R1208 vss.n853 vss.n852 5.47239
R1209 vss.n928 vss.n927 5.47239
R1210 vss.n777 vss.n124 5.47239
R1211 vss.n648 vss.n647 5.47239
R1212 vss.n614 vss.n613 5.47239
R1213 vss.n179 vss.n39 5.47239
R1214 vss.n388 vss.n252 5.47239
R1215 vss.n511 vss.n510 5.03414
R1216 vss.n225 vss.n224 5.03414
R1217 vss.n312 vss.n311 5.03414
R1218 vss.n324 vss.n323 5.03414
R1219 vss.n406 vss.n400 5.03414
R1220 vss.n423 vss.n422 5.03414
R1221 vss.n430 vss.n429 5.03414
R1222 vss.n456 vss.n455 5.03414
R1223 vss.n532 vss.n174 5.03414
R1224 vss.n523 vss.n522 5.03414
R1225 vss.n541 vss.n540 5.03414
R1226 vss.n605 vss.n604 5.03414
R1227 vss.n570 vss.n569 5.03414
R1228 vss.n550 vss.n549 5.03414
R1229 vss.n598 vss.n597 5.03414
R1230 vss.n794 vss.n793 5.03414
R1231 vss.n803 vss.n802 5.03414
R1232 vss.n552 vss.n551 5.03414
R1233 vss.n714 vss.n713 5.03414
R1234 vss.n807 vss.n806 5.03414
R1235 vss.n723 vss.n722 5.03414
R1236 vss.n696 vss.n695 5.03414
R1237 vss.n836 vss.n835 5.03414
R1238 vss.n843 vss.n842 5.03414
R1239 vss.n861 vss.n860 5.03414
R1240 vss.n726 vss.n725 5.03414
R1241 vss.n114 vss.n113 5.03414
R1242 vss.n487 vss.n486 5.03414
R1243 vss.n355 vss.n354 5.03414
R1244 vss.n14 vss.n13 5.03414
R1245 vss.n588 vss.n587 5.03414
R1246 vss.n2 vss.n1 5.03414
R1247 vss.n472 vss.n471 5.03414
R1248 vss.n379 vss.n11 5.03414
R1249 vss.n330 vss.n329 5.03414
R1250 vss.n248 vss.n247 5.03414
R1251 vss.n370 vss.n369 5.03414
R1252 vss.n266 vss.n265 5.03414
R1253 vss.n352 vss.n351 5.03414
R1254 vss.n258 vss.n257 5.03414
R1255 vss.n500 vss.n481 5.03414
R1256 vss.n900 vss.n42 5.03414
R1257 vss.n482 vss.n155 5.03414
R1258 vss.n295 vss.n294 5.03414
R1259 vss.n269 vss.n33 5.03414
R1260 vss.n31 vss.n30 5.03414
R1261 vss.n286 vss.n284 5.03414
R1262 vss.n656 vss.n655 5.03414
R1263 vss.n897 vss.n45 5.03414
R1264 vss.n641 vss.n640 5.03414
R1265 vss.n894 vss.n49 5.03414
R1266 vss.n637 vss.n636 5.03414
R1267 vss.n668 vss.n667 5.03414
R1268 vss.n662 vss.n661 5.03414
R1269 vss.n682 vss.n681 5.03414
R1270 vss.n768 vss.n767 5.03414
R1271 vss.n760 vss.n759 5.03414
R1272 vss.n689 vss.n688 5.03414
R1273 vss.n738 vss.n737 5.03414
R1274 vss.n888 vss.n887 5.03414
R1275 vss.n745 vss.n744 5.03414
R1276 vss.n626 vss.n625 5.03414
R1277 vss.n828 vss.n827 5.03414
R1278 vss.n874 vss.n873 5.03414
R1279 vss.n62 vss.n61 5.03414
R1280 vss.n866 vss.n865 5.03414
R1281 vss.n790 vss.n107 5.03414
R1282 vss.n176 vss.n175 5.03414
R1283 vss.n507 vss.n218 5.03414
R1284 vss.n520 vss.n519 5.03414
R1285 vss.n443 vss.t23 4.7885
R1286 vss.n511 vss.t44 4.7885
R1287 vss.n225 vss.t143 4.7885
R1288 vss.n311 vss.t248 4.7885
R1289 vss.n323 vss.t250 4.7885
R1290 vss.n400 vss.t138 4.7885
R1291 vss.n422 vss.t334 4.7885
R1292 vss.n415 vss.t61 4.7885
R1293 vss.n430 vss.t125 4.7885
R1294 vss.n252 vss.t336 4.7885
R1295 vss.n451 vss.t70 4.7885
R1296 vss.n455 vss.t223 4.7885
R1297 vss.n532 vss.t163 4.7885
R1298 vss.n195 vss.t35 4.7885
R1299 vss.n522 vss.t320 4.7885
R1300 vss.n540 vss.t128 4.7885
R1301 vss.n605 vss.t136 4.7885
R1302 vss.n558 vss.t84 4.7885
R1303 vss.n569 vss.t165 4.7885
R1304 vss.n549 vss.t10 4.7885
R1305 vss.n598 vss.t156 4.7885
R1306 vss.n794 vss.t195 4.7885
R1307 vss.n815 vss.t318 4.7885
R1308 vss.n802 vss.t87 4.7885
R1309 vss.n552 vss.t20 4.7885
R1310 vss.n714 vss.t115 4.7885
R1311 vss.n706 vss.t140 4.7885
R1312 vss.n806 vss.t82 4.7885
R1313 vss.n722 vss.t18 4.7885
R1314 vss.n696 vss.t190 4.7885
R1315 vss.n836 vss.t237 4.7885
R1316 vss.n842 vss.t326 4.7885
R1317 vss.n852 vss.t330 4.7885
R1318 vss.n860 vss.t201 4.7885
R1319 vss.n725 vss.t74 4.7885
R1320 vss.n114 vss.t183 4.7885
R1321 vss.n486 vss.t154 4.7885
R1322 vss.n355 vss.t104 4.7885
R1323 vss.n179 vss.t122 4.7885
R1324 vss.n14 vss.t322 4.7885
R1325 vss.n587 vss.t147 4.7885
R1326 vss.n927 vss.t169 4.7885
R1327 vss.n2 vss.t63 4.7885
R1328 vss.n472 vss.t188 4.7885
R1329 vss.n379 vss.t98 4.7885
R1330 vss.n330 vss.t13 4.7885
R1331 vss.n247 vss.t15 4.7885
R1332 vss.n369 vss.t308 4.7885
R1333 vss.n265 vss.t32 4.7885
R1334 vss.n351 vss.t311 4.7885
R1335 vss.n257 vss.t235 4.7885
R1336 vss.n481 vss.t57 4.7885
R1337 vss.n614 vss.t244 4.7885
R1338 vss.n42 vss.t221 4.7885
R1339 vss.n482 vss.t52 4.7885
R1340 vss.n294 vss.t107 4.7885
R1341 vss.n269 vss.t50 4.7885
R1342 vss.n30 vss.t95 4.7885
R1343 vss.n284 vss.t117 4.7885
R1344 vss.n655 vss.t40 4.7885
R1345 vss.n647 vss.t175 4.7885
R1346 vss.n45 vss.t257 4.7885
R1347 vss.n641 vss.t47 4.7885
R1348 vss.n124 vss.t38 4.7885
R1349 vss.n49 vss.t4 4.7885
R1350 vss.n636 vss.t229 4.7885
R1351 vss.n667 vss.t254 4.7885
R1352 vss.n662 vss.t239 4.7885
R1353 vss.n681 vss.t241 4.7885
R1354 vss.n767 vss.t77 4.7885
R1355 vss.n760 vss.t66 4.7885
R1356 vss.n689 vss.t79 4.7885
R1357 vss.n737 vss.t131 4.7885
R1358 vss.n887 vss.t206 4.7885
R1359 vss.n744 vss.t186 4.7885
R1360 vss.n625 vss.t152 4.7885
R1361 vss.n828 vss.t283 4.7885
R1362 vss.n873 vss.t173 4.7885
R1363 vss.n61 vss.t277 4.7885
R1364 vss.n866 vss.t1 4.7885
R1365 vss.n107 vss.t158 4.7885
R1366 vss.n176 vss.t150 4.7885
R1367 vss.n218 vss.t145 4.7885
R1368 vss.n519 vss.t339 4.7885
R1369 vss.n414 vss.n413 4.28213
R1370 vss.n389 vss.n388 4.28213
R1371 vss.n903 vss.n39 4.28213
R1372 vss.n613 vss.n37 4.28213
R1373 vss.n648 vss.n46 4.28213
R1374 vss.n777 vss.n776 4.28213
R1375 vss.n853 vss.n851 4.28213
R1376 vss.n707 vss.n86 4.28213
R1377 vss.n817 vss.n816 4.28213
R1378 vss.n928 vss.n926 4.28213
R1379 vss.n445 vss.n444 4.28213
R1380 vss.n453 vss.n452 4.28213
R1381 vss.n196 vss.n190 4.28213
R1382 vss.n557 vss.n189 4.28213
R1383 vss.n403 dffrs_12.nand3_6.B 2.17818
R1384 vss.n839 vss.n79 2.06007
R1385 vss.n334 vss.n7 2.02164
R1386 vss.n918 vss.n917 2.02164
R1387 vss.n911 vss.n28 2.02164
R1388 vss.n652 vss.n150 2.02164
R1389 vss.n717 vss.n122 2.02164
R1390 vss.n797 vss.n99 2.02164
R1391 vss.n609 vss.n608 2.02164
R1392 vss.n535 vss.n19 2.02164
R1393 vss.n514 vss.n8 2.02164
R1394 vss.n397 vss.n396 2.02164
R1395 vss.n403 dffrs_12.nand3_1.A 1.34729
R1396 vss.n419 vss.n236 1.3005
R1397 vss.n422 vss.n421 1.3005
R1398 vss.n421 vss.n420 1.3005
R1399 vss.n416 vss.n415 1.3005
R1400 vss.n417 vss.n416 1.3005
R1401 vss.n307 vss.n238 1.3005
R1402 vss.n459 vss.n458 1.3005
R1403 vss.n455 vss.n437 1.3005
R1404 vss.n437 vss.n209 1.3005
R1405 vss.n204 vss.n192 1.3005
R1406 vss.n540 vss.n539 1.3005
R1407 vss.n539 vss.n538 1.3005
R1408 vss.n526 vss.n525 1.3005
R1409 vss.n522 vss.n205 1.3005
R1410 vss.n205 vss.n193 1.3005
R1411 vss.n544 vss.n185 1.3005
R1412 vss.n549 vss.n548 1.3005
R1413 vss.n548 vss.n547 1.3005
R1414 vss.n573 vss.n572 1.3005
R1415 vss.n569 vss.n186 1.3005
R1416 vss.n545 vss.n186 1.3005
R1417 vss.n564 vss.n563 1.3005
R1418 vss.n553 vss.n552 1.3005
R1419 vss.n553 vss.n97 1.3005
R1420 vss.n554 vss.n96 1.3005
R1421 vss.n802 vss.n801 1.3005
R1422 vss.n801 vss.n800 1.3005
R1423 vss.n703 vss.n92 1.3005
R1424 vss.n722 vss.n721 1.3005
R1425 vss.n721 vss.n720 1.3005
R1426 vss.n810 vss.n809 1.3005
R1427 vss.n806 vss.n93 1.3005
R1428 vss.n704 vss.n93 1.3005
R1429 vss.n729 vss.n728 1.3005
R1430 vss.n725 vss.n701 1.3005
R1431 vss.n701 vss.n78 1.3005
R1432 vss.n730 vss.n77 1.3005
R1433 vss.n860 vss.n859 1.3005
R1434 vss.n859 vss.n858 1.3005
R1435 vss.n784 vss.n783 1.3005
R1436 vss.n115 vss.n114 1.3005
R1437 vss.n782 vss.n115 1.3005
R1438 vss.n490 vss.n489 1.3005
R1439 vss.n486 vss.n485 1.3005
R1440 vss.n485 vss.n484 1.3005
R1441 vss.n585 vss.n584 1.3005
R1442 vss.n587 vss.n586 1.3005
R1443 vss.n586 vss.n17 1.3005
R1444 vss.n923 vss.n922 1.3005
R1445 vss.n15 vss.n14 1.3005
R1446 vss.n921 vss.n15 1.3005
R1447 vss.n383 vss.n382 1.3005
R1448 vss.n380 vss.n379 1.3005
R1449 vss.n380 vss.n5 1.3005
R1450 vss.n475 vss.n474 1.3005
R1451 vss.n473 vss.n472 1.3005
R1452 vss.n473 vss.n6 1.3005
R1453 vss.n935 vss.n934 1.3005
R1454 vss.n3 vss.n2 1.3005
R1455 vss.n933 vss.n3 1.3005
R1456 vss.n351 vss.n350 1.3005
R1457 vss.n350 vss.n349 1.3005
R1458 vss.n348 vss.n346 1.3005
R1459 vss.n339 vss.n338 1.3005
R1460 vss.n331 vss.n330 1.3005
R1461 vss.n337 vss.n331 1.3005
R1462 vss.n333 vss.n262 1.3005
R1463 vss.n369 vss.n368 1.3005
R1464 vss.n368 vss.n367 1.3005
R1465 vss.n365 vss.n364 1.3005
R1466 vss.n265 vss.n264 1.3005
R1467 vss.n264 vss.n21 1.3005
R1468 vss.n930 vss.n929 1.3005
R1469 vss.n927 vss.n9 1.3005
R1470 vss.n200 vss.n9 1.3005
R1471 vss.n481 vss.n480 1.3005
R1472 vss.n480 vss.n18 1.3005
R1473 vss.n479 vss.n478 1.3005
R1474 vss.n491 vss.n42 1.3005
R1475 vss.n492 vss.n491 1.3005
R1476 vss.n493 vss.n41 1.3005
R1477 vss.n483 vss.n482 1.3005
R1478 vss.n495 vss.n483 1.3005
R1479 vss.n497 vss.n496 1.3005
R1480 vss.n284 vss.n283 1.3005
R1481 vss.n283 vss.n282 1.3005
R1482 vss.n279 vss.n278 1.3005
R1483 vss.n118 vss.n49 1.3005
R1484 vss.n119 vss.n118 1.3005
R1485 vss.n117 vss.n48 1.3005
R1486 vss.n636 vss.n635 1.3005
R1487 vss.n635 vss.n120 1.3005
R1488 vss.n634 vss.n633 1.3005
R1489 vss.n663 vss.n662 1.3005
R1490 vss.n664 vss.n663 1.3005
R1491 vss.n149 vss.n141 1.3005
R1492 vss.n681 vss.n680 1.3005
R1493 vss.n680 vss.n679 1.3005
R1494 vss.n675 vss.n138 1.3005
R1495 vss.n767 vss.n766 1.3005
R1496 vss.n766 vss.n765 1.3005
R1497 vss.n133 vss.n131 1.3005
R1498 vss.n737 vss.n736 1.3005
R1499 vss.n736 vss.n735 1.3005
R1500 vss.n741 vss.n740 1.3005
R1501 vss.n744 vss.n743 1.3005
R1502 vss.n743 vss.n742 1.3005
R1503 vss.n750 vss.n749 1.3005
R1504 vss.n358 vss.n22 1.3005
R1505 vss.n357 vss.n355 1.3005
R1506 vss.n357 vss.n356 1.3005
R1507 vss.n273 vss.n272 1.3005
R1508 vss.n270 vss.n269 1.3005
R1509 vss.n271 vss.n270 1.3005
R1510 vss.n178 vss.n20 1.3005
R1511 vss.n180 vss.n179 1.3005
R1512 vss.n181 vss.n180 1.3005
R1513 vss.n291 vss.n25 1.3005
R1514 vss.n294 vss.n293 1.3005
R1515 vss.n293 vss.n26 1.3005
R1516 vss.n910 vss.n909 1.3005
R1517 vss.n30 vss.n29 1.3005
R1518 vss.n160 vss.n29 1.3005
R1519 vss.n161 vss.n148 1.3005
R1520 vss.n655 vss.n654 1.3005
R1521 vss.n654 vss.n653 1.3005
R1522 vss.n612 vss.n611 1.3005
R1523 vss.n615 vss.n614 1.3005
R1524 vss.n616 vss.n615 1.3005
R1525 vss.n619 vss.n44 1.3005
R1526 vss.n151 vss.n45 1.3005
R1527 vss.n152 vss.n151 1.3005
R1528 vss.n622 vss.n621 1.3005
R1529 vss.n625 vss.n624 1.3005
R1530 vss.n624 vss.n153 1.3005
R1531 vss.n618 vss.n154 1.3005
R1532 vss.n642 vss.n641 1.3005
R1533 vss.n643 vss.n642 1.3005
R1534 vss.n650 vss.n649 1.3005
R1535 vss.n647 vss.n646 1.3005
R1536 vss.n646 vss.n645 1.3005
R1537 vss.n671 vss.n670 1.3005
R1538 vss.n667 vss.n666 1.3005
R1539 vss.n666 vss.n665 1.3005
R1540 vss.n676 vss.n135 1.3005
R1541 vss.n690 vss.n689 1.3005
R1542 vss.n691 vss.n690 1.3005
R1543 vss.n756 vss.n755 1.3005
R1544 vss.n761 vss.n760 1.3005
R1545 vss.n762 vss.n761 1.3005
R1546 vss.n779 vss.n778 1.3005
R1547 vss.n124 vss.n123 1.3005
R1548 vss.n734 vss.n123 1.3005
R1549 vss.n751 vss.n54 1.3005
R1550 vss.n887 vss.n886 1.3005
R1551 vss.n886 vss.n885 1.3005
R1552 vss.n832 vss.n831 1.3005
R1553 vss.n829 vss.n828 1.3005
R1554 vss.n830 vss.n829 1.3005
R1555 vss.n881 vss.n880 1.3005
R1556 vss.n61 vss.n60 1.3005
R1557 vss.n60 vss.n59 1.3005
R1558 vss.n68 vss.n67 1.3005
R1559 vss.n873 vss.n872 1.3005
R1560 vss.n872 vss.n871 1.3005
R1561 vss.n855 vss.n854 1.3005
R1562 vss.n852 vss.n850 1.3005
R1563 vss.n850 vss.n849 1.3005
R1564 vss.n846 vss.n845 1.3005
R1565 vss.n842 vss.n841 1.3005
R1566 vss.n841 vss.n69 1.3005
R1567 vss.n867 vss.n866 1.3005
R1568 vss.n868 vss.n867 1.3005
R1569 vss.n840 vss.n70 1.3005
R1570 vss.n693 vss.n692 1.3005
R1571 vss.n697 vss.n696 1.3005
R1572 vss.n698 vss.n697 1.3005
R1573 vss.n699 vss.n80 1.3005
R1574 vss.n837 vss.n836 1.3005
R1575 vss.n838 vss.n837 1.3005
R1576 vss.n709 vss.n708 1.3005
R1577 vss.n706 vss.n705 1.3005
R1578 vss.n705 vss.n700 1.3005
R1579 vss.n711 vss.n710 1.3005
R1580 vss.n715 vss.n714 1.3005
R1581 vss.n716 vss.n715 1.3005
R1582 vss.n98 vss.n90 1.3005
R1583 vss.n815 vss.n814 1.3005
R1584 vss.n814 vss.n813 1.3005
R1585 vss.n107 vss.n106 1.3005
R1586 vss.n106 vss.n105 1.3005
R1587 vss.n104 vss.n103 1.3005
R1588 vss.n601 vss.n166 1.3005
R1589 vss.n600 vss.n598 1.3005
R1590 vss.n600 vss.n599 1.3005
R1591 vss.n163 vss.n100 1.3005
R1592 vss.n795 vss.n794 1.3005
R1593 vss.n796 vss.n795 1.3005
R1594 vss.n556 vss.n555 1.3005
R1595 vss.n559 vss.n558 1.3005
R1596 vss.n560 vss.n559 1.3005
R1597 vss.n579 vss.n578 1.3005
R1598 vss.n177 vss.n176 1.3005
R1599 vss.n577 vss.n177 1.3005
R1600 vss.n183 vss.n168 1.3005
R1601 vss.n606 vss.n605 1.3005
R1602 vss.n607 vss.n606 1.3005
R1603 vss.n198 vss.n197 1.3005
R1604 vss.n195 vss.n194 1.3005
R1605 vss.n194 vss.n184 1.3005
R1606 vss.n531 vss.n530 1.3005
R1607 vss.n533 vss.n532 1.3005
R1608 vss.n534 vss.n533 1.3005
R1609 vss.n449 vss.n210 1.3005
R1610 vss.n451 vss.n450 1.3005
R1611 vss.n450 vss.n203 1.3005
R1612 vss.n218 vss.n217 1.3005
R1613 vss.n217 vss.n202 1.3005
R1614 vss.n216 vss.n215 1.3005
R1615 vss.n315 vss.n314 1.3005
R1616 vss.n311 vss.n309 1.3005
R1617 vss.n309 vss.n308 1.3005
R1618 vss.n244 vss.n243 1.3005
R1619 vss.n400 vss.n399 1.3005
R1620 vss.n399 vss.n398 1.3005
R1621 vss.n318 vss.n303 1.3005
R1622 vss.n323 vss.n322 1.3005
R1623 vss.n322 vss.n321 1.3005
R1624 vss.n395 vss.n394 1.3005
R1625 vss.n247 vss.n246 1.3005
R1626 vss.n254 vss.n246 1.3005
R1627 vss.n377 vss.n376 1.3005
R1628 vss.n257 vss.n256 1.3005
R1629 vss.n256 vss.n255 1.3005
R1630 vss.n387 vss.n229 1.3005
R1631 vss.n386 vss.n252 1.3005
R1632 vss.n386 vss.n385 1.3005
R1633 vss.n305 vss.n230 1.3005
R1634 vss.n431 vss.n430 1.3005
R1635 vss.n432 vss.n431 1.3005
R1636 vss.n466 vss.n465 1.3005
R1637 vss.n226 vss.n225 1.3005
R1638 vss.n464 vss.n226 1.3005
R1639 vss.n435 vss.n211 1.3005
R1640 vss.n512 vss.n511 1.3005
R1641 vss.n513 vss.n512 1.3005
R1642 vss.n441 vss.n440 1.3005
R1643 vss.n443 vss.n442 1.3005
R1644 vss.n442 vss.n436 1.3005
R1645 vss.n519 vss.n518 1.3005
R1646 vss.n518 vss.n517 1.3005
R1647 vss.n460 vss.n208 1.3005
R1648 vss.n510 vss.n212 0.92075
R1649 vss.n467 vss.n224 0.92075
R1650 vss.n324 vss.n302 0.92075
R1651 vss.n407 vss.n406 0.92075
R1652 vss.n423 vss.n235 0.92075
R1653 vss.n429 vss.n231 0.92075
R1654 vss.n457 vss.n456 0.92075
R1655 vss.n199 vss.n174 0.92075
R1656 vss.n524 vss.n523 0.92075
R1657 vss.n541 vss.n191 0.92075
R1658 vss.n604 vss.n169 0.92075
R1659 vss.n571 vss.n570 0.92075
R1660 vss.n550 vss.n543 0.92075
R1661 vss.n793 vss.n101 0.92075
R1662 vss.n803 vss.n95 0.92075
R1663 vss.n565 vss.n551 0.92075
R1664 vss.n713 vss.n712 0.92075
R1665 vss.n808 vss.n807 0.92075
R1666 vss.n723 vss.n702 0.92075
R1667 vss.n835 vss.n81 0.92075
R1668 vss.n844 vss.n843 0.92075
R1669 vss.n861 vss.n76 0.92075
R1670 vss.n727 vss.n726 0.92075
R1671 vss.n785 vss.n113 0.92075
R1672 vss.n488 vss.n487 0.92075
R1673 vss.n924 vss.n13 0.92075
R1674 vss.n588 vss.n583 0.92075
R1675 vss.n936 vss.n1 0.92075
R1676 vss.n476 vss.n471 0.92075
R1677 vss.n381 vss.n11 0.92075
R1678 vss.n393 vss.n248 0.92075
R1679 vss.n363 vss.n266 0.92075
R1680 vss.n352 vss.n345 0.92075
R1681 vss.n371 vss.n370 0.92075
R1682 vss.n375 vss.n258 0.92075
R1683 vss.n340 vss.n329 0.92075
R1684 vss.n501 vss.n500 0.92075
R1685 vss.n901 vss.n900 0.92075
R1686 vss.n498 vss.n155 0.92075
R1687 vss.n296 vss.n295 0.92075
R1688 vss.n274 vss.n33 0.92075
R1689 vss.n908 vss.n31 0.92075
R1690 vss.n287 vss.n286 0.92075
R1691 vss.n656 vss.n147 0.92075
R1692 vss.n898 vss.n897 0.92075
R1693 vss.n640 vss.n632 0.92075
R1694 vss.n895 vss.n894 0.92075
R1695 vss.n638 vss.n637 0.92075
R1696 vss.n669 vss.n668 0.92075
R1697 vss.n661 vss.n142 0.92075
R1698 vss.n682 vss.n137 0.92075
R1699 vss.n769 vss.n768 0.92075
R1700 vss.n759 vss.n757 0.92075
R1701 vss.n688 vss.n687 0.92075
R1702 vss.n739 vss.n738 0.92075
R1703 vss.n889 vss.n888 0.92075
R1704 vss.n748 vss.n745 0.92075
R1705 vss.n627 vss.n626 0.92075
R1706 vss.n359 vss.n354 0.92075
R1707 vss.n874 vss.n66 0.92075
R1708 vss.n879 vss.n62 0.92075
R1709 vss.n833 vss.n827 0.92075
R1710 vss.n865 vss.n71 0.92075
R1711 vss.n695 vss.n694 0.92075
R1712 vss.n791 vss.n790 0.92075
R1713 vss.n602 vss.n597 0.92075
R1714 vss.n580 vss.n175 0.92075
R1715 vss.n508 vss.n507 0.92075
R1716 vss.n313 vss.n312 0.92075
R1717 vss.n520 vss.n207 0.92075
R1718 dffrs_12.d dffrs_12.nand3_8.A 0.784786
R1719 dffrs_13.d dffrs_13.nand3_8.A 0.784786
R1720 vss.n746 vss.n52 0.779467
R1721 dffrs_12.clk vss.n403 0.611214
R1722 vss.n327 vss.n300 0.52742
R1723 vss.n327 vss.n326 0.195855
R1724 vss.n892 vss.n51 0.143322
R1725 vss.n326 vss.n249 0.140365
R1726 vss.n240 vss.n239 0.122607
R1727 vss.n470 vss.n469 0.122607
R1728 vss.n392 vss.n249 0.118169
R1729 vss.n863 vss.n74 0.115241
R1730 vss.n774 vss.n125 0.10457
R1731 vss.n876 vss.n64 0.10457
R1732 vss.n110 dffrs_14.vss 0.102612
R1733 dffrs_7.vss vss.n109 0.102537
R1734 dffrs_8.vss vss.n630 0.102537
R1735 vss.n590 dffrs_9.vss 0.102537
R1736 vss.n503 dffrs_10.vss 0.102537
R1737 vss.n404 vss.n234 0.078611
R1738 vss.n392 vss.n391 0.0781858
R1739 vss.n426 vss.n425 0.0660086
R1740 vss.n425 vss.n0 0.0655096
R1741 vss.n412 vss.n232 0.0645882
R1742 vss.n439 vss.n438 0.0645882
R1743 vss.n823 vss.n82 0.0625376
R1744 vss.n469 vss.n222 0.0622481
R1745 vss.n410 vss.n239 0.0622481
R1746 vss.n373 vss.n260 0.0616538
R1747 vss.n285 vss.n143 0.0616538
R1748 vss.n292 vss.n32 0.0616538
R1749 vss.n361 vss.n353 0.0616538
R1750 vss.n112 vss.n111 0.0616538
R1751 vss.n623 vss.n102 0.0616538
R1752 vss.n219 vss.n213 0.0616538
R1753 vss.n589 vss.n582 0.0616538
R1754 vss.n594 vss.n156 0.0616538
R1755 vss.n684 vss.n683 0.0615256
R1756 vss.n326 vss.n242 0.0551896
R1757 vss.n774 vss.n51 0.054837
R1758 vss.n74 vss.n64 0.054837
R1759 vss.n771 vss.n129 0.0478906
R1760 vss.n343 vss.n342 0.0478478
R1761 vss.n328 vss.n327 0.0478478
R1762 vss.n277 vss.n145 0.0478478
R1763 vss.n110 vss.n83 0.0478478
R1764 vss.n290 vss.n289 0.0478478
R1765 vss.n299 vss.n298 0.0478478
R1766 vss.n630 vss.n629 0.0478478
R1767 vss.n746 vss.n63 0.0478478
R1768 vss.n787 vss.n109 0.0478478
R1769 vss.n504 vss.n503 0.0478478
R1770 vss.n591 vss.n590 0.0478478
R1771 vss.n130 vss.n125 0.0466843
R1772 vss.n877 vss.n876 0.0466843
R1773 vss.n325 vss.n300 0.0465106
R1774 vss.n405 vss.n242 0.0465106
R1775 vss.n424 vss.n234 0.0465106
R1776 vss.n896 vss.n47 0.0465022
R1777 vss.n899 vss.n43 0.0465022
R1778 vss.n902 vss.n40 0.0465022
R1779 vss.n925 vss.n12 0.0465022
R1780 vss.n893 vss.n892 0.0464521
R1781 vss.n411 vss.n410 0.0415307
R1782 vss.n446 vss.n222 0.0415307
R1783 vss.n758 vss.n128 0.0405109
R1784 vss.n770 vss.n130 0.0405109
R1785 vss.n878 vss.n877 0.0405109
R1786 vss.n875 vss.n65 0.0405109
R1787 vss.n310 vss.n241 0.0405109
R1788 vss.n468 vss.n223 0.0405109
R1789 vss.n391 vss.n390 0.040346
R1790 vss.n863 vss.n75 0.0368083
R1791 vss.n724 vss.n73 0.036505
R1792 vss.n94 vss.n89 0.036505
R1793 vss.n454 vss.n206 0.036505
R1794 vss.n542 vss.n188 0.036505
R1795 vss.n567 vss.n566 0.036505
R1796 vss.n373 vss.n259 0.0361576
R1797 vss.n250 vss.n249 0.0361576
R1798 vss.n361 vss.n268 0.0361576
R1799 vss.n660 vss.n143 0.0361576
R1800 vss.n684 vss.n127 0.0361576
R1801 vss.n34 vss.n32 0.0361576
R1802 vss.n826 vss.n823 0.0361576
R1803 vss.n111 vss.n84 0.0361576
R1804 vss.n789 vss.n102 0.0361576
R1805 vss.n596 vss.n594 0.0361576
R1806 vss.n506 vss.n213 0.0361576
R1807 vss.n582 vss.n171 0.0361576
R1808 vss.n413 vss.n411 0.0349747
R1809 vss.n446 vss.n445 0.0349747
R1810 vss.n834 vss.n823 0.0340549
R1811 vss.n390 vss.n389 0.0339793
R1812 vss.n342 vss.n260 0.0335769
R1813 vss.n373 vss.n372 0.0335769
R1814 vss.n683 vss.n129 0.0335769
R1815 vss.n285 vss.n277 0.0335769
R1816 vss.n657 vss.n143 0.0335769
R1817 vss.n292 vss.n290 0.0335769
R1818 vss.n907 vss.n32 0.0335769
R1819 vss.n353 vss.n299 0.0335769
R1820 vss.n361 vss.n360 0.0335769
R1821 vss.n111 vss.n85 0.0335769
R1822 vss.n792 vss.n102 0.0335769
R1823 vss.n509 vss.n213 0.0335769
R1824 vss.n582 vss.n581 0.0335769
R1825 vss.n603 vss.n594 0.0335769
R1826 vss.n686 vss.n685 0.0334487
R1827 vss.n592 vss.n170 0.0322085
R1828 vss.n788 vss.n88 0.0322085
R1829 vss.n391 vss.n251 0.0322085
R1830 vss.n343 vss.n267 0.0322085
R1831 vss.n267 vss.n261 0.0322085
R1832 vss.n328 vss.n251 0.0322085
R1833 vss.n276 vss.n38 0.0322085
R1834 vss.n298 vss.n276 0.0322085
R1835 vss.n659 vss.n145 0.0322085
R1836 vss.n659 vss.n658 0.0322085
R1837 vss.n772 vss.n771 0.0322085
R1838 vss.n773 vss.n772 0.0322085
R1839 vss.n821 vss.n83 0.0322085
R1840 vss.n289 vss.n35 0.0322085
R1841 vss.n906 vss.n35 0.0322085
R1842 vss.n629 vss.n159 0.0322085
R1843 vss.n825 vss.n824 0.0322085
R1844 vss.n825 vss.n63 0.0322085
R1845 vss.n788 vss.n787 0.0322085
R1846 vss.n821 vss.n820 0.0322085
R1847 vss.n505 vss.n504 0.0322085
R1848 vss.n409 vss.n240 0.0322085
R1849 vss.n410 vss.n409 0.0322085
R1850 vss.n470 vss.n221 0.0322085
R1851 vss.n222 vss.n221 0.0322085
R1852 vss.n505 vss.n214 0.0322085
R1853 vss.n592 vss.n591 0.0322085
R1854 vss.n595 vss.n159 0.0322085
R1855 vss.n326 vss.n325 0.0308765
R1856 vss.n344 vss.n299 0.0268641
R1857 vss.n362 vss.n361 0.0268641
R1858 vss.n374 vss.n373 0.0268641
R1859 vss.n342 vss.n341 0.0268641
R1860 vss.n275 vss.n32 0.0268641
R1861 vss.n144 vss.n129 0.0268641
R1862 vss.n685 vss.n136 0.0268641
R1863 vss.n747 vss.n746 0.0268641
R1864 vss.n146 vss.n143 0.0268641
R1865 vss.n288 vss.n277 0.0268641
R1866 vss.n297 vss.n290 0.0268641
R1867 vss.n628 vss.n109 0.0268641
R1868 vss.n823 vss.n822 0.0268641
R1869 vss.n111 vss.n108 0.0268641
R1870 vss.n786 vss.n110 0.0268641
R1871 vss.n158 vss.n102 0.0268641
R1872 vss.n582 vss.n173 0.0268641
R1873 vss.n590 vss.n172 0.0268641
R1874 vss.n301 vss.n300 0.0268641
R1875 vss.n408 vss.n242 0.0268641
R1876 vss.n220 vss.n213 0.0268641
R1877 vss.n503 vss.n477 0.0268641
R1878 vss.n594 vss.n593 0.0268641
R1879 vss.n630 vss.n157 0.0268641
R1880 vss.n892 vss.n52 0.0263346
R1881 vss.n824 vss.n64 0.0237454
R1882 vss.n774 vss.n773 0.0235512
R1883 vss.n658 vss.n36 0.0235512
R1884 vss.n906 vss.n905 0.0235512
R1885 vss.n904 vss.n38 0.0235512
R1886 vss.n820 vss.n819 0.0235512
R1887 vss.n818 vss.n88 0.0235512
R1888 vss.n261 vss.n10 0.0235512
R1889 vss.n448 vss.n214 0.0235512
R1890 vss.n447 vss.n170 0.0235512
R1891 vss.n595 vss.n87 0.0235512
R1892 vss.n834 vss.n824 0.0226532
R1893 vss.n411 vss.n234 0.0225109
R1894 vss.n775 vss.n36 0.0225109
R1895 vss.n905 vss.n36 0.0225109
R1896 vss.n905 vss.n904 0.0225109
R1897 vss.n904 vss.n10 0.0225109
R1898 vss.n819 vss.n64 0.0225109
R1899 vss.n819 vss.n818 0.0225109
R1900 vss.n818 vss.n87 0.0225109
R1901 vss.n390 vss.n10 0.0225109
R1902 vss.n448 vss.n446 0.0225109
R1903 vss.n447 vss.n87 0.0225109
R1904 vss.n448 vss.n447 0.0225109
R1905 vss.n567 vss.n188 0.0223682
R1906 vss.n206 vss.n188 0.0223682
R1907 vss.n426 vss.n232 0.0223682
R1908 vss.n567 vss.n94 0.0223682
R1909 vss.n94 vss.n73 0.0223682
R1910 vss.n863 vss.n73 0.0223682
R1911 vss.n438 vss.n206 0.0223682
R1912 vss.n372 vss.n261 0.0223376
R1913 vss.n658 vss.n657 0.0223376
R1914 vss.n907 vss.n906 0.0223376
R1915 vss.n360 vss.n38 0.0223376
R1916 vss.n820 vss.n85 0.0223376
R1917 vss.n792 vss.n88 0.0223376
R1918 vss.n509 vss.n214 0.0223376
R1919 vss.n581 vss.n170 0.0223376
R1920 vss.n603 vss.n595 0.0223376
R1921 vss.n773 vss.n126 0.0222094
R1922 vss.n344 vss.n343 0.0214837
R1923 vss.n362 vss.n267 0.0214837
R1924 vss.n374 vss.n251 0.0214837
R1925 vss.n341 vss.n328 0.0214837
R1926 vss.n276 vss.n275 0.0214837
R1927 vss.n145 vss.n144 0.0214837
R1928 vss.n659 vss.n136 0.0214837
R1929 vss.n772 vss.n128 0.0214837
R1930 vss.n771 vss.n770 0.0214837
R1931 vss.n747 vss.n83 0.0214837
R1932 vss.n146 vss.n35 0.0214837
R1933 vss.n289 vss.n288 0.0214837
R1934 vss.n298 vss.n297 0.0214837
R1935 vss.n629 vss.n628 0.0214837
R1936 vss.n878 vss.n63 0.0214837
R1937 vss.n825 vss.n65 0.0214837
R1938 vss.n822 vss.n821 0.0214837
R1939 vss.n788 vss.n108 0.0214837
R1940 vss.n787 vss.n786 0.0214837
R1941 vss.n159 vss.n158 0.0214837
R1942 vss.n505 vss.n173 0.0214837
R1943 vss.n504 vss.n172 0.0214837
R1944 vss.n301 vss.n240 0.0214837
R1945 vss.n409 vss.n408 0.0214837
R1946 vss.n221 vss.n220 0.0214837
R1947 vss.n477 vss.n470 0.0214837
R1948 vss.n593 vss.n592 0.0214837
R1949 vss.n591 vss.n157 0.0214837
R1950 vss.n425 vss.n424 0.0204141
R1951 vss.n851 vss.n64 0.0200312
R1952 vss.n863 vss.n862 0.0199048
R1953 vss.n46 vss.n36 0.019868
R1954 vss.n905 vss.n37 0.019868
R1955 vss.n904 vss.n903 0.019868
R1956 vss.n819 vss.n86 0.019868
R1957 vss.n818 vss.n817 0.019868
R1958 vss.n926 vss.n10 0.019868
R1959 vss.n453 vss.n448 0.019868
R1960 vss.n447 vss.n190 0.019868
R1961 vss.n189 vss.n87 0.019868
R1962 vss.n776 vss.n775 0.0197929
R1963 vss.n805 vss.n73 0.0197428
R1964 vss.n804 vss.n94 0.0197428
R1965 vss.n521 vss.n206 0.0197428
R1966 vss.n188 vss.n187 0.0197428
R1967 vss.n568 vss.n567 0.0197428
R1968 vss.n937 vss.n0 0.0164817
R1969 vss.n12 vss.n0 0.0157888
R1970 vss.n40 vss.n12 0.0157888
R1971 vss.n43 vss.n40 0.0157888
R1972 vss.n47 vss.n43 0.0157888
R1973 vss.n891 vss.n47 0.0157888
R1974 vss.n425 vss.n233 0.0150091
R1975 vss.n746 vss.n82 0.0142428
R1976 vss.n112 vss.n110 0.014047
R1977 vss.n623 vss.n109 0.014047
R1978 vss.n503 vss.n219 0.014047
R1979 vss.n590 vss.n589 0.014047
R1980 vss.n630 vss.n156 0.014047
R1981 vss.n267 vss.n259 0.0121902
R1982 vss.n251 vss.n250 0.0121902
R1983 vss.n276 vss.n268 0.0121902
R1984 vss.n660 vss.n659 0.0121902
R1985 vss.n772 vss.n127 0.0121902
R1986 vss.n35 vss.n34 0.0121902
R1987 vss.n826 vss.n825 0.0121902
R1988 vss.n821 vss.n84 0.0121902
R1989 vss.n789 vss.n788 0.0121902
R1990 vss.n596 vss.n159 0.0121902
R1991 vss.n506 vss.n505 0.0121902
R1992 vss.n409 vss.n241 0.0121902
R1993 vss.n223 vss.n221 0.0121902
R1994 vss.n592 vss.n171 0.0121902
R1995 vss.n864 vss.n863 0.0102582
R1996 vss.n639 vss.n47 0.00974555
R1997 vss.n631 vss.n43 0.00974555
R1998 vss.n499 vss.n40 0.00974555
R1999 vss.n502 vss.n12 0.00974555
R2000 vss.n891 vss.n890 0.00967038
R2001 vss.n310 vss.n239 0.00915761
R2002 vss.n469 vss.n468 0.00915761
R2003 vss.n405 vss.n404 0.00745509
R2004 dffrs_11.vss vss.n937 0.00734312
R2005 vss.n758 vss.n125 0.00720109
R2006 vss.n876 vss.n875 0.00720109
R2007 vss.n428 vss.n426 0.00638507
R2008 vss.n639 dffrs_7.vss 0.0044588
R2009 vss.n631 dffrs_8.vss 0.0044588
R2010 vss.n499 dffrs_9.vss 0.0044588
R2011 dffrs_10.vss vss.n502 0.0044588
R2012 vss.n568 vss 0.0044588
R2013 dffrs_14.vss vss.n53 0.00438363
R2014 vss.n685 vss.n684 0.000628205
R2015 vss.n686 vss.n126 0.000628205
R2016 vss.n775 vss.n774 0.000575167
R2017 vss.n893 vss.n50 0.000575167
R2018 vss.n890 vss.n53 0.000575167
R2019 vss.n892 vss.n891 0.000550111
R2020 vss.n413 vss.n412 0.000544599
R2021 vss.n445 vss.n439 0.000544599
R2022 vss.n389 vss.n233 0.000543311
R2023 vss.n851 vss.n75 0.000525267
R2024 vss.n776 vss.n50 0.000525056
R2025 vss.n896 vss.n46 0.000525056
R2026 vss.n899 vss.n37 0.000525056
R2027 vss.n903 vss.n902 0.000525056
R2028 vss.n724 vss.n86 0.000525056
R2029 vss.n817 vss.n89 0.000525056
R2030 vss.n926 vss.n925 0.000525056
R2031 vss.n454 vss.n453 0.000525056
R2032 vss.n542 vss.n190 0.000525056
R2033 vss.n566 vss.n189 0.000525056
R2034 dffrs_13.nand3_8.Z.n0 dffrs_13.nand3_8.Z.t5 41.0041
R2035 dffrs_13.nand3_8.Z.n1 dffrs_13.nand3_8.Z.t6 40.8177
R2036 dffrs_13.nand3_8.Z.n1 dffrs_13.nand3_8.Z.t4 27.1302
R2037 dffrs_13.nand3_8.Z.n0 dffrs_13.nand3_8.Z.t7 26.9438
R2038 dffrs_13.nand3_6.A dffrs_13.nand3_0.B 17.0041
R2039 dffrs_13.nand3_8.Z dffrs_13.nand3_8.Z.n2 14.8493
R2040 dffrs_13.nand3_8.Z.n5 dffrs_13.nand3_8.Z.t3 10.0473
R2041 dffrs_13.nand3_8.Z.n4 dffrs_13.nand3_8.Z.t2 6.51042
R2042 dffrs_13.nand3_8.Z.n4 dffrs_13.nand3_8.Z.n3 6.04952
R2043 dffrs_13.nand3_8.Z.n2 dffrs_13.nand3_8.Z.n0 5.7305
R2044 dffrs_13.nand3_0.B dffrs_13.nand3_8.Z.n1 5.47979
R2045 dffrs_13.nand3_8.Z dffrs_13.nand3_8.Z.n5 4.72925
R2046 dffrs_13.nand3_8.Z.n5 dffrs_13.nand3_8.Z.n4 0.732092
R2047 dffrs_13.nand3_8.Z.n3 dffrs_13.nand3_8.Z.t1 0.7285
R2048 dffrs_13.nand3_8.Z.n3 dffrs_13.nand3_8.Z.t0 0.7285
R2049 dffrs_13.nand3_8.Z.n2 dffrs_13.nand3_6.A 0.0455
R2050 vdd.t225 vdd.n482 250.9
R2051 vdd.n483 vdd.t149 250.9
R2052 vdd.t6 vdd.n367 250.9
R2053 vdd.n368 vdd.t70 250.9
R2054 vdd.t261 vdd.n299 250.9
R2055 vdd.n300 vdd.t167 250.9
R2056 vdd.t323 vdd.n231 250.9
R2057 vdd.n232 vdd.t179 250.9
R2058 vdd.t467 vdd.n163 250.9
R2059 vdd.n164 vdd.t463 250.9
R2060 vdd.t197 vdd.n95 250.9
R2061 vdd.n96 vdd.t501 250.9
R2062 vdd.t371 vdd.n400 250.9
R2063 vdd.n401 vdd.t82 250.9
R2064 vdd.t207 vdd.n394 250.9
R2065 vdd.n395 vdd.t147 250.9
R2066 vdd.t349 vdd.n332 250.9
R2067 vdd.n333 vdd.t361 250.9
R2068 vdd.t40 vdd.n326 250.9
R2069 vdd.n327 vdd.t68 250.9
R2070 vdd.t513 vdd.n264 250.9
R2071 vdd.n265 vdd.t44 250.9
R2072 vdd.t32 vdd.n258 250.9
R2073 vdd.n259 vdd.t205 250.9
R2074 vdd.t295 vdd.n196 250.9
R2075 vdd.n197 vdd.t62 250.9
R2076 vdd.t34 vdd.n190 250.9
R2077 vdd.n191 vdd.t177 250.9
R2078 vdd.t511 vdd.n128 250.9
R2079 vdd.n129 vdd.t36 250.9
R2080 vdd.t341 vdd.n122 250.9
R2081 vdd.n123 vdd.t329 250.9
R2082 vdd.t76 vdd.n60 250.9
R2083 vdd.n61 vdd.t343 250.9
R2084 vdd.t2 vdd.n54 250.9
R2085 vdd.n55 vdd.t12 250.9
R2086 vdd.t327 vdd.n477 250.9
R2087 vdd.n478 vdd.t223 250.9
R2088 vdd.t391 vdd.n379 250.9
R2089 vdd.n380 vdd.t42 250.9
R2090 vdd.t48 vdd.n362 250.9
R2091 vdd.n363 vdd.t461 250.9
R2092 vdd.t433 vdd.n311 250.9
R2093 vdd.n312 vdd.t369 250.9
R2094 vdd.t267 vdd.n294 250.9
R2095 vdd.n295 vdd.t259 250.9
R2096 vdd.t379 vdd.n243 250.9
R2097 vdd.n244 vdd.t239 250.9
R2098 vdd.t129 vdd.n226 250.9
R2099 vdd.n227 vdd.t319 250.9
R2100 vdd.t429 vdd.n175 250.9
R2101 vdd.n176 vdd.t515 250.9
R2102 vdd.t281 vdd.n158 250.9
R2103 vdd.n159 vdd.t469 250.9
R2104 vdd.t447 vdd.n107 250.9
R2105 vdd.n108 vdd.t245 250.9
R2106 vdd.t273 vdd.n90 250.9
R2107 vdd.n91 vdd.t199 250.9
R2108 vdd.t413 vdd.n39 250.9
R2109 vdd.n40 vdd.t507 250.9
R2110 vdd.t337 vdd.n405 250.9
R2111 vdd.n406 vdd.t301 250.9
R2112 vdd.t26 vdd.n337 250.9
R2113 vdd.n338 vdd.t331 250.9
R2114 vdd.t333 vdd.n269 250.9
R2115 vdd.n270 vdd.t60 250.9
R2116 vdd.t335 vdd.n201 250.9
R2117 vdd.n202 vdd.t74 250.9
R2118 vdd.t339 vdd.n133 250.9
R2119 vdd.n134 vdd.t155 250.9
R2120 vdd.t28 vdd.n65 250.9
R2121 vdd.n66 vdd.t473 250.9
R2122 vdd.t141 vdd.n472 250.9
R2123 vdd.n473 vdd.t91 250.9
R2124 vdd.t171 vdd.n410 250.9
R2125 vdd.n411 vdd.t345 250.9
R2126 vdd.t457 vdd.n357 250.9
R2127 vdd.n358 vdd.t97 250.9
R2128 vdd.t347 vdd.n389 250.9
R2129 vdd.n390 vdd.t85 250.9
R2130 vdd.t481 vdd.n342 250.9
R2131 vdd.n343 vdd.t201 250.9
R2132 vdd.t8 vdd.n289 250.9
R2133 vdd.n290 vdd.t115 250.9
R2134 vdd.t203 vdd.n321 250.9
R2135 vdd.n322 vdd.t103 250.9
R2136 vdd.t165 vdd.n274 250.9
R2137 vdd.n275 vdd.t287 250.9
R2138 vdd.t50 vdd.n221 250.9
R2139 vdd.n222 vdd.t112 250.9
R2140 vdd.t181 vdd.n253 250.9
R2141 vdd.n254 vdd.t106 250.9
R2142 vdd.t163 vdd.n206 250.9
R2143 vdd.n207 vdd.t227 250.9
R2144 vdd.t217 vdd.n153 250.9
R2145 vdd.n154 vdd.t124 250.9
R2146 vdd.t465 vdd.n185 250.9
R2147 vdd.n186 vdd.t109 250.9
R2148 vdd.t191 vdd.n138 250.9
R2149 vdd.n139 vdd.t243 250.9
R2150 vdd.t317 vdd.n85 250.9
R2151 vdd.n86 vdd.t88 250.9
R2152 vdd.t14 vdd.n117 250.9
R2153 vdd.n118 vdd.t121 250.9
R2154 vdd.t175 vdd.n70 250.9
R2155 vdd.n71 vdd.t56 250.9
R2156 vdd.t353 vdd.n49 250.9
R2157 vdd.n50 vdd.t127 250.9
R2158 vdd.t365 vdd.n467 250.9
R2159 vdd.n468 vdd.t139 250.9
R2160 vdd.t411 vdd.n384 250.9
R2161 vdd.n385 vdd.t235 250.9
R2162 vdd.t251 vdd.n352 250.9
R2163 vdd.n353 vdd.t459 250.9
R2164 vdd.t435 vdd.n316 250.9
R2165 vdd.n317 vdd.t475 250.9
R2166 vdd.t277 vdd.n284 250.9
R2167 vdd.n285 vdd.t4 250.9
R2168 vdd.t381 vdd.n248 250.9
R2169 vdd.n249 vdd.t297 250.9
R2170 vdd.t289 vdd.n216 250.9
R2171 vdd.n217 vdd.t24 250.9
R2172 vdd.t385 vdd.n180 250.9
R2173 vdd.n181 vdd.t38 250.9
R2174 vdd.t357 vdd.n148 250.9
R2175 vdd.n149 vdd.t219 250.9
R2176 vdd.t399 vdd.n112 250.9
R2177 vdd.n113 vdd.t133 250.9
R2178 vdd.t283 vdd.n80 250.9
R2179 vdd.n81 vdd.t315 250.9
R2180 vdd.t405 vdd.n44 250.9
R2181 vdd.n45 vdd.t20 250.9
R2182 vdd.t151 vdd.n415 250.9
R2183 vdd.n416 vdd.t189 250.9
R2184 vdd.t233 vdd.n347 250.9
R2185 vdd.n348 vdd.t183 250.9
R2186 vdd.t477 vdd.n279 250.9
R2187 vdd.n280 vdd.t54 250.9
R2188 vdd.t299 vdd.n211 250.9
R2189 vdd.n212 vdd.t249 250.9
R2190 vdd.t229 vdd.n143 250.9
R2191 vdd.n144 vdd.t363 250.9
R2192 vdd.t135 vdd.n75 250.9
R2193 vdd.n76 vdd.t143 250.9
R2194 vdd.t491 vdd.n420 250.9
R2195 vdd.n421 vdd.t439 250.9
R2196 vdd.t193 vdd.n436 250.9
R2197 vdd.n437 vdd.t263 250.9
R2198 vdd.t145 vdd.n431 250.9
R2199 vdd.n432 vdd.t443 250.9
R2200 vdd.t257 vdd.n454 250.9
R2201 vdd.n455 vdd.t493 250.9
R2202 vdd.t94 vdd.n460 250.9
R2203 vdd.n461 vdd.t497 250.9
R2204 vdd.t311 vdd.n448 250.9
R2205 vdd.n449 vdd.t30 250.9
R2206 vdd.t64 vdd.n25 250.9
R2207 vdd.n26 vdd.t505 250.9
R2208 vdd.t415 vdd.n19 250.9
R2209 vdd.n20 vdd.t78 250.9
R2210 vdd.t309 vdd.n32 250.9
R2211 vdd.n33 vdd.t211 250.9
R2212 vdd.t503 vdd.n2 250.9
R2213 vdd.n3 vdd.t351 250.9
R2214 vdd.t305 vdd.n13 250.9
R2215 vdd.n14 vdd.t231 250.9
R2216 vdd.t269 vdd.n8 250.9
R2217 vdd.n9 vdd.t355 250.9
R2218 vdd.t325 vdd.t225 200
R2219 vdd.t149 vdd.t325 200
R2220 vdd.t46 vdd.t6 200
R2221 vdd.t70 vdd.t46 200
R2222 vdd.t265 vdd.t261 200
R2223 vdd.t167 vdd.t265 200
R2224 vdd.t131 vdd.t323 200
R2225 vdd.t179 vdd.t131 200
R2226 vdd.t279 vdd.t467 200
R2227 vdd.t463 vdd.t279 200
R2228 vdd.t271 vdd.t197 200
R2229 vdd.t501 vdd.t271 200
R2230 vdd.t401 vdd.t371 200
R2231 vdd.t82 vdd.t401 200
R2232 vdd.t221 vdd.t207 200
R2233 vdd.t147 vdd.t221 200
R2234 vdd.t377 vdd.t349 200
R2235 vdd.t361 vdd.t377 200
R2236 vdd.t455 vdd.t40 200
R2237 vdd.t68 vdd.t455 200
R2238 vdd.t407 vdd.t513 200
R2239 vdd.t44 vdd.t407 200
R2240 vdd.t237 vdd.t32 200
R2241 vdd.t205 vdd.t237 200
R2242 vdd.t437 vdd.t295 200
R2243 vdd.t62 vdd.t437 200
R2244 vdd.t321 vdd.t34 200
R2245 vdd.t177 vdd.t321 200
R2246 vdd.t393 vdd.t511 200
R2247 vdd.t36 vdd.t393 200
R2248 vdd.t471 vdd.t341 200
R2249 vdd.t329 vdd.t471 200
R2250 vdd.t453 vdd.t76 200
R2251 vdd.t343 vdd.t453 200
R2252 vdd.t195 vdd.t2 200
R2253 vdd.t12 vdd.t195 200
R2254 vdd.t159 vdd.t327 200
R2255 vdd.t223 vdd.t159 200
R2256 vdd.t303 vdd.t391 200
R2257 vdd.t42 vdd.t303 200
R2258 vdd.t241 vdd.t48 200
R2259 vdd.t461 vdd.t241 200
R2260 vdd.t499 vdd.t433 200
R2261 vdd.t369 vdd.t499 200
R2262 vdd.t209 vdd.t267 200
R2263 vdd.t259 vdd.t209 200
R2264 vdd.t58 vdd.t379 200
R2265 vdd.t239 vdd.t58 200
R2266 vdd.t253 vdd.t129 200
R2267 vdd.t319 vdd.t253 200
R2268 vdd.t72 vdd.t429 200
R2269 vdd.t515 vdd.t72 200
R2270 vdd.t509 vdd.t281 200
R2271 vdd.t469 vdd.t509 200
R2272 vdd.t153 vdd.t447 200
R2273 vdd.t245 vdd.t153 200
R2274 vdd.t157 vdd.t273 200
R2275 vdd.t199 vdd.t157 200
R2276 vdd.t80 vdd.t413 200
R2277 vdd.t507 vdd.t80 200
R2278 vdd.t431 vdd.t337 200
R2279 vdd.t301 vdd.t431 200
R2280 vdd.t403 vdd.t26 200
R2281 vdd.t331 vdd.t403 200
R2282 vdd.t445 vdd.t333 200
R2283 vdd.t60 vdd.t445 200
R2284 vdd.t383 vdd.t335 200
R2285 vdd.t74 vdd.t383 200
R2286 vdd.t425 vdd.t339 200
R2287 vdd.t155 vdd.t425 200
R2288 vdd.t397 vdd.t28 200
R2289 vdd.t473 vdd.t397 200
R2290 vdd.t367 vdd.t141 200
R2291 vdd.t91 vdd.t367 200
R2292 vdd.t427 vdd.t171 200
R2293 vdd.t345 vdd.t427 200
R2294 vdd.t293 vdd.t457 200
R2295 vdd.t97 vdd.t293 200
R2296 vdd.t137 vdd.t347 200
R2297 vdd.t85 vdd.t137 200
R2298 vdd.t375 vdd.t481 200
R2299 vdd.t201 vdd.t375 200
R2300 vdd.t275 vdd.t8 200
R2301 vdd.t115 vdd.t275 200
R2302 vdd.t16 vdd.t203 200
R2303 vdd.t103 vdd.t16 200
R2304 vdd.t387 vdd.t165 200
R2305 vdd.t287 vdd.t387 200
R2306 vdd.t291 vdd.t50 200
R2307 vdd.t112 vdd.t291 200
R2308 vdd.t18 vdd.t181 200
R2309 vdd.t106 vdd.t18 200
R2310 vdd.t421 vdd.t163 200
R2311 vdd.t227 vdd.t421 200
R2312 vdd.t359 vdd.t217 200
R2313 vdd.t124 vdd.t359 200
R2314 vdd.t22 vdd.t465 200
R2315 vdd.t109 vdd.t22 200
R2316 vdd.t409 vdd.t191 200
R2317 vdd.t243 vdd.t409 200
R2318 vdd.t285 vdd.t317 200
R2319 vdd.t88 vdd.t285 200
R2320 vdd.t215 vdd.t14 200
R2321 vdd.t121 vdd.t215 200
R2322 vdd.t419 vdd.t175 200
R2323 vdd.t56 vdd.t419 200
R2324 vdd.t313 vdd.t353 200
R2325 vdd.t127 vdd.t313 200
R2326 vdd.t495 vdd.t365 200
R2327 vdd.t139 vdd.t495 200
R2328 vdd.t187 vdd.t411 200
R2329 vdd.t235 vdd.t187 200
R2330 vdd.t161 vdd.t251 200
R2331 vdd.t459 vdd.t161 200
R2332 vdd.t185 vdd.t435 200
R2333 vdd.t475 vdd.t185 200
R2334 vdd.t173 vdd.t277 200
R2335 vdd.t4 vdd.t173 200
R2336 vdd.t52 vdd.t381 200
R2337 vdd.t297 vdd.t52 200
R2338 vdd.t483 vdd.t289 200
R2339 vdd.t24 vdd.t483 200
R2340 vdd.t247 vdd.t385 200
R2341 vdd.t38 vdd.t247 200
R2342 vdd.t487 vdd.t357 200
R2343 vdd.t219 vdd.t487 200
R2344 vdd.t479 vdd.t399 200
R2345 vdd.t133 vdd.t479 200
R2346 vdd.t485 vdd.t283 200
R2347 vdd.t315 vdd.t485 200
R2348 vdd.t517 vdd.t405 200
R2349 vdd.t20 vdd.t517 200
R2350 vdd.t373 vdd.t151 200
R2351 vdd.t189 vdd.t373 200
R2352 vdd.t395 vdd.t233 200
R2353 vdd.t183 vdd.t395 200
R2354 vdd.t417 vdd.t477 200
R2355 vdd.t54 vdd.t417 200
R2356 vdd.t451 vdd.t299 200
R2357 vdd.t249 vdd.t451 200
R2358 vdd.t441 vdd.t229 200
R2359 vdd.t363 vdd.t441 200
R2360 vdd.t449 vdd.t135 200
R2361 vdd.t143 vdd.t449 200
R2362 vdd.t255 vdd.t491 200
R2363 vdd.t439 vdd.t255 200
R2364 vdd.t100 vdd.t193 200
R2365 vdd.t263 vdd.t100 200
R2366 vdd.t10 vdd.t145 200
R2367 vdd.t443 vdd.t10 200
R2368 vdd.t489 vdd.t257 200
R2369 vdd.t493 vdd.t489 200
R2370 vdd.t0 vdd.t94 200
R2371 vdd.t497 vdd.t0 200
R2372 vdd.t118 vdd.t311 200
R2373 vdd.t30 vdd.t118 200
R2374 vdd.t307 vdd.t64 200
R2375 vdd.t505 vdd.t307 200
R2376 vdd.t213 vdd.t415 200
R2377 vdd.t78 vdd.t213 200
R2378 vdd.t423 vdd.t309 200
R2379 vdd.t211 vdd.t423 200
R2380 vdd.t66 vdd.t503 200
R2381 vdd.t351 vdd.t66 200
R2382 vdd.t389 vdd.t305 200
R2383 vdd.t231 vdd.t389 200
R2384 vdd.t169 vdd.t269 200
R2385 vdd.t355 vdd.t169 200
R2386 vdd.n483 vdd.n482 68.0765
R2387 vdd.n368 vdd.n367 68.0765
R2388 vdd.n300 vdd.n299 68.0765
R2389 vdd.n232 vdd.n231 68.0765
R2390 vdd.n164 vdd.n163 68.0765
R2391 vdd.n96 vdd.n95 68.0765
R2392 vdd.n401 vdd.n400 68.0765
R2393 vdd.n395 vdd.n394 68.0765
R2394 vdd.n333 vdd.n332 68.0765
R2395 vdd.n327 vdd.n326 68.0765
R2396 vdd.n265 vdd.n264 68.0765
R2397 vdd.n259 vdd.n258 68.0765
R2398 vdd.n197 vdd.n196 68.0765
R2399 vdd.n191 vdd.n190 68.0765
R2400 vdd.n129 vdd.n128 68.0765
R2401 vdd.n123 vdd.n122 68.0765
R2402 vdd.n61 vdd.n60 68.0765
R2403 vdd.n55 vdd.n54 68.0765
R2404 vdd.n478 vdd.n477 68.0765
R2405 vdd.n380 vdd.n379 68.0765
R2406 vdd.n363 vdd.n362 68.0765
R2407 vdd.n312 vdd.n311 68.0765
R2408 vdd.n295 vdd.n294 68.0765
R2409 vdd.n244 vdd.n243 68.0765
R2410 vdd.n227 vdd.n226 68.0765
R2411 vdd.n176 vdd.n175 68.0765
R2412 vdd.n159 vdd.n158 68.0765
R2413 vdd.n108 vdd.n107 68.0765
R2414 vdd.n91 vdd.n90 68.0765
R2415 vdd.n40 vdd.n39 68.0765
R2416 vdd.n406 vdd.n405 68.0765
R2417 vdd.n338 vdd.n337 68.0765
R2418 vdd.n270 vdd.n269 68.0765
R2419 vdd.n202 vdd.n201 68.0765
R2420 vdd.n134 vdd.n133 68.0765
R2421 vdd.n66 vdd.n65 68.0765
R2422 vdd.n473 vdd.n472 68.0765
R2423 vdd.n411 vdd.n410 68.0765
R2424 vdd.n358 vdd.n357 68.0765
R2425 vdd.n390 vdd.n389 68.0765
R2426 vdd.n343 vdd.n342 68.0765
R2427 vdd.n290 vdd.n289 68.0765
R2428 vdd.n322 vdd.n321 68.0765
R2429 vdd.n275 vdd.n274 68.0765
R2430 vdd.n222 vdd.n221 68.0765
R2431 vdd.n254 vdd.n253 68.0765
R2432 vdd.n207 vdd.n206 68.0765
R2433 vdd.n154 vdd.n153 68.0765
R2434 vdd.n186 vdd.n185 68.0765
R2435 vdd.n139 vdd.n138 68.0765
R2436 vdd.n86 vdd.n85 68.0765
R2437 vdd.n118 vdd.n117 68.0765
R2438 vdd.n71 vdd.n70 68.0765
R2439 vdd.n50 vdd.n49 68.0765
R2440 vdd.n468 vdd.n467 68.0765
R2441 vdd.n385 vdd.n384 68.0765
R2442 vdd.n353 vdd.n352 68.0765
R2443 vdd.n317 vdd.n316 68.0765
R2444 vdd.n285 vdd.n284 68.0765
R2445 vdd.n249 vdd.n248 68.0765
R2446 vdd.n217 vdd.n216 68.0765
R2447 vdd.n181 vdd.n180 68.0765
R2448 vdd.n149 vdd.n148 68.0765
R2449 vdd.n113 vdd.n112 68.0765
R2450 vdd.n81 vdd.n80 68.0765
R2451 vdd.n45 vdd.n44 68.0765
R2452 vdd.n416 vdd.n415 68.0765
R2453 vdd.n348 vdd.n347 68.0765
R2454 vdd.n280 vdd.n279 68.0765
R2455 vdd.n212 vdd.n211 68.0765
R2456 vdd.n144 vdd.n143 68.0765
R2457 vdd.n76 vdd.n75 68.0765
R2458 vdd.n421 vdd.n420 68.0765
R2459 vdd.n437 vdd.n436 68.0765
R2460 vdd.n432 vdd.n431 68.0765
R2461 vdd.n455 vdd.n454 68.0765
R2462 vdd.n461 vdd.n460 68.0765
R2463 vdd.n449 vdd.n448 68.0765
R2464 vdd.n26 vdd.n25 68.0765
R2465 vdd.n20 vdd.n19 68.0765
R2466 vdd.n33 vdd.n32 68.0765
R2467 vdd.n3 vdd.n2 68.0765
R2468 vdd.n14 vdd.n13 68.0765
R2469 vdd.n9 vdd.n8 68.0765
R2470 vdd.n30 vdd.n0 66.7247
R2471 vdd.n6 vdd.n0 54.3605
R2472 vdd.n441 vdd.t93 41.0041
R2473 vdd.n444 vdd.t117 40.8177
R2474 vdd.n443 vdd.t99 40.8177
R2475 vdd.n374 vdd.t96 40.6313
R2476 vdd.n372 vdd.t102 40.6313
R2477 vdd.n306 vdd.t114 40.6313
R2478 vdd.n304 vdd.t105 40.6313
R2479 vdd.n238 vdd.t111 40.6313
R2480 vdd.n236 vdd.t108 40.6313
R2481 vdd.n170 vdd.t123 40.6313
R2482 vdd.n168 vdd.t120 40.6313
R2483 vdd.n102 vdd.t87 40.6313
R2484 vdd.n100 vdd.t126 40.6313
R2485 vdd.n426 vdd.t90 40.6313
R2486 vdd.n424 vdd.t84 40.6313
R2487 vdd.n374 vdd.t519 27.3166
R2488 vdd.n372 vdd.t532 27.3166
R2489 vdd.n306 vdd.t529 27.3166
R2490 vdd.n304 vdd.t531 27.3166
R2491 vdd.n238 vdd.t530 27.3166
R2492 vdd.n236 vdd.t528 27.3166
R2493 vdd.n170 vdd.t526 27.3166
R2494 vdd.n168 vdd.t525 27.3166
R2495 vdd.n102 vdd.t522 27.3166
R2496 vdd.n100 vdd.t524 27.3166
R2497 vdd.n426 vdd.t521 27.3166
R2498 vdd.n424 vdd.t523 27.3166
R2499 vdd.n444 vdd.t527 27.1302
R2500 vdd.n443 vdd.t533 27.1302
R2501 vdd.n441 vdd.t520 26.9438
R2502 vdd.n452 dffrs_13.resetb 18.2673
R2503 vdd.n377 vdd.n376 18.0005
R2504 vdd.n309 vdd.n308 18.0005
R2505 vdd.n241 vdd.n240 18.0005
R2506 vdd.n173 vdd.n172 18.0005
R2507 vdd.n105 vdd.n104 18.0005
R2508 vdd.n429 vdd.n428 18.0005
R2509 vdd.n6 vdd.n5 13.533
R2510 vdd.n429 vdd.n423 13.5152
R2511 vdd.n486 vdd.n485 13.5005
R2512 vdd.n371 vdd.n370 13.5005
R2513 vdd.n303 vdd.n302 13.5005
R2514 vdd.n235 vdd.n234 13.5005
R2515 vdd.n167 vdd.n166 13.5005
R2516 vdd.n99 vdd.n98 13.5005
R2517 vdd.n486 vdd.n403 13.5005
R2518 vdd.n398 vdd.n397 13.5005
R2519 vdd.n371 vdd.n335 13.5005
R2520 vdd.n330 vdd.n329 13.5005
R2521 vdd.n303 vdd.n267 13.5005
R2522 vdd.n262 vdd.n261 13.5005
R2523 vdd.n235 vdd.n199 13.5005
R2524 vdd.n194 vdd.n193 13.5005
R2525 vdd.n167 vdd.n131 13.5005
R2526 vdd.n126 vdd.n125 13.5005
R2527 vdd.n99 vdd.n63 13.5005
R2528 vdd.n58 vdd.n57 13.5005
R2529 vdd.n486 vdd.n480 13.5005
R2530 vdd.n398 vdd.n382 13.5005
R2531 vdd.n371 vdd.n365 13.5005
R2532 vdd.n330 vdd.n314 13.5005
R2533 vdd.n303 vdd.n297 13.5005
R2534 vdd.n262 vdd.n246 13.5005
R2535 vdd.n235 vdd.n229 13.5005
R2536 vdd.n194 vdd.n178 13.5005
R2537 vdd.n167 vdd.n161 13.5005
R2538 vdd.n126 vdd.n110 13.5005
R2539 vdd.n99 vdd.n93 13.5005
R2540 vdd.n58 vdd.n42 13.5005
R2541 vdd.n486 vdd.n408 13.5005
R2542 vdd.n371 vdd.n340 13.5005
R2543 vdd.n303 vdd.n272 13.5005
R2544 vdd.n235 vdd.n204 13.5005
R2545 vdd.n167 vdd.n136 13.5005
R2546 vdd.n99 vdd.n68 13.5005
R2547 vdd.n486 vdd.n475 13.5005
R2548 vdd.n486 vdd.n413 13.5005
R2549 vdd.n371 vdd.n360 13.5005
R2550 vdd.n398 vdd.n392 13.5005
R2551 vdd.n371 vdd.n345 13.5005
R2552 vdd.n303 vdd.n292 13.5005
R2553 vdd.n330 vdd.n324 13.5005
R2554 vdd.n303 vdd.n277 13.5005
R2555 vdd.n235 vdd.n224 13.5005
R2556 vdd.n262 vdd.n256 13.5005
R2557 vdd.n235 vdd.n209 13.5005
R2558 vdd.n167 vdd.n156 13.5005
R2559 vdd.n194 vdd.n188 13.5005
R2560 vdd.n167 vdd.n141 13.5005
R2561 vdd.n99 vdd.n88 13.5005
R2562 vdd.n126 vdd.n120 13.5005
R2563 vdd.n99 vdd.n73 13.5005
R2564 vdd.n58 vdd.n52 13.5005
R2565 vdd.n486 vdd.n470 13.5005
R2566 vdd.n398 vdd.n387 13.5005
R2567 vdd.n371 vdd.n355 13.5005
R2568 vdd.n330 vdd.n319 13.5005
R2569 vdd.n303 vdd.n287 13.5005
R2570 vdd.n262 vdd.n251 13.5005
R2571 vdd.n235 vdd.n219 13.5005
R2572 vdd.n194 vdd.n183 13.5005
R2573 vdd.n167 vdd.n151 13.5005
R2574 vdd.n126 vdd.n115 13.5005
R2575 vdd.n99 vdd.n83 13.5005
R2576 vdd.n58 vdd.n47 13.5005
R2577 vdd.n486 vdd.n418 13.5005
R2578 vdd.n371 vdd.n350 13.5005
R2579 vdd.n303 vdd.n282 13.5005
R2580 vdd.n235 vdd.n214 13.5005
R2581 vdd.n167 vdd.n146 13.5005
R2582 vdd.n99 vdd.n78 13.5005
R2583 vdd.n440 vdd.n439 13.5005
R2584 vdd.n440 vdd.n434 13.5005
R2585 vdd.n458 vdd.n457 13.5005
R2586 vdd.n464 vdd.n463 13.5005
R2587 vdd.n452 vdd.n451 13.5005
R2588 vdd.n29 vdd.n28 13.5005
R2589 vdd.n23 vdd.n22 13.5005
R2590 vdd.n36 vdd.n35 13.5005
R2591 vdd.n17 vdd.n16 13.5005
R2592 vdd.n17 vdd.n11 13.5005
R2593 vdd.n445 dffrs_13.nand3_1.B 12.1571
R2594 vdd.n375 vdd.n373 9.22229
R2595 vdd.n307 vdd.n305 9.22229
R2596 vdd.n239 vdd.n237 9.22229
R2597 vdd.n171 vdd.n169 9.22229
R2598 vdd.n103 vdd.n101 9.22229
R2599 vdd.n427 vdd.n425 9.22229
R2600 vdd.n446 vdd.n442 7.75389
R2601 vdd.n485 vdd.n482 6.4802
R2602 vdd.n370 vdd.n367 6.4802
R2603 vdd.n302 vdd.n299 6.4802
R2604 vdd.n234 vdd.n231 6.4802
R2605 vdd.n166 vdd.n163 6.4802
R2606 vdd.n98 vdd.n95 6.4802
R2607 vdd.n403 vdd.n400 6.4802
R2608 vdd.n397 vdd.n394 6.4802
R2609 vdd.n335 vdd.n332 6.4802
R2610 vdd.n329 vdd.n326 6.4802
R2611 vdd.n267 vdd.n264 6.4802
R2612 vdd.n261 vdd.n258 6.4802
R2613 vdd.n199 vdd.n196 6.4802
R2614 vdd.n193 vdd.n190 6.4802
R2615 vdd.n131 vdd.n128 6.4802
R2616 vdd.n125 vdd.n122 6.4802
R2617 vdd.n63 vdd.n60 6.4802
R2618 vdd.n57 vdd.n54 6.4802
R2619 vdd.n480 vdd.n477 6.4802
R2620 vdd.n382 vdd.n379 6.4802
R2621 vdd.n365 vdd.n362 6.4802
R2622 vdd.n314 vdd.n311 6.4802
R2623 vdd.n297 vdd.n294 6.4802
R2624 vdd.n246 vdd.n243 6.4802
R2625 vdd.n229 vdd.n226 6.4802
R2626 vdd.n178 vdd.n175 6.4802
R2627 vdd.n161 vdd.n158 6.4802
R2628 vdd.n110 vdd.n107 6.4802
R2629 vdd.n93 vdd.n90 6.4802
R2630 vdd.n42 vdd.n39 6.4802
R2631 vdd.n408 vdd.n405 6.4802
R2632 vdd.n340 vdd.n337 6.4802
R2633 vdd.n272 vdd.n269 6.4802
R2634 vdd.n204 vdd.n201 6.4802
R2635 vdd.n136 vdd.n133 6.4802
R2636 vdd.n68 vdd.n65 6.4802
R2637 vdd.n475 vdd.n472 6.4802
R2638 vdd.n413 vdd.n410 6.4802
R2639 vdd.n360 vdd.n357 6.4802
R2640 vdd.n392 vdd.n389 6.4802
R2641 vdd.n345 vdd.n342 6.4802
R2642 vdd.n292 vdd.n289 6.4802
R2643 vdd.n324 vdd.n321 6.4802
R2644 vdd.n277 vdd.n274 6.4802
R2645 vdd.n224 vdd.n221 6.4802
R2646 vdd.n256 vdd.n253 6.4802
R2647 vdd.n209 vdd.n206 6.4802
R2648 vdd.n156 vdd.n153 6.4802
R2649 vdd.n188 vdd.n185 6.4802
R2650 vdd.n141 vdd.n138 6.4802
R2651 vdd.n88 vdd.n85 6.4802
R2652 vdd.n120 vdd.n117 6.4802
R2653 vdd.n73 vdd.n70 6.4802
R2654 vdd.n52 vdd.n49 6.4802
R2655 vdd.n470 vdd.n467 6.4802
R2656 vdd.n387 vdd.n384 6.4802
R2657 vdd.n355 vdd.n352 6.4802
R2658 vdd.n319 vdd.n316 6.4802
R2659 vdd.n287 vdd.n284 6.4802
R2660 vdd.n251 vdd.n248 6.4802
R2661 vdd.n219 vdd.n216 6.4802
R2662 vdd.n183 vdd.n180 6.4802
R2663 vdd.n151 vdd.n148 6.4802
R2664 vdd.n115 vdd.n112 6.4802
R2665 vdd.n83 vdd.n80 6.4802
R2666 vdd.n47 vdd.n44 6.4802
R2667 vdd.n418 vdd.n415 6.4802
R2668 vdd.n350 vdd.n347 6.4802
R2669 vdd.n282 vdd.n279 6.4802
R2670 vdd.n214 vdd.n211 6.4802
R2671 vdd.n146 vdd.n143 6.4802
R2672 vdd.n78 vdd.n75 6.4802
R2673 vdd.n423 vdd.n420 6.4802
R2674 vdd.n439 vdd.n436 6.4802
R2675 vdd.n434 vdd.n431 6.4802
R2676 vdd.n457 vdd.n454 6.4802
R2677 vdd.n463 vdd.n460 6.4802
R2678 vdd.n451 vdd.n448 6.4802
R2679 vdd.n28 vdd.n25 6.4802
R2680 vdd.n22 vdd.n19 6.4802
R2681 vdd.n35 vdd.n32 6.4802
R2682 vdd.n5 vdd.n2 6.4802
R2683 vdd.n16 vdd.n13 6.4802
R2684 vdd.n11 vdd.n8 6.4802
R2685 vdd.n485 vdd.n481 6.25878
R2686 vdd.n370 vdd.n366 6.25878
R2687 vdd.n302 vdd.n298 6.25878
R2688 vdd.n234 vdd.n230 6.25878
R2689 vdd.n166 vdd.n162 6.25878
R2690 vdd.n98 vdd.n94 6.25878
R2691 vdd.n403 vdd.n399 6.25878
R2692 vdd.n397 vdd.n393 6.25878
R2693 vdd.n335 vdd.n331 6.25878
R2694 vdd.n329 vdd.n325 6.25878
R2695 vdd.n267 vdd.n263 6.25878
R2696 vdd.n261 vdd.n257 6.25878
R2697 vdd.n199 vdd.n195 6.25878
R2698 vdd.n193 vdd.n189 6.25878
R2699 vdd.n131 vdd.n127 6.25878
R2700 vdd.n125 vdd.n121 6.25878
R2701 vdd.n63 vdd.n59 6.25878
R2702 vdd.n57 vdd.n53 6.25878
R2703 vdd.n480 vdd.n476 6.25878
R2704 vdd.n382 vdd.n378 6.25878
R2705 vdd.n365 vdd.n361 6.25878
R2706 vdd.n314 vdd.n310 6.25878
R2707 vdd.n297 vdd.n293 6.25878
R2708 vdd.n246 vdd.n242 6.25878
R2709 vdd.n229 vdd.n225 6.25878
R2710 vdd.n178 vdd.n174 6.25878
R2711 vdd.n161 vdd.n157 6.25878
R2712 vdd.n110 vdd.n106 6.25878
R2713 vdd.n93 vdd.n89 6.25878
R2714 vdd.n42 vdd.n38 6.25878
R2715 vdd.n408 vdd.n404 6.25878
R2716 vdd.n340 vdd.n336 6.25878
R2717 vdd.n272 vdd.n268 6.25878
R2718 vdd.n204 vdd.n200 6.25878
R2719 vdd.n136 vdd.n132 6.25878
R2720 vdd.n68 vdd.n64 6.25878
R2721 vdd.n475 vdd.n471 6.25878
R2722 vdd.n413 vdd.n409 6.25878
R2723 vdd.n360 vdd.n356 6.25878
R2724 vdd.n392 vdd.n388 6.25878
R2725 vdd.n345 vdd.n341 6.25878
R2726 vdd.n292 vdd.n288 6.25878
R2727 vdd.n324 vdd.n320 6.25878
R2728 vdd.n277 vdd.n273 6.25878
R2729 vdd.n224 vdd.n220 6.25878
R2730 vdd.n256 vdd.n252 6.25878
R2731 vdd.n209 vdd.n205 6.25878
R2732 vdd.n156 vdd.n152 6.25878
R2733 vdd.n188 vdd.n184 6.25878
R2734 vdd.n141 vdd.n137 6.25878
R2735 vdd.n88 vdd.n84 6.25878
R2736 vdd.n120 vdd.n116 6.25878
R2737 vdd.n73 vdd.n69 6.25878
R2738 vdd.n52 vdd.n48 6.25878
R2739 vdd.n470 vdd.n466 6.25878
R2740 vdd.n387 vdd.n383 6.25878
R2741 vdd.n355 vdd.n351 6.25878
R2742 vdd.n319 vdd.n315 6.25878
R2743 vdd.n287 vdd.n283 6.25878
R2744 vdd.n251 vdd.n247 6.25878
R2745 vdd.n219 vdd.n215 6.25878
R2746 vdd.n183 vdd.n179 6.25878
R2747 vdd.n151 vdd.n147 6.25878
R2748 vdd.n115 vdd.n111 6.25878
R2749 vdd.n83 vdd.n79 6.25878
R2750 vdd.n47 vdd.n43 6.25878
R2751 vdd.n418 vdd.n414 6.25878
R2752 vdd.n350 vdd.n346 6.25878
R2753 vdd.n282 vdd.n278 6.25878
R2754 vdd.n214 vdd.n210 6.25878
R2755 vdd.n146 vdd.n142 6.25878
R2756 vdd.n78 vdd.n74 6.25878
R2757 vdd.n423 vdd.n419 6.25878
R2758 vdd.n439 vdd.n435 6.25878
R2759 vdd.n434 vdd.n430 6.25878
R2760 vdd.n457 vdd.n453 6.25878
R2761 vdd.n463 vdd.n459 6.25878
R2762 vdd.n451 vdd.n447 6.25878
R2763 vdd.n28 vdd.n24 6.25878
R2764 vdd.n22 vdd.n18 6.25878
R2765 vdd.n35 vdd.n31 6.25878
R2766 vdd.n5 vdd.n1 6.25878
R2767 vdd.n16 vdd.n12 6.25878
R2768 vdd.n11 vdd.n7 6.25878
R2769 vdd.n446 vdd.n445 5.93546
R2770 vdd.n442 vdd.n441 5.7305
R2771 dffrs_13.nand3_8.B vdd.n444 5.47979
R2772 dffrs_13.nand3_1.B vdd.n443 5.47979
R2773 vdd.n485 vdd.n484 5.44497
R2774 vdd.n370 vdd.n369 5.44497
R2775 vdd.n302 vdd.n301 5.44497
R2776 vdd.n234 vdd.n233 5.44497
R2777 vdd.n166 vdd.n165 5.44497
R2778 vdd.n98 vdd.n97 5.44497
R2779 vdd.n403 vdd.n402 5.44497
R2780 vdd.n397 vdd.n396 5.44497
R2781 vdd.n335 vdd.n334 5.44497
R2782 vdd.n329 vdd.n328 5.44497
R2783 vdd.n267 vdd.n266 5.44497
R2784 vdd.n261 vdd.n260 5.44497
R2785 vdd.n199 vdd.n198 5.44497
R2786 vdd.n193 vdd.n192 5.44497
R2787 vdd.n131 vdd.n130 5.44497
R2788 vdd.n125 vdd.n124 5.44497
R2789 vdd.n63 vdd.n62 5.44497
R2790 vdd.n57 vdd.n56 5.44497
R2791 vdd.n480 vdd.n479 5.44497
R2792 vdd.n382 vdd.n381 5.44497
R2793 vdd.n365 vdd.n364 5.44497
R2794 vdd.n314 vdd.n313 5.44497
R2795 vdd.n297 vdd.n296 5.44497
R2796 vdd.n246 vdd.n245 5.44497
R2797 vdd.n229 vdd.n228 5.44497
R2798 vdd.n178 vdd.n177 5.44497
R2799 vdd.n161 vdd.n160 5.44497
R2800 vdd.n110 vdd.n109 5.44497
R2801 vdd.n93 vdd.n92 5.44497
R2802 vdd.n42 vdd.n41 5.44497
R2803 vdd.n408 vdd.n407 5.44497
R2804 vdd.n340 vdd.n339 5.44497
R2805 vdd.n272 vdd.n271 5.44497
R2806 vdd.n204 vdd.n203 5.44497
R2807 vdd.n136 vdd.n135 5.44497
R2808 vdd.n68 vdd.n67 5.44497
R2809 vdd.n475 vdd.n474 5.44497
R2810 vdd.n413 vdd.n412 5.44497
R2811 vdd.n360 vdd.n359 5.44497
R2812 vdd.n392 vdd.n391 5.44497
R2813 vdd.n345 vdd.n344 5.44497
R2814 vdd.n292 vdd.n291 5.44497
R2815 vdd.n324 vdd.n323 5.44497
R2816 vdd.n277 vdd.n276 5.44497
R2817 vdd.n224 vdd.n223 5.44497
R2818 vdd.n256 vdd.n255 5.44497
R2819 vdd.n209 vdd.n208 5.44497
R2820 vdd.n156 vdd.n155 5.44497
R2821 vdd.n188 vdd.n187 5.44497
R2822 vdd.n141 vdd.n140 5.44497
R2823 vdd.n88 vdd.n87 5.44497
R2824 vdd.n120 vdd.n119 5.44497
R2825 vdd.n73 vdd.n72 5.44497
R2826 vdd.n52 vdd.n51 5.44497
R2827 vdd.n470 vdd.n469 5.44497
R2828 vdd.n387 vdd.n386 5.44497
R2829 vdd.n355 vdd.n354 5.44497
R2830 vdd.n319 vdd.n318 5.44497
R2831 vdd.n287 vdd.n286 5.44497
R2832 vdd.n251 vdd.n250 5.44497
R2833 vdd.n219 vdd.n218 5.44497
R2834 vdd.n183 vdd.n182 5.44497
R2835 vdd.n151 vdd.n150 5.44497
R2836 vdd.n115 vdd.n114 5.44497
R2837 vdd.n83 vdd.n82 5.44497
R2838 vdd.n47 vdd.n46 5.44497
R2839 vdd.n418 vdd.n417 5.44497
R2840 vdd.n350 vdd.n349 5.44497
R2841 vdd.n282 vdd.n281 5.44497
R2842 vdd.n214 vdd.n213 5.44497
R2843 vdd.n146 vdd.n145 5.44497
R2844 vdd.n78 vdd.n77 5.44497
R2845 vdd.n423 vdd.n422 5.44497
R2846 vdd.n439 vdd.n438 5.44497
R2847 vdd.n434 vdd.n433 5.44497
R2848 vdd.n457 vdd.n456 5.44497
R2849 vdd.n463 vdd.n462 5.44497
R2850 vdd.n451 vdd.n450 5.44497
R2851 vdd.n28 vdd.n27 5.44497
R2852 vdd.n22 vdd.n21 5.44497
R2853 vdd.n35 vdd.n34 5.44497
R2854 vdd.n5 vdd.n4 5.44497
R2855 vdd.n16 vdd.n15 5.44497
R2856 vdd.n11 vdd.n10 5.44497
R2857 vdd.n375 vdd.n374 5.14711
R2858 vdd.n307 vdd.n306 5.14711
R2859 vdd.n239 vdd.n238 5.14711
R2860 vdd.n171 vdd.n170 5.14711
R2861 vdd.n103 vdd.n102 5.14711
R2862 vdd.n427 vdd.n426 5.14711
R2863 vdd.n373 vdd.n372 5.13907
R2864 vdd.n305 vdd.n304 5.13907
R2865 vdd.n237 vdd.n236 5.13907
R2866 vdd.n169 vdd.n168 5.13907
R2867 vdd.n101 vdd.n100 5.13907
R2868 vdd.n425 vdd.n424 5.13907
R2869 vdd.n445 dffrs_13.nand3_8.B 5.09593
R2870 vdd.n484 vdd.t150 1.85637
R2871 vdd.n369 vdd.t71 1.85637
R2872 vdd.n301 vdd.t168 1.85637
R2873 vdd.n233 vdd.t180 1.85637
R2874 vdd.n165 vdd.t464 1.85637
R2875 vdd.n97 vdd.t502 1.85637
R2876 vdd.n402 vdd.t83 1.85637
R2877 vdd.n396 vdd.t148 1.85637
R2878 vdd.n334 vdd.t362 1.85637
R2879 vdd.n328 vdd.t69 1.85637
R2880 vdd.n266 vdd.t45 1.85637
R2881 vdd.n260 vdd.t206 1.85637
R2882 vdd.n198 vdd.t63 1.85637
R2883 vdd.n192 vdd.t178 1.85637
R2884 vdd.n130 vdd.t37 1.85637
R2885 vdd.n124 vdd.t330 1.85637
R2886 vdd.n62 vdd.t344 1.85637
R2887 vdd.n56 vdd.t13 1.85637
R2888 vdd.n479 vdd.t224 1.85637
R2889 vdd.n381 vdd.t43 1.85637
R2890 vdd.n364 vdd.t462 1.85637
R2891 vdd.n313 vdd.t370 1.85637
R2892 vdd.n296 vdd.t260 1.85637
R2893 vdd.n245 vdd.t240 1.85637
R2894 vdd.n228 vdd.t320 1.85637
R2895 vdd.n177 vdd.t516 1.85637
R2896 vdd.n160 vdd.t470 1.85637
R2897 vdd.n109 vdd.t246 1.85637
R2898 vdd.n92 vdd.t200 1.85637
R2899 vdd.n41 vdd.t508 1.85637
R2900 vdd.n407 vdd.t302 1.85637
R2901 vdd.n339 vdd.t332 1.85637
R2902 vdd.n271 vdd.t61 1.85637
R2903 vdd.n203 vdd.t75 1.85637
R2904 vdd.n135 vdd.t156 1.85637
R2905 vdd.n67 vdd.t474 1.85637
R2906 vdd.n474 vdd.t92 1.85637
R2907 vdd.n412 vdd.t346 1.85637
R2908 vdd.n359 vdd.t98 1.85637
R2909 vdd.n391 vdd.t86 1.85637
R2910 vdd.n344 vdd.t202 1.85637
R2911 vdd.n291 vdd.t116 1.85637
R2912 vdd.n323 vdd.t104 1.85637
R2913 vdd.n276 vdd.t288 1.85637
R2914 vdd.n223 vdd.t113 1.85637
R2915 vdd.n255 vdd.t107 1.85637
R2916 vdd.n208 vdd.t228 1.85637
R2917 vdd.n155 vdd.t125 1.85637
R2918 vdd.n187 vdd.t110 1.85637
R2919 vdd.n140 vdd.t244 1.85637
R2920 vdd.n87 vdd.t89 1.85637
R2921 vdd.n119 vdd.t122 1.85637
R2922 vdd.n72 vdd.t57 1.85637
R2923 vdd.n51 vdd.t128 1.85637
R2924 vdd.n469 vdd.t140 1.85637
R2925 vdd.n386 vdd.t236 1.85637
R2926 vdd.n354 vdd.t460 1.85637
R2927 vdd.n318 vdd.t476 1.85637
R2928 vdd.n286 vdd.t5 1.85637
R2929 vdd.n250 vdd.t298 1.85637
R2930 vdd.n218 vdd.t25 1.85637
R2931 vdd.n182 vdd.t39 1.85637
R2932 vdd.n150 vdd.t220 1.85637
R2933 vdd.n114 vdd.t134 1.85637
R2934 vdd.n82 vdd.t316 1.85637
R2935 vdd.n46 vdd.t21 1.85637
R2936 vdd.n417 vdd.t190 1.85637
R2937 vdd.n349 vdd.t184 1.85637
R2938 vdd.n281 vdd.t55 1.85637
R2939 vdd.n213 vdd.t250 1.85637
R2940 vdd.n145 vdd.t364 1.85637
R2941 vdd.n77 vdd.t144 1.85637
R2942 vdd.n422 vdd.t440 1.85637
R2943 vdd.n438 vdd.t264 1.85637
R2944 vdd.n433 vdd.t444 1.85637
R2945 vdd.n456 vdd.t494 1.85637
R2946 vdd.n462 vdd.t498 1.85637
R2947 vdd.n450 vdd.t31 1.85637
R2948 vdd.n27 vdd.t506 1.85637
R2949 vdd.n21 vdd.t79 1.85637
R2950 vdd.n34 vdd.t212 1.85637
R2951 vdd.n4 vdd.t352 1.85637
R2952 vdd.n15 vdd.t232 1.85637
R2953 vdd.n10 vdd.t356 1.85637
R2954 vdd.n484 vdd.n483 1.04105
R2955 vdd.n369 vdd.n368 1.04105
R2956 vdd.n301 vdd.n300 1.04105
R2957 vdd.n233 vdd.n232 1.04105
R2958 vdd.n165 vdd.n164 1.04105
R2959 vdd.n97 vdd.n96 1.04105
R2960 vdd.n402 vdd.n401 1.04105
R2961 vdd.n396 vdd.n395 1.04105
R2962 vdd.n334 vdd.n333 1.04105
R2963 vdd.n328 vdd.n327 1.04105
R2964 vdd.n266 vdd.n265 1.04105
R2965 vdd.n260 vdd.n259 1.04105
R2966 vdd.n198 vdd.n197 1.04105
R2967 vdd.n192 vdd.n191 1.04105
R2968 vdd.n130 vdd.n129 1.04105
R2969 vdd.n124 vdd.n123 1.04105
R2970 vdd.n62 vdd.n61 1.04105
R2971 vdd.n56 vdd.n55 1.04105
R2972 vdd.n479 vdd.n478 1.04105
R2973 vdd.n381 vdd.n380 1.04105
R2974 vdd.n364 vdd.n363 1.04105
R2975 vdd.n313 vdd.n312 1.04105
R2976 vdd.n296 vdd.n295 1.04105
R2977 vdd.n245 vdd.n244 1.04105
R2978 vdd.n228 vdd.n227 1.04105
R2979 vdd.n177 vdd.n176 1.04105
R2980 vdd.n160 vdd.n159 1.04105
R2981 vdd.n109 vdd.n108 1.04105
R2982 vdd.n92 vdd.n91 1.04105
R2983 vdd.n41 vdd.n40 1.04105
R2984 vdd.n407 vdd.n406 1.04105
R2985 vdd.n339 vdd.n338 1.04105
R2986 vdd.n271 vdd.n270 1.04105
R2987 vdd.n203 vdd.n202 1.04105
R2988 vdd.n135 vdd.n134 1.04105
R2989 vdd.n67 vdd.n66 1.04105
R2990 vdd.n474 vdd.n473 1.04105
R2991 vdd.n412 vdd.n411 1.04105
R2992 vdd.n359 vdd.n358 1.04105
R2993 vdd.n391 vdd.n390 1.04105
R2994 vdd.n344 vdd.n343 1.04105
R2995 vdd.n291 vdd.n290 1.04105
R2996 vdd.n323 vdd.n322 1.04105
R2997 vdd.n276 vdd.n275 1.04105
R2998 vdd.n223 vdd.n222 1.04105
R2999 vdd.n255 vdd.n254 1.04105
R3000 vdd.n208 vdd.n207 1.04105
R3001 vdd.n155 vdd.n154 1.04105
R3002 vdd.n187 vdd.n186 1.04105
R3003 vdd.n140 vdd.n139 1.04105
R3004 vdd.n87 vdd.n86 1.04105
R3005 vdd.n119 vdd.n118 1.04105
R3006 vdd.n72 vdd.n71 1.04105
R3007 vdd.n51 vdd.n50 1.04105
R3008 vdd.n469 vdd.n468 1.04105
R3009 vdd.n386 vdd.n385 1.04105
R3010 vdd.n354 vdd.n353 1.04105
R3011 vdd.n318 vdd.n317 1.04105
R3012 vdd.n286 vdd.n285 1.04105
R3013 vdd.n250 vdd.n249 1.04105
R3014 vdd.n218 vdd.n217 1.04105
R3015 vdd.n182 vdd.n181 1.04105
R3016 vdd.n150 vdd.n149 1.04105
R3017 vdd.n114 vdd.n113 1.04105
R3018 vdd.n82 vdd.n81 1.04105
R3019 vdd.n46 vdd.n45 1.04105
R3020 vdd.n417 vdd.n416 1.04105
R3021 vdd.n349 vdd.n348 1.04105
R3022 vdd.n281 vdd.n280 1.04105
R3023 vdd.n213 vdd.n212 1.04105
R3024 vdd.n145 vdd.n144 1.04105
R3025 vdd.n77 vdd.n76 1.04105
R3026 vdd.n422 vdd.n421 1.04105
R3027 vdd.n438 vdd.n437 1.04105
R3028 vdd.n433 vdd.n432 1.04105
R3029 vdd.n456 vdd.n455 1.04105
R3030 vdd.n462 vdd.n461 1.04105
R3031 vdd.n450 vdd.n449 1.04105
R3032 vdd.n27 vdd.n26 1.04105
R3033 vdd.n21 vdd.n20 1.04105
R3034 vdd.n34 vdd.n33 1.04105
R3035 vdd.n4 vdd.n3 1.04105
R3036 vdd.n15 vdd.n14 1.04105
R3037 vdd.n10 vdd.n9 1.04105
R3038 vdd.n37 vdd.n36 0.839436
R3039 vdd.n481 vdd.t226 0.7285
R3040 vdd.n481 vdd.t326 0.7285
R3041 vdd.n366 vdd.t7 0.7285
R3042 vdd.n366 vdd.t47 0.7285
R3043 vdd.n298 vdd.t262 0.7285
R3044 vdd.n298 vdd.t266 0.7285
R3045 vdd.n230 vdd.t324 0.7285
R3046 vdd.n230 vdd.t132 0.7285
R3047 vdd.n162 vdd.t468 0.7285
R3048 vdd.n162 vdd.t280 0.7285
R3049 vdd.n94 vdd.t198 0.7285
R3050 vdd.n94 vdd.t272 0.7285
R3051 vdd.n399 vdd.t372 0.7285
R3052 vdd.n399 vdd.t402 0.7285
R3053 vdd.n393 vdd.t208 0.7285
R3054 vdd.n393 vdd.t222 0.7285
R3055 vdd.n331 vdd.t350 0.7285
R3056 vdd.n331 vdd.t378 0.7285
R3057 vdd.n325 vdd.t41 0.7285
R3058 vdd.n325 vdd.t456 0.7285
R3059 vdd.n263 vdd.t514 0.7285
R3060 vdd.n263 vdd.t408 0.7285
R3061 vdd.n257 vdd.t33 0.7285
R3062 vdd.n257 vdd.t238 0.7285
R3063 vdd.n195 vdd.t296 0.7285
R3064 vdd.n195 vdd.t438 0.7285
R3065 vdd.n189 vdd.t35 0.7285
R3066 vdd.n189 vdd.t322 0.7285
R3067 vdd.n127 vdd.t512 0.7285
R3068 vdd.n127 vdd.t394 0.7285
R3069 vdd.n121 vdd.t342 0.7285
R3070 vdd.n121 vdd.t472 0.7285
R3071 vdd.n59 vdd.t77 0.7285
R3072 vdd.n59 vdd.t454 0.7285
R3073 vdd.n53 vdd.t3 0.7285
R3074 vdd.n53 vdd.t196 0.7285
R3075 vdd.n476 vdd.t328 0.7285
R3076 vdd.n476 vdd.t160 0.7285
R3077 vdd.n378 vdd.t392 0.7285
R3078 vdd.n378 vdd.t304 0.7285
R3079 vdd.n361 vdd.t49 0.7285
R3080 vdd.n361 vdd.t242 0.7285
R3081 vdd.n310 vdd.t434 0.7285
R3082 vdd.n310 vdd.t500 0.7285
R3083 vdd.n293 vdd.t268 0.7285
R3084 vdd.n293 vdd.t210 0.7285
R3085 vdd.n242 vdd.t380 0.7285
R3086 vdd.n242 vdd.t59 0.7285
R3087 vdd.n225 vdd.t130 0.7285
R3088 vdd.n225 vdd.t254 0.7285
R3089 vdd.n174 vdd.t430 0.7285
R3090 vdd.n174 vdd.t73 0.7285
R3091 vdd.n157 vdd.t282 0.7285
R3092 vdd.n157 vdd.t510 0.7285
R3093 vdd.n106 vdd.t448 0.7285
R3094 vdd.n106 vdd.t154 0.7285
R3095 vdd.n89 vdd.t274 0.7285
R3096 vdd.n89 vdd.t158 0.7285
R3097 vdd.n38 vdd.t414 0.7285
R3098 vdd.n38 vdd.t81 0.7285
R3099 vdd.n404 vdd.t338 0.7285
R3100 vdd.n404 vdd.t432 0.7285
R3101 vdd.n336 vdd.t27 0.7285
R3102 vdd.n336 vdd.t404 0.7285
R3103 vdd.n268 vdd.t334 0.7285
R3104 vdd.n268 vdd.t446 0.7285
R3105 vdd.n200 vdd.t336 0.7285
R3106 vdd.n200 vdd.t384 0.7285
R3107 vdd.n132 vdd.t340 0.7285
R3108 vdd.n132 vdd.t426 0.7285
R3109 vdd.n64 vdd.t29 0.7285
R3110 vdd.n64 vdd.t398 0.7285
R3111 vdd.n471 vdd.t142 0.7285
R3112 vdd.n471 vdd.t368 0.7285
R3113 vdd.n409 vdd.t172 0.7285
R3114 vdd.n409 vdd.t428 0.7285
R3115 vdd.n356 vdd.t458 0.7285
R3116 vdd.n356 vdd.t294 0.7285
R3117 vdd.n388 vdd.t348 0.7285
R3118 vdd.n388 vdd.t138 0.7285
R3119 vdd.n341 vdd.t482 0.7285
R3120 vdd.n341 vdd.t376 0.7285
R3121 vdd.n288 vdd.t9 0.7285
R3122 vdd.n288 vdd.t276 0.7285
R3123 vdd.n320 vdd.t204 0.7285
R3124 vdd.n320 vdd.t17 0.7285
R3125 vdd.n273 vdd.t166 0.7285
R3126 vdd.n273 vdd.t388 0.7285
R3127 vdd.n220 vdd.t51 0.7285
R3128 vdd.n220 vdd.t292 0.7285
R3129 vdd.n252 vdd.t182 0.7285
R3130 vdd.n252 vdd.t19 0.7285
R3131 vdd.n205 vdd.t164 0.7285
R3132 vdd.n205 vdd.t422 0.7285
R3133 vdd.n152 vdd.t218 0.7285
R3134 vdd.n152 vdd.t360 0.7285
R3135 vdd.n184 vdd.t466 0.7285
R3136 vdd.n184 vdd.t23 0.7285
R3137 vdd.n137 vdd.t192 0.7285
R3138 vdd.n137 vdd.t410 0.7285
R3139 vdd.n84 vdd.t318 0.7285
R3140 vdd.n84 vdd.t286 0.7285
R3141 vdd.n116 vdd.t15 0.7285
R3142 vdd.n116 vdd.t216 0.7285
R3143 vdd.n69 vdd.t176 0.7285
R3144 vdd.n69 vdd.t420 0.7285
R3145 vdd.n48 vdd.t354 0.7285
R3146 vdd.n48 vdd.t314 0.7285
R3147 vdd.n466 vdd.t366 0.7285
R3148 vdd.n466 vdd.t496 0.7285
R3149 vdd.n383 vdd.t412 0.7285
R3150 vdd.n383 vdd.t188 0.7285
R3151 vdd.n351 vdd.t252 0.7285
R3152 vdd.n351 vdd.t162 0.7285
R3153 vdd.n315 vdd.t436 0.7285
R3154 vdd.n315 vdd.t186 0.7285
R3155 vdd.n283 vdd.t278 0.7285
R3156 vdd.n283 vdd.t174 0.7285
R3157 vdd.n247 vdd.t382 0.7285
R3158 vdd.n247 vdd.t53 0.7285
R3159 vdd.n215 vdd.t290 0.7285
R3160 vdd.n215 vdd.t484 0.7285
R3161 vdd.n179 vdd.t386 0.7285
R3162 vdd.n179 vdd.t248 0.7285
R3163 vdd.n147 vdd.t358 0.7285
R3164 vdd.n147 vdd.t488 0.7285
R3165 vdd.n111 vdd.t400 0.7285
R3166 vdd.n111 vdd.t480 0.7285
R3167 vdd.n79 vdd.t284 0.7285
R3168 vdd.n79 vdd.t486 0.7285
R3169 vdd.n43 vdd.t406 0.7285
R3170 vdd.n43 vdd.t518 0.7285
R3171 vdd.n414 vdd.t152 0.7285
R3172 vdd.n414 vdd.t374 0.7285
R3173 vdd.n346 vdd.t234 0.7285
R3174 vdd.n346 vdd.t396 0.7285
R3175 vdd.n278 vdd.t478 0.7285
R3176 vdd.n278 vdd.t418 0.7285
R3177 vdd.n210 vdd.t300 0.7285
R3178 vdd.n210 vdd.t452 0.7285
R3179 vdd.n142 vdd.t230 0.7285
R3180 vdd.n142 vdd.t442 0.7285
R3181 vdd.n74 vdd.t136 0.7285
R3182 vdd.n74 vdd.t450 0.7285
R3183 vdd.n419 vdd.t492 0.7285
R3184 vdd.n419 vdd.t256 0.7285
R3185 vdd.n435 vdd.t194 0.7285
R3186 vdd.n435 vdd.t101 0.7285
R3187 vdd.n430 vdd.t146 0.7285
R3188 vdd.n430 vdd.t11 0.7285
R3189 vdd.n453 vdd.t258 0.7285
R3190 vdd.n453 vdd.t490 0.7285
R3191 vdd.n459 vdd.t95 0.7285
R3192 vdd.n459 vdd.t1 0.7285
R3193 vdd.n447 vdd.t312 0.7285
R3194 vdd.n447 vdd.t119 0.7285
R3195 vdd.n24 vdd.t65 0.7285
R3196 vdd.n24 vdd.t308 0.7285
R3197 vdd.n18 vdd.t416 0.7285
R3198 vdd.n18 vdd.t214 0.7285
R3199 vdd.n31 vdd.t310 0.7285
R3200 vdd.n31 vdd.t424 0.7285
R3201 vdd.n1 vdd.t504 0.7285
R3202 vdd.n1 vdd.t67 0.7285
R3203 vdd.n12 vdd.t306 0.7285
R3204 vdd.n12 vdd.t390 0.7285
R3205 vdd.n7 vdd.t270 0.7285
R3206 vdd.n7 vdd.t170 0.7285
R3207 vdd.n376 dffrs_1.nand3_0.C 0.717607
R3208 vdd.n308 dffrs_2.nand3_0.C 0.717607
R3209 vdd.n240 dffrs_3.nand3_0.C 0.717607
R3210 vdd.n172 dffrs_4.nand3_0.C 0.717607
R3211 vdd.n104 dffrs_5.nand3_0.C 0.717607
R3212 vdd.n428 dffrs_0.nand3_0.C 0.717607
R3213 vdd.n486 vdd.n465 0.403945
R3214 vdd.n58 vdd.n37 0.400984
R3215 dffrs_13.resetb vdd.n446 0.136036
R3216 vdd.n37 vdd.n0 0.0817571
R3217 vdd.n373 dffrs_1.nand3_2.C 0.0455
R3218 vdd.n305 dffrs_2.nand3_2.C 0.0455
R3219 vdd.n237 dffrs_3.nand3_2.C 0.0455
R3220 vdd.n169 dffrs_4.nand3_2.C 0.0455
R3221 vdd.n101 dffrs_5.nand3_2.C 0.0455
R3222 vdd.n425 dffrs_0.nand3_2.C 0.0455
R3223 vdd.n442 dffrs_13.nand3_7.A 0.0455
R3224 dffrs_1.nand3_0.C vdd.n375 0.0374643
R3225 dffrs_2.nand3_0.C vdd.n307 0.0374643
R3226 dffrs_3.nand3_0.C vdd.n239 0.0374643
R3227 dffrs_4.nand3_0.C vdd.n171 0.0374643
R3228 dffrs_5.nand3_0.C vdd.n103 0.0374643
R3229 dffrs_0.nand3_0.C vdd.n427 0.0374643
R3230 vdd.n23 vdd.n17 0.0373206
R3231 vdd.n458 vdd.n452 0.0339767
R3232 vdd.n376 dffrs_1.setb 0.032
R3233 vdd.n308 dffrs_2.setb 0.032
R3234 vdd.n240 dffrs_3.setb 0.032
R3235 vdd.n172 dffrs_4.setb 0.032
R3236 vdd.n104 dffrs_5.setb 0.032
R3237 vdd.n428 dffrs_0.setb 0.032
R3238 vdd.n465 vdd.n440 0.0316083
R3239 vdd.n30 vdd.n29 0.0286958
R3240 vdd.n440 vdd.n429 0.0192652
R3241 vdd.n36 vdd.n30 0.0113078
R3242 vdd.n126 vdd.n105 0.00505026
R3243 vdd.n262 vdd.n241 0.00505026
R3244 vdd.n330 vdd.n309 0.00505026
R3245 vdd.n398 vdd.n377 0.00505026
R3246 vdd.n17 vdd.n6 0.00441736
R3247 vdd.n105 vdd.n99 0.00430496
R3248 vdd.n173 vdd.n167 0.00430496
R3249 vdd.n241 vdd.n235 0.00430496
R3250 vdd.n309 vdd.n303 0.00430496
R3251 vdd.n377 vdd.n371 0.00430496
R3252 vdd.n99 dffrs_5.vdd 0.00349428
R3253 vdd.n167 dffrs_4.vdd 0.00349428
R3254 vdd.n235 dffrs_3.vdd 0.00349428
R3255 vdd.n303 dffrs_2.vdd 0.00349428
R3256 vdd.n371 dffrs_1.vdd 0.00349428
R3257 dffrs_0.vdd vdd.n486 0.00349428
R3258 vdd.n194 vdd 0.00312817
R3259 vdd.n465 vdd.n464 0.00285324
R3260 vdd vdd.n173 0.00242209
R3261 dffrs_5.vdd vdd.n58 0.00236325
R3262 dffrs_4.vdd vdd.n126 0.00236325
R3263 dffrs_3.vdd vdd.n194 0.00236325
R3264 dffrs_2.vdd vdd.n262 0.00236325
R3265 dffrs_1.vdd vdd.n330 0.00236325
R3266 dffrs_0.vdd vdd.n398 0.00236325
R3267 vdd.n29 vdd.n23 0.000517689
R3268 vdd.n464 vdd.n458 0.000515182
R3269 dffrs_5.nand3_6.C.n1 dffrs_5.nand3_6.C.t7 41.0041
R3270 dffrs_5.nand3_6.C.n0 dffrs_5.nand3_6.C.t5 40.8177
R3271 dffrs_5.nand3_6.C.n3 dffrs_5.nand3_6.C.t6 40.6313
R3272 dffrs_5.nand3_6.C.n3 dffrs_5.nand3_6.C.t9 27.3166
R3273 dffrs_5.nand3_6.C.n0 dffrs_5.nand3_6.C.t8 27.1302
R3274 dffrs_5.nand3_6.C.n1 dffrs_5.nand3_6.C.t4 26.9438
R3275 dffrs_5.nand3_6.C.n9 dffrs_5.nand3_6.C.t1 10.0473
R3276 dffrs_5.nand3_6.C.n5 dffrs_5.nand3_6.C.n4 9.90747
R3277 dffrs_5.nand3_6.C.n5 dffrs_5.nand3_6.C.n2 9.90116
R3278 dffrs_5.nand3_6.C.n8 dffrs_5.nand3_6.C.t2 6.51042
R3279 dffrs_5.nand3_6.C.n8 dffrs_5.nand3_6.C.n7 6.04952
R3280 dffrs_5.nand3_6.C.n2 dffrs_5.nand3_6.C.n1 5.7305
R3281 dffrs_5.nand3_2.B dffrs_5.nand3_6.C.n0 5.47979
R3282 dffrs_5.nand3_6.C.n4 dffrs_5.nand3_6.C.n3 5.13907
R3283 dffrs_5.nand3_1.Z dffrs_5.nand3_6.C.n9 4.72925
R3284 dffrs_5.nand3_6.C.n6 dffrs_5.nand3_6.C.n5 4.5005
R3285 dffrs_5.nand3_6.C.n9 dffrs_5.nand3_6.C.n8 0.732092
R3286 dffrs_5.nand3_6.C.n7 dffrs_5.nand3_6.C.t3 0.7285
R3287 dffrs_5.nand3_6.C.n7 dffrs_5.nand3_6.C.t0 0.7285
R3288 dffrs_5.nand3_1.Z dffrs_5.nand3_6.C.n6 0.449758
R3289 dffrs_5.nand3_6.C.n6 dffrs_5.nand3_2.B 0.166901
R3290 dffrs_5.nand3_6.C.n2 dffrs_5.nand3_0.A 0.0455
R3291 dffrs_5.nand3_6.C.n4 dffrs_5.nand3_6.C 0.0455
R3292 dffrs_5.nand3_1.C.n0 dffrs_5.nand3_1.C.t5 40.6313
R3293 dffrs_5.nand3_1.C.n0 dffrs_5.nand3_1.C.t4 27.3166
R3294 dffrs_5.nand3_0.Z dffrs_5.nand3_1.C.n1 14.2854
R3295 dffrs_5.nand3_1.C.n4 dffrs_5.nand3_1.C.t1 10.0473
R3296 dffrs_5.nand3_1.C.n3 dffrs_5.nand3_1.C.t0 6.51042
R3297 dffrs_5.nand3_1.C.n3 dffrs_5.nand3_1.C.n2 6.04952
R3298 dffrs_5.nand3_1.C.n1 dffrs_5.nand3_1.C.n0 5.13907
R3299 dffrs_5.nand3_0.Z dffrs_5.nand3_1.C.n4 4.72925
R3300 dffrs_5.nand3_1.C.n4 dffrs_5.nand3_1.C.n3 0.732092
R3301 dffrs_5.nand3_1.C.n2 dffrs_5.nand3_1.C.t3 0.7285
R3302 dffrs_5.nand3_1.C.n2 dffrs_5.nand3_1.C.t2 0.7285
R3303 dffrs_5.nand3_1.C.n1 dffrs_5.nand3_1.C 0.0455
R3304 dffrs_8.nand3_8.C.n0 dffrs_8.nand3_8.C.t7 40.8177
R3305 dffrs_8.nand3_8.C.n1 dffrs_8.nand3_8.C.t5 40.6313
R3306 dffrs_8.nand3_8.C.n1 dffrs_8.nand3_8.C.t6 27.3166
R3307 dffrs_8.nand3_8.C.n0 dffrs_8.nand3_8.C.t4 27.1302
R3308 dffrs_8.nand3_8.C.n3 dffrs_8.nand3_8.C.n2 14.119
R3309 dffrs_8.nand3_8.C.n6 dffrs_8.nand3_8.C.t3 10.0473
R3310 dffrs_8.nand3_8.C.n5 dffrs_8.nand3_8.C.t2 6.51042
R3311 dffrs_8.nand3_8.C.n5 dffrs_8.nand3_8.C.n4 6.04952
R3312 dffrs_8.nand3_7.B dffrs_8.nand3_8.C.n0 5.47979
R3313 dffrs_8.nand3_8.C.n2 dffrs_8.nand3_8.C.n1 5.13907
R3314 dffrs_8.nand3_6.Z dffrs_8.nand3_8.C.n6 4.72925
R3315 dffrs_8.nand3_8.C.n6 dffrs_8.nand3_8.C.n5 0.732092
R3316 dffrs_8.nand3_8.C.n4 dffrs_8.nand3_8.C.t0 0.7285
R3317 dffrs_8.nand3_8.C.n4 dffrs_8.nand3_8.C.t1 0.7285
R3318 dffrs_8.nand3_8.C.n3 dffrs_8.nand3_7.B 0.438233
R3319 dffrs_8.nand3_6.Z dffrs_8.nand3_8.C.n3 0.166901
R3320 dffrs_8.nand3_8.C.n2 dffrs_8.nand3_8.C 0.0455
R3321 dffrs_10.nand3_8.C.n0 dffrs_10.nand3_8.C.t4 40.8177
R3322 dffrs_10.nand3_8.C.n1 dffrs_10.nand3_8.C.t6 40.6313
R3323 dffrs_10.nand3_8.C.n1 dffrs_10.nand3_8.C.t7 27.3166
R3324 dffrs_10.nand3_8.C.n0 dffrs_10.nand3_8.C.t5 27.1302
R3325 dffrs_10.nand3_8.C.n3 dffrs_10.nand3_8.C.n2 14.119
R3326 dffrs_10.nand3_8.C.n6 dffrs_10.nand3_8.C.t1 10.0473
R3327 dffrs_10.nand3_8.C.n5 dffrs_10.nand3_8.C.t0 6.51042
R3328 dffrs_10.nand3_8.C.n5 dffrs_10.nand3_8.C.n4 6.04952
R3329 dffrs_10.nand3_7.B dffrs_10.nand3_8.C.n0 5.47979
R3330 dffrs_10.nand3_8.C.n2 dffrs_10.nand3_8.C.n1 5.13907
R3331 dffrs_10.nand3_6.Z dffrs_10.nand3_8.C.n6 4.72925
R3332 dffrs_10.nand3_8.C.n6 dffrs_10.nand3_8.C.n5 0.732092
R3333 dffrs_10.nand3_8.C.n4 dffrs_10.nand3_8.C.t3 0.7285
R3334 dffrs_10.nand3_8.C.n4 dffrs_10.nand3_8.C.t2 0.7285
R3335 dffrs_10.nand3_8.C.n3 dffrs_10.nand3_7.B 0.438233
R3336 dffrs_10.nand3_6.Z dffrs_10.nand3_8.C.n3 0.166901
R3337 dffrs_10.nand3_8.C.n2 dffrs_10.nand3_8.C 0.0455
R3338 dffrs_12.Q.n5 dffrs_11.clk 44.4671
R3339 dffrs_12.Q.n0 dffrs_12.Q.t5 41.0041
R3340 dffrs_12.Q.n1 dffrs_12.Q.t4 40.8177
R3341 dffrs_12.Q.n3 dffrs_12.Q.t8 40.6313
R3342 dffrs_12.Q.n3 dffrs_12.Q.t9 27.3166
R3343 dffrs_12.Q.n1 dffrs_12.Q.t6 27.1302
R3344 dffrs_12.Q.n0 dffrs_12.Q.t7 26.9438
R3345 dffrs_12.Q.n5 dffrs_12.Q.n4 14.0582
R3346 dffrs_12.Q.n8 dffrs_12.Q.t2 10.0473
R3347 dffrs_12.Q.n7 dffrs_12.Q.t1 6.51042
R3348 dffrs_12.Q.n7 dffrs_12.Q.n6 6.04952
R3349 dffrs_11.nand3_1.A dffrs_12.Q.n0 5.7755
R3350 dffrs_11.nand3_6.B dffrs_12.Q.n1 5.47979
R3351 dffrs_12.Q.n4 dffrs_12.Q.n3 5.13907
R3352 dffrs_12.nand3_2.Z dffrs_12.Q.n8 4.72925
R3353 dffrs_12.Q.n2 dffrs_11.nand3_6.B 2.17818
R3354 dffrs_12.Q.n2 dffrs_11.nand3_1.A 1.34729
R3355 dffrs_12.Q.n8 dffrs_12.Q.n7 0.732092
R3356 dffrs_12.Q.n6 dffrs_12.Q.t0 0.7285
R3357 dffrs_12.Q.n6 dffrs_12.Q.t3 0.7285
R3358 dffrs_11.clk dffrs_12.Q.n2 0.610571
R3359 dffrs_12.nand3_2.Z dffrs_12.Q.n5 0.166901
R3360 dffrs_12.Q.n4 dffrs_12.nand3_7.C 0.0455
R3361 dffrs_11.nand3_8.C.n0 dffrs_11.nand3_8.C.t6 40.8177
R3362 dffrs_11.nand3_8.C.n1 dffrs_11.nand3_8.C.t4 40.6313
R3363 dffrs_11.nand3_8.C.n1 dffrs_11.nand3_8.C.t5 27.3166
R3364 dffrs_11.nand3_8.C.n0 dffrs_11.nand3_8.C.t7 27.1302
R3365 dffrs_11.nand3_8.C.n3 dffrs_11.nand3_8.C.n2 14.119
R3366 dffrs_11.nand3_8.C.n6 dffrs_11.nand3_8.C.t2 10.0473
R3367 dffrs_11.nand3_8.C.n5 dffrs_11.nand3_8.C.t3 6.51042
R3368 dffrs_11.nand3_8.C.n5 dffrs_11.nand3_8.C.n4 6.04952
R3369 dffrs_11.nand3_7.B dffrs_11.nand3_8.C.n0 5.47979
R3370 dffrs_11.nand3_8.C.n2 dffrs_11.nand3_8.C.n1 5.13907
R3371 dffrs_11.nand3_6.Z dffrs_11.nand3_8.C.n6 4.72925
R3372 dffrs_11.nand3_8.C.n6 dffrs_11.nand3_8.C.n5 0.732092
R3373 dffrs_11.nand3_8.C.n4 dffrs_11.nand3_8.C.t0 0.7285
R3374 dffrs_11.nand3_8.C.n4 dffrs_11.nand3_8.C.t1 0.7285
R3375 dffrs_11.nand3_8.C.n3 dffrs_11.nand3_7.B 0.438233
R3376 dffrs_11.nand3_6.Z dffrs_11.nand3_8.C.n3 0.166901
R3377 dffrs_11.nand3_8.C.n2 dffrs_11.nand3_8.C 0.0455
R3378 dffrs_1.nand3_1.C.n0 dffrs_1.nand3_1.C.t5 40.6313
R3379 dffrs_1.nand3_1.C.n0 dffrs_1.nand3_1.C.t4 27.3166
R3380 dffrs_1.nand3_0.Z dffrs_1.nand3_1.C.n1 14.2854
R3381 dffrs_1.nand3_1.C.n4 dffrs_1.nand3_1.C.t0 10.0473
R3382 dffrs_1.nand3_1.C.n3 dffrs_1.nand3_1.C.t3 6.51042
R3383 dffrs_1.nand3_1.C.n3 dffrs_1.nand3_1.C.n2 6.04952
R3384 dffrs_1.nand3_1.C.n1 dffrs_1.nand3_1.C.n0 5.13907
R3385 dffrs_1.nand3_0.Z dffrs_1.nand3_1.C.n4 4.72925
R3386 dffrs_1.nand3_1.C.n4 dffrs_1.nand3_1.C.n3 0.732092
R3387 dffrs_1.nand3_1.C.n2 dffrs_1.nand3_1.C.t2 0.7285
R3388 dffrs_1.nand3_1.C.n2 dffrs_1.nand3_1.C.t1 0.7285
R3389 dffrs_1.nand3_1.C.n1 dffrs_1.nand3_1.C 0.0455
R3390 dffrs_2.Qb.n0 dffrs_2.Qb.t9 41.0041
R3391 dffrs_2.Qb.n4 dffrs_2.Qb.t7 40.6313
R3392 dffrs_2.Qb.n2 dffrs_2.Qb.t4 40.6313
R3393 dffrs_2.Qb dffrs_9.setb 28.021
R3394 dffrs_2.Qb.n4 dffrs_2.Qb.t8 27.3166
R3395 dffrs_2.Qb.n2 dffrs_2.Qb.t5 27.3166
R3396 dffrs_2.Qb.n0 dffrs_2.Qb.t6 26.9438
R3397 dffrs_2.Qb.n9 dffrs_2.Qb.t2 10.0473
R3398 dffrs_2.Qb.n6 dffrs_2.Qb.n1 9.84255
R3399 dffrs_2.Qb.n5 dffrs_2.Qb.n3 9.22229
R3400 dffrs_2.Qb.n8 dffrs_2.Qb.t3 6.51042
R3401 dffrs_2.Qb.n8 dffrs_2.Qb.n7 6.04952
R3402 dffrs_2.Qb.n1 dffrs_2.Qb.n0 5.7305
R3403 dffrs_2.Qb.n5 dffrs_2.Qb.n4 5.14711
R3404 dffrs_2.Qb.n3 dffrs_2.Qb.n2 5.13907
R3405 dffrs_2.nand3_7.Z dffrs_2.Qb.n6 4.94976
R3406 dffrs_2.nand3_7.Z dffrs_2.Qb.n9 4.72925
R3407 dffrs_9.setb dffrs_9.nand3_0.C 0.784786
R3408 dffrs_2.Qb.n9 dffrs_2.Qb.n8 0.732092
R3409 dffrs_2.Qb.n7 dffrs_2.Qb.t0 0.7285
R3410 dffrs_2.Qb.n7 dffrs_2.Qb.t1 0.7285
R3411 dffrs_2.Qb.n6 dffrs_2.Qb 0.175225
R3412 dffrs_2.Qb.n1 dffrs_2.nand3_2.A 0.0455
R3413 dffrs_2.Qb.n3 dffrs_9.nand3_2.C 0.0455
R3414 dffrs_9.nand3_0.C dffrs_2.Qb.n5 0.0374643
R3415 d2.n0 d2.t4 41.0041
R3416 d2.n1 d2.t6 40.8177
R3417 d2.n4 d2.t5 40.6313
R3418 d2.n3 dffrs_8.clk 34.1594
R3419 d2.n4 d2.t8 27.3166
R3420 d2.n1 d2.t9 27.1302
R3421 d2.n0 d2.t7 26.9438
R3422 d2.n6 d2.n5 14.0582
R3423 d2.n6 d2.n3 12.0118
R3424 d2.n9 d2.t0 10.0473
R3425 d2.n8 d2.t1 6.51042
R3426 d2.n8 d2.n7 6.04952
R3427 dffrs_8.nand3_1.A d2.n0 5.7755
R3428 dffrs_8.nand3_6.B d2.n1 5.47979
R3429 d2.n5 d2.n4 5.13907
R3430 dffrs_9.nand3_2.Z d2.n9 4.72925
R3431 d2.n2 dffrs_8.nand3_6.B 2.17818
R3432 d2.n2 dffrs_8.nand3_1.A 1.34729
R3433 d2.n9 d2.n8 0.732092
R3434 d2.n7 d2.t3 0.7285
R3435 d2.n7 d2.t2 0.7285
R3436 d2.n3 d2 0.698
R3437 dffrs_8.clk d2.n2 0.610571
R3438 dffrs_9.nand3_2.Z d2.n6 0.166901
R3439 d2.n5 dffrs_9.nand3_7.C 0.0455
R3440 dffrs_9.nand3_6.C.n1 dffrs_9.nand3_6.C.t9 41.0041
R3441 dffrs_9.nand3_6.C.n0 dffrs_9.nand3_6.C.t8 40.8177
R3442 dffrs_9.nand3_6.C.n3 dffrs_9.nand3_6.C.t5 40.6313
R3443 dffrs_9.nand3_6.C.n3 dffrs_9.nand3_6.C.t7 27.3166
R3444 dffrs_9.nand3_6.C.n0 dffrs_9.nand3_6.C.t4 27.1302
R3445 dffrs_9.nand3_6.C.n1 dffrs_9.nand3_6.C.t6 26.9438
R3446 dffrs_9.nand3_6.C.n9 dffrs_9.nand3_6.C.t2 10.0473
R3447 dffrs_9.nand3_6.C.n5 dffrs_9.nand3_6.C.n4 9.90747
R3448 dffrs_9.nand3_6.C.n5 dffrs_9.nand3_6.C.n2 9.90116
R3449 dffrs_9.nand3_6.C.n8 dffrs_9.nand3_6.C.t1 6.51042
R3450 dffrs_9.nand3_6.C.n8 dffrs_9.nand3_6.C.n7 6.04952
R3451 dffrs_9.nand3_6.C.n2 dffrs_9.nand3_6.C.n1 5.7305
R3452 dffrs_9.nand3_2.B dffrs_9.nand3_6.C.n0 5.47979
R3453 dffrs_9.nand3_6.C.n4 dffrs_9.nand3_6.C.n3 5.13907
R3454 dffrs_9.nand3_1.Z dffrs_9.nand3_6.C.n9 4.72925
R3455 dffrs_9.nand3_6.C.n6 dffrs_9.nand3_6.C.n5 4.5005
R3456 dffrs_9.nand3_6.C.n9 dffrs_9.nand3_6.C.n8 0.732092
R3457 dffrs_9.nand3_6.C.n7 dffrs_9.nand3_6.C.t3 0.7285
R3458 dffrs_9.nand3_6.C.n7 dffrs_9.nand3_6.C.t0 0.7285
R3459 dffrs_9.nand3_1.Z dffrs_9.nand3_6.C.n6 0.449758
R3460 dffrs_9.nand3_6.C.n6 dffrs_9.nand3_2.B 0.166901
R3461 dffrs_9.nand3_6.C.n2 dffrs_9.nand3_0.A 0.0455
R3462 dffrs_9.nand3_6.C.n4 dffrs_9.nand3_6.C 0.0455
R3463 d0.n0 d0.t8 41.0041
R3464 d0.n1 d0.t6 40.8177
R3465 d0.n4 d0.t5 40.6313
R3466 d0.n3 dffrs_10.clk 33.5936
R3467 d0.n4 d0.t7 27.3166
R3468 d0.n1 d0.t9 27.1302
R3469 d0.n0 d0.t4 26.9438
R3470 d0.n6 d0.n5 14.0582
R3471 d0.n6 d0.n3 11.4461
R3472 d0.n9 d0.t1 10.0473
R3473 d0.n8 d0.t0 6.51042
R3474 d0.n8 d0.n7 6.04952
R3475 dffrs_10.nand3_1.A d0.n0 5.7755
R3476 dffrs_10.nand3_6.B d0.n1 5.47979
R3477 d0.n5 d0.n4 5.13907
R3478 dffrs_11.nand3_2.Z d0.n9 4.72925
R3479 d0.n2 dffrs_10.nand3_6.B 2.17818
R3480 d0.n2 dffrs_10.nand3_1.A 1.34729
R3481 d0.n3 d0 1.26371
R3482 d0.n9 d0.n8 0.732092
R3483 d0.n7 d0.t3 0.7285
R3484 d0.n7 d0.t2 0.7285
R3485 dffrs_10.clk d0.n2 0.610571
R3486 dffrs_11.nand3_2.Z d0.n6 0.166901
R3487 d0.n5 dffrs_11.nand3_7.C 0.0455
R3488 dffrs_10.nand3_6.C.n1 dffrs_10.nand3_6.C.t5 41.0041
R3489 dffrs_10.nand3_6.C.n0 dffrs_10.nand3_6.C.t9 40.8177
R3490 dffrs_10.nand3_6.C.n3 dffrs_10.nand3_6.C.t8 40.6313
R3491 dffrs_10.nand3_6.C.n3 dffrs_10.nand3_6.C.t4 27.3166
R3492 dffrs_10.nand3_6.C.n0 dffrs_10.nand3_6.C.t6 27.1302
R3493 dffrs_10.nand3_6.C.n1 dffrs_10.nand3_6.C.t7 26.9438
R3494 dffrs_10.nand3_6.C.n9 dffrs_10.nand3_6.C.t1 10.0473
R3495 dffrs_10.nand3_6.C.n5 dffrs_10.nand3_6.C.n4 9.90747
R3496 dffrs_10.nand3_6.C.n5 dffrs_10.nand3_6.C.n2 9.90116
R3497 dffrs_10.nand3_6.C.n8 dffrs_10.nand3_6.C.t2 6.51042
R3498 dffrs_10.nand3_6.C.n8 dffrs_10.nand3_6.C.n7 6.04952
R3499 dffrs_10.nand3_6.C.n2 dffrs_10.nand3_6.C.n1 5.7305
R3500 dffrs_10.nand3_2.B dffrs_10.nand3_6.C.n0 5.47979
R3501 dffrs_10.nand3_6.C.n4 dffrs_10.nand3_6.C.n3 5.13907
R3502 dffrs_10.nand3_1.Z dffrs_10.nand3_6.C.n9 4.72925
R3503 dffrs_10.nand3_6.C.n6 dffrs_10.nand3_6.C.n5 4.5005
R3504 dffrs_10.nand3_6.C.n9 dffrs_10.nand3_6.C.n8 0.732092
R3505 dffrs_10.nand3_6.C.n7 dffrs_10.nand3_6.C.t3 0.7285
R3506 dffrs_10.nand3_6.C.n7 dffrs_10.nand3_6.C.t0 0.7285
R3507 dffrs_10.nand3_1.Z dffrs_10.nand3_6.C.n6 0.449758
R3508 dffrs_10.nand3_6.C.n6 dffrs_10.nand3_2.B 0.166901
R3509 dffrs_10.nand3_6.C.n2 dffrs_10.nand3_0.A 0.0455
R3510 dffrs_10.nand3_6.C.n4 dffrs_10.nand3_6.C 0.0455
R3511 dffrs_3.Qb.n0 dffrs_3.Qb.t8 41.0041
R3512 dffrs_3.Qb.n4 dffrs_3.Qb.t5 40.6313
R3513 dffrs_3.Qb.n2 dffrs_3.Qb.t9 40.6313
R3514 dffrs_3.Qb dffrs_10.setb 28.021
R3515 dffrs_3.Qb.n4 dffrs_3.Qb.t7 27.3166
R3516 dffrs_3.Qb.n2 dffrs_3.Qb.t4 27.3166
R3517 dffrs_3.Qb.n0 dffrs_3.Qb.t6 26.9438
R3518 dffrs_3.Qb.n9 dffrs_3.Qb.t3 10.0473
R3519 dffrs_3.Qb.n6 dffrs_3.Qb.n1 9.84255
R3520 dffrs_3.Qb.n5 dffrs_3.Qb.n3 9.22229
R3521 dffrs_3.Qb.n8 dffrs_3.Qb.t2 6.51042
R3522 dffrs_3.Qb.n8 dffrs_3.Qb.n7 6.04952
R3523 dffrs_3.Qb.n1 dffrs_3.Qb.n0 5.7305
R3524 dffrs_3.Qb.n5 dffrs_3.Qb.n4 5.14711
R3525 dffrs_3.Qb.n3 dffrs_3.Qb.n2 5.13907
R3526 dffrs_3.nand3_7.Z dffrs_3.Qb.n6 4.94976
R3527 dffrs_3.nand3_7.Z dffrs_3.Qb.n9 4.72925
R3528 dffrs_10.setb dffrs_10.nand3_0.C 0.784786
R3529 dffrs_3.Qb.n9 dffrs_3.Qb.n8 0.732092
R3530 dffrs_3.Qb.n7 dffrs_3.Qb.t1 0.7285
R3531 dffrs_3.Qb.n7 dffrs_3.Qb.t0 0.7285
R3532 dffrs_3.Qb.n6 dffrs_3.Qb 0.175225
R3533 dffrs_3.Qb.n1 dffrs_3.nand3_2.A 0.0455
R3534 dffrs_3.Qb.n3 dffrs_10.nand3_2.C 0.0455
R3535 dffrs_10.nand3_0.C dffrs_3.Qb.n5 0.0374643
R3536 dffrs_11.nand3_6.C.n1 dffrs_11.nand3_6.C.t5 41.0041
R3537 dffrs_11.nand3_6.C.n0 dffrs_11.nand3_6.C.t4 40.8177
R3538 dffrs_11.nand3_6.C.n3 dffrs_11.nand3_6.C.t7 40.6313
R3539 dffrs_11.nand3_6.C.n3 dffrs_11.nand3_6.C.t9 27.3166
R3540 dffrs_11.nand3_6.C.n0 dffrs_11.nand3_6.C.t6 27.1302
R3541 dffrs_11.nand3_6.C.n1 dffrs_11.nand3_6.C.t8 26.9438
R3542 dffrs_11.nand3_6.C.n9 dffrs_11.nand3_6.C.t0 10.0473
R3543 dffrs_11.nand3_6.C.n5 dffrs_11.nand3_6.C.n4 9.90747
R3544 dffrs_11.nand3_6.C.n5 dffrs_11.nand3_6.C.n2 9.90116
R3545 dffrs_11.nand3_6.C.n8 dffrs_11.nand3_6.C.t1 6.51042
R3546 dffrs_11.nand3_6.C.n8 dffrs_11.nand3_6.C.n7 6.04952
R3547 dffrs_11.nand3_6.C.n2 dffrs_11.nand3_6.C.n1 5.7305
R3548 dffrs_11.nand3_2.B dffrs_11.nand3_6.C.n0 5.47979
R3549 dffrs_11.nand3_6.C.n4 dffrs_11.nand3_6.C.n3 5.13907
R3550 dffrs_11.nand3_1.Z dffrs_11.nand3_6.C.n9 4.72925
R3551 dffrs_11.nand3_6.C.n6 dffrs_11.nand3_6.C.n5 4.5005
R3552 dffrs_11.nand3_6.C.n9 dffrs_11.nand3_6.C.n8 0.732092
R3553 dffrs_11.nand3_6.C.n7 dffrs_11.nand3_6.C.t3 0.7285
R3554 dffrs_11.nand3_6.C.n7 dffrs_11.nand3_6.C.t2 0.7285
R3555 dffrs_11.nand3_1.Z dffrs_11.nand3_6.C.n6 0.449758
R3556 dffrs_11.nand3_6.C.n6 dffrs_11.nand3_2.B 0.166901
R3557 dffrs_11.nand3_6.C.n2 dffrs_11.nand3_0.A 0.0455
R3558 dffrs_11.nand3_6.C.n4 dffrs_11.nand3_6.C 0.0455
R3559 clk.n3 clk.t19 41.0041
R3560 clk.n7 clk.t9 41.0041
R3561 clk.n11 clk.t3 41.0041
R3562 clk.n15 clk.t2 41.0041
R3563 clk.n19 clk.t26 41.0041
R3564 clk.n23 clk.t16 41.0041
R3565 clk.n0 clk.t13 41.0041
R3566 clk.n4 clk.t8 40.8177
R3567 clk.n8 clk.t27 40.8177
R3568 clk.n12 clk.t22 40.8177
R3569 clk.n16 clk.t10 40.8177
R3570 clk.n20 clk.t4 40.8177
R3571 clk.n24 clk.t7 40.8177
R3572 clk.n1 clk.t5 40.8177
R3573 clk.n4 clk.t21 27.1302
R3574 clk.n8 clk.t12 27.1302
R3575 clk.n12 clk.t6 27.1302
R3576 clk.n16 clk.t24 27.1302
R3577 clk.n20 clk.t17 27.1302
R3578 clk.n24 clk.t20 27.1302
R3579 clk.n1 clk.t18 27.1302
R3580 clk.n3 clk.t1 26.9438
R3581 clk.n7 clk.t23 26.9438
R3582 clk.n11 clk.t15 26.9438
R3583 clk.n15 clk.t14 26.9438
R3584 clk.n19 clk.t11 26.9438
R3585 clk.n23 clk.t0 26.9438
R3586 clk.n0 clk.t25 26.9438
R3587 dffrs_5.clk clk.n26 20.5278
R3588 clk.n14 dffrs_1.clk 16.89
R3589 clk.n18 dffrs_2.clk 16.89
R3590 clk.n22 dffrs_3.clk 16.89
R3591 clk.n26 dffrs_4.clk 16.89
R3592 clk.n10 dffrs_0.clk 16.8417
R3593 clk.n6 dffrs_13.clk 12.2453
R3594 clk.n10 clk.n6 8.1113
R3595 dffrs_13.nand3_1.A clk.n3 5.7755
R3596 dffrs_0.nand3_1.A clk.n7 5.7755
R3597 dffrs_1.nand3_1.A clk.n11 5.7755
R3598 dffrs_2.nand3_1.A clk.n15 5.7755
R3599 dffrs_3.nand3_1.A clk.n19 5.7755
R3600 dffrs_4.nand3_1.A clk.n23 5.7755
R3601 dffrs_5.nand3_1.A clk.n0 5.7755
R3602 dffrs_13.nand3_6.B clk.n4 5.47979
R3603 dffrs_0.nand3_6.B clk.n8 5.47979
R3604 dffrs_1.nand3_6.B clk.n12 5.47979
R3605 dffrs_2.nand3_6.B clk.n16 5.47979
R3606 dffrs_3.nand3_6.B clk.n20 5.47979
R3607 dffrs_4.nand3_6.B clk.n24 5.47979
R3608 dffrs_5.nand3_6.B clk.n1 5.47979
R3609 clk.n26 clk.n22 3.6383
R3610 clk.n22 clk.n18 3.6383
R3611 clk.n18 clk.n14 3.6383
R3612 clk.n14 clk.n10 3.6113
R3613 clk.n5 dffrs_13.nand3_6.B 2.17818
R3614 clk.n9 dffrs_0.nand3_6.B 2.17818
R3615 clk.n13 dffrs_1.nand3_6.B 2.17818
R3616 clk.n17 dffrs_2.nand3_6.B 2.17818
R3617 clk.n21 dffrs_3.nand3_6.B 2.17818
R3618 clk.n25 dffrs_4.nand3_6.B 2.17818
R3619 clk.n2 dffrs_5.nand3_6.B 2.17818
R3620 clk.n5 dffrs_13.nand3_1.A 1.34729
R3621 clk.n9 dffrs_0.nand3_1.A 1.34729
R3622 clk.n13 dffrs_1.nand3_1.A 1.34729
R3623 clk.n17 dffrs_2.nand3_1.A 1.34729
R3624 clk.n21 dffrs_3.nand3_1.A 1.34729
R3625 clk.n25 dffrs_4.nand3_1.A 1.34729
R3626 clk.n2 dffrs_5.nand3_1.A 1.34729
R3627 dffrs_13.clk clk.n5 0.611214
R3628 dffrs_0.clk clk.n9 0.611214
R3629 dffrs_1.clk clk.n13 0.611214
R3630 dffrs_2.clk clk.n17 0.611214
R3631 dffrs_3.clk clk.n21 0.611214
R3632 dffrs_4.clk clk.n25 0.611214
R3633 dffrs_5.clk clk.n2 0.611214
R3634 clk.n6 clk 0.13775
R3635 dffrs_4.nand3_6.C.n1 dffrs_4.nand3_6.C.t7 41.0041
R3636 dffrs_4.nand3_6.C.n0 dffrs_4.nand3_6.C.t5 40.8177
R3637 dffrs_4.nand3_6.C.n3 dffrs_4.nand3_6.C.t9 40.6313
R3638 dffrs_4.nand3_6.C.n3 dffrs_4.nand3_6.C.t6 27.3166
R3639 dffrs_4.nand3_6.C.n0 dffrs_4.nand3_6.C.t8 27.1302
R3640 dffrs_4.nand3_6.C.n1 dffrs_4.nand3_6.C.t4 26.9438
R3641 dffrs_4.nand3_6.C.n9 dffrs_4.nand3_6.C.t1 10.0473
R3642 dffrs_4.nand3_6.C.n5 dffrs_4.nand3_6.C.n4 9.90747
R3643 dffrs_4.nand3_6.C.n5 dffrs_4.nand3_6.C.n2 9.90116
R3644 dffrs_4.nand3_6.C.n8 dffrs_4.nand3_6.C.t0 6.51042
R3645 dffrs_4.nand3_6.C.n8 dffrs_4.nand3_6.C.n7 6.04952
R3646 dffrs_4.nand3_6.C.n2 dffrs_4.nand3_6.C.n1 5.7305
R3647 dffrs_4.nand3_2.B dffrs_4.nand3_6.C.n0 5.47979
R3648 dffrs_4.nand3_6.C.n4 dffrs_4.nand3_6.C.n3 5.13907
R3649 dffrs_4.nand3_1.Z dffrs_4.nand3_6.C.n9 4.72925
R3650 dffrs_4.nand3_6.C.n6 dffrs_4.nand3_6.C.n5 4.5005
R3651 dffrs_4.nand3_6.C.n9 dffrs_4.nand3_6.C.n8 0.732092
R3652 dffrs_4.nand3_6.C.n7 dffrs_4.nand3_6.C.t3 0.7285
R3653 dffrs_4.nand3_6.C.n7 dffrs_4.nand3_6.C.t2 0.7285
R3654 dffrs_4.nand3_1.Z dffrs_4.nand3_6.C.n6 0.449758
R3655 dffrs_4.nand3_6.C.n6 dffrs_4.nand3_2.B 0.166901
R3656 dffrs_4.nand3_6.C.n2 dffrs_4.nand3_0.A 0.0455
R3657 dffrs_4.nand3_6.C.n4 dffrs_4.nand3_6.C 0.0455
R3658 dffrs_1.Qb.n0 dffrs_1.Qb.t5 41.0041
R3659 dffrs_1.Qb.n4 dffrs_1.Qb.t8 40.6313
R3660 dffrs_1.Qb.n2 dffrs_1.Qb.t6 40.6313
R3661 dffrs_1.Qb dffrs_8.setb 28.021
R3662 dffrs_1.Qb.n4 dffrs_1.Qb.t4 27.3166
R3663 dffrs_1.Qb.n2 dffrs_1.Qb.t9 27.3166
R3664 dffrs_1.Qb.n0 dffrs_1.Qb.t7 26.9438
R3665 dffrs_1.Qb.n9 dffrs_1.Qb.t2 10.0473
R3666 dffrs_1.Qb.n6 dffrs_1.Qb.n1 9.84255
R3667 dffrs_1.Qb.n5 dffrs_1.Qb.n3 9.22229
R3668 dffrs_1.Qb.n8 dffrs_1.Qb.t1 6.51042
R3669 dffrs_1.Qb.n8 dffrs_1.Qb.n7 6.04952
R3670 dffrs_1.Qb.n1 dffrs_1.Qb.n0 5.7305
R3671 dffrs_1.Qb.n5 dffrs_1.Qb.n4 5.14711
R3672 dffrs_1.Qb.n3 dffrs_1.Qb.n2 5.13907
R3673 dffrs_1.nand3_7.Z dffrs_1.Qb.n6 4.94976
R3674 dffrs_1.nand3_7.Z dffrs_1.Qb.n9 4.72925
R3675 dffrs_8.setb dffrs_8.nand3_0.C 0.784786
R3676 dffrs_1.Qb.n9 dffrs_1.Qb.n8 0.732092
R3677 dffrs_1.Qb.n7 dffrs_1.Qb.t0 0.7285
R3678 dffrs_1.Qb.n7 dffrs_1.Qb.t3 0.7285
R3679 dffrs_1.Qb.n6 dffrs_1.Qb 0.175225
R3680 dffrs_1.Qb.n1 dffrs_1.nand3_2.A 0.0455
R3681 dffrs_1.Qb.n3 dffrs_8.nand3_2.C 0.0455
R3682 dffrs_8.nand3_0.C dffrs_1.Qb.n5 0.0374643
R3683 dffrs_12.nand3_8.C.n0 dffrs_12.nand3_8.C.t5 40.8177
R3684 dffrs_12.nand3_8.C.n1 dffrs_12.nand3_8.C.t4 40.6313
R3685 dffrs_12.nand3_8.C.n1 dffrs_12.nand3_8.C.t6 27.3166
R3686 dffrs_12.nand3_8.C.n0 dffrs_12.nand3_8.C.t7 27.1302
R3687 dffrs_12.nand3_8.C.n3 dffrs_12.nand3_8.C.n2 14.119
R3688 dffrs_12.nand3_8.C.n6 dffrs_12.nand3_8.C.t0 10.0473
R3689 dffrs_12.nand3_8.C.n5 dffrs_12.nand3_8.C.t1 6.51042
R3690 dffrs_12.nand3_8.C.n5 dffrs_12.nand3_8.C.n4 6.04952
R3691 dffrs_12.nand3_7.B dffrs_12.nand3_8.C.n0 5.47979
R3692 dffrs_12.nand3_8.C.n2 dffrs_12.nand3_8.C.n1 5.13907
R3693 dffrs_12.nand3_6.Z dffrs_12.nand3_8.C.n6 4.72925
R3694 dffrs_12.nand3_8.C.n6 dffrs_12.nand3_8.C.n5 0.732092
R3695 dffrs_12.nand3_8.C.n4 dffrs_12.nand3_8.C.t2 0.7285
R3696 dffrs_12.nand3_8.C.n4 dffrs_12.nand3_8.C.t3 0.7285
R3697 dffrs_12.nand3_8.C.n3 dffrs_12.nand3_7.B 0.438233
R3698 dffrs_12.nand3_6.Z dffrs_12.nand3_8.C.n3 0.166901
R3699 dffrs_12.nand3_8.C.n2 dffrs_12.nand3_8.C 0.0455
R3700 dffrs_14.nand3_6.C.n1 dffrs_14.nand3_6.C.t6 41.0041
R3701 dffrs_14.nand3_6.C.n0 dffrs_14.nand3_6.C.t8 40.8177
R3702 dffrs_14.nand3_6.C.n3 dffrs_14.nand3_6.C.t5 40.6313
R3703 dffrs_14.nand3_6.C.n3 dffrs_14.nand3_6.C.t7 27.3166
R3704 dffrs_14.nand3_6.C.n0 dffrs_14.nand3_6.C.t4 27.1302
R3705 dffrs_14.nand3_6.C.n1 dffrs_14.nand3_6.C.t9 26.9438
R3706 dffrs_14.nand3_6.C.n9 dffrs_14.nand3_6.C.t1 10.0473
R3707 dffrs_14.nand3_6.C.n5 dffrs_14.nand3_6.C.n4 9.90747
R3708 dffrs_14.nand3_6.C.n5 dffrs_14.nand3_6.C.n2 9.90116
R3709 dffrs_14.nand3_6.C.n8 dffrs_14.nand3_6.C.t2 6.51042
R3710 dffrs_14.nand3_6.C.n8 dffrs_14.nand3_6.C.n7 6.04952
R3711 dffrs_14.nand3_6.C.n2 dffrs_14.nand3_6.C.n1 5.7305
R3712 dffrs_14.nand3_2.B dffrs_14.nand3_6.C.n0 5.47979
R3713 dffrs_14.nand3_6.C.n4 dffrs_14.nand3_6.C.n3 5.13907
R3714 dffrs_14.nand3_1.Z dffrs_14.nand3_6.C.n9 4.72925
R3715 dffrs_14.nand3_6.C.n6 dffrs_14.nand3_6.C.n5 4.5005
R3716 dffrs_14.nand3_6.C.n9 dffrs_14.nand3_6.C.n8 0.732092
R3717 dffrs_14.nand3_6.C.n7 dffrs_14.nand3_6.C.t3 0.7285
R3718 dffrs_14.nand3_6.C.n7 dffrs_14.nand3_6.C.t0 0.7285
R3719 dffrs_14.nand3_1.Z dffrs_14.nand3_6.C.n6 0.449758
R3720 dffrs_14.nand3_6.C.n6 dffrs_14.nand3_2.B 0.166901
R3721 dffrs_14.nand3_6.C.n2 dffrs_14.nand3_0.A 0.0455
R3722 dffrs_14.nand3_6.C.n4 dffrs_14.nand3_6.C 0.0455
R3723 dffrs_13.nand3_6.C.n1 dffrs_13.nand3_6.C.t7 41.0041
R3724 dffrs_13.nand3_6.C.n0 dffrs_13.nand3_6.C.t5 40.8177
R3725 dffrs_13.nand3_6.C.n3 dffrs_13.nand3_6.C.t9 40.6313
R3726 dffrs_13.nand3_6.C.n3 dffrs_13.nand3_6.C.t6 27.3166
R3727 dffrs_13.nand3_6.C.n0 dffrs_13.nand3_6.C.t8 27.1302
R3728 dffrs_13.nand3_6.C.n1 dffrs_13.nand3_6.C.t4 26.9438
R3729 dffrs_13.nand3_6.C.n9 dffrs_13.nand3_6.C.t1 10.0473
R3730 dffrs_13.nand3_6.C.n5 dffrs_13.nand3_6.C.n4 9.90747
R3731 dffrs_13.nand3_6.C.n5 dffrs_13.nand3_6.C.n2 9.90116
R3732 dffrs_13.nand3_6.C.n8 dffrs_13.nand3_6.C.t0 6.51042
R3733 dffrs_13.nand3_6.C.n8 dffrs_13.nand3_6.C.n7 6.04952
R3734 dffrs_13.nand3_6.C.n2 dffrs_13.nand3_6.C.n1 5.7305
R3735 dffrs_13.nand3_2.B dffrs_13.nand3_6.C.n0 5.47979
R3736 dffrs_13.nand3_6.C.n4 dffrs_13.nand3_6.C.n3 5.13907
R3737 dffrs_13.nand3_1.Z dffrs_13.nand3_6.C.n9 4.72925
R3738 dffrs_13.nand3_6.C.n6 dffrs_13.nand3_6.C.n5 4.5005
R3739 dffrs_13.nand3_6.C.n9 dffrs_13.nand3_6.C.n8 0.732092
R3740 dffrs_13.nand3_6.C.n7 dffrs_13.nand3_6.C.t2 0.7285
R3741 dffrs_13.nand3_6.C.n7 dffrs_13.nand3_6.C.t3 0.7285
R3742 dffrs_13.nand3_1.Z dffrs_13.nand3_6.C.n6 0.449758
R3743 dffrs_13.nand3_6.C.n6 dffrs_13.nand3_2.B 0.166901
R3744 dffrs_13.nand3_6.C.n2 dffrs_13.nand3_0.A 0.0455
R3745 dffrs_13.nand3_6.C.n4 dffrs_13.nand3_6.C 0.0455
R3746 dffrs_12.nand3_6.C.n1 dffrs_12.nand3_6.C.t5 41.0041
R3747 dffrs_12.nand3_6.C.n0 dffrs_12.nand3_6.C.t4 40.8177
R3748 dffrs_12.nand3_6.C.n3 dffrs_12.nand3_6.C.t8 40.6313
R3749 dffrs_12.nand3_6.C.n3 dffrs_12.nand3_6.C.t9 27.3166
R3750 dffrs_12.nand3_6.C.n0 dffrs_12.nand3_6.C.t6 27.1302
R3751 dffrs_12.nand3_6.C.n1 dffrs_12.nand3_6.C.t7 26.9438
R3752 dffrs_12.nand3_6.C.n9 dffrs_12.nand3_6.C.t1 10.0473
R3753 dffrs_12.nand3_6.C.n5 dffrs_12.nand3_6.C.n4 9.90747
R3754 dffrs_12.nand3_6.C.n5 dffrs_12.nand3_6.C.n2 9.90116
R3755 dffrs_12.nand3_6.C.n8 dffrs_12.nand3_6.C.t2 6.51042
R3756 dffrs_12.nand3_6.C.n8 dffrs_12.nand3_6.C.n7 6.04952
R3757 dffrs_12.nand3_6.C.n2 dffrs_12.nand3_6.C.n1 5.7305
R3758 dffrs_12.nand3_2.B dffrs_12.nand3_6.C.n0 5.47979
R3759 dffrs_12.nand3_6.C.n4 dffrs_12.nand3_6.C.n3 5.13907
R3760 dffrs_12.nand3_1.Z dffrs_12.nand3_6.C.n9 4.72925
R3761 dffrs_12.nand3_6.C.n6 dffrs_12.nand3_6.C.n5 4.5005
R3762 dffrs_12.nand3_6.C.n9 dffrs_12.nand3_6.C.n8 0.732092
R3763 dffrs_12.nand3_6.C.n7 dffrs_12.nand3_6.C.t3 0.7285
R3764 dffrs_12.nand3_6.C.n7 dffrs_12.nand3_6.C.t0 0.7285
R3765 dffrs_12.nand3_1.Z dffrs_12.nand3_6.C.n6 0.449758
R3766 dffrs_12.nand3_6.C.n6 dffrs_12.nand3_2.B 0.166901
R3767 dffrs_12.nand3_6.C.n2 dffrs_12.nand3_0.A 0.0455
R3768 dffrs_12.nand3_6.C.n4 dffrs_12.nand3_6.C 0.0455
R3769 dffrs_4.Qb.n0 dffrs_4.Qb.t8 41.0041
R3770 dffrs_4.Qb.n4 dffrs_4.Qb.t9 40.6313
R3771 dffrs_4.Qb.n2 dffrs_4.Qb.t6 40.6313
R3772 dffrs_4.Qb dffrs_11.setb 28.021
R3773 dffrs_4.Qb.n4 dffrs_4.Qb.t5 27.3166
R3774 dffrs_4.Qb.n2 dffrs_4.Qb.t7 27.3166
R3775 dffrs_4.Qb.n0 dffrs_4.Qb.t4 26.9438
R3776 dffrs_4.Qb.n9 dffrs_4.Qb.t1 10.0473
R3777 dffrs_4.Qb.n6 dffrs_4.Qb.n1 9.84255
R3778 dffrs_4.Qb.n5 dffrs_4.Qb.n3 9.22229
R3779 dffrs_4.Qb.n8 dffrs_4.Qb.t2 6.51042
R3780 dffrs_4.Qb.n8 dffrs_4.Qb.n7 6.04952
R3781 dffrs_4.Qb.n1 dffrs_4.Qb.n0 5.7305
R3782 dffrs_4.Qb.n5 dffrs_4.Qb.n4 5.14711
R3783 dffrs_4.Qb.n3 dffrs_4.Qb.n2 5.13907
R3784 dffrs_4.nand3_7.Z dffrs_4.Qb.n6 4.94976
R3785 dffrs_4.nand3_7.Z dffrs_4.Qb.n9 4.72925
R3786 dffrs_11.setb dffrs_11.nand3_0.C 0.784786
R3787 dffrs_4.Qb.n9 dffrs_4.Qb.n8 0.732092
R3788 dffrs_4.Qb.n7 dffrs_4.Qb.t3 0.7285
R3789 dffrs_4.Qb.n7 dffrs_4.Qb.t0 0.7285
R3790 dffrs_4.Qb.n6 dffrs_4.Qb 0.175225
R3791 dffrs_4.Qb.n1 dffrs_4.nand3_2.A 0.0455
R3792 dffrs_4.Qb.n3 dffrs_11.nand3_2.C 0.0455
R3793 dffrs_11.nand3_0.C dffrs_4.Qb.n5 0.0374643
R3794 dffrs_4.Q.n0 dffrs_4.Q.t5 41.0041
R3795 dffrs_4.Q.n1 dffrs_4.Q.t6 40.6313
R3796 dffrs_4.Q.n1 dffrs_4.Q.t7 27.3166
R3797 dffrs_4.Q.n0 dffrs_4.Q.t4 26.9438
R3798 dffrs_4.Q.n3 dffrs_5.d 17.5382
R3799 dffrs_4.Q.n3 dffrs_4.Q.n2 14.0582
R3800 dffrs_4.Q.n6 dffrs_4.Q.t3 10.0473
R3801 dffrs_4.Q.n5 dffrs_4.Q.t2 6.51042
R3802 dffrs_4.Q.n5 dffrs_4.Q.n4 6.04952
R3803 dffrs_5.nand3_8.A dffrs_4.Q.n0 5.7755
R3804 dffrs_4.Q.n2 dffrs_4.Q.n1 5.13907
R3805 dffrs_4.nand3_2.Z dffrs_4.Q.n6 4.72925
R3806 dffrs_5.d dffrs_5.nand3_8.A 0.784786
R3807 dffrs_4.Q.n6 dffrs_4.Q.n5 0.732092
R3808 dffrs_4.Q.n4 dffrs_4.Q.t0 0.7285
R3809 dffrs_4.Q.n4 dffrs_4.Q.t1 0.7285
R3810 dffrs_4.nand3_2.Z dffrs_4.Q.n3 0.166901
R3811 dffrs_4.Q.n2 dffrs_4.nand3_7.C 0.0455
R3812 comp_in.n1 comp_in.t3 41.0041
R3813 comp_in.n3 comp_in.t7 41.0041
R3814 comp_in.n5 comp_in.t11 41.0041
R3815 comp_in.n7 comp_in.t2 41.0041
R3816 comp_in.n9 comp_in.t4 41.0041
R3817 comp_in.n0 comp_in.t9 41.0041
R3818 comp_in.n1 comp_in.t6 26.9438
R3819 comp_in.n3 comp_in.t10 26.9438
R3820 comp_in.n5 comp_in.t1 26.9438
R3821 comp_in.n7 comp_in.t5 26.9438
R3822 comp_in.n9 comp_in.t8 26.9438
R3823 comp_in.n0 comp_in.t0 26.9438
R3824 dffrs_11.d comp_in.n10 15.3544
R3825 comp_in.n4 dffrs_7.d 11.7166
R3826 comp_in.n6 dffrs_8.d 11.7166
R3827 comp_in.n8 dffrs_9.d 11.7166
R3828 comp_in.n10 dffrs_10.d 11.7166
R3829 comp_in.n2 dffrs_14.d 11.6732
R3830 comp_in.n2 comp_in 7.63655
R3831 dffrs_14.nand3_8.A comp_in.n1 5.7755
R3832 dffrs_7.nand3_8.A comp_in.n3 5.7755
R3833 dffrs_8.nand3_8.A comp_in.n5 5.7755
R3834 dffrs_9.nand3_8.A comp_in.n7 5.7755
R3835 dffrs_10.nand3_8.A comp_in.n9 5.7755
R3836 dffrs_11.nand3_8.A comp_in.n0 5.7755
R3837 comp_in.n10 comp_in.n8 3.6383
R3838 comp_in.n8 comp_in.n6 3.6383
R3839 comp_in.n6 comp_in.n4 3.6383
R3840 comp_in.n4 comp_in.n2 3.6113
R3841 dffrs_14.d dffrs_14.nand3_8.A 0.784786
R3842 dffrs_7.d dffrs_7.nand3_8.A 0.784786
R3843 dffrs_8.d dffrs_8.nand3_8.A 0.784786
R3844 dffrs_9.d dffrs_9.nand3_8.A 0.784786
R3845 dffrs_10.d dffrs_10.nand3_8.A 0.784786
R3846 dffrs_11.d dffrs_11.nand3_8.A 0.784786
R3847 dffrs_7.nand3_8.C.n0 dffrs_7.nand3_8.C.t4 40.8177
R3848 dffrs_7.nand3_8.C.n1 dffrs_7.nand3_8.C.t5 40.6313
R3849 dffrs_7.nand3_8.C.n1 dffrs_7.nand3_8.C.t7 27.3166
R3850 dffrs_7.nand3_8.C.n0 dffrs_7.nand3_8.C.t6 27.1302
R3851 dffrs_7.nand3_8.C.n3 dffrs_7.nand3_8.C.n2 14.119
R3852 dffrs_7.nand3_8.C.n6 dffrs_7.nand3_8.C.t1 10.0473
R3853 dffrs_7.nand3_8.C.n5 dffrs_7.nand3_8.C.t0 6.51042
R3854 dffrs_7.nand3_8.C.n5 dffrs_7.nand3_8.C.n4 6.04952
R3855 dffrs_7.nand3_7.B dffrs_7.nand3_8.C.n0 5.47979
R3856 dffrs_7.nand3_8.C.n2 dffrs_7.nand3_8.C.n1 5.13907
R3857 dffrs_7.nand3_6.Z dffrs_7.nand3_8.C.n6 4.72925
R3858 dffrs_7.nand3_8.C.n6 dffrs_7.nand3_8.C.n5 0.732092
R3859 dffrs_7.nand3_8.C.n4 dffrs_7.nand3_8.C.t2 0.7285
R3860 dffrs_7.nand3_8.C.n4 dffrs_7.nand3_8.C.t3 0.7285
R3861 dffrs_7.nand3_8.C.n3 dffrs_7.nand3_7.B 0.438233
R3862 dffrs_7.nand3_6.Z dffrs_7.nand3_8.C.n3 0.166901
R3863 dffrs_7.nand3_8.C.n2 dffrs_7.nand3_8.C 0.0455
R3864 dffrs_13.Qb.n0 dffrs_13.Qb.t6 41.0041
R3865 dffrs_13.Qb.n4 dffrs_13.Qb.t8 40.6313
R3866 dffrs_13.Qb.n2 dffrs_13.Qb.t7 40.6313
R3867 dffrs_13.Qb dffrs_14.setb 27.9776
R3868 dffrs_13.Qb.n4 dffrs_13.Qb.t5 27.3166
R3869 dffrs_13.Qb.n2 dffrs_13.Qb.t9 27.3166
R3870 dffrs_13.Qb.n0 dffrs_13.Qb.t4 26.9438
R3871 dffrs_13.Qb.n9 dffrs_13.Qb.t2 10.0473
R3872 dffrs_13.Qb.n6 dffrs_13.Qb.n1 9.84255
R3873 dffrs_13.Qb.n5 dffrs_13.Qb.n3 9.22229
R3874 dffrs_13.Qb.n8 dffrs_13.Qb.t1 6.51042
R3875 dffrs_13.Qb.n8 dffrs_13.Qb.n7 6.04952
R3876 dffrs_13.Qb.n1 dffrs_13.Qb.n0 5.7305
R3877 dffrs_13.Qb.n5 dffrs_13.Qb.n4 5.14711
R3878 dffrs_13.Qb.n3 dffrs_13.Qb.n2 5.13907
R3879 dffrs_13.nand3_7.Z dffrs_13.Qb.n6 4.94976
R3880 dffrs_13.nand3_7.Z dffrs_13.Qb.n9 4.72925
R3881 dffrs_14.setb dffrs_14.nand3_0.C 0.784786
R3882 dffrs_13.Qb.n9 dffrs_13.Qb.n8 0.732092
R3883 dffrs_13.Qb.n7 dffrs_13.Qb.t0 0.7285
R3884 dffrs_13.Qb.n7 dffrs_13.Qb.t3 0.7285
R3885 dffrs_13.Qb.n6 dffrs_13.Qb 0.175225
R3886 dffrs_13.Qb.n1 dffrs_13.nand3_2.A 0.0455
R3887 dffrs_13.Qb.n3 dffrs_14.nand3_2.C 0.0455
R3888 dffrs_14.nand3_0.C dffrs_13.Qb.n5 0.0374643
R3889 dffrs_0.d.n0 dffrs_0.d.t4 41.0041
R3890 dffrs_0.d.n1 dffrs_0.d.t5 40.6313
R3891 dffrs_0.d.n1 dffrs_0.d.t7 27.3166
R3892 dffrs_0.d.n0 dffrs_0.d.t6 26.9438
R3893 dffrs_0.d.n3 dffrs_0.d 17.5022
R3894 dffrs_0.d.n3 dffrs_0.d.n2 14.0582
R3895 dffrs_0.d.n6 dffrs_0.d.t0 10.0473
R3896 dffrs_0.d.n5 dffrs_0.d.t1 6.51042
R3897 dffrs_0.d.n5 dffrs_0.d.n4 6.04952
R3898 dffrs_0.nand3_8.A dffrs_0.d.n0 5.7755
R3899 dffrs_0.d.n2 dffrs_0.d.n1 5.13907
R3900 dffrs_13.nand3_2.Z dffrs_0.d.n6 4.72925
R3901 dffrs_0.d dffrs_0.nand3_8.A 0.783821
R3902 dffrs_0.d.n6 dffrs_0.d.n5 0.732092
R3903 dffrs_0.d.n4 dffrs_0.d.t2 0.7285
R3904 dffrs_0.d.n4 dffrs_0.d.t3 0.7285
R3905 dffrs_13.nand3_2.Z dffrs_0.d.n3 0.166901
R3906 dffrs_0.d.n2 dffrs_13.nand3_7.C 0.0455
R3907 dffrs_9.nand3_8.C.n0 dffrs_9.nand3_8.C.t4 40.8177
R3908 dffrs_9.nand3_8.C.n1 dffrs_9.nand3_8.C.t6 40.6313
R3909 dffrs_9.nand3_8.C.n1 dffrs_9.nand3_8.C.t7 27.3166
R3910 dffrs_9.nand3_8.C.n0 dffrs_9.nand3_8.C.t5 27.1302
R3911 dffrs_9.nand3_8.C.n3 dffrs_9.nand3_8.C.n2 14.119
R3912 dffrs_9.nand3_8.C.n6 dffrs_9.nand3_8.C.t1 10.0473
R3913 dffrs_9.nand3_8.C.n5 dffrs_9.nand3_8.C.t0 6.51042
R3914 dffrs_9.nand3_8.C.n5 dffrs_9.nand3_8.C.n4 6.04952
R3915 dffrs_9.nand3_7.B dffrs_9.nand3_8.C.n0 5.47979
R3916 dffrs_9.nand3_8.C.n2 dffrs_9.nand3_8.C.n1 5.13907
R3917 dffrs_9.nand3_6.Z dffrs_9.nand3_8.C.n6 4.72925
R3918 dffrs_9.nand3_8.C.n6 dffrs_9.nand3_8.C.n5 0.732092
R3919 dffrs_9.nand3_8.C.n4 dffrs_9.nand3_8.C.t2 0.7285
R3920 dffrs_9.nand3_8.C.n4 dffrs_9.nand3_8.C.t3 0.7285
R3921 dffrs_9.nand3_8.C.n3 dffrs_9.nand3_7.B 0.438233
R3922 dffrs_9.nand3_6.Z dffrs_9.nand3_8.C.n3 0.166901
R3923 dffrs_9.nand3_8.C.n2 dffrs_9.nand3_8.C 0.0455
R3924 dffrs_0.nand3_6.C.n1 dffrs_0.nand3_6.C.t6 41.0041
R3925 dffrs_0.nand3_6.C.n0 dffrs_0.nand3_6.C.t4 40.8177
R3926 dffrs_0.nand3_6.C.n3 dffrs_0.nand3_6.C.t5 40.6313
R3927 dffrs_0.nand3_6.C.n3 dffrs_0.nand3_6.C.t8 27.3166
R3928 dffrs_0.nand3_6.C.n0 dffrs_0.nand3_6.C.t7 27.1302
R3929 dffrs_0.nand3_6.C.n1 dffrs_0.nand3_6.C.t9 26.9438
R3930 dffrs_0.nand3_6.C.n9 dffrs_0.nand3_6.C.t1 10.0473
R3931 dffrs_0.nand3_6.C.n5 dffrs_0.nand3_6.C.n4 9.90747
R3932 dffrs_0.nand3_6.C.n5 dffrs_0.nand3_6.C.n2 9.90116
R3933 dffrs_0.nand3_6.C.n8 dffrs_0.nand3_6.C.t0 6.51042
R3934 dffrs_0.nand3_6.C.n8 dffrs_0.nand3_6.C.n7 6.04952
R3935 dffrs_0.nand3_6.C.n2 dffrs_0.nand3_6.C.n1 5.7305
R3936 dffrs_0.nand3_2.B dffrs_0.nand3_6.C.n0 5.47979
R3937 dffrs_0.nand3_6.C.n4 dffrs_0.nand3_6.C.n3 5.13907
R3938 dffrs_0.nand3_1.Z dffrs_0.nand3_6.C.n9 4.72925
R3939 dffrs_0.nand3_6.C.n6 dffrs_0.nand3_6.C.n5 4.5005
R3940 dffrs_0.nand3_6.C.n9 dffrs_0.nand3_6.C.n8 0.732092
R3941 dffrs_0.nand3_6.C.n7 dffrs_0.nand3_6.C.t3 0.7285
R3942 dffrs_0.nand3_6.C.n7 dffrs_0.nand3_6.C.t2 0.7285
R3943 dffrs_0.nand3_1.Z dffrs_0.nand3_6.C.n6 0.449758
R3944 dffrs_0.nand3_6.C.n6 dffrs_0.nand3_2.B 0.166901
R3945 dffrs_0.nand3_6.C.n2 dffrs_0.nand3_0.A 0.0455
R3946 dffrs_0.nand3_6.C.n4 dffrs_0.nand3_6.C 0.0455
R3947 dffrs_0.Q.n0 dffrs_0.Q.t6 41.0041
R3948 dffrs_0.Q.n1 dffrs_0.Q.t7 40.6313
R3949 dffrs_0.Q.n1 dffrs_0.Q.t5 27.3166
R3950 dffrs_0.Q.n0 dffrs_0.Q.t4 26.9438
R3951 dffrs_0.Q.n3 dffrs_1.d 17.5382
R3952 dffrs_0.Q.n3 dffrs_0.Q.n2 14.0582
R3953 dffrs_0.Q.n6 dffrs_0.Q.t3 10.0473
R3954 dffrs_0.Q.n5 dffrs_0.Q.t1 6.51042
R3955 dffrs_0.Q.n5 dffrs_0.Q.n4 6.04952
R3956 dffrs_1.nand3_8.A dffrs_0.Q.n0 5.7755
R3957 dffrs_0.Q.n2 dffrs_0.Q.n1 5.13907
R3958 dffrs_0.nand3_2.Z dffrs_0.Q.n6 4.72925
R3959 dffrs_1.d dffrs_1.nand3_8.A 0.784786
R3960 dffrs_0.Q.n6 dffrs_0.Q.n5 0.732092
R3961 dffrs_0.Q.n4 dffrs_0.Q.t2 0.7285
R3962 dffrs_0.Q.n4 dffrs_0.Q.t0 0.7285
R3963 dffrs_0.nand3_2.Z dffrs_0.Q.n3 0.166901
R3964 dffrs_0.Q.n2 dffrs_0.nand3_7.C 0.0455
R3965 d3.n0 d3.t4 41.0041
R3966 d3.n1 d3.t9 40.8177
R3967 d3.n4 d3.t8 40.6313
R3968 d3.n3 dffrs_7.clk 33.3108
R3969 d3.n4 d3.t5 27.3166
R3970 d3.n1 d3.t6 27.1302
R3971 d3.n0 d3.t7 26.9438
R3972 d3.n6 d3.n5 14.0582
R3973 d3.n6 d3.n3 11.1633
R3974 d3.n9 d3.t1 10.0473
R3975 d3.n8 d3.t0 6.51042
R3976 d3.n8 d3.n7 6.04952
R3977 dffrs_7.nand3_1.A d3.n0 5.7755
R3978 dffrs_7.nand3_6.B d3.n1 5.47979
R3979 d3.n5 d3.n4 5.13907
R3980 dffrs_8.nand3_2.Z d3.n9 4.72925
R3981 d3.n2 dffrs_7.nand3_6.B 2.17818
R3982 d3.n3 d3 1.54657
R3983 d3.n2 dffrs_7.nand3_1.A 1.34729
R3984 d3.n9 d3.n8 0.732092
R3985 d3.n7 d3.t2 0.7285
R3986 d3.n7 d3.t3 0.7285
R3987 dffrs_7.clk d3.n2 0.610571
R3988 dffrs_8.nand3_2.Z d3.n6 0.166901
R3989 d3.n5 dffrs_8.nand3_7.C 0.0455
R3990 dffrs_7.nand3_6.C.n1 dffrs_7.nand3_6.C.t7 41.0041
R3991 dffrs_7.nand3_6.C.n0 dffrs_7.nand3_6.C.t4 40.8177
R3992 dffrs_7.nand3_6.C.n3 dffrs_7.nand3_6.C.t9 40.6313
R3993 dffrs_7.nand3_6.C.n3 dffrs_7.nand3_6.C.t5 27.3166
R3994 dffrs_7.nand3_6.C.n0 dffrs_7.nand3_6.C.t6 27.1302
R3995 dffrs_7.nand3_6.C.n1 dffrs_7.nand3_6.C.t8 26.9438
R3996 dffrs_7.nand3_6.C.n9 dffrs_7.nand3_6.C.t1 10.0473
R3997 dffrs_7.nand3_6.C.n5 dffrs_7.nand3_6.C.n4 9.90747
R3998 dffrs_7.nand3_6.C.n5 dffrs_7.nand3_6.C.n2 9.90116
R3999 dffrs_7.nand3_6.C.n8 dffrs_7.nand3_6.C.t0 6.51042
R4000 dffrs_7.nand3_6.C.n8 dffrs_7.nand3_6.C.n7 6.04952
R4001 dffrs_7.nand3_6.C.n2 dffrs_7.nand3_6.C.n1 5.7305
R4002 dffrs_7.nand3_2.B dffrs_7.nand3_6.C.n0 5.47979
R4003 dffrs_7.nand3_6.C.n4 dffrs_7.nand3_6.C.n3 5.13907
R4004 dffrs_7.nand3_1.Z dffrs_7.nand3_6.C.n9 4.72925
R4005 dffrs_7.nand3_6.C.n6 dffrs_7.nand3_6.C.n5 4.5005
R4006 dffrs_7.nand3_6.C.n9 dffrs_7.nand3_6.C.n8 0.732092
R4007 dffrs_7.nand3_6.C.n7 dffrs_7.nand3_6.C.t3 0.7285
R4008 dffrs_7.nand3_6.C.n7 dffrs_7.nand3_6.C.t2 0.7285
R4009 dffrs_7.nand3_1.Z dffrs_7.nand3_6.C.n6 0.449758
R4010 dffrs_7.nand3_6.C.n6 dffrs_7.nand3_2.B 0.166901
R4011 dffrs_7.nand3_6.C.n2 dffrs_7.nand3_0.A 0.0455
R4012 dffrs_7.nand3_6.C.n4 dffrs_7.nand3_6.C 0.0455
R4013 dffrs_5.Q.n0 dffrs_5.Q.t4 40.6313
R4014 dffrs_5.Q.n0 dffrs_5.Q.t5 27.3166
R4015 dffrs_5.nand3_2.Z dffrs_5.Q.n1 14.2246
R4016 dffrs_5.Q.n4 dffrs_5.Q.t3 10.0473
R4017 dffrs_5.Q.n3 dffrs_5.Q.t2 6.51042
R4018 dffrs_5.Q.n3 dffrs_5.Q.n2 6.04952
R4019 dffrs_5.Q.n1 dffrs_5.Q.n0 5.13907
R4020 dffrs_5.nand3_2.Z dffrs_5.Q.n4 4.72925
R4021 dffrs_5.Q.n4 dffrs_5.Q.n3 0.732092
R4022 dffrs_5.Q.n2 dffrs_5.Q.t0 0.7285
R4023 dffrs_5.Q.n2 dffrs_5.Q.t1 0.7285
R4024 dffrs_5.Q.n1 dffrs_5.nand3_7.C 0.0455
R4025 dffrs_2.nand3_6.C.n1 dffrs_2.nand3_6.C.t4 41.0041
R4026 dffrs_2.nand3_6.C.n0 dffrs_2.nand3_6.C.t8 40.8177
R4027 dffrs_2.nand3_6.C.n3 dffrs_2.nand3_6.C.t9 40.6313
R4028 dffrs_2.nand3_6.C.n3 dffrs_2.nand3_6.C.t6 27.3166
R4029 dffrs_2.nand3_6.C.n0 dffrs_2.nand3_6.C.t5 27.1302
R4030 dffrs_2.nand3_6.C.n1 dffrs_2.nand3_6.C.t7 26.9438
R4031 dffrs_2.nand3_6.C.n9 dffrs_2.nand3_6.C.t1 10.0473
R4032 dffrs_2.nand3_6.C.n5 dffrs_2.nand3_6.C.n4 9.90747
R4033 dffrs_2.nand3_6.C.n5 dffrs_2.nand3_6.C.n2 9.90116
R4034 dffrs_2.nand3_6.C.n8 dffrs_2.nand3_6.C.t0 6.51042
R4035 dffrs_2.nand3_6.C.n8 dffrs_2.nand3_6.C.n7 6.04952
R4036 dffrs_2.nand3_6.C.n2 dffrs_2.nand3_6.C.n1 5.7305
R4037 dffrs_2.nand3_2.B dffrs_2.nand3_6.C.n0 5.47979
R4038 dffrs_2.nand3_6.C.n4 dffrs_2.nand3_6.C.n3 5.13907
R4039 dffrs_2.nand3_1.Z dffrs_2.nand3_6.C.n9 4.72925
R4040 dffrs_2.nand3_6.C.n6 dffrs_2.nand3_6.C.n5 4.5005
R4041 dffrs_2.nand3_6.C.n9 dffrs_2.nand3_6.C.n8 0.732092
R4042 dffrs_2.nand3_6.C.n7 dffrs_2.nand3_6.C.t3 0.7285
R4043 dffrs_2.nand3_6.C.n7 dffrs_2.nand3_6.C.t2 0.7285
R4044 dffrs_2.nand3_1.Z dffrs_2.nand3_6.C.n6 0.449758
R4045 dffrs_2.nand3_6.C.n6 dffrs_2.nand3_2.B 0.166901
R4046 dffrs_2.nand3_6.C.n2 dffrs_2.nand3_0.A 0.0455
R4047 dffrs_2.nand3_6.C.n4 dffrs_2.nand3_6.C 0.0455
R4048 dffrs_1.nand3_6.C.n1 dffrs_1.nand3_6.C.t4 41.0041
R4049 dffrs_1.nand3_6.C.n0 dffrs_1.nand3_6.C.t9 40.8177
R4050 dffrs_1.nand3_6.C.n3 dffrs_1.nand3_6.C.t5 40.6313
R4051 dffrs_1.nand3_6.C.n3 dffrs_1.nand3_6.C.t8 27.3166
R4052 dffrs_1.nand3_6.C.n0 dffrs_1.nand3_6.C.t6 27.1302
R4053 dffrs_1.nand3_6.C.n1 dffrs_1.nand3_6.C.t7 26.9438
R4054 dffrs_1.nand3_6.C.n9 dffrs_1.nand3_6.C.t1 10.0473
R4055 dffrs_1.nand3_6.C.n5 dffrs_1.nand3_6.C.n4 9.90747
R4056 dffrs_1.nand3_6.C.n5 dffrs_1.nand3_6.C.n2 9.90116
R4057 dffrs_1.nand3_6.C.n8 dffrs_1.nand3_6.C.t0 6.51042
R4058 dffrs_1.nand3_6.C.n8 dffrs_1.nand3_6.C.n7 6.04952
R4059 dffrs_1.nand3_6.C.n2 dffrs_1.nand3_6.C.n1 5.7305
R4060 dffrs_1.nand3_2.B dffrs_1.nand3_6.C.n0 5.47979
R4061 dffrs_1.nand3_6.C.n4 dffrs_1.nand3_6.C.n3 5.13907
R4062 dffrs_1.nand3_1.Z dffrs_1.nand3_6.C.n9 4.72925
R4063 dffrs_1.nand3_6.C.n6 dffrs_1.nand3_6.C.n5 4.5005
R4064 dffrs_1.nand3_6.C.n9 dffrs_1.nand3_6.C.n8 0.732092
R4065 dffrs_1.nand3_6.C.n7 dffrs_1.nand3_6.C.t3 0.7285
R4066 dffrs_1.nand3_6.C.n7 dffrs_1.nand3_6.C.t2 0.7285
R4067 dffrs_1.nand3_1.Z dffrs_1.nand3_6.C.n6 0.449758
R4068 dffrs_1.nand3_6.C.n6 dffrs_1.nand3_2.B 0.166901
R4069 dffrs_1.nand3_6.C.n2 dffrs_1.nand3_0.A 0.0455
R4070 dffrs_1.nand3_6.C.n4 dffrs_1.nand3_6.C 0.0455
R4071 dffrs_13.nand3_8.C.n0 dffrs_13.nand3_8.C.t5 40.8177
R4072 dffrs_13.nand3_8.C.n1 dffrs_13.nand3_8.C.t7 40.6313
R4073 dffrs_13.nand3_8.C.n1 dffrs_13.nand3_8.C.t4 27.3166
R4074 dffrs_13.nand3_8.C.n0 dffrs_13.nand3_8.C.t6 27.1302
R4075 dffrs_13.nand3_8.C.n3 dffrs_13.nand3_8.C.n2 14.119
R4076 dffrs_13.nand3_8.C.n6 dffrs_13.nand3_8.C.t3 10.0473
R4077 dffrs_13.nand3_8.C.n5 dffrs_13.nand3_8.C.t2 6.51042
R4078 dffrs_13.nand3_8.C.n5 dffrs_13.nand3_8.C.n4 6.04952
R4079 dffrs_13.nand3_7.B dffrs_13.nand3_8.C.n0 5.47979
R4080 dffrs_13.nand3_8.C.n2 dffrs_13.nand3_8.C.n1 5.13907
R4081 dffrs_13.nand3_6.Z dffrs_13.nand3_8.C.n6 4.72925
R4082 dffrs_13.nand3_8.C.n6 dffrs_13.nand3_8.C.n5 0.732092
R4083 dffrs_13.nand3_8.C.n4 dffrs_13.nand3_8.C.t0 0.7285
R4084 dffrs_13.nand3_8.C.n4 dffrs_13.nand3_8.C.t1 0.7285
R4085 dffrs_13.nand3_8.C.n3 dffrs_13.nand3_7.B 0.438233
R4086 dffrs_13.nand3_6.Z dffrs_13.nand3_8.C.n3 0.166901
R4087 dffrs_13.nand3_8.C.n2 dffrs_13.nand3_8.C 0.0455
R4088 dffrs_14.nand3_8.C.n0 dffrs_14.nand3_8.C.t7 40.8177
R4089 dffrs_14.nand3_8.C.n1 dffrs_14.nand3_8.C.t5 40.6313
R4090 dffrs_14.nand3_8.C.n1 dffrs_14.nand3_8.C.t6 27.3166
R4091 dffrs_14.nand3_8.C.n0 dffrs_14.nand3_8.C.t4 27.1302
R4092 dffrs_14.nand3_8.C.n3 dffrs_14.nand3_8.C.n2 14.119
R4093 dffrs_14.nand3_8.C.n6 dffrs_14.nand3_8.C.t2 10.0473
R4094 dffrs_14.nand3_8.C.n5 dffrs_14.nand3_8.C.t3 6.51042
R4095 dffrs_14.nand3_8.C.n5 dffrs_14.nand3_8.C.n4 6.04952
R4096 dffrs_14.nand3_7.B dffrs_14.nand3_8.C.n0 5.47979
R4097 dffrs_14.nand3_8.C.n2 dffrs_14.nand3_8.C.n1 5.13907
R4098 dffrs_14.nand3_6.Z dffrs_14.nand3_8.C.n6 4.72925
R4099 dffrs_14.nand3_8.C.n6 dffrs_14.nand3_8.C.n5 0.732092
R4100 dffrs_14.nand3_8.C.n4 dffrs_14.nand3_8.C.t1 0.7285
R4101 dffrs_14.nand3_8.C.n4 dffrs_14.nand3_8.C.t0 0.7285
R4102 dffrs_14.nand3_8.C.n3 dffrs_14.nand3_7.B 0.438233
R4103 dffrs_14.nand3_6.Z dffrs_14.nand3_8.C.n3 0.166901
R4104 dffrs_14.nand3_8.C.n2 dffrs_14.nand3_8.C 0.0455
R4105 dffrs_0.nand3_8.Z.n0 dffrs_0.nand3_8.Z.t4 41.0041
R4106 dffrs_0.nand3_8.Z.n1 dffrs_0.nand3_8.Z.t5 40.8177
R4107 dffrs_0.nand3_8.Z.n1 dffrs_0.nand3_8.Z.t7 27.1302
R4108 dffrs_0.nand3_8.Z.n0 dffrs_0.nand3_8.Z.t6 26.9438
R4109 dffrs_0.nand3_6.A dffrs_0.nand3_0.B 17.0041
R4110 dffrs_0.nand3_8.Z dffrs_0.nand3_8.Z.n2 14.8493
R4111 dffrs_0.nand3_8.Z.n5 dffrs_0.nand3_8.Z.t2 10.0473
R4112 dffrs_0.nand3_8.Z.n4 dffrs_0.nand3_8.Z.t1 6.51042
R4113 dffrs_0.nand3_8.Z.n4 dffrs_0.nand3_8.Z.n3 6.04952
R4114 dffrs_0.nand3_8.Z.n2 dffrs_0.nand3_8.Z.n0 5.7305
R4115 dffrs_0.nand3_0.B dffrs_0.nand3_8.Z.n1 5.47979
R4116 dffrs_0.nand3_8.Z dffrs_0.nand3_8.Z.n5 4.72925
R4117 dffrs_0.nand3_8.Z.n5 dffrs_0.nand3_8.Z.n4 0.732092
R4118 dffrs_0.nand3_8.Z.n3 dffrs_0.nand3_8.Z.t3 0.7285
R4119 dffrs_0.nand3_8.Z.n3 dffrs_0.nand3_8.Z.t0 0.7285
R4120 dffrs_0.nand3_8.Z.n2 dffrs_0.nand3_6.A 0.0455
R4121 dffrs_2.nand3_1.C.n0 dffrs_2.nand3_1.C.t4 40.6313
R4122 dffrs_2.nand3_1.C.n0 dffrs_2.nand3_1.C.t5 27.3166
R4123 dffrs_2.nand3_0.Z dffrs_2.nand3_1.C.n1 14.2854
R4124 dffrs_2.nand3_1.C.n4 dffrs_2.nand3_1.C.t1 10.0473
R4125 dffrs_2.nand3_1.C.n3 dffrs_2.nand3_1.C.t2 6.51042
R4126 dffrs_2.nand3_1.C.n3 dffrs_2.nand3_1.C.n2 6.04952
R4127 dffrs_2.nand3_1.C.n1 dffrs_2.nand3_1.C.n0 5.13907
R4128 dffrs_2.nand3_0.Z dffrs_2.nand3_1.C.n4 4.72925
R4129 dffrs_2.nand3_1.C.n4 dffrs_2.nand3_1.C.n3 0.732092
R4130 dffrs_2.nand3_1.C.n2 dffrs_2.nand3_1.C.t3 0.7285
R4131 dffrs_2.nand3_1.C.n2 dffrs_2.nand3_1.C.t0 0.7285
R4132 dffrs_2.nand3_1.C.n1 dffrs_2.nand3_1.C 0.0455
R4133 dffrs_3.nand3_8.Z.n0 dffrs_3.nand3_8.Z.t6 41.0041
R4134 dffrs_3.nand3_8.Z.n1 dffrs_3.nand3_8.Z.t5 40.8177
R4135 dffrs_3.nand3_8.Z.n1 dffrs_3.nand3_8.Z.t7 27.1302
R4136 dffrs_3.nand3_8.Z.n0 dffrs_3.nand3_8.Z.t4 26.9438
R4137 dffrs_3.nand3_6.A dffrs_3.nand3_0.B 17.0041
R4138 dffrs_3.nand3_8.Z dffrs_3.nand3_8.Z.n2 14.8493
R4139 dffrs_3.nand3_8.Z.n5 dffrs_3.nand3_8.Z.t2 10.0473
R4140 dffrs_3.nand3_8.Z.n4 dffrs_3.nand3_8.Z.t1 6.51042
R4141 dffrs_3.nand3_8.Z.n4 dffrs_3.nand3_8.Z.n3 6.04952
R4142 dffrs_3.nand3_8.Z.n2 dffrs_3.nand3_8.Z.n0 5.7305
R4143 dffrs_3.nand3_0.B dffrs_3.nand3_8.Z.n1 5.47979
R4144 dffrs_3.nand3_8.Z dffrs_3.nand3_8.Z.n5 4.72925
R4145 dffrs_3.nand3_8.Z.n5 dffrs_3.nand3_8.Z.n4 0.732092
R4146 dffrs_3.nand3_8.Z.n3 dffrs_3.nand3_8.Z.t3 0.7285
R4147 dffrs_3.nand3_8.Z.n3 dffrs_3.nand3_8.Z.t0 0.7285
R4148 dffrs_3.nand3_8.Z.n2 dffrs_3.nand3_6.A 0.0455
R4149 dffrs_5.nand3_8.Z.n0 dffrs_5.nand3_8.Z.t4 41.0041
R4150 dffrs_5.nand3_8.Z.n1 dffrs_5.nand3_8.Z.t5 40.8177
R4151 dffrs_5.nand3_8.Z.n1 dffrs_5.nand3_8.Z.t7 27.1302
R4152 dffrs_5.nand3_8.Z.n0 dffrs_5.nand3_8.Z.t6 26.9438
R4153 dffrs_5.nand3_6.A dffrs_5.nand3_0.B 17.0041
R4154 dffrs_5.nand3_8.Z dffrs_5.nand3_8.Z.n2 14.8493
R4155 dffrs_5.nand3_8.Z.n5 dffrs_5.nand3_8.Z.t1 10.0473
R4156 dffrs_5.nand3_8.Z.n4 dffrs_5.nand3_8.Z.t2 6.51042
R4157 dffrs_5.nand3_8.Z.n4 dffrs_5.nand3_8.Z.n3 6.04952
R4158 dffrs_5.nand3_8.Z.n2 dffrs_5.nand3_8.Z.n0 5.7305
R4159 dffrs_5.nand3_0.B dffrs_5.nand3_8.Z.n1 5.47979
R4160 dffrs_5.nand3_8.Z dffrs_5.nand3_8.Z.n5 4.72925
R4161 dffrs_5.nand3_8.Z.n5 dffrs_5.nand3_8.Z.n4 0.732092
R4162 dffrs_5.nand3_8.Z.n3 dffrs_5.nand3_8.Z.t3 0.7285
R4163 dffrs_5.nand3_8.Z.n3 dffrs_5.nand3_8.Z.t0 0.7285
R4164 dffrs_5.nand3_8.Z.n2 dffrs_5.nand3_6.A 0.0455
R4165 dffrs_0.nand3_8.C.n0 dffrs_0.nand3_8.C.t4 40.8177
R4166 dffrs_0.nand3_8.C.n1 dffrs_0.nand3_8.C.t5 40.6313
R4167 dffrs_0.nand3_8.C.n1 dffrs_0.nand3_8.C.t6 27.3166
R4168 dffrs_0.nand3_8.C.n0 dffrs_0.nand3_8.C.t7 27.1302
R4169 dffrs_0.nand3_8.C.n3 dffrs_0.nand3_8.C.n2 14.119
R4170 dffrs_0.nand3_8.C.n6 dffrs_0.nand3_8.C.t2 10.0473
R4171 dffrs_0.nand3_8.C.n5 dffrs_0.nand3_8.C.t1 6.51042
R4172 dffrs_0.nand3_8.C.n5 dffrs_0.nand3_8.C.n4 6.04952
R4173 dffrs_0.nand3_7.B dffrs_0.nand3_8.C.n0 5.47979
R4174 dffrs_0.nand3_8.C.n2 dffrs_0.nand3_8.C.n1 5.13907
R4175 dffrs_0.nand3_6.Z dffrs_0.nand3_8.C.n6 4.72925
R4176 dffrs_0.nand3_8.C.n6 dffrs_0.nand3_8.C.n5 0.732092
R4177 dffrs_0.nand3_8.C.n4 dffrs_0.nand3_8.C.t0 0.7285
R4178 dffrs_0.nand3_8.C.n4 dffrs_0.nand3_8.C.t3 0.7285
R4179 dffrs_0.nand3_8.C.n3 dffrs_0.nand3_7.B 0.438233
R4180 dffrs_0.nand3_6.Z dffrs_0.nand3_8.C.n3 0.166901
R4181 dffrs_0.nand3_8.C.n2 dffrs_0.nand3_8.C 0.0455
R4182 dffrs_3.nand3_8.C.n0 dffrs_3.nand3_8.C.t5 40.8177
R4183 dffrs_3.nand3_8.C.n1 dffrs_3.nand3_8.C.t7 40.6313
R4184 dffrs_3.nand3_8.C.n1 dffrs_3.nand3_8.C.t6 27.3166
R4185 dffrs_3.nand3_8.C.n0 dffrs_3.nand3_8.C.t4 27.1302
R4186 dffrs_3.nand3_8.C.n3 dffrs_3.nand3_8.C.n2 14.119
R4187 dffrs_3.nand3_8.C.n6 dffrs_3.nand3_8.C.t2 10.0473
R4188 dffrs_3.nand3_8.C.n5 dffrs_3.nand3_8.C.t1 6.51042
R4189 dffrs_3.nand3_8.C.n5 dffrs_3.nand3_8.C.n4 6.04952
R4190 dffrs_3.nand3_7.B dffrs_3.nand3_8.C.n0 5.47979
R4191 dffrs_3.nand3_8.C.n2 dffrs_3.nand3_8.C.n1 5.13907
R4192 dffrs_3.nand3_6.Z dffrs_3.nand3_8.C.n6 4.72925
R4193 dffrs_3.nand3_8.C.n6 dffrs_3.nand3_8.C.n5 0.732092
R4194 dffrs_3.nand3_8.C.n4 dffrs_3.nand3_8.C.t3 0.7285
R4195 dffrs_3.nand3_8.C.n4 dffrs_3.nand3_8.C.t0 0.7285
R4196 dffrs_3.nand3_8.C.n3 dffrs_3.nand3_7.B 0.438233
R4197 dffrs_3.nand3_6.Z dffrs_3.nand3_8.C.n3 0.166901
R4198 dffrs_3.nand3_8.C.n2 dffrs_3.nand3_8.C 0.0455
R4199 dffrs_0.nand3_1.C.n0 dffrs_0.nand3_1.C.t5 40.6313
R4200 dffrs_0.nand3_1.C.n0 dffrs_0.nand3_1.C.t4 27.3166
R4201 dffrs_0.nand3_0.Z dffrs_0.nand3_1.C.n1 14.2854
R4202 dffrs_0.nand3_1.C.n4 dffrs_0.nand3_1.C.t3 10.0473
R4203 dffrs_0.nand3_1.C.n3 dffrs_0.nand3_1.C.t2 6.51042
R4204 dffrs_0.nand3_1.C.n3 dffrs_0.nand3_1.C.n2 6.04952
R4205 dffrs_0.nand3_1.C.n1 dffrs_0.nand3_1.C.n0 5.13907
R4206 dffrs_0.nand3_0.Z dffrs_0.nand3_1.C.n4 4.72925
R4207 dffrs_0.nand3_1.C.n4 dffrs_0.nand3_1.C.n3 0.732092
R4208 dffrs_0.nand3_1.C.n2 dffrs_0.nand3_1.C.t1 0.7285
R4209 dffrs_0.nand3_1.C.n2 dffrs_0.nand3_1.C.t0 0.7285
R4210 dffrs_0.nand3_1.C.n1 dffrs_0.nand3_1.C 0.0455
R4211 dffrs_5.nand3_8.C.n0 dffrs_5.nand3_8.C.t5 40.8177
R4212 dffrs_5.nand3_8.C.n1 dffrs_5.nand3_8.C.t6 40.6313
R4213 dffrs_5.nand3_8.C.n1 dffrs_5.nand3_8.C.t4 27.3166
R4214 dffrs_5.nand3_8.C.n0 dffrs_5.nand3_8.C.t7 27.1302
R4215 dffrs_5.nand3_8.C.n3 dffrs_5.nand3_8.C.n2 14.119
R4216 dffrs_5.nand3_8.C.n6 dffrs_5.nand3_8.C.t3 10.0473
R4217 dffrs_5.nand3_8.C.n5 dffrs_5.nand3_8.C.t2 6.51042
R4218 dffrs_5.nand3_8.C.n5 dffrs_5.nand3_8.C.n4 6.04952
R4219 dffrs_5.nand3_7.B dffrs_5.nand3_8.C.n0 5.47979
R4220 dffrs_5.nand3_8.C.n2 dffrs_5.nand3_8.C.n1 5.13907
R4221 dffrs_5.nand3_6.Z dffrs_5.nand3_8.C.n6 4.72925
R4222 dffrs_5.nand3_8.C.n6 dffrs_5.nand3_8.C.n5 0.732092
R4223 dffrs_5.nand3_8.C.n4 dffrs_5.nand3_8.C.t1 0.7285
R4224 dffrs_5.nand3_8.C.n4 dffrs_5.nand3_8.C.t0 0.7285
R4225 dffrs_5.nand3_8.C.n3 dffrs_5.nand3_7.B 0.438233
R4226 dffrs_5.nand3_6.Z dffrs_5.nand3_8.C.n3 0.166901
R4227 dffrs_5.nand3_8.C.n2 dffrs_5.nand3_8.C 0.0455
R4228 dffrs_4.nand3_1.C.n0 dffrs_4.nand3_1.C.t4 40.6313
R4229 dffrs_4.nand3_1.C.n0 dffrs_4.nand3_1.C.t5 27.3166
R4230 dffrs_4.nand3_0.Z dffrs_4.nand3_1.C.n1 14.2854
R4231 dffrs_4.nand3_1.C.n4 dffrs_4.nand3_1.C.t0 10.0473
R4232 dffrs_4.nand3_1.C.n3 dffrs_4.nand3_1.C.t1 6.51042
R4233 dffrs_4.nand3_1.C.n3 dffrs_4.nand3_1.C.n2 6.04952
R4234 dffrs_4.nand3_1.C.n1 dffrs_4.nand3_1.C.n0 5.13907
R4235 dffrs_4.nand3_0.Z dffrs_4.nand3_1.C.n4 4.72925
R4236 dffrs_4.nand3_1.C.n4 dffrs_4.nand3_1.C.n3 0.732092
R4237 dffrs_4.nand3_1.C.n2 dffrs_4.nand3_1.C.t3 0.7285
R4238 dffrs_4.nand3_1.C.n2 dffrs_4.nand3_1.C.t2 0.7285
R4239 dffrs_4.nand3_1.C.n1 dffrs_4.nand3_1.C 0.0455
R4240 dffrs_0.Qb.n0 dffrs_0.Qb.t6 41.0041
R4241 dffrs_0.Qb.n4 dffrs_0.Qb.t5 40.6313
R4242 dffrs_0.Qb.n2 dffrs_0.Qb.t4 40.6313
R4243 dffrs_0.Qb dffrs_7.setb 28.021
R4244 dffrs_0.Qb.n4 dffrs_0.Qb.t8 27.3166
R4245 dffrs_0.Qb.n2 dffrs_0.Qb.t7 27.3166
R4246 dffrs_0.Qb.n0 dffrs_0.Qb.t9 26.9438
R4247 dffrs_0.Qb.n9 dffrs_0.Qb.t1 10.0473
R4248 dffrs_0.Qb.n6 dffrs_0.Qb.n1 9.84255
R4249 dffrs_0.Qb.n5 dffrs_0.Qb.n3 9.22229
R4250 dffrs_0.Qb.n8 dffrs_0.Qb.t2 6.51042
R4251 dffrs_0.Qb.n8 dffrs_0.Qb.n7 6.04952
R4252 dffrs_0.Qb.n1 dffrs_0.Qb.n0 5.7305
R4253 dffrs_0.Qb.n5 dffrs_0.Qb.n4 5.14711
R4254 dffrs_0.Qb.n3 dffrs_0.Qb.n2 5.13907
R4255 dffrs_0.nand3_7.Z dffrs_0.Qb.n6 4.94976
R4256 dffrs_0.nand3_7.Z dffrs_0.Qb.n9 4.72925
R4257 dffrs_7.setb dffrs_7.nand3_0.C 0.784786
R4258 dffrs_0.Qb.n9 dffrs_0.Qb.n8 0.732092
R4259 dffrs_0.Qb.n7 dffrs_0.Qb.t0 0.7285
R4260 dffrs_0.Qb.n7 dffrs_0.Qb.t3 0.7285
R4261 dffrs_0.Qb.n6 dffrs_0.Qb 0.175225
R4262 dffrs_0.Qb.n1 dffrs_0.nand3_2.A 0.0455
R4263 dffrs_0.Qb.n3 dffrs_7.nand3_2.C 0.0455
R4264 dffrs_7.nand3_0.C dffrs_0.Qb.n5 0.0374643
R4265 dffrs_13.nand3_1.C.n0 dffrs_13.nand3_1.C.t4 40.6313
R4266 dffrs_13.nand3_1.C.n0 dffrs_13.nand3_1.C.t5 27.3166
R4267 dffrs_13.nand3_0.Z dffrs_13.nand3_1.C.n1 14.2854
R4268 dffrs_13.nand3_1.C.n4 dffrs_13.nand3_1.C.t0 10.0473
R4269 dffrs_13.nand3_1.C.n3 dffrs_13.nand3_1.C.t1 6.51042
R4270 dffrs_13.nand3_1.C.n3 dffrs_13.nand3_1.C.n2 6.04952
R4271 dffrs_13.nand3_1.C.n1 dffrs_13.nand3_1.C.n0 5.13907
R4272 dffrs_13.nand3_0.Z dffrs_13.nand3_1.C.n4 4.72925
R4273 dffrs_13.nand3_1.C.n4 dffrs_13.nand3_1.C.n3 0.732092
R4274 dffrs_13.nand3_1.C.n2 dffrs_13.nand3_1.C.t2 0.7285
R4275 dffrs_13.nand3_1.C.n2 dffrs_13.nand3_1.C.t3 0.7285
R4276 dffrs_13.nand3_1.C.n1 dffrs_13.nand3_1.C 0.0455
R4277 d4.n0 d4.t7 41.0041
R4278 d4.n1 d4.t4 40.8177
R4279 d4.n4 d4.t6 40.6313
R4280 d4.n3 dffrs_14.clk 33.675
R4281 d4.n4 d4.t8 27.3166
R4282 d4.n1 d4.t5 27.1302
R4283 d4.n0 d4.t9 26.9438
R4284 d4.n6 d4.n5 14.0582
R4285 d4.n6 d4.n3 11.3593
R4286 d4.n9 d4.t1 10.0473
R4287 d4.n8 d4.t0 6.51042
R4288 d4.n8 d4.n7 6.04952
R4289 dffrs_14.nand3_1.A d4.n0 5.7755
R4290 dffrs_14.nand3_6.B d4.n1 5.47979
R4291 d4.n5 d4.n4 5.13907
R4292 dffrs_7.nand3_2.Z d4.n9 4.72925
R4293 d4.n2 dffrs_14.nand3_6.B 2.17818
R4294 d4.n2 dffrs_14.nand3_1.A 1.34729
R4295 d4.n3 d4 1.26371
R4296 d4.n9 d4.n8 0.732092
R4297 d4.n7 d4.t3 0.7285
R4298 d4.n7 d4.t2 0.7285
R4299 dffrs_14.clk d4.n2 0.611214
R4300 dffrs_7.nand3_2.Z d4.n6 0.166901
R4301 d4.n5 dffrs_7.nand3_7.C 0.0455
R4302 dffrs_1.nand3_8.C.n0 dffrs_1.nand3_8.C.t7 40.8177
R4303 dffrs_1.nand3_8.C.n1 dffrs_1.nand3_8.C.t5 40.6313
R4304 dffrs_1.nand3_8.C.n1 dffrs_1.nand3_8.C.t4 27.3166
R4305 dffrs_1.nand3_8.C.n0 dffrs_1.nand3_8.C.t6 27.1302
R4306 dffrs_1.nand3_8.C.n3 dffrs_1.nand3_8.C.n2 14.119
R4307 dffrs_1.nand3_8.C.n6 dffrs_1.nand3_8.C.t1 10.0473
R4308 dffrs_1.nand3_8.C.n5 dffrs_1.nand3_8.C.t2 6.51042
R4309 dffrs_1.nand3_8.C.n5 dffrs_1.nand3_8.C.n4 6.04952
R4310 dffrs_1.nand3_7.B dffrs_1.nand3_8.C.n0 5.47979
R4311 dffrs_1.nand3_8.C.n2 dffrs_1.nand3_8.C.n1 5.13907
R4312 dffrs_1.nand3_6.Z dffrs_1.nand3_8.C.n6 4.72925
R4313 dffrs_1.nand3_8.C.n6 dffrs_1.nand3_8.C.n5 0.732092
R4314 dffrs_1.nand3_8.C.n4 dffrs_1.nand3_8.C.t0 0.7285
R4315 dffrs_1.nand3_8.C.n4 dffrs_1.nand3_8.C.t3 0.7285
R4316 dffrs_1.nand3_8.C.n3 dffrs_1.nand3_7.B 0.438233
R4317 dffrs_1.nand3_6.Z dffrs_1.nand3_8.C.n3 0.166901
R4318 dffrs_1.nand3_8.C.n2 dffrs_1.nand3_8.C 0.0455
R4319 dffrs_1.nand3_8.Z.n0 dffrs_1.nand3_8.Z.t6 41.0041
R4320 dffrs_1.nand3_8.Z.n1 dffrs_1.nand3_8.Z.t7 40.8177
R4321 dffrs_1.nand3_8.Z.n1 dffrs_1.nand3_8.Z.t5 27.1302
R4322 dffrs_1.nand3_8.Z.n0 dffrs_1.nand3_8.Z.t4 26.9438
R4323 dffrs_1.nand3_6.A dffrs_1.nand3_0.B 17.0041
R4324 dffrs_1.nand3_8.Z dffrs_1.nand3_8.Z.n2 14.8493
R4325 dffrs_1.nand3_8.Z.n5 dffrs_1.nand3_8.Z.t3 10.0473
R4326 dffrs_1.nand3_8.Z.n4 dffrs_1.nand3_8.Z.t2 6.51042
R4327 dffrs_1.nand3_8.Z.n4 dffrs_1.nand3_8.Z.n3 6.04952
R4328 dffrs_1.nand3_8.Z.n2 dffrs_1.nand3_8.Z.n0 5.7305
R4329 dffrs_1.nand3_0.B dffrs_1.nand3_8.Z.n1 5.47979
R4330 dffrs_1.nand3_8.Z dffrs_1.nand3_8.Z.n5 4.72925
R4331 dffrs_1.nand3_8.Z.n5 dffrs_1.nand3_8.Z.n4 0.732092
R4332 dffrs_1.nand3_8.Z.n3 dffrs_1.nand3_8.Z.t1 0.7285
R4333 dffrs_1.nand3_8.Z.n3 dffrs_1.nand3_8.Z.t0 0.7285
R4334 dffrs_1.nand3_8.Z.n2 dffrs_1.nand3_6.A 0.0455
R4335 d1.n0 d1.t8 41.0041
R4336 d1.n1 d1.t5 40.8177
R4337 d1.n4 d1.t4 40.6313
R4338 d1.n3 dffrs_9.clk 33.8765
R4339 d1.n4 d1.t6 27.3166
R4340 d1.n1 d1.t7 27.1302
R4341 d1.n0 d1.t9 26.9438
R4342 d1.n6 d1.n5 14.0582
R4343 d1.n6 d1.n3 11.729
R4344 d1.n9 d1.t2 10.0473
R4345 d1.n8 d1.t3 6.51042
R4346 d1.n8 d1.n7 6.04952
R4347 dffrs_9.nand3_1.A d1.n0 5.7755
R4348 dffrs_9.nand3_6.B d1.n1 5.47979
R4349 d1.n5 d1.n4 5.13907
R4350 dffrs_10.nand3_2.Z d1.n9 4.72925
R4351 d1.n2 dffrs_9.nand3_6.B 2.17818
R4352 d1.n2 dffrs_9.nand3_1.A 1.34729
R4353 d1.n3 d1 0.985679
R4354 d1.n9 d1.n8 0.732092
R4355 d1.n7 d1.t1 0.7285
R4356 d1.n7 d1.t0 0.7285
R4357 dffrs_9.clk d1.n2 0.610571
R4358 dffrs_10.nand3_2.Z d1.n6 0.166901
R4359 d1.n5 dffrs_10.nand3_7.C 0.0455
R4360 dffrs_3.nand3_6.C.n1 dffrs_3.nand3_6.C.t9 41.0041
R4361 dffrs_3.nand3_6.C.n0 dffrs_3.nand3_6.C.t7 40.8177
R4362 dffrs_3.nand3_6.C.n3 dffrs_3.nand3_6.C.t8 40.6313
R4363 dffrs_3.nand3_6.C.n3 dffrs_3.nand3_6.C.t5 27.3166
R4364 dffrs_3.nand3_6.C.n0 dffrs_3.nand3_6.C.t4 27.1302
R4365 dffrs_3.nand3_6.C.n1 dffrs_3.nand3_6.C.t6 26.9438
R4366 dffrs_3.nand3_6.C.n9 dffrs_3.nand3_6.C.t1 10.0473
R4367 dffrs_3.nand3_6.C.n5 dffrs_3.nand3_6.C.n4 9.90747
R4368 dffrs_3.nand3_6.C.n5 dffrs_3.nand3_6.C.n2 9.90116
R4369 dffrs_3.nand3_6.C.n8 dffrs_3.nand3_6.C.t0 6.51042
R4370 dffrs_3.nand3_6.C.n8 dffrs_3.nand3_6.C.n7 6.04952
R4371 dffrs_3.nand3_6.C.n2 dffrs_3.nand3_6.C.n1 5.7305
R4372 dffrs_3.nand3_2.B dffrs_3.nand3_6.C.n0 5.47979
R4373 dffrs_3.nand3_6.C.n4 dffrs_3.nand3_6.C.n3 5.13907
R4374 dffrs_3.nand3_1.Z dffrs_3.nand3_6.C.n9 4.72925
R4375 dffrs_3.nand3_6.C.n6 dffrs_3.nand3_6.C.n5 4.5005
R4376 dffrs_3.nand3_6.C.n9 dffrs_3.nand3_6.C.n8 0.732092
R4377 dffrs_3.nand3_6.C.n7 dffrs_3.nand3_6.C.t3 0.7285
R4378 dffrs_3.nand3_6.C.n7 dffrs_3.nand3_6.C.t2 0.7285
R4379 dffrs_3.nand3_1.Z dffrs_3.nand3_6.C.n6 0.449758
R4380 dffrs_3.nand3_6.C.n6 dffrs_3.nand3_2.B 0.166901
R4381 dffrs_3.nand3_6.C.n2 dffrs_3.nand3_0.A 0.0455
R4382 dffrs_3.nand3_6.C.n4 dffrs_3.nand3_6.C 0.0455
R4383 dffrs_2.d.n0 dffrs_2.d.t6 41.0041
R4384 dffrs_2.d.n1 dffrs_2.d.t5 40.6313
R4385 dffrs_2.d.n1 dffrs_2.d.t7 27.3166
R4386 dffrs_2.d.n0 dffrs_2.d.t4 26.9438
R4387 dffrs_2.d.n3 dffrs_2.d 17.5382
R4388 dffrs_2.d.n3 dffrs_2.d.n2 14.0582
R4389 dffrs_2.d.n6 dffrs_2.d.t3 10.0473
R4390 dffrs_2.d.n5 dffrs_2.d.t2 6.51042
R4391 dffrs_2.d.n5 dffrs_2.d.n4 6.04952
R4392 dffrs_2.nand3_8.A dffrs_2.d.n0 5.7755
R4393 dffrs_2.d.n2 dffrs_2.d.n1 5.13907
R4394 dffrs_1.nand3_2.Z dffrs_2.d.n6 4.72925
R4395 dffrs_2.d dffrs_2.nand3_8.A 0.784786
R4396 dffrs_2.d.n6 dffrs_2.d.n5 0.732092
R4397 dffrs_2.d.n4 dffrs_2.d.t1 0.7285
R4398 dffrs_2.d.n4 dffrs_2.d.t0 0.7285
R4399 dffrs_1.nand3_2.Z dffrs_2.d.n3 0.166901
R4400 dffrs_2.d.n2 dffrs_1.nand3_7.C 0.0455
R4401 dffrs_4.nand3_8.Z.n0 dffrs_4.nand3_8.Z.t4 41.0041
R4402 dffrs_4.nand3_8.Z.n1 dffrs_4.nand3_8.Z.t5 40.8177
R4403 dffrs_4.nand3_8.Z.n1 dffrs_4.nand3_8.Z.t7 27.1302
R4404 dffrs_4.nand3_8.Z.n0 dffrs_4.nand3_8.Z.t6 26.9438
R4405 dffrs_4.nand3_6.A dffrs_4.nand3_0.B 17.0041
R4406 dffrs_4.nand3_8.Z dffrs_4.nand3_8.Z.n2 14.8493
R4407 dffrs_4.nand3_8.Z.n5 dffrs_4.nand3_8.Z.t0 10.0473
R4408 dffrs_4.nand3_8.Z.n4 dffrs_4.nand3_8.Z.t1 6.51042
R4409 dffrs_4.nand3_8.Z.n4 dffrs_4.nand3_8.Z.n3 6.04952
R4410 dffrs_4.nand3_8.Z.n2 dffrs_4.nand3_8.Z.n0 5.7305
R4411 dffrs_4.nand3_0.B dffrs_4.nand3_8.Z.n1 5.47979
R4412 dffrs_4.nand3_8.Z dffrs_4.nand3_8.Z.n5 4.72925
R4413 dffrs_4.nand3_8.Z.n5 dffrs_4.nand3_8.Z.n4 0.732092
R4414 dffrs_4.nand3_8.Z.n3 dffrs_4.nand3_8.Z.t3 0.7285
R4415 dffrs_4.nand3_8.Z.n3 dffrs_4.nand3_8.Z.t2 0.7285
R4416 dffrs_4.nand3_8.Z.n2 dffrs_4.nand3_6.A 0.0455
R4417 dffrs_4.nand3_8.C.n0 dffrs_4.nand3_8.C.t4 40.8177
R4418 dffrs_4.nand3_8.C.n1 dffrs_4.nand3_8.C.t7 40.6313
R4419 dffrs_4.nand3_8.C.n1 dffrs_4.nand3_8.C.t5 27.3166
R4420 dffrs_4.nand3_8.C.n0 dffrs_4.nand3_8.C.t6 27.1302
R4421 dffrs_4.nand3_8.C.n3 dffrs_4.nand3_8.C.n2 14.119
R4422 dffrs_4.nand3_8.C.n6 dffrs_4.nand3_8.C.t3 10.0473
R4423 dffrs_4.nand3_8.C.n5 dffrs_4.nand3_8.C.t2 6.51042
R4424 dffrs_4.nand3_8.C.n5 dffrs_4.nand3_8.C.n4 6.04952
R4425 dffrs_4.nand3_7.B dffrs_4.nand3_8.C.n0 5.47979
R4426 dffrs_4.nand3_8.C.n2 dffrs_4.nand3_8.C.n1 5.13907
R4427 dffrs_4.nand3_6.Z dffrs_4.nand3_8.C.n6 4.72925
R4428 dffrs_4.nand3_8.C.n6 dffrs_4.nand3_8.C.n5 0.732092
R4429 dffrs_4.nand3_8.C.n4 dffrs_4.nand3_8.C.t1 0.7285
R4430 dffrs_4.nand3_8.C.n4 dffrs_4.nand3_8.C.t0 0.7285
R4431 dffrs_4.nand3_8.C.n3 dffrs_4.nand3_7.B 0.438233
R4432 dffrs_4.nand3_6.Z dffrs_4.nand3_8.C.n3 0.166901
R4433 dffrs_4.nand3_8.C.n2 dffrs_4.nand3_8.C 0.0455
R4434 dffrs_4.d.n0 dffrs_4.d.t4 41.0041
R4435 dffrs_4.d.n1 dffrs_4.d.t5 40.6313
R4436 dffrs_4.d.n1 dffrs_4.d.t7 27.3166
R4437 dffrs_4.d.n0 dffrs_4.d.t6 26.9438
R4438 dffrs_4.d.n3 dffrs_4.d 17.5382
R4439 dffrs_4.d.n3 dffrs_4.d.n2 14.0582
R4440 dffrs_4.d.n6 dffrs_4.d.t0 10.0473
R4441 dffrs_4.d.n5 dffrs_4.d.t1 6.51042
R4442 dffrs_4.d.n5 dffrs_4.d.n4 6.04952
R4443 dffrs_4.nand3_8.A dffrs_4.d.n0 5.7755
R4444 dffrs_4.d.n2 dffrs_4.d.n1 5.13907
R4445 dffrs_3.nand3_2.Z dffrs_4.d.n6 4.72925
R4446 dffrs_4.d dffrs_4.nand3_8.A 0.784786
R4447 dffrs_4.d.n6 dffrs_4.d.n5 0.732092
R4448 dffrs_4.d.n4 dffrs_4.d.t2 0.7285
R4449 dffrs_4.d.n4 dffrs_4.d.t3 0.7285
R4450 dffrs_3.nand3_2.Z dffrs_4.d.n3 0.166901
R4451 dffrs_4.d.n2 dffrs_3.nand3_7.C 0.0455
R4452 dffrs_2.nand3_8.Z.n0 dffrs_2.nand3_8.Z.t7 41.0041
R4453 dffrs_2.nand3_8.Z.n1 dffrs_2.nand3_8.Z.t6 40.8177
R4454 dffrs_2.nand3_8.Z.n1 dffrs_2.nand3_8.Z.t5 27.1302
R4455 dffrs_2.nand3_8.Z.n0 dffrs_2.nand3_8.Z.t4 26.9438
R4456 dffrs_2.nand3_6.A dffrs_2.nand3_0.B 17.0041
R4457 dffrs_2.nand3_8.Z dffrs_2.nand3_8.Z.n2 14.8493
R4458 dffrs_2.nand3_8.Z.n5 dffrs_2.nand3_8.Z.t1 10.0473
R4459 dffrs_2.nand3_8.Z.n4 dffrs_2.nand3_8.Z.t2 6.51042
R4460 dffrs_2.nand3_8.Z.n4 dffrs_2.nand3_8.Z.n3 6.04952
R4461 dffrs_2.nand3_8.Z.n2 dffrs_2.nand3_8.Z.n0 5.7305
R4462 dffrs_2.nand3_0.B dffrs_2.nand3_8.Z.n1 5.47979
R4463 dffrs_2.nand3_8.Z dffrs_2.nand3_8.Z.n5 4.72925
R4464 dffrs_2.nand3_8.Z.n5 dffrs_2.nand3_8.Z.n4 0.732092
R4465 dffrs_2.nand3_8.Z.n3 dffrs_2.nand3_8.Z.t3 0.7285
R4466 dffrs_2.nand3_8.Z.n3 dffrs_2.nand3_8.Z.t0 0.7285
R4467 dffrs_2.nand3_8.Z.n2 dffrs_2.nand3_6.A 0.0455
R4468 dffrs_2.nand3_8.C.n0 dffrs_2.nand3_8.C.t6 40.8177
R4469 dffrs_2.nand3_8.C.n1 dffrs_2.nand3_8.C.t7 40.6313
R4470 dffrs_2.nand3_8.C.n1 dffrs_2.nand3_8.C.t5 27.3166
R4471 dffrs_2.nand3_8.C.n0 dffrs_2.nand3_8.C.t4 27.1302
R4472 dffrs_2.nand3_8.C.n3 dffrs_2.nand3_8.C.n2 14.119
R4473 dffrs_2.nand3_8.C.n6 dffrs_2.nand3_8.C.t3 10.0473
R4474 dffrs_2.nand3_8.C.n5 dffrs_2.nand3_8.C.t2 6.51042
R4475 dffrs_2.nand3_8.C.n5 dffrs_2.nand3_8.C.n4 6.04952
R4476 dffrs_2.nand3_7.B dffrs_2.nand3_8.C.n0 5.47979
R4477 dffrs_2.nand3_8.C.n2 dffrs_2.nand3_8.C.n1 5.13907
R4478 dffrs_2.nand3_6.Z dffrs_2.nand3_8.C.n6 4.72925
R4479 dffrs_2.nand3_8.C.n6 dffrs_2.nand3_8.C.n5 0.732092
R4480 dffrs_2.nand3_8.C.n4 dffrs_2.nand3_8.C.t0 0.7285
R4481 dffrs_2.nand3_8.C.n4 dffrs_2.nand3_8.C.t1 0.7285
R4482 dffrs_2.nand3_8.C.n3 dffrs_2.nand3_7.B 0.438233
R4483 dffrs_2.nand3_6.Z dffrs_2.nand3_8.C.n3 0.166901
R4484 dffrs_2.nand3_8.C.n2 dffrs_2.nand3_8.C 0.0455
R4485 dffrs_2.Q.n0 dffrs_2.Q.t5 41.0041
R4486 dffrs_2.Q.n1 dffrs_2.Q.t4 40.6313
R4487 dffrs_2.Q.n1 dffrs_2.Q.t7 27.3166
R4488 dffrs_2.Q.n0 dffrs_2.Q.t6 26.9438
R4489 dffrs_2.Q.n3 dffrs_3.d 17.5382
R4490 dffrs_2.Q.n3 dffrs_2.Q.n2 14.0582
R4491 dffrs_2.Q.n6 dffrs_2.Q.t2 10.0473
R4492 dffrs_2.Q.n5 dffrs_2.Q.t1 6.51042
R4493 dffrs_2.Q.n5 dffrs_2.Q.n4 6.04952
R4494 dffrs_3.nand3_8.A dffrs_2.Q.n0 5.7755
R4495 dffrs_2.Q.n2 dffrs_2.Q.n1 5.13907
R4496 dffrs_2.nand3_2.Z dffrs_2.Q.n6 4.72925
R4497 dffrs_3.d dffrs_3.nand3_8.A 0.784786
R4498 dffrs_2.Q.n6 dffrs_2.Q.n5 0.732092
R4499 dffrs_2.Q.n4 dffrs_2.Q.t3 0.7285
R4500 dffrs_2.Q.n4 dffrs_2.Q.t0 0.7285
R4501 dffrs_2.nand3_2.Z dffrs_2.Q.n3 0.166901
R4502 dffrs_2.Q.n2 dffrs_2.nand3_7.C 0.0455
R4503 dffrs_3.nand3_1.C.n0 dffrs_3.nand3_1.C.t4 40.6313
R4504 dffrs_3.nand3_1.C.n0 dffrs_3.nand3_1.C.t5 27.3166
R4505 dffrs_3.nand3_0.Z dffrs_3.nand3_1.C.n1 14.2854
R4506 dffrs_3.nand3_1.C.n4 dffrs_3.nand3_1.C.t1 10.0473
R4507 dffrs_3.nand3_1.C.n3 dffrs_3.nand3_1.C.t0 6.51042
R4508 dffrs_3.nand3_1.C.n3 dffrs_3.nand3_1.C.n2 6.04952
R4509 dffrs_3.nand3_1.C.n1 dffrs_3.nand3_1.C.n0 5.13907
R4510 dffrs_3.nand3_0.Z dffrs_3.nand3_1.C.n4 4.72925
R4511 dffrs_3.nand3_1.C.n4 dffrs_3.nand3_1.C.n3 0.732092
R4512 dffrs_3.nand3_1.C.n2 dffrs_3.nand3_1.C.t2 0.7285
R4513 dffrs_3.nand3_1.C.n2 dffrs_3.nand3_1.C.t3 0.7285
R4514 dffrs_3.nand3_1.C.n1 dffrs_3.nand3_1.C 0.0455
R4515 dffrs_8.nand3_6.C.n1 dffrs_8.nand3_6.C.t6 41.0041
R4516 dffrs_8.nand3_6.C.n0 dffrs_8.nand3_6.C.t4 40.8177
R4517 dffrs_8.nand3_6.C.n3 dffrs_8.nand3_6.C.t5 40.6313
R4518 dffrs_8.nand3_6.C.n3 dffrs_8.nand3_6.C.t8 27.3166
R4519 dffrs_8.nand3_6.C.n0 dffrs_8.nand3_6.C.t7 27.1302
R4520 dffrs_8.nand3_6.C.n1 dffrs_8.nand3_6.C.t9 26.9438
R4521 dffrs_8.nand3_6.C.n9 dffrs_8.nand3_6.C.t2 10.0473
R4522 dffrs_8.nand3_6.C.n5 dffrs_8.nand3_6.C.n4 9.90747
R4523 dffrs_8.nand3_6.C.n5 dffrs_8.nand3_6.C.n2 9.90116
R4524 dffrs_8.nand3_6.C.n8 dffrs_8.nand3_6.C.t1 6.51042
R4525 dffrs_8.nand3_6.C.n8 dffrs_8.nand3_6.C.n7 6.04952
R4526 dffrs_8.nand3_6.C.n2 dffrs_8.nand3_6.C.n1 5.7305
R4527 dffrs_8.nand3_2.B dffrs_8.nand3_6.C.n0 5.47979
R4528 dffrs_8.nand3_6.C.n4 dffrs_8.nand3_6.C.n3 5.13907
R4529 dffrs_8.nand3_1.Z dffrs_8.nand3_6.C.n9 4.72925
R4530 dffrs_8.nand3_6.C.n6 dffrs_8.nand3_6.C.n5 4.5005
R4531 dffrs_8.nand3_6.C.n9 dffrs_8.nand3_6.C.n8 0.732092
R4532 dffrs_8.nand3_6.C.n7 dffrs_8.nand3_6.C.t3 0.7285
R4533 dffrs_8.nand3_6.C.n7 dffrs_8.nand3_6.C.t0 0.7285
R4534 dffrs_8.nand3_1.Z dffrs_8.nand3_6.C.n6 0.449758
R4535 dffrs_8.nand3_6.C.n6 dffrs_8.nand3_2.B 0.166901
R4536 dffrs_8.nand3_6.C.n2 dffrs_8.nand3_0.A 0.0455
R4537 dffrs_8.nand3_6.C.n4 dffrs_8.nand3_6.C 0.0455
R4538 d5.n0 d5.t4 40.6313
R4539 d5.n0 d5.t5 27.3166
R4540 d5.n2 d5.n1 14.0582
R4541 d5.n2 d5 12.6306
R4542 d5.n5 d5.t3 10.0473
R4543 d5.n4 d5.t2 6.51042
R4544 d5.n4 d5.n3 6.04952
R4545 d5.n1 d5.n0 5.13907
R4546 dffrs_14.nand3_2.Z d5.n5 4.72925
R4547 d5.n5 d5.n4 0.732092
R4548 d5.n3 d5.t1 0.7285
R4549 d5.n3 d5.t0 0.7285
R4550 dffrs_14.nand3_2.Z d5.n2 0.166901
R4551 d5.n1 dffrs_14.nand3_7.C 0.0455
.ends

