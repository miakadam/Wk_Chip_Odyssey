magic
tech gf180mcuD
magscale 1 10
timestamp 1757708813
<< metal1 >>
rect 5565 1279 5659 1291
rect 7675 1279 7747 1281
rect 5565 1203 5577 1279
rect 5657 1203 6695 1279
rect 6823 1203 7677 1279
rect 7733 1203 7747 1279
rect 5565 1201 5659 1203
rect 7675 1191 7747 1203
rect 8123 1279 8195 1281
rect 10201 1279 10305 1291
rect 8123 1203 8137 1279
rect 8193 1203 8979 1279
rect 9175 1203 10213 1279
rect 10293 1203 10305 1279
rect 8123 1191 8195 1203
rect 10201 1201 10305 1203
rect 1470 -3350 6470 -3275
rect 1470 -3675 6470 -3600
rect 1565 -5180 7841 -5100
<< via1 >>
rect 5577 1203 5657 1279
rect 7677 1203 7733 1279
rect 8137 1203 8193 1279
rect 10213 1203 10293 1279
<< metal2 >>
rect 1725 2783 5325 2843
rect 5909 2527 7276 2579
rect 5985 2523 7276 2527
rect 7220 2136 7276 2523
rect 5565 1279 5659 1291
rect 7677 1281 7733 1302
rect 8137 1281 8193 1648
rect 5565 1203 5577 1279
rect 5657 1203 5659 1279
rect 5565 1201 5659 1203
rect 7675 1279 7747 1281
rect 7675 1203 7677 1279
rect 7733 1203 7747 1279
rect 5577 -924 5657 1201
rect 7675 1191 7747 1203
rect 8123 1279 8195 1281
rect 8123 1203 8137 1279
rect 8193 1203 8195 1279
rect 8123 1191 8195 1203
rect 10201 1279 10305 1291
rect 10201 1203 10213 1279
rect 10293 1203 10305 1279
rect 10201 1201 10305 1203
rect 10213 100 10293 1201
use lvsclean_SAlatch  x1 /foss/designs/comparator/final_magic/fullcomp
timestamp 1757676563
transform 1 0 -9053 0 1 -1780
box 11023 -3410 22953 2129
use rslatch  x2 /foss/designs/comparator/final_magic/fullcomp
timestamp 1757675171
transform 1 0 5355 0 1 3480
box 1870 -2178 3290 -420
use inv_mia  x3 /foss/designs/comparator/final_magic/fullcomp
timestamp 1757680375
transform 1 0 1295 0 1 2105
box 5150 -1650 5730 322
use osu_sc_buf_4  x4 /foss/designs/comparator/final_magic/fullcomp
timestamp 1757675583
transform -1 0 6205 0 1 2073
box 0 -10 1140 1260
use inv_mia  x5
timestamp 1757680375
transform -1 0 14575 0 1 2105
box 5150 -1650 5730 322
<< labels >>
rlabel metal1 1470 -3310 1470 -3310 7 Vin1
port 6 w
rlabel metal1 1470 -3638 1470 -3638 7 Vin2
port 8 w
rlabel space 3494 -2927 3494 -2927 5 off3
port 5 s
rlabel space 1992 -2918 1992 -2918 5 off4
port 7 s
rlabel space 3392 -1380 3392 -1380 1 off2
port 3 n
rlabel space 4035 -1380 4035 -1380 1 off1
port 0 n
rlabel space 11850 -1380 11850 -1380 1 off5
port 9 n
rlabel space 12501 -1380 12501 -1380 1 off6
port 11 n
rlabel space 13866 -2918 13866 -2918 5 off8
port 13 s
rlabel space 12405 -2927 12405 -2927 5 off7
port 12 s
rlabel metal2 5577 172 5577 172 7 out1
rlabel metal2 10293 152 10293 152 3 out2
rlabel via1 8161 1233 8161 1233 7 out
port 3 w
rlabel metal2 5618 192 5618 192 1 Vout2
port 6 n
rlabel via1 5645 1229 5645 1229 3 in
port 2 w
rlabel metal1 1565 -5144 1565 -5144 7 CLK
port 4 w
rlabel metal2 1725 2811 1725 2811 7 Vout
port 10 w
rlabel metal1 7231 1279 7231 1279 1 inv1
rlabel metal1 8411 1279 8411 1279 1 inv2
rlabel metal2 6801 2579 6801 2579 1 latch
rlabel space 5523 3333 5523 3333 1 VDD
port 1 n
rlabel space 7660 3060 7660 3060 1 VDD
rlabel space 6535 2389 6535 2389 1 VDD
rlabel space 9317 2389 9317 2389 1 VDD
rlabel space 7953 146 7953 146 1 VDD
rlabel space 5790 -4801 5790 -4801 7 VSS
rlabel space 6775 481 6775 481 5 VSS
rlabel space 9203 481 9203 481 5 VSS
rlabel space 7897 1460 7897 1460 5 VSS
rlabel space 5543 2063 5543 2063 5 VSS
port 2 s
<< end >>
