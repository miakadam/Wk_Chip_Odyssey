magic
tech gf180mcuD
magscale 1 5
timestamp 1755275691
<< checkpaint >>
rect 1238 22530 4192 39774
rect 6614 22530 11332 28240
rect 1238 12392 11332 22530
rect -1030 9722 11332 12392
rect -1030 428 11752 9722
rect -1030 -342 13958 428
rect -1030 -500 17052 -342
rect -1030 -530 17724 -500
rect -1030 -644 18396 -530
rect -1030 -2630 18868 -644
rect -106 -2660 18868 -2630
rect 566 -2690 18868 -2660
rect 1238 -2720 18868 -2690
rect 2162 -2750 18868 -2720
rect 3086 -2780 18868 -2750
rect 3506 -2810 18868 -2780
rect 3926 -2840 18868 -2810
rect 6614 -2870 18868 -2840
rect 9302 -2900 18868 -2870
rect 9722 -2930 18868 -2900
rect 11928 -2960 18868 -2930
rect 12400 -2990 18868 -2960
rect 12872 -3020 18868 -2990
rect 13344 -3050 18868 -3020
rect 13816 -3080 18868 -3050
rect 15022 -3110 18868 -3080
rect 15694 -3140 18868 -3110
rect 16366 -3170 18868 -3140
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
use pfet_03v3_6Z3D7A  M1
timestamp 0
transform 1 0 13179 0 1 -1697
box -251 -263 251 263
use pfet_03v3_6Z3D7A  M2
timestamp 0
transform 1 0 13651 0 1 -1727
box -251 -263 251 263
use nfet_03v3_5MQYYT  M3
timestamp 0
transform 1 0 14123 0 1 -1865
box -251 -155 251 155
use nfet_03v3_5MQYYT  M4
timestamp 0
transform 1 0 14595 0 1 -1895
box -251 -155 251 155
use pfet_03v3_6Z3D7A  M5
timestamp 0
transform 1 0 17617 0 1 -1907
box -251 -263 251 263
use nfet_03v3_M5KWLQ  M6
timestamp 0
transform 1 0 16373 0 1 -1805
box -351 -305 351 305
use nfet_03v3_M5KWLQ  M7
timestamp 0
transform 1 0 17045 0 1 -1835
box -351 -305 351 305
use nfet_03v3_JSLSQ7  MN_CD
timestamp 0
transform 1 0 8973 0 1 12685
box -1359 -14555 1359 14555
use nfet_03v3_M2CYLQ  MN_CD_LOAD
timestamp 0
transform 1 0 10527 0 1 3411
box -225 -5311 225 5311
use nfet_03v3_BU4HR4  MN_CS
timestamp 0
transform 1 0 6285 0 1 9845
box -1359 -11685 1359 11685
use nfet_03v3_M2DZKQ  MN_LOAD_L
timestamp 0
transform 1 0 4731 0 1 -1105
box -225 -705 225 705
use nfet_03v3_M2DZKQ  MN_LOAD_R
timestamp 0
transform 1 0 4311 0 1 -1075
box -225 -705 225 705
use pfet_03v3_DA6X4Y  MP_CS_LOAD
timestamp 0
transform 1 0 2715 0 1 18527
box -477 -20247 477 20247
use pfet_03v3_DA94CY  MP_DIFF_L
timestamp 0
transform 1 0 1245 0 1 3967
box -351 -5627 351 5627
use pfet_03v3_DA94CY  MP_DIFF_R
timestamp 0
transform 1 0 1917 0 1 3937
box -351 -5627 351 5627
use pfet_03v3_4ZM98G  MP_MIRROR
timestamp 0
transform 1 0 3639 0 1 -895
box -477 -855 477 855
use pfet_03v3_4Z5NAG  MP_TAIL
timestamp 0
transform 1 0 447 0 1 4881
box -477 -6511 477 6511
use ppolyf_u_1k_MSK24U  XR1
timestamp 0
transform 1 0 15434 0 1 -1711
box -618 -369 618 369
use ppolyf_u_1k_XXBPKD  XR2
timestamp 0
transform 1 0 11840 0 1 -1251
box -1118 -679 1118 679
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 A_VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 IN_N
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 IN_P
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 640 0 0 0 A_VSS
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 640 0 0 0 I_REF
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 640 0 0 0 OUT
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 640 0 0 0 I_REF
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 640 0 0 0 A_VSS
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 640 0 0 0 A_VDD
port 8 nsew
<< end >>
