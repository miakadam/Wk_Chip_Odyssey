magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -702 -610 702 610
<< nmos >>
rect -452 -400 -52 400
rect 52 -400 452 400
<< ndiff >>
rect -540 387 -452 400
rect -540 -387 -527 387
rect -481 -387 -452 387
rect -540 -400 -452 -387
rect -52 387 52 400
rect -52 -387 -23 387
rect 23 -387 52 387
rect -52 -400 52 -387
rect 452 387 540 400
rect 452 -387 481 387
rect 527 -387 540 387
rect 452 -400 540 -387
<< ndiffc >>
rect -527 -387 -481 387
rect -23 -387 23 387
rect 481 -387 527 387
<< psubdiff >>
rect -678 514 678 586
rect -678 470 -606 514
rect -678 -470 -665 470
rect -619 -470 -606 470
rect 606 470 678 514
rect -678 -514 -606 -470
rect 606 -470 619 470
rect 665 -470 678 470
rect 606 -514 678 -470
rect -678 -586 678 -514
<< psubdiffcont >>
rect -665 -470 -619 470
rect 619 -470 665 470
<< polysilicon >>
rect -452 479 -52 492
rect -452 433 -439 479
rect -65 433 -52 479
rect -452 400 -52 433
rect 52 479 452 492
rect 52 433 65 479
rect 439 433 452 479
rect 52 400 452 433
rect -452 -433 -52 -400
rect -452 -479 -439 -433
rect -65 -479 -52 -433
rect -452 -492 -52 -479
rect 52 -433 452 -400
rect 52 -479 65 -433
rect 439 -479 452 -433
rect 52 -492 452 -479
<< polycontact >>
rect -439 433 -65 479
rect 65 433 439 479
rect -439 -479 -65 -433
rect 65 -479 439 -433
<< metal1 >>
rect -665 527 665 573
rect -665 470 -619 527
rect -450 433 -439 479
rect -65 433 -54 479
rect 54 433 65 479
rect 439 433 450 479
rect 619 470 665 527
rect -527 387 -481 398
rect -527 -398 -481 -387
rect -23 387 23 398
rect -23 -398 23 -387
rect 481 387 527 398
rect 481 -398 527 -387
rect -665 -527 -619 -470
rect -450 -479 -439 -433
rect -65 -479 -54 -433
rect 54 -479 65 -433
rect 439 -479 450 -433
rect 619 -527 665 -470
rect -665 -573 665 -527
<< properties >>
string FIXED_BBOX -642 -550 642 550
string gencell nfet_03v3
string library gf180mcu
string parameters w 4.0 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
