magic
tech gf180mcuD
magscale 1 10
timestamp 1758007907
<< metal1 >>
rect -800 1940 96 2140
rect 2062 1940 4290 2140
rect -800 720 -200 1940
rect 2322 967 4290 1940
rect 2412 804 2422 944
rect 4190 804 4200 944
rect 1352 30 1362 170
rect 1962 30 1972 170
rect 1352 -370 1362 -230
rect 1962 -370 1972 -230
rect 2412 -1156 2422 -1016
rect 4190 -1156 4200 -1016
rect -800 -2140 -200 -1420
rect 2322 -2140 4290 -1179
rect -800 -2340 96 -2140
rect 2062 -2340 4290 -2140
<< via1 >>
rect 2422 804 4190 944
rect 1362 30 1962 170
rect 1362 -370 1962 -230
rect 2422 -1156 4190 -1016
<< metal2 >>
rect -1024 920 0 976
rect 2410 944 4202 956
rect 2069 842 2181 898
rect -1024 764 0 820
rect -912 -522 -856 764
rect 1350 170 1974 182
rect 1350 30 1362 170
rect 1962 30 1974 170
rect 1350 18 1974 30
rect 2125 -200 2181 842
rect 2410 804 2422 944
rect 4190 804 4202 944
rect 2410 792 4202 804
rect 1350 -230 1974 -218
rect 1350 -370 1362 -230
rect 1962 -370 1974 -230
rect 2125 -256 2318 -200
rect 4294 -334 4350 -278
rect 1350 -382 1974 -370
rect 2125 -412 2263 -356
rect -912 -578 -800 -522
rect -200 -578 0 -522
rect -56 -1420 0 -578
rect 2125 -1442 2181 -412
rect 2410 -1016 4202 -1004
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
rect 2069 -1498 2181 -1442
rect -1024 -1576 0 -1520
<< via2 >>
rect 1362 30 1962 170
rect 2422 804 4190 944
rect 1362 -370 1962 -230
rect 2422 -1156 4190 -1016
<< metal3 >>
rect 2410 944 4202 956
rect 2410 804 2422 944
rect 4190 804 4202 944
rect 1350 170 1974 182
rect 1350 30 1362 170
rect 1962 30 1974 170
rect 1350 18 1974 30
rect 2410 -218 4202 804
rect 1350 -230 4202 -218
rect 1350 -370 1362 -230
rect 1962 -370 4202 -230
rect 1350 -382 4202 -370
rect 2410 -1016 4202 -1004
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
<< via3 >>
rect 1362 30 1962 170
rect 2422 -1156 4190 -1016
<< metal4 >>
rect 1350 170 4202 182
rect 1350 30 1362 170
rect 1962 30 4202 170
rect 1350 18 4202 30
rect 2410 -1016 4202 18
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
use and2  and2_0
timestamp 1758005944
transform 1 0 1647 0 1 10
box -1647 -10 422 2130
use and2  and2_1
timestamp 1758005944
transform 1 0 1647 0 1 -2330
box -1647 -10 422 2130
use inv2  inv2_0
timestamp 1757998295
transform 1 0 -2050 0 1 -50
box 1250 -1370 1850 770
use or2  or2_0
timestamp 1758004169
transform 1 0 2216 0 1 -1436
box 46 257 2078 2403
<< labels >>
rlabel metal2 -1024 947 -1024 947 7 Bit
port 0 w
rlabel metal2 -1024 791 -1024 791 7 Load
port 1 w
rlabel metal1 -469 2140 -469 2140 1 VDD
port 2 n
rlabel metal2 4350 -306 4350 -306 3 OUT
port 3 e
rlabel metal1 -500 -2340 -500 -2340 5 VSS
port 4 s
rlabel metal2 -1024 -1549 -1024 -1549 7 In
port 5 w
<< end >>
