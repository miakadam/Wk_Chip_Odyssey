magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< nwell >>
rect -502 -526 502 526
<< pmos >>
rect -252 116 -52 316
rect 52 116 252 316
rect -252 -316 -52 -116
rect 52 -316 252 -116
<< pdiff >>
rect -340 303 -252 316
rect -340 129 -327 303
rect -281 129 -252 303
rect -340 116 -252 129
rect -52 303 52 316
rect -52 129 -23 303
rect 23 129 52 303
rect -52 116 52 129
rect 252 303 340 316
rect 252 129 281 303
rect 327 129 340 303
rect 252 116 340 129
rect -340 -129 -252 -116
rect -340 -303 -327 -129
rect -281 -303 -252 -129
rect -340 -316 -252 -303
rect -52 -129 52 -116
rect -52 -303 -23 -129
rect 23 -303 52 -129
rect -52 -316 52 -303
rect 252 -129 340 -116
rect 252 -303 281 -129
rect 327 -303 340 -129
rect 252 -316 340 -303
<< pdiffc >>
rect -327 129 -281 303
rect -23 129 23 303
rect 281 129 327 303
rect -327 -303 -281 -129
rect -23 -303 23 -129
rect 281 -303 327 -129
<< nsubdiff >>
rect -478 430 478 502
rect -478 386 -406 430
rect -478 -386 -465 386
rect -419 -386 -406 386
rect 406 386 478 430
rect -478 -430 -406 -386
rect 406 -386 419 386
rect 465 -386 478 386
rect 406 -430 478 -386
rect -478 -502 478 -430
<< nsubdiffcont >>
rect -465 -386 -419 386
rect 419 -386 465 386
<< polysilicon >>
rect -252 395 -52 408
rect -252 349 -239 395
rect -65 349 -52 395
rect -252 316 -52 349
rect 52 395 252 408
rect 52 349 65 395
rect 239 349 252 395
rect 52 316 252 349
rect -252 83 -52 116
rect -252 37 -239 83
rect -65 37 -52 83
rect -252 24 -52 37
rect 52 83 252 116
rect 52 37 65 83
rect 239 37 252 83
rect 52 24 252 37
rect -252 -37 -52 -24
rect -252 -83 -239 -37
rect -65 -83 -52 -37
rect -252 -116 -52 -83
rect 52 -37 252 -24
rect 52 -83 65 -37
rect 239 -83 252 -37
rect 52 -116 252 -83
rect -252 -349 -52 -316
rect -252 -395 -239 -349
rect -65 -395 -52 -349
rect -252 -408 -52 -395
rect 52 -349 252 -316
rect 52 -395 65 -349
rect 239 -395 252 -349
rect 52 -408 252 -395
<< polycontact >>
rect -239 349 -65 395
rect 65 349 239 395
rect -239 37 -65 83
rect 65 37 239 83
rect -239 -83 -65 -37
rect 65 -83 239 -37
rect -239 -395 -65 -349
rect 65 -395 239 -349
<< metal1 >>
rect -465 443 465 489
rect -465 386 -419 443
rect -250 349 -239 395
rect -65 349 -54 395
rect 54 349 65 395
rect 239 349 250 395
rect 419 386 465 443
rect -327 303 -281 314
rect -327 118 -281 129
rect -23 303 23 314
rect -23 118 23 129
rect 281 303 327 314
rect 281 118 327 129
rect -250 37 -239 83
rect -65 37 -54 83
rect 54 37 65 83
rect 239 37 250 83
rect -250 -83 -239 -37
rect -65 -83 -54 -37
rect 54 -83 65 -37
rect 239 -83 250 -37
rect -327 -129 -281 -118
rect -327 -314 -281 -303
rect -23 -129 23 -118
rect -23 -314 23 -303
rect 281 -129 327 -118
rect 281 -314 327 -303
rect -465 -443 -419 -386
rect -250 -395 -239 -349
rect -65 -395 -54 -349
rect 54 -395 65 -349
rect 239 -395 250 -349
rect 419 -443 465 -386
rect -465 -489 465 -443
<< properties >>
string FIXED_BBOX -442 -466 442 466
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
