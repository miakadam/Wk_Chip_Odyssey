magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 1165 -23 1211
rect 23 1165 34 1176
rect -103 1054 -57 1130
rect 57 1054 103 1130
rect -34 973 -23 1019
rect -34 853 -23 899
rect 23 853 34 864
rect -103 742 -57 818
rect 57 742 103 818
rect -34 661 -23 707
rect -34 541 -23 587
rect 23 541 34 552
rect -103 430 -57 506
rect 57 430 103 506
rect -34 349 -23 395
rect -34 229 -23 275
rect 23 229 34 240
rect -103 118 -57 194
rect 57 118 103 194
rect -34 37 -23 83
rect -34 -83 -23 -37
rect 23 -83 34 -72
rect -103 -194 -57 -118
rect 57 -194 103 -118
rect -34 -275 -23 -229
rect -34 -395 -23 -349
rect 23 -395 34 -384
rect -103 -506 -57 -430
rect 57 -506 103 -430
rect -34 -587 -23 -541
rect -34 -707 -23 -661
rect 23 -707 34 -696
rect -103 -818 -57 -742
rect 57 -818 103 -742
rect -34 -899 -23 -853
rect -34 -1019 -23 -973
rect 23 -1019 34 -1008
rect -103 -1130 -57 -1054
rect 57 -1130 103 -1054
rect -34 -1211 -23 -1165
<< nwell >>
rect -278 -1342 278 1342
<< pmos >>
rect -28 1052 28 1132
rect -28 740 28 820
rect -28 428 28 508
rect -28 116 28 196
rect -28 -196 28 -116
rect -28 -508 28 -428
rect -28 -820 28 -740
rect -28 -1132 28 -1052
<< pdiff >>
rect -116 1119 -28 1132
rect -116 1065 -103 1119
rect -57 1065 -28 1119
rect -116 1052 -28 1065
rect 28 1119 116 1132
rect 28 1065 57 1119
rect 103 1065 116 1119
rect 28 1052 116 1065
rect -116 807 -28 820
rect -116 753 -103 807
rect -57 753 -28 807
rect -116 740 -28 753
rect 28 807 116 820
rect 28 753 57 807
rect 103 753 116 807
rect 28 740 116 753
rect -116 495 -28 508
rect -116 441 -103 495
rect -57 441 -28 495
rect -116 428 -28 441
rect 28 495 116 508
rect 28 441 57 495
rect 103 441 116 495
rect 28 428 116 441
rect -116 183 -28 196
rect -116 129 -103 183
rect -57 129 -28 183
rect -116 116 -28 129
rect 28 183 116 196
rect 28 129 57 183
rect 103 129 116 183
rect 28 116 116 129
rect -116 -129 -28 -116
rect -116 -183 -103 -129
rect -57 -183 -28 -129
rect -116 -196 -28 -183
rect 28 -129 116 -116
rect 28 -183 57 -129
rect 103 -183 116 -129
rect 28 -196 116 -183
rect -116 -441 -28 -428
rect -116 -495 -103 -441
rect -57 -495 -28 -441
rect -116 -508 -28 -495
rect 28 -441 116 -428
rect 28 -495 57 -441
rect 103 -495 116 -441
rect 28 -508 116 -495
rect -116 -753 -28 -740
rect -116 -807 -103 -753
rect -57 -807 -28 -753
rect -116 -820 -28 -807
rect 28 -753 116 -740
rect 28 -807 57 -753
rect 103 -807 116 -753
rect 28 -820 116 -807
rect -116 -1065 -28 -1052
rect -116 -1119 -103 -1065
rect -57 -1119 -28 -1065
rect -116 -1132 -28 -1119
rect 28 -1065 116 -1052
rect 28 -1119 57 -1065
rect 103 -1119 116 -1065
rect 28 -1132 116 -1119
<< pdiffc >>
rect -103 1065 -57 1119
rect 57 1065 103 1119
rect -103 753 -57 807
rect 57 753 103 807
rect -103 441 -57 495
rect 57 441 103 495
rect -103 129 -57 183
rect 57 129 103 183
rect -103 -183 -57 -129
rect 57 -183 103 -129
rect -103 -495 -57 -441
rect 57 -495 103 -441
rect -103 -807 -57 -753
rect 57 -807 103 -753
rect -103 -1119 -57 -1065
rect 57 -1119 103 -1065
<< nsubdiff >>
rect -254 1246 254 1318
rect -254 1202 -182 1246
rect -254 -1202 -241 1202
rect -195 -1202 -182 1202
rect 182 1202 254 1246
rect -254 -1246 -182 -1202
rect 182 -1202 195 1202
rect 241 -1202 254 1202
rect 182 -1246 254 -1202
rect -254 -1318 254 -1246
<< nsubdiffcont >>
rect -241 -1202 -195 1202
rect 195 -1202 241 1202
<< polysilicon >>
rect -36 1211 36 1224
rect -36 1165 -23 1211
rect 23 1165 36 1211
rect -36 1152 36 1165
rect -28 1132 28 1152
rect -28 1032 28 1052
rect -36 1019 36 1032
rect -36 973 -23 1019
rect 23 973 36 1019
rect -36 960 36 973
rect -36 899 36 912
rect -36 853 -23 899
rect 23 853 36 899
rect -36 840 36 853
rect -28 820 28 840
rect -28 720 28 740
rect -36 707 36 720
rect -36 661 -23 707
rect 23 661 36 707
rect -36 648 36 661
rect -36 587 36 600
rect -36 541 -23 587
rect 23 541 36 587
rect -36 528 36 541
rect -28 508 28 528
rect -28 408 28 428
rect -36 395 36 408
rect -36 349 -23 395
rect 23 349 36 395
rect -36 336 36 349
rect -36 275 36 288
rect -36 229 -23 275
rect 23 229 36 275
rect -36 216 36 229
rect -28 196 28 216
rect -28 96 28 116
rect -36 83 36 96
rect -36 37 -23 83
rect 23 37 36 83
rect -36 24 36 37
rect -36 -37 36 -24
rect -36 -83 -23 -37
rect 23 -83 36 -37
rect -36 -96 36 -83
rect -28 -116 28 -96
rect -28 -216 28 -196
rect -36 -229 36 -216
rect -36 -275 -23 -229
rect 23 -275 36 -229
rect -36 -288 36 -275
rect -36 -349 36 -336
rect -36 -395 -23 -349
rect 23 -395 36 -349
rect -36 -408 36 -395
rect -28 -428 28 -408
rect -28 -528 28 -508
rect -36 -541 36 -528
rect -36 -587 -23 -541
rect 23 -587 36 -541
rect -36 -600 36 -587
rect -36 -661 36 -648
rect -36 -707 -23 -661
rect 23 -707 36 -661
rect -36 -720 36 -707
rect -28 -740 28 -720
rect -28 -840 28 -820
rect -36 -853 36 -840
rect -36 -899 -23 -853
rect 23 -899 36 -853
rect -36 -912 36 -899
rect -36 -973 36 -960
rect -36 -1019 -23 -973
rect 23 -1019 36 -973
rect -36 -1032 36 -1019
rect -28 -1052 28 -1032
rect -28 -1152 28 -1132
rect -36 -1165 36 -1152
rect -36 -1211 -23 -1165
rect 23 -1211 36 -1165
rect -36 -1224 36 -1211
<< polycontact >>
rect -23 1165 23 1211
rect -23 973 23 1019
rect -23 853 23 899
rect -23 661 23 707
rect -23 541 23 587
rect -23 349 23 395
rect -23 229 23 275
rect -23 37 23 83
rect -23 -83 23 -37
rect -23 -275 23 -229
rect -23 -395 23 -349
rect -23 -587 23 -541
rect -23 -707 23 -661
rect -23 -899 23 -853
rect -23 -1019 23 -973
rect -23 -1211 23 -1165
<< metal1 >>
rect -241 1259 241 1305
rect -241 1202 -195 1259
rect -34 1165 -23 1211
rect 23 1165 34 1211
rect 195 1202 241 1259
rect -103 1119 -57 1130
rect -103 1054 -57 1065
rect 57 1119 103 1130
rect 57 1054 103 1065
rect -34 973 -23 1019
rect 23 973 34 1019
rect -34 853 -23 899
rect 23 853 34 899
rect -103 807 -57 818
rect -103 742 -57 753
rect 57 807 103 818
rect 57 742 103 753
rect -34 661 -23 707
rect 23 661 34 707
rect -34 541 -23 587
rect 23 541 34 587
rect -103 495 -57 506
rect -103 430 -57 441
rect 57 495 103 506
rect 57 430 103 441
rect -34 349 -23 395
rect 23 349 34 395
rect -34 229 -23 275
rect 23 229 34 275
rect -103 183 -57 194
rect -103 118 -57 129
rect 57 183 103 194
rect 57 118 103 129
rect -34 37 -23 83
rect 23 37 34 83
rect -34 -83 -23 -37
rect 23 -83 34 -37
rect -103 -129 -57 -118
rect -103 -194 -57 -183
rect 57 -129 103 -118
rect 57 -194 103 -183
rect -34 -275 -23 -229
rect 23 -275 34 -229
rect -34 -395 -23 -349
rect 23 -395 34 -349
rect -103 -441 -57 -430
rect -103 -506 -57 -495
rect 57 -441 103 -430
rect 57 -506 103 -495
rect -34 -587 -23 -541
rect 23 -587 34 -541
rect -34 -707 -23 -661
rect 23 -707 34 -661
rect -103 -753 -57 -742
rect -103 -818 -57 -807
rect 57 -753 103 -742
rect 57 -818 103 -807
rect -34 -899 -23 -853
rect 23 -899 34 -853
rect -34 -1019 -23 -973
rect 23 -1019 34 -973
rect -103 -1065 -57 -1054
rect -103 -1130 -57 -1119
rect 57 -1065 103 -1054
rect 57 -1130 103 -1119
rect -241 -1259 -195 -1202
rect -34 -1211 -23 -1165
rect 23 -1211 34 -1165
rect 195 -1259 241 -1202
rect -241 -1305 241 -1259
<< properties >>
string FIXED_BBOX -218 -1282 218 1282
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.4 l 0.28 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
