magic
tech gf180mcuD
magscale 1 10
timestamp 1755256602
<< error_s >>
rect 954 -2247 965 -2201
rect 1011 -2247 1022 -2236
rect 3234 -2357 3245 -2311
rect 3291 -2357 3302 -2346
rect 184 -2417 195 -2371
rect 241 -2417 252 -2406
rect 1714 -2467 1725 -2421
rect 1771 -2467 1782 -2456
rect 3924 -2457 3935 -2411
rect 3981 -2457 3992 -2446
rect 2474 -2507 2485 -2461
rect 4694 -2487 4705 -2441
rect 4751 -2487 4762 -2476
rect 2531 -2507 2542 -2496
rect 5424 -2567 5435 -2521
rect 5481 -2567 5492 -2556
rect 6224 -2637 6235 -2591
rect 6281 -2637 6292 -2626
rect 138 -2648 161 -2637
rect 275 -2648 298 -2637
rect 908 -2678 931 -2667
rect 1045 -2678 1068 -2667
rect 184 -2729 195 -2683
rect 1668 -2698 1691 -2687
rect 1805 -2698 1828 -2687
rect 954 -2759 965 -2713
rect 1714 -2779 1725 -2733
rect 2428 -2738 2451 -2727
rect 2565 -2738 2588 -2727
rect 2474 -2819 2485 -2773
rect 3188 -2788 3211 -2777
rect 3325 -2788 3348 -2777
rect 3234 -2869 3245 -2823
rect 3878 -2888 3901 -2877
rect 4015 -2888 4038 -2877
rect 4648 -2918 4671 -2907
rect 4785 -2918 4808 -2907
rect 3924 -2969 3935 -2923
rect 4694 -2999 4705 -2953
rect 5380 -2998 5401 -2987
rect 5515 -2998 5538 -2987
rect 5424 -3079 5435 -3033
rect 6178 -3068 6201 -3057
rect 6315 -3068 6338 -3057
rect 6224 -3149 6235 -3103
rect 174 -3547 185 -3501
rect 231 -3547 242 -3536
rect 964 -3567 975 -3521
rect 1021 -3567 1032 -3556
rect 1794 -3717 1805 -3671
rect 2494 -3687 2505 -3641
rect 2551 -3687 2562 -3676
rect 1851 -3717 1862 -3706
rect 3234 -3727 3245 -3681
rect 3291 -3727 3302 -3716
rect 2448 -3918 2471 -3907
rect 2585 -3918 2608 -3907
rect 1748 -3948 1771 -3937
rect 1885 -3948 1908 -3937
rect 128 -3978 151 -3967
rect 265 -3978 288 -3967
rect 918 -3998 941 -3987
rect 1055 -3998 1078 -3987
rect 174 -4059 185 -4013
rect 1794 -4029 1805 -3983
rect 2494 -3999 2505 -3953
rect 3964 -3997 3975 -3951
rect 4021 -3997 4032 -3986
rect 4644 -4017 4655 -3971
rect 5444 -3997 5455 -3951
rect 5501 -3997 5512 -3986
rect 4701 -4017 4712 -4006
rect 964 -4079 975 -4033
rect 6184 -4057 6195 -4011
rect 6241 -4057 6252 -4046
rect 3188 -4158 3211 -4147
rect 3325 -4158 3348 -4147
rect 3234 -4239 3245 -4193
rect 3918 -4228 3941 -4217
rect 4055 -4228 4078 -4217
rect 5398 -4228 5421 -4217
rect 5535 -4228 5558 -4217
rect 4598 -4248 4621 -4237
rect 4735 -4248 4758 -4237
rect 3964 -4309 3975 -4263
rect 4644 -4329 4655 -4283
rect 5444 -4309 5455 -4263
rect 6138 -4288 6161 -4277
rect 6275 -4288 6298 -4277
rect 6184 -4369 6195 -4323
<< metal1 >>
rect 10 -1620 210 -1420
rect 470 -1640 670 -1440
rect 1180 -1590 1380 -1390
rect 1610 -1650 1810 -1450
rect 2150 -1670 2350 -1470
rect 2710 -1750 2910 -1550
rect 3450 -1660 3650 -1460
rect 3980 -1830 4180 -1630
use nfet_03v3_NRMGVU  XM1
timestamp 1755256602
transform 1 0 218 0 1 -2550
box -278 -310 278 310
use pfet_03v3_NE88KN  XM2
timestamp 1755256602
transform 1 0 208 0 1 -3780
box -278 -410 278 410
use pfet_03v3_NE88KN  XM3
timestamp 1755256602
transform 1 0 988 0 1 -2480
box -278 -410 278 410
use pfet_03v3_NE88KN  XM4
timestamp 1755256602
transform 1 0 998 0 1 -3800
box -278 -410 278 410
use nfet_03v3_NRMGVU  XM5
timestamp 1755256602
transform 1 0 1748 0 1 -2600
box -278 -310 278 310
use nfet_03v3_NRMGVU  XM6
timestamp 1755256602
transform 1 0 1828 0 1 -3850
box -278 -310 278 310
use nfet_03v3_NRMGVU  XM7
timestamp 1755256602
transform 1 0 2508 0 1 -2640
box -278 -310 278 310
use nfet_03v3_NRMGVU  XM8
timestamp 1755256602
transform 1 0 2528 0 1 -3820
box -278 -310 278 310
use pfet_03v3_NE88KN  XM9
timestamp 1755256602
transform 1 0 3268 0 1 -2590
box -278 -410 278 410
use pfet_03v3_NE88KN  XM10
timestamp 1755256602
transform 1 0 3268 0 1 -3960
box -278 -410 278 410
use pfet_03v3_NE88KN  XM11
timestamp 1755256602
transform 1 0 3958 0 1 -2690
box -278 -410 278 410
use nfet_03v3_NRMGVU  XM12
timestamp 1755256602
transform 1 0 3998 0 1 -4130
box -278 -310 278 310
use pfet_03v3_NE88KN  XM13
timestamp 1755256602
transform 1 0 4728 0 1 -2720
box -278 -410 278 410
use nfet_03v3_NRMGVU  XM14
timestamp 1755256602
transform 1 0 4678 0 1 -4150
box -278 -310 278 310
use pfet_03v3_NE88KN  XM15
timestamp 1755256602
transform 1 0 5458 0 1 -2800
box -278 -410 278 410
use nfet_03v3_NRMGVU  XM16
timestamp 1755256602
transform 1 0 5478 0 1 -4130
box -278 -310 278 310
use pfet_03v3_NE88KN  XM17
timestamp 1755256602
transform 1 0 6258 0 1 -2870
box -278 -410 278 410
use nfet_03v3_NRMGVU  XM18
timestamp 1755256602
transform 1 0 6218 0 1 -4190
box -278 -310 278 310
<< labels >>
flabel metal1 2710 -1750 2910 -1550 0 FreeSans 1280 0 0 0 clk
port 3 nsew
flabel metal1 2150 -1670 2350 -1470 0 FreeSans 1280 0 0 0 set
port 4 nsew
flabel metal1 1610 -1650 1810 -1450 0 FreeSans 1280 0 0 0 q
port 6 nsew
flabel metal1 3450 -1660 3650 -1460 0 FreeSans 1280 0 0 0 reset
port 5 nsew
flabel metal1 3980 -1830 4180 -1630 0 FreeSans 1280 0 0 0 qb
port 7 nsew
flabel metal1 10 -1620 210 -1420 0 FreeSans 1280 0 0 0 vdd
port 0 nsew
flabel metal1 470 -1640 670 -1440 0 FreeSans 1280 0 0 0 vss
port 1 nsew
flabel metal1 1180 -1590 1380 -1390 0 FreeSans 1280 0 0 0 d
port 2 nsew
<< end >>
