magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -502 -310 502 310
<< nmos >>
rect -252 -100 -52 100
rect 52 -100 252 100
<< ndiff >>
rect -340 87 -252 100
rect -340 -87 -327 87
rect -281 -87 -252 87
rect -340 -100 -252 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 252 87 340 100
rect 252 -87 281 87
rect 327 -87 340 87
rect 252 -100 340 -87
<< ndiffc >>
rect -327 -87 -281 87
rect -23 -87 23 87
rect 281 -87 327 87
<< psubdiff >>
rect -478 214 478 286
rect -478 170 -406 214
rect -478 -170 -465 170
rect -419 -170 -406 170
rect 406 170 478 214
rect -478 -214 -406 -170
rect 406 -170 419 170
rect 465 -170 478 170
rect 406 -214 478 -170
rect -478 -286 478 -214
<< psubdiffcont >>
rect -465 -170 -419 170
rect 419 -170 465 170
<< polysilicon >>
rect -252 179 -52 192
rect -252 133 -239 179
rect -65 133 -52 179
rect -252 100 -52 133
rect 52 179 252 192
rect 52 133 65 179
rect 239 133 252 179
rect 52 100 252 133
rect -252 -133 -52 -100
rect -252 -179 -239 -133
rect -65 -179 -52 -133
rect -252 -192 -52 -179
rect 52 -133 252 -100
rect 52 -179 65 -133
rect 239 -179 252 -133
rect 52 -192 252 -179
<< polycontact >>
rect -239 133 -65 179
rect 65 133 239 179
rect -239 -179 -65 -133
rect 65 -179 239 -133
<< metal1 >>
rect -465 227 465 273
rect -465 170 -419 227
rect -250 133 -239 179
rect -65 133 -54 179
rect 54 133 65 179
rect 239 133 250 179
rect 419 170 465 227
rect -327 87 -281 98
rect -327 -98 -281 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 281 87 327 98
rect 281 -98 327 -87
rect -465 -227 -419 -170
rect -250 -179 -239 -133
rect -65 -179 -54 -133
rect 54 -179 65 -133
rect 239 -179 250 -133
rect 419 -227 465 -170
rect -465 -273 465 -227
<< properties >>
string FIXED_BBOX -442 -250 442 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
