* NGSPICE file created from dffrs.ext - technology: gf180mcuD

.subckt nfet_03v3_EPF4UP a_n224_n192# a_n40_n192# a_n450_n286# a_224_n100# a_n312_n100#
+ a_144_n192#
X0 a_224_n100# a_144_n192# a_40_n100# a_n450_n286# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.4u
X1 a_n144_n100# a_n224_n192# a_n312_n100# a_n450_n286# nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.4u
X2 a_40_n100# a_n40_n192# a_n144_n100# a_n450_n286# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.4u
.ends

.subckt pfet_03v3_54RA84 a_224_n250# a_n40_n342# a_n224_n342# a_40_n250# a_n312_n250#
+ a_n144_n250# w_n474_n460# a_144_n342#
X0 a_n144_n250# a_n224_n342# a_n312_n250# w_n474_n460# pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.4u
X1 a_40_n250# a_n40_n342# a_n144_n250# w_n474_n460# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.4u
X2 a_224_n250# a_144_n342# a_40_n250# w_n474_n460# pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.4u
.ends

.subckt nand3 VDD Z A B C VSS
XM1 C B VSS Z VSS A nfet_03v3_EPF4UP
XM3 Z B C VDD VDD Z VDD A pfet_03v3_54RA84
.ends

.subckt dffrs vdd vss d clk setb resetb Q Qb
Xnand3_0 vdd nand3_1/C nand3_6/C nand3_8/Z setb vss nand3
Xnand3_1 vdd nand3_6/C clk resetb nand3_1/C vss nand3
Xnand3_2 vdd Q Qb nand3_6/C setb vss nand3
Xnand3_7 vdd Qb resetb nand3_8/C Q vss nand3
Xnand3_6 vdd nand3_8/C nand3_8/Z clk nand3_6/C vss nand3
Xnand3_8 vdd nand3_8/Z d resetb nand3_8/C vss nand3
.ends

