* NGSPICE file created from v2comparator_no_offsetcal.ext - technology: gf180mcuD

.subckt comparator_no_offsetcal VDD VSS CLK Vin1 Vin2 Vout
X0 VDD a_5265_2223# Vout VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 VDD a_6467_n692# a_6379_n600# VDD pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=1u
X2 lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X3 VSS a_7711_n4982# a_7623_n4890# VSS nfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.4u
X4 VDD a_5265_2223# Vout VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VDD lvsclean_SAlatch_0.Vout2 x5.out VDD pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.4u
X6 lvsclean_SAlatch_0.Vp CLK VDD VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X7 a_9403_n600# a_9203_n692# VDD VDD pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=1u
X8 VDD CLK lvsclean_SAlatch_0.Vout2 VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X9 lvsclean_SAlatch_0.Vout2 a_8125_n1848# a_8037_n1756# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X10 lvsclean_SAlatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X11 a_6667_n4104# Vin1 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X12 VDD lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X13 lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X14 lvsclean_SAlatch_0.Vp a_6163_n3233# a_6075_n3141# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X15 lvsclean_SAlatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X16 a_6667_n4104# Vin2 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X17 a_6667_n4104# Vin1 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X18 a_9707_n4104# a_9507_n4196# lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
X19 Vout a_5265_2223# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X20 lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X21 VDD CLK lvsclean_SAlatch_0.Vq VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X22 a_7745_n1756# a_7545_n1848# lvsclean_SAlatch_0.Vout1 VSS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X23 a_5265_2223# x4.A VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X24 lvsclean_SAlatch_0.Vq lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X25 x4.A x2.Vout2 VDD VDD pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X26 x4.A x3.out VSS VSS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X27 lvsclean_SAlatch_0.Vq a_6163_n4196# a_6075_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X28 lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X29 a_6667_n4104# Vin2 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X30 a_6667_n4104# Vin2 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X31 Vout a_5265_2223# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X32 Vout a_5265_2223# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X33 lvsclean_SAlatch_0.Vout1 CLK VDD VDD pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.4u
X34 lvsclean_SAlatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X35 lvsclean_SAlatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X36 a_5265_2223# x4.A VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X37 VDD lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X38 lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X39 lvsclean_SAlatch_0.Vp lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X40 a_6667_n4104# Vin1 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X41 Vout a_5265_2223# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X42 lvsclean_SAlatch_0.Vq lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X43 a_9541_n1756# a_9341_n1848# lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X44 lvsclean_SAlatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X45 VDD x4.A x2.Vout2 VDD pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X46 VSS x5.out x2.Vout2 VSS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.4u
X47 a_6667_n4104# Vin1 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X48 lvsclean_SAlatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X49 lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X50 lvsclean_SAlatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X51 x3.out lvsclean_SAlatch_0.Vout1 VSS VSS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.4u
X52 lvsclean_SAlatch_0.Vp a_6329_n1848# a_6241_n1756# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X53 a_6667_n4104# CLK VSS VSS nfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.4u
X54 a_8159_n4890# a_8079_n4982# a_6667_n4104# VSS nfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.4u
X55 VSS a_5265_2223# Vout VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X56 VSS lvsclean_SAlatch_0.Vout2 x5.out VSS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.4u
X57 x3.out lvsclean_SAlatch_0.Vout1 VDD VDD pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.4u
X58 VDD lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X59 lvsclean_SAlatch_0.Vout2 lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X60 a_6667_n4104# Vin2 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X61 a_6667_n4104# Vin2 lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X62 VSS a_5265_2223# Vout VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X63 lvsclean_SAlatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X64 lvsclean_SAlatch_0.Vp Vin1 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X65 lvsclean_SAlatch_0.Vq Vin2 a_6667_n4104# VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X66 a_6667_n4104# Vin1 lvsclean_SAlatch_0.Vp VSS nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X67 VDD lvsclean_SAlatch_0.Vout1 lvsclean_SAlatch_0.Vout2 VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X68 a_9707_n3141# a_9507_n3233# lvsclean_SAlatch_0.Vq VSS nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
.ends

