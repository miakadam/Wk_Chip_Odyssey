magic
tech gf180mcuD
magscale 1 10
timestamp 1756985263
<< error_s >>
rect 451 423 483 469
rect 192 343 203 389
rect 449 320 483 368
rect 497 320 529 423
rect 971 403 1003 423
rect 192 71 203 117
rect 497 80 531 320
rect 712 283 723 329
rect 969 300 1003 320
rect 1017 300 1049 403
rect 2219 343 2251 389
rect 497 -23 529 80
rect 712 11 723 57
rect 1017 20 1051 300
rect 2217 240 2251 288
rect 2265 240 2297 343
rect 3467 243 3499 289
rect 1017 -83 1049 20
rect 2265 -40 2299 240
rect 3465 140 3499 188
rect 3513 140 3545 243
rect 3987 183 4019 229
rect 4516 183 4576 200
rect 2265 -143 2297 -40
rect 3513 -100 3547 140
rect 3728 103 3739 149
rect 3985 80 4019 128
rect 4033 80 4065 183
rect 4507 163 4576 183
rect 3513 -203 3545 -100
rect 3728 -169 3739 -123
rect 4033 -160 4067 80
rect 4248 43 4259 89
rect 4516 80 4585 163
rect 6363 103 6395 149
rect 4505 60 4585 80
rect 4033 -263 4065 -160
rect 4248 -229 4259 -183
rect 4516 -220 4587 60
rect 6361 0 6395 48
rect 6409 0 6441 103
rect 4516 -323 4585 -220
rect 6409 -280 6443 0
rect 12451 -140 12483 -131
rect 12451 -177 12520 -140
rect 12192 -257 12203 -211
rect 12460 -232 12529 -177
rect 12449 -280 12529 -232
rect 12971 -237 13003 -191
rect 4516 -360 4576 -323
rect 6409 -383 6441 -280
rect 12192 -529 12203 -483
rect 12460 -520 12531 -280
rect 12712 -317 12723 -271
rect 12969 -340 13003 -292
rect 13017 -340 13049 -237
rect 13675 -297 13707 -251
rect 12460 -623 12529 -520
rect 12712 -589 12723 -543
rect 13017 -580 13051 -340
rect 13232 -377 13243 -331
rect 13416 -377 13427 -331
rect 13673 -400 13707 -352
rect 13721 -400 13753 -297
rect 14747 -357 14779 -311
rect 12460 -660 12520 -623
rect 13017 -683 13049 -580
rect 13232 -649 13243 -603
rect 13416 -649 13427 -603
rect 13721 -640 13755 -400
rect 13936 -437 13947 -391
rect 14120 -437 14131 -391
rect 14304 -437 14315 -391
rect 14488 -437 14499 -391
rect 14745 -460 14779 -412
rect 14793 -460 14825 -357
rect 15819 -417 15851 -371
rect 13721 -743 13753 -640
rect 13936 -709 13947 -663
rect 14120 -709 14131 -663
rect 14304 -709 14315 -663
rect 14488 -709 14499 -663
rect 14793 -700 14827 -460
rect 15008 -497 15019 -451
rect 15192 -497 15203 -451
rect 15376 -497 15387 -451
rect 15560 -497 15571 -451
rect 15817 -520 15851 -472
rect 15865 -520 15897 -417
rect 16339 -477 16371 -431
rect 14793 -803 14825 -700
rect 15008 -769 15019 -723
rect 15192 -769 15203 -723
rect 15376 -769 15387 -723
rect 15560 -769 15571 -723
rect 15865 -760 15899 -520
rect 16080 -557 16091 -511
rect 16337 -580 16371 -532
rect 16385 -580 16417 -477
rect 17043 -537 17075 -491
rect 15865 -863 15897 -760
rect 16080 -829 16091 -783
rect 16385 -820 16419 -580
rect 16600 -617 16611 -571
rect 16784 -617 16795 -571
rect 17041 -640 17075 -592
rect 17089 -640 17121 -537
rect 18115 -597 18147 -551
rect 16385 -923 16417 -820
rect 16600 -889 16611 -843
rect 16784 -889 16795 -843
rect 17089 -880 17123 -640
rect 17304 -677 17315 -631
rect 17488 -677 17499 -631
rect 17672 -677 17683 -631
rect 17856 -677 17867 -631
rect 18113 -700 18147 -652
rect 18161 -700 18193 -597
rect 17089 -983 17121 -880
rect 17304 -949 17315 -903
rect 17488 -949 17499 -903
rect 17672 -949 17683 -903
rect 17856 -949 17867 -903
rect 18161 -940 18195 -700
rect 18376 -737 18387 -691
rect 18560 -737 18571 -691
rect 18744 -737 18755 -691
rect 18928 -737 18939 -691
rect 23971 -837 24003 -791
rect 23160 -917 23171 -871
rect 23344 -917 23355 -871
rect 23528 -917 23539 -871
rect 23712 -917 23723 -871
rect 23969 -940 24003 -892
rect 24017 -940 24049 -837
rect 18161 -1043 18193 -940
rect 18376 -1009 18387 -963
rect 18560 -1009 18571 -963
rect 18744 -1009 18755 -963
rect 18928 -1009 18939 -963
rect 23160 -1189 23171 -1143
rect 23344 -1189 23355 -1143
rect 23528 -1189 23539 -1143
rect 23712 -1189 23723 -1143
rect 24017 -1180 24051 -940
rect 24232 -977 24243 -931
rect 24416 -977 24427 -931
rect 24600 -977 24611 -931
rect 24784 -977 24795 -931
rect 24017 -1283 24049 -1180
rect 24232 -1249 24243 -1203
rect 24416 -1249 24427 -1203
rect 24600 -1249 24611 -1203
rect 24784 -1249 24795 -1203
<< pwell >>
rect 9945 3495 10040 3814
rect 13040 3485 13135 3804
rect 13055 3235 13120 3250
rect 10430 3135 10520 3205
rect 10430 3125 10520 3130
rect 10588 2140 10668 2235
<< polysilicon >>
rect 10430 3135 10520 3205
rect 10430 3125 10520 3130
<< metal1 >>
rect 10588 3486 10668 3496
rect 9900 3260 9960 3485
rect 10025 3260 10035 3485
rect 9900 3255 10035 3260
rect 10284 3402 10364 3412
rect 10284 3241 10296 3402
rect 10352 3241 10364 3402
rect 10588 3269 10600 3486
rect 10656 3269 10668 3486
rect 11196 3486 11276 3496
rect 11196 3430 11208 3486
rect 11264 3430 11276 3486
rect 11196 3420 11276 3430
rect 11804 3486 11884 3496
rect 11804 3430 11816 3486
rect 11872 3430 11884 3486
rect 11804 3420 11884 3430
rect 12412 3486 12492 3496
rect 10588 3261 10668 3269
rect 10892 3402 10972 3412
rect 10284 3231 10364 3241
rect 10892 3241 10904 3402
rect 10960 3241 10972 3402
rect 10892 3231 10972 3241
rect 11500 3402 11580 3412
rect 11500 3241 11512 3402
rect 11568 3241 11580 3402
rect 11500 3231 11580 3241
rect 12108 3402 12188 3412
rect 12108 3241 12120 3402
rect 12176 3241 12188 3402
rect 12108 3231 12188 3241
rect 12412 3241 12424 3486
rect 12480 3241 12492 3486
rect 12412 3231 12492 3241
rect 12716 3402 12796 3412
rect 12716 3241 12728 3402
rect 12784 3241 12796 3402
rect 13045 3260 13055 3485
rect 13120 3260 13180 3485
rect 13045 3255 13180 3260
rect 12716 3231 12796 3241
rect 10425 3140 10440 3195
rect 10075 3085 10270 3140
rect 10380 3135 10440 3140
rect 10510 3140 10525 3195
rect 10510 3135 10565 3140
rect 10730 3135 10745 3195
rect 10815 3135 10830 3195
rect 10985 3085 11180 3140
rect 11290 3085 11485 3140
rect 11640 3135 11655 3195
rect 11725 3135 11740 3195
rect 11945 3135 11960 3195
rect 12030 3135 12045 3195
rect 12205 3085 12400 3140
rect 12505 3085 12700 3140
rect 12860 3135 12875 3195
rect 12945 3135 12960 3195
rect 10075 3070 13670 3085
rect 10075 3010 13190 3070
rect 13250 3010 13670 3070
rect 10075 2700 13450 2760
rect 13510 2700 13670 2760
rect 10075 2685 13670 2700
rect 10075 2635 10270 2685
rect 10985 2635 11180 2685
rect 11290 2635 11485 2685
rect 12200 2635 12395 2685
rect 12505 2635 12700 2685
rect 10430 2590 10440 2635
rect 10425 2575 10440 2590
rect 10510 2590 10520 2635
rect 10735 2590 10745 2635
rect 10510 2575 10525 2590
rect 10730 2575 10745 2590
rect 10815 2590 10825 2635
rect 11645 2590 11655 2635
rect 10815 2575 10830 2590
rect 11640 2575 11655 2590
rect 11725 2590 11735 2635
rect 11950 2590 11960 2635
rect 11725 2575 11740 2590
rect 11945 2575 11960 2590
rect 12030 2590 12040 2635
rect 12865 2590 12875 2635
rect 12030 2575 12045 2590
rect 12860 2575 12875 2590
rect 12945 2590 12955 2635
rect 12945 2575 12960 2590
rect 10284 2531 10364 2541
rect 10284 2370 10296 2531
rect 10352 2370 10364 2531
rect 10892 2531 10972 2541
rect 10284 2360 10364 2370
rect 10588 2497 10668 2507
rect 9980 2342 10060 2352
rect 9980 2286 9992 2342
rect 10048 2286 10060 2342
rect 9980 2276 10060 2286
rect 10588 2286 10600 2497
rect 10656 2286 10668 2497
rect 10892 2370 10904 2531
rect 10960 2370 10972 2531
rect 10892 2360 10972 2370
rect 11196 2531 11276 2541
rect 10588 2276 10668 2286
rect 11196 2286 11208 2531
rect 11264 2286 11276 2531
rect 11500 2531 11580 2541
rect 11500 2370 11512 2531
rect 11568 2370 11580 2531
rect 12108 2531 12188 2541
rect 11500 2360 11580 2370
rect 11804 2497 11884 2507
rect 11196 2276 11276 2286
rect 11804 2286 11816 2497
rect 11872 2286 11884 2497
rect 12108 2370 12120 2531
rect 12176 2370 12188 2531
rect 12108 2360 12188 2370
rect 12412 2531 12492 2541
rect 11804 2276 11884 2286
rect 12412 2286 12424 2531
rect 12480 2286 12492 2531
rect 12412 2276 12492 2286
rect 12716 2531 12796 2541
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2276 12796 2286
rect 13020 2343 13100 2353
rect 13020 2286 13032 2343
rect 13088 2286 13100 2343
rect 13020 2276 13100 2286
<< via1 >>
rect 9960 3260 10025 3485
rect 10296 3241 10352 3402
rect 10600 3269 10656 3486
rect 11208 3430 11264 3486
rect 11816 3430 11872 3486
rect 10904 3241 10960 3402
rect 11512 3241 11568 3402
rect 12120 3241 12176 3402
rect 12424 3241 12480 3486
rect 12728 3241 12784 3402
rect 13055 3260 13120 3485
rect 10440 3135 10510 3195
rect 10745 3135 10815 3195
rect 11655 3135 11725 3195
rect 11960 3135 12030 3195
rect 12875 3135 12945 3195
rect 13190 3010 13250 3070
rect 13450 2700 13510 2760
rect 10440 2575 10510 2635
rect 10745 2575 10815 2635
rect 11655 2575 11725 2635
rect 11960 2575 12030 2635
rect 12875 2575 12945 2635
rect 10296 2370 10352 2531
rect 9992 2286 10048 2342
rect 10600 2286 10656 2497
rect 10904 2370 10960 2531
rect 11208 2286 11264 2531
rect 11512 2370 11568 2531
rect 11816 2286 11872 2497
rect 12120 2370 12176 2531
rect 12424 2286 12480 2531
rect 12728 2286 12784 2531
rect 13032 2286 13088 2343
<< metal2 >>
rect 9945 3485 10040 3814
rect 13040 3688 13135 3804
rect 9945 3260 9960 3485
rect 10025 3260 10040 3485
rect 10588 3632 13135 3688
rect 10588 3486 10668 3632
rect 9945 3255 10040 3260
rect 10284 3402 10364 3412
rect 10284 3241 10296 3402
rect 10352 3241 10364 3402
rect 10588 3269 10600 3486
rect 10656 3269 10668 3486
rect 11196 3486 11276 3496
rect 11196 3430 11208 3486
rect 11264 3430 11276 3486
rect 11196 3420 11276 3430
rect 11804 3486 11884 3632
rect 11804 3430 11816 3486
rect 11872 3430 11884 3486
rect 11804 3420 11884 3430
rect 12412 3486 12492 3496
rect 10588 3261 10668 3269
rect 10892 3402 10972 3412
rect 10284 2911 10364 3241
rect 10892 3241 10904 3402
rect 10960 3241 10972 3402
rect 10425 3195 10830 3205
rect 10425 3135 10440 3195
rect 10510 3135 10745 3195
rect 10815 3135 10830 3195
rect 10425 3125 10830 3135
rect 10892 2911 10972 3241
rect 11500 3402 11580 3412
rect 11500 3241 11512 3402
rect 11568 3241 11580 3402
rect 11500 2911 11580 3241
rect 12108 3402 12188 3412
rect 12108 3241 12120 3402
rect 12176 3241 12188 3402
rect 11640 3195 12045 3205
rect 11640 3135 11655 3195
rect 11725 3135 11960 3195
rect 12030 3135 12045 3195
rect 11640 3125 12045 3135
rect 12108 2911 12188 3241
rect 12412 3241 12424 3486
rect 12480 3241 12492 3486
rect 13040 3485 13135 3632
rect 12412 3231 12492 3241
rect 12716 3402 12796 3412
rect 12716 3241 12728 3402
rect 12784 3241 12796 3402
rect 13040 3260 13055 3485
rect 13120 3260 13135 3485
rect 13040 3255 13135 3260
rect 12716 2911 12796 3241
rect 12860 3195 12960 3205
rect 13154 3195 13380 3196
rect 12860 3135 12875 3195
rect 12945 3136 13380 3195
rect 12945 3135 13119 3136
rect 12860 3125 12960 3135
rect 13175 3070 13260 3080
rect 13175 3010 13190 3070
rect 13250 3010 13260 3070
rect 13175 2995 13260 3010
rect 10284 2855 12796 2911
rect 10284 2531 10364 2855
rect 10425 2635 10830 2645
rect 10425 2575 10440 2635
rect 10510 2575 10745 2635
rect 10815 2575 10830 2635
rect 10425 2565 10830 2575
rect 10284 2370 10296 2531
rect 10352 2370 10364 2531
rect 10892 2531 10972 2855
rect 9980 2342 10060 2352
rect 9980 2286 9992 2342
rect 10048 2286 10060 2342
rect 9980 2276 10060 2286
rect 10284 2024 10364 2370
rect 10588 2497 10668 2507
rect 10588 2286 10600 2497
rect 10656 2286 10668 2497
rect 10892 2370 10904 2531
rect 10960 2370 10972 2531
rect 10892 2360 10972 2370
rect 11196 2531 11276 2541
rect 10588 2140 10668 2286
rect 11196 2286 11208 2531
rect 11264 2286 11276 2531
rect 11500 2531 11580 2855
rect 11640 2635 12045 2645
rect 11640 2575 11655 2635
rect 11725 2575 11960 2635
rect 12030 2575 12045 2635
rect 11640 2565 12045 2575
rect 11500 2370 11512 2531
rect 11568 2370 11580 2531
rect 12108 2531 12188 2855
rect 11500 2360 11580 2370
rect 11804 2497 11884 2507
rect 11196 2276 11276 2286
rect 11804 2286 11816 2497
rect 11872 2286 11884 2497
rect 12108 2370 12120 2531
rect 12176 2370 12188 2531
rect 12108 2360 12188 2370
rect 12412 2531 12492 2541
rect 11804 2140 11884 2286
rect 12412 2286 12424 2531
rect 12480 2286 12492 2531
rect 12412 2276 12492 2286
rect 12716 2531 12796 2855
rect 13190 2855 13250 2995
rect 13320 2975 13380 3136
rect 13320 2915 13510 2975
rect 13190 2795 13380 2855
rect 12860 2635 12960 2645
rect 13320 2635 13380 2795
rect 13450 2770 13510 2915
rect 13440 2760 13520 2770
rect 13440 2700 13450 2760
rect 13510 2700 13520 2760
rect 13440 2690 13520 2700
rect 12860 2575 12875 2635
rect 12945 2575 13380 2635
rect 12860 2565 12960 2575
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2276 12796 2286
rect 13020 2343 13100 2353
rect 13020 2286 13032 2343
rect 13088 2286 13100 2343
rect 13020 2140 13100 2286
rect 10588 2084 13100 2140
rect 10284 2013 12806 2024
rect 10284 1957 12716 2013
rect 12796 1957 12806 2013
rect 10284 1947 12806 1957
<< via2 >>
rect 9960 3260 10025 3485
rect 10600 3269 10656 3325
rect 11208 3430 11264 3486
rect 12424 3241 12480 3486
rect 13055 3260 13120 3485
rect 9992 2286 10048 2342
rect 10600 2441 10656 2497
rect 11208 2286 11264 2531
rect 11816 2441 11872 2497
rect 12424 2286 12480 2531
rect 12728 2286 12784 2531
rect 12716 1957 12796 2013
<< metal3 >>
rect 10035 3486 12492 3496
rect 10035 3485 11208 3486
rect 9950 3260 9960 3485
rect 10025 3430 11208 3485
rect 11264 3430 12424 3486
rect 10025 3420 12424 3430
rect 10025 3260 10035 3420
rect 10588 3325 10668 3335
rect 10588 3269 10600 3325
rect 10656 3269 10668 3325
rect 9960 2855 10025 3260
rect 10588 2971 10668 3269
rect 12412 3241 12424 3420
rect 12480 3241 12492 3486
rect 13045 3260 13055 3485
rect 13120 3260 13130 3485
rect 13045 3255 13130 3260
rect 12412 2971 12492 3241
rect 10588 2911 11276 2971
rect 9960 2795 10668 2855
rect 10588 2497 10668 2795
rect 10588 2441 10600 2497
rect 10656 2441 10668 2497
rect 10588 2431 10668 2441
rect 11196 2531 11276 2911
rect 11196 2352 11208 2531
rect 9980 2342 11208 2352
rect 9980 2286 9992 2342
rect 10048 2286 11208 2342
rect 11264 2352 11276 2531
rect 11804 2911 12492 2971
rect 11804 2497 11884 2911
rect 13055 2855 13120 3255
rect 11804 2441 11816 2497
rect 11872 2441 11884 2497
rect 11804 2431 11884 2441
rect 12412 2795 13120 2855
rect 12412 2531 12492 2795
rect 12412 2352 12424 2531
rect 11264 2286 12424 2352
rect 12480 2286 12492 2531
rect 9980 2276 12492 2286
rect 12716 2531 12796 2541
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2024 12796 2286
rect 12706 2013 12806 2024
rect 12706 1957 12716 2013
rect 12796 1957 12806 2013
rect 12706 1947 12806 1957
use nfet_03v3_RPTYYZ  nfet_03v3_RPTYYZ_0
timestamp 1756981609
transform 1 0 12300 0 1 3366
box -820 -266 820 266
use pfet_03v3_PQ9NUS  XM1
timestamp 1756981609
transform 1 0 230 0 1 230
box -290 -290 290 290
use pfet_03v3_PQ9NUS  XM2
timestamp 1756981609
transform 1 0 750 0 1 170
box -290 -290 290 290
use pfet_03v3_V5CHCW  XM3
timestamp 1756981609
transform 1 0 1634 0 1 130
box -654 -310 654 310
use pfet_03v3_V5CHCW  XM4
timestamp 1756981609
transform 1 0 2882 0 1 70
box -654 -310 654 310
use pfet_03v3_PQ9NUS  XM5
timestamp 1756981609
transform 1 0 3766 0 1 -10
box -290 -290 290 290
use pfet_03v3_PQ9NUS  XM6
timestamp 1756981609
transform 1 0 4286 0 1 -70
box -290 -290 290 290
use nfet_03v3_KVLVYL  XM7
timestamp 1756981609
transform 1 0 5474 0 1 -110
box -958 -310 958 310
use nfet_03v3_KVLVYL  XM8
timestamp 1756981609
transform 1 0 7330 0 1 -170
box -958 -310 958 310
use nfet_03v3_RPTYYZ  XM9
timestamp 1756981609
transform 1 0 10780 0 1 2406
box -820 -266 820 266
use nfet_03v3_RPTYYZ  XM10
timestamp 1756981609
transform 1 0 12300 0 1 2406
box -820 -266 820 266
use nfet_03v3_KTKMNW  XM11
timestamp 1756981609
transform 1 0 12230 0 1 -370
box -290 -290 290 290
use pfet_03v3_PQ9NUS  XM12
timestamp 1756981609
transform 1 0 12750 0 1 -430
box -290 -290 290 290
use pfet_03v3_75ANUS  XM13
timestamp 1756981609
transform 1 0 13362 0 1 -490
box -382 -290 382 290
use pfet_03v3_9LZZ5X  XM14
timestamp 1756981609
transform 1 0 14250 0 1 -550
box -566 -290 566 290
use pfet_03v3_9LZZ5X  XM15
timestamp 1756981609
transform 1 0 15322 0 1 -610
box -566 -290 566 290
use pfet_03v3_PQ9NUS  XM16
timestamp 1756981609
transform 1 0 16118 0 1 -670
box -290 -290 290 290
use pfet_03v3_75ANUS  XM17
timestamp 1756981609
transform 1 0 16730 0 1 -730
box -382 -290 382 290
use pfet_03v3_9LZZ5X  XM18
timestamp 1756981609
transform 1 0 17618 0 1 -790
box -566 -290 566 290
use pfet_03v3_9LZZ5X  XM19
timestamp 1756981609
transform 1 0 18690 0 1 -850
box -566 -290 566 290
use nfet_03v3_RPTYYZ  XM20
timestamp 1756981609
transform 1 0 10780 0 1 3366
box -820 -266 820 266
use pfet_03v3_9LZZ5X  XM22
timestamp 1756981609
transform 1 0 23474 0 1 -1030
box -566 -290 566 290
use pfet_03v3_9LZZ5X  XM23
timestamp 1756981609
transform 1 0 24546 0 1 -1090
box -566 -290 566 290
<< end >>
