* NGSPICE file created from nor2.ext - technology: (null)

.subckt nor2 VDD VSS OUT A B
X0 a_2130_n110 A.t0 VDD.t5 VDD.t4 pfet_03v3
**devattr s=52800,1376 d=31200,704
X1 OUT.t2 B.t0 VSS.t1 VSS.t0 nfet_03v3
**devattr s=17600,576 d=17600,576
X2 VSS.t3 A.t1 OUT.t3 VSS.t2 nfet_03v3
**devattr s=17600,576 d=17600,576
X3 OUT.t1 B.t1 a_2130_n110 VDD.t1 pfet_03v3
**devattr s=31200,704 d=52800,1376
X4 VDD.t3 A.t2 a_2130_n110 VDD.t2 pfet_03v3
**devattr s=31200,704 d=52800,1376
X5 a_2130_n110 B.t2 OUT.t0 VDD.t0 pfet_03v3
**devattr s=52800,1376 d=31200,704
R0 A.n0 A.t2 34.2311
R1 A.n0 A.t0 34.011
R2 A.n1 A.t1 19.6529
R3 A A.n1 5.0495
R4 A.n1 A.n0 0.096125
R5 VDD.t1 VDD.n3 236.083
R6 VDD.n6 VDD.t4 236.083
R7 VDD.n5 VDD.t0 235.294
R8 VDD.t2 VDD.n5 235.294
R9 VDD.t0 VDD.t1 200
R10 VDD.t4 VDD.t2 200
R11 VDD.n3 VDD.n1 96.0755
R12 VDD.n6 VDD.n1 96.0755
R13 VDD.n6 VDD.n2 96.0755
R14 VDD.n3 VDD.n2 96.0755
R15 VDD.n4 VDD.n1 36.2255
R16 VDD.n4 VDD.n2 36.2255
R17 VDD.n3 VDD 2.09318
R18 VDD.n7 VDD.t5 1.47383
R19 VDD.n0 VDD.t3 1.47383
R20 VDD.n8 VDD.n7 0.868843
R21 VDD.n4 VDD.n0 0.788
R22 VDD.n5 VDD.n4 0.788
R23 VDD.n7 VDD.n6 0.788
R24 VDD.n8 VDD.n0 0.561043
R25 VDD.n8 VDD 0.00095
R26 B.n0 B.t1 34.2311
R27 B.n0 B.t2 34.011
R28 B.n1 B.t0 19.5066
R29 B B.n1 6.15163
R30 B.n1 B.n0 0.242375
R31 VSS.n2 VSS.t0 849.126
R32 VSS.n9 VSS.t2 849.126
R33 VSS.n7 VSS.t0 847.827
R34 VSS.t2 VSS.n8 847.827
R35 VSS.n8 VSS.n7 720.653
R36 VSS.n6 VSS.n2 44.1404
R37 VSS.n9 VSS.n1 44.1404
R38 VSS.n3 VSS.t3 4.84702
R39 VSS.n5 VSS.t1 4.84702
R40 VSS.n2 VSS.n0 2.16892
R41 VSS VSS.n9 2.16712
R42 VSS.n6 VSS.n5 1.3005
R43 VSS.n7 VSS.n6 1.3005
R44 VSS.n3 VSS.n1 1.3005
R45 VSS.n8 VSS.n1 1.3005
R46 VSS.n4 VSS.n0 0.073981
R47 VSS.n5 VSS.n4 0.0258591
R48 VSS.n4 VSS.n3 0.0258591
R49 VSS VSS.n0 0.0023
R50 OUT.n1 OUT.t3 10.3401
R51 OUT.n1 OUT.t2 9.2885
R52 OUT.n0 OUT.t0 4.09202
R53 OUT.n0 OUT.t1 3.95079
R54 OUT.n2 OUT.n1 0.599711
R55 OUT.n2 OUT.n0 0.296375
R56 OUT OUT.n2 0.254429
.ends

