magic
tech gf180mcuD
magscale 1 10
timestamp 1755272603
<< checkpaint >>
rect -1974 1160 2582 2500
rect -2810 1040 2582 1160
rect -2810 980 2738 1040
rect -2810 920 3234 980
rect -2870 -3840 3234 920
rect -2870 -3900 3174 -3840
rect -2374 -3960 3174 -3900
rect -1878 -4020 3174 -3960
rect -1382 -4080 3174 -4020
<< error_s >>
rect 109 417 196 446
rect 26 268 86 360
rect 270 323 281 369
rect 327 323 338 334
rect -226 183 -215 229
rect -169 183 -158 194
rect -96 0 -89 46
rect -272 -48 -249 -37
rect -135 -48 -112 -37
rect -50 -48 -43 0
rect -226 -129 -215 -83
rect 26 -120 97 268
rect 201 0 246 246
rect 224 -108 247 -97
rect 361 -108 384 -97
rect 26 -260 86 -120
rect 270 -189 281 -143
rect -323 -937 -291 -891
rect -566 -1017 -555 -971
rect -509 -1017 -498 -1006
rect -325 -1040 -291 -992
rect -277 -1040 -245 -937
rect -46 -983 159 -954
rect 173 -960 205 -951
rect 173 -997 242 -960
rect -612 -1448 -589 -1437
rect -475 -1448 -452 -1437
rect -566 -1529 -555 -1483
rect -277 -1520 -243 -1040
rect -70 -1077 -59 -1031
rect 0 -1077 44 -1000
rect 182 -1052 251 -997
rect 171 -1100 251 -1052
rect 669 -1057 701 -1011
rect -116 -1508 -93 -1497
rect -277 -1623 -245 -1520
rect -70 -1589 -59 -1543
rect 0 -1589 44 -1497
rect 182 -1580 253 -1100
rect 426 -1137 437 -1091
rect 483 -1137 494 -1126
rect 667 -1160 701 -1112
rect 715 -1160 747 -1057
rect 380 -1568 403 -1557
rect 517 -1568 540 -1557
rect 0 -1600 159 -1591
rect 182 -1683 251 -1580
rect 426 -1649 437 -1603
rect 715 -1640 749 -1160
rect 922 -1197 933 -1151
rect 979 -1197 990 -1186
rect 876 -1628 899 -1617
rect 1013 -1628 1036 -1617
rect 182 -1720 242 -1683
rect 715 -1743 747 -1640
rect 922 -1709 933 -1663
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
<< metal2 >>
rect -750 1430 570 1540
rect -750 520 -630 1430
rect 480 1270 570 1430
rect 1060 610 1150 810
rect 470 540 1150 610
rect 470 520 550 540
rect -750 410 -100 520
rect -40 410 550 520
rect -750 -370 -630 410
rect 480 310 550 410
rect 1060 -370 1150 -160
rect -750 -450 1160 -370
use inv_test  x1
timestamp 1755272338
transform 1 0 -50 0 1 1000
box -420 -1320 632 246
use nfet_03v3_AUBTWU  XM1
timestamp 1755271904
transform 1 0 -592 0 1 -1490
box -278 -410 278 410
use pfet_03v3_NE88KN  XM2
timestamp 1755271904
transform 1 0 896 0 1 -1670
box -278 -410 278 410
use nfet_03v3_AUBTWU  XM3
timestamp 1755271904
transform 1 0 -96 0 1 -1550
box -278 -410 278 410
use pfet_03v3_NE88KN  XM4
timestamp 1755271904
transform 1 0 400 0 1 -1610
box -278 -410 278 410
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 sw_vout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 sw_bit
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 sw_Vref
port 4 nsew
<< end >>
