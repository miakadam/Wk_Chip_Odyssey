magic
tech gf180mcuD
magscale 1 10
timestamp 1758003743
<< nwell >>
rect 1780 -320 3268 700
<< pwell >>
rect 1780 -1040 2380 -420
rect 2464 -510 3064 -420
rect 2464 -768 3110 -510
rect 2464 -1040 3064 -768
<< nmos >>
rect 2030 -830 2130 -630
rect 2714 -830 2814 -630
<< pmos >>
rect 2030 -110 2130 490
rect 2234 -110 2334 490
rect 2714 -110 2814 490
rect 2918 -110 3018 490
<< ndiff >>
rect 1942 -643 2030 -630
rect 1942 -817 1955 -643
rect 2001 -817 2030 -643
rect 1942 -830 2030 -817
rect 2130 -643 2218 -630
rect 2130 -817 2159 -643
rect 2205 -817 2218 -643
rect 2130 -830 2218 -817
rect 2626 -643 2714 -630
rect 2626 -817 2639 -643
rect 2685 -817 2714 -643
rect 2626 -830 2714 -817
rect 2814 -643 2902 -630
rect 2814 -817 2843 -643
rect 2889 -817 2902 -643
rect 2814 -830 2902 -817
<< pdiff >>
rect 1942 477 2030 490
rect 1942 -97 1955 477
rect 2001 -97 2030 477
rect 1942 -110 2030 -97
rect 2130 477 2234 490
rect 2130 -97 2159 477
rect 2205 -97 2234 477
rect 2130 -110 2234 -97
rect 2334 477 2422 490
rect 2334 -97 2363 477
rect 2409 -97 2422 477
rect 2334 -110 2422 -97
rect 2626 477 2714 490
rect 2626 -97 2639 477
rect 2685 -97 2714 477
rect 2626 -110 2714 -97
rect 2814 477 2918 490
rect 2814 -97 2843 477
rect 2889 -97 2918 477
rect 2814 -110 2918 -97
rect 3018 477 3106 490
rect 3018 -97 3047 477
rect 3093 -97 3106 477
rect 3018 -110 3106 -97
<< ndiffc >>
rect 1955 -817 2001 -643
rect 2159 -817 2205 -643
rect 2639 -817 2685 -643
rect 2843 -817 2889 -643
<< pdiffc >>
rect 1955 -97 2001 477
rect 2159 -97 2205 477
rect 2363 -97 2409 477
rect 2639 -97 2685 477
rect 2843 -97 2889 477
rect 3047 -97 3093 477
<< psubdiff >>
rect 1804 -516 2356 -444
rect 1804 -560 1876 -516
rect 1804 -900 1817 -560
rect 1863 -900 1876 -560
rect 2284 -560 2356 -516
rect 1804 -944 1876 -900
rect 2284 -900 2297 -560
rect 2343 -900 2356 -560
rect 2284 -944 2356 -900
rect 1804 -1016 2356 -944
rect 2488 -516 3040 -444
rect 2488 -560 2560 -516
rect 2488 -900 2501 -560
rect 2547 -900 2560 -560
rect 2968 -560 3040 -516
rect 2488 -944 2560 -900
rect 2968 -900 2981 -560
rect 3027 -900 3040 -560
rect 2968 -944 3040 -900
rect 2488 -1016 3040 -944
<< nsubdiff >>
rect 1804 604 3244 676
rect 1804 560 1876 604
rect 1804 -180 1817 560
rect 1863 -180 1876 560
rect 2488 560 2560 604
rect 1804 -224 1876 -180
rect 2488 -180 2501 560
rect 2547 -180 2560 560
rect 3172 560 3244 604
rect 2488 -224 2560 -180
rect 3172 -180 3185 560
rect 3231 -180 3244 560
rect 3172 -224 3244 -180
rect 1804 -296 3244 -224
<< psubdiffcont >>
rect 1817 -900 1863 -560
rect 2297 -900 2343 -560
rect 2501 -900 2547 -560
rect 2981 -900 3027 -560
<< nsubdiffcont >>
rect 1817 -180 1863 560
rect 2501 -180 2547 560
rect 3185 -180 3231 560
<< polysilicon >>
rect 2030 569 2130 582
rect 2030 523 2043 569
rect 2117 523 2130 569
rect 2030 490 2130 523
rect 2234 569 2334 582
rect 2234 523 2247 569
rect 2321 523 2334 569
rect 2234 490 2334 523
rect 2030 -143 2130 -110
rect 2030 -189 2043 -143
rect 2117 -189 2130 -143
rect 2030 -202 2130 -189
rect 2234 -143 2334 -110
rect 2234 -189 2247 -143
rect 2321 -189 2334 -143
rect 2234 -202 2334 -189
rect 2714 569 2814 582
rect 2714 523 2727 569
rect 2801 523 2814 569
rect 2714 490 2814 523
rect 2918 569 3018 582
rect 2918 523 2931 569
rect 3005 523 3018 569
rect 2918 490 3018 523
rect 2714 -143 2814 -110
rect 2714 -189 2727 -143
rect 2801 -189 2814 -143
rect 2714 -202 2814 -189
rect 2918 -143 3018 -110
rect 2918 -189 2931 -143
rect 3005 -189 3018 -143
rect 2918 -202 3018 -189
rect 2030 -551 2130 -538
rect 2030 -597 2043 -551
rect 2117 -597 2130 -551
rect 2030 -630 2130 -597
rect 2030 -863 2130 -830
rect 2030 -909 2043 -863
rect 2117 -909 2130 -863
rect 2030 -922 2130 -909
rect 2714 -551 2814 -538
rect 2714 -597 2727 -551
rect 2801 -597 2814 -551
rect 2714 -630 2814 -597
rect 2714 -863 2814 -830
rect 2714 -909 2727 -863
rect 2801 -909 2814 -863
rect 2714 -922 2814 -909
<< polycontact >>
rect 2043 523 2117 569
rect 2247 523 2321 569
rect 2043 -189 2117 -143
rect 2247 -189 2321 -143
rect 2727 523 2801 569
rect 2931 523 3005 569
rect 2727 -189 2801 -143
rect 2931 -189 3005 -143
rect 2043 -597 2117 -551
rect 2043 -909 2117 -863
rect 2727 -597 2801 -551
rect 2727 -909 2801 -863
<< metal1 >>
rect 1780 700 3268 900
rect 1817 560 1863 700
rect 2032 569 2128 600
rect 2032 523 2043 569
rect 2117 523 2128 569
rect 2236 569 2332 600
rect 2236 523 2247 569
rect 2321 523 2332 569
rect 2501 560 2547 700
rect 1863 477 2001 488
rect 2159 477 2205 488
rect 2363 477 2501 488
rect 1863 -97 1955 477
rect 2142 237 2154 477
rect 2210 237 2222 477
rect 1863 -108 2001 -97
rect 2159 -108 2205 -97
rect 2409 -97 2501 477
rect 2363 -108 2501 -97
rect 1817 -191 1863 -180
rect 2032 -189 2043 -143
rect 2117 -163 2128 -143
rect 2236 -163 2247 -143
rect 2117 -189 2247 -163
rect 2321 -189 2332 -143
rect 2032 -216 2332 -189
rect 2716 569 2812 600
rect 2716 523 2727 569
rect 2801 523 2812 569
rect 2920 569 3016 600
rect 2920 523 2931 569
rect 3005 523 3016 569
rect 3185 560 3231 700
rect 2639 477 2685 488
rect 2843 477 2889 488
rect 3047 477 3093 488
rect 2826 237 2838 477
rect 2894 237 2906 477
rect 2622 -97 2634 143
rect 2690 -97 2702 143
rect 3030 -97 3042 143
rect 3098 -97 3110 143
rect 2639 -108 2685 -97
rect 2843 -108 2889 -97
rect 3047 -108 3093 -97
rect 2501 -191 2547 -180
rect 2716 -189 2727 -143
rect 2801 -163 2812 -143
rect 2920 -163 2931 -143
rect 2801 -189 2931 -163
rect 3005 -189 3016 -143
rect 2716 -216 3016 -189
rect 3185 -191 3231 -180
rect 2032 -264 2128 -216
rect 2032 -320 2052 -264
rect 2108 -320 2128 -264
rect 1817 -560 1863 -549
rect 2032 -551 2128 -320
rect 2716 -420 2812 -216
rect 2716 -476 2736 -420
rect 2792 -476 2812 -420
rect 2032 -597 2043 -551
rect 2117 -597 2128 -551
rect 2297 -560 2547 -549
rect 1955 -643 2001 -632
rect 1938 -702 1955 -692
rect 2159 -643 2297 -632
rect 2001 -702 2018 -692
rect 1938 -758 1950 -702
rect 2006 -758 2018 -702
rect 1938 -768 1955 -758
rect 2001 -768 2018 -758
rect 1955 -828 2001 -817
rect 2205 -817 2297 -643
rect 2159 -828 2297 -817
rect 1817 -1040 1863 -900
rect 2032 -909 2043 -863
rect 2117 -909 2128 -863
rect 2032 -940 2128 -909
rect 2343 -900 2501 -560
rect 2716 -551 2812 -476
rect 2716 -597 2727 -551
rect 2801 -597 2812 -551
rect 2981 -560 3027 -549
rect 2547 -643 2685 -632
rect 2547 -817 2639 -643
rect 2843 -643 2889 -632
rect 2826 -702 2843 -692
rect 2889 -702 2906 -692
rect 2826 -758 2838 -702
rect 2894 -758 2906 -702
rect 2826 -768 2843 -758
rect 2547 -828 2685 -817
rect 2889 -768 2906 -758
rect 2843 -828 2889 -817
rect 2297 -911 2547 -900
rect 2716 -909 2727 -863
rect 2801 -909 2812 -863
rect 2343 -1040 2501 -911
rect 2716 -940 2812 -909
rect 2981 -1040 3027 -900
rect 1780 -1240 3064 -1040
<< via1 >>
rect 2154 237 2159 477
rect 2159 237 2205 477
rect 2205 237 2210 477
rect 2838 237 2843 477
rect 2843 237 2889 477
rect 2889 237 2894 477
rect 2634 -97 2639 143
rect 2639 -97 2685 143
rect 2685 -97 2690 143
rect 3042 -97 3047 143
rect 3047 -97 3093 143
rect 3093 -97 3098 143
rect 2052 -320 2108 -264
rect 2736 -476 2792 -420
rect 1950 -758 1955 -702
rect 1955 -758 2001 -702
rect 2001 -758 2006 -702
rect 2838 -758 2843 -702
rect 2843 -758 2889 -702
rect 2889 -758 2894 -702
<< metal2 >>
rect 2142 477 2906 487
rect 2142 237 2154 477
rect 2210 237 2838 477
rect 2894 237 2906 477
rect 2142 227 2906 237
rect 2622 143 3110 153
rect 2622 -97 2634 143
rect 2690 -97 3042 143
rect 3098 -97 3110 143
rect 2622 -107 3110 -97
rect 2032 -264 2128 -252
rect 1724 -320 2052 -264
rect 2108 -320 2128 -264
rect 2032 -332 2128 -320
rect 3030 -342 3110 -107
rect 3030 -398 3268 -342
rect 2716 -420 2812 -410
rect 1724 -476 2736 -420
rect 2792 -476 2812 -420
rect 2716 -486 2812 -476
rect 3030 -692 3110 -398
rect 1938 -702 3110 -692
rect 1938 -758 1950 -702
rect 2006 -758 2838 -702
rect 2894 -758 3110 -702
rect 1938 -768 3110 -758
<< labels >>
rlabel metal1 2525 900 2525 900 1 VDD
port 0 n
rlabel metal1 2418 -1240 2418 -1240 5 VSS
port 1 s
rlabel metal2 3268 -371 3268 -371 3 OUT
port 2 e
rlabel metal2 1724 -291 1724 -291 7 A
port 3 w
rlabel metal2 1724 -448 1724 -448 7 B
port 4 w
<< end >>
