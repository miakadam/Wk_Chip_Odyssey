* NGSPICE file created from nand2.ext - technology: (null)

.subckt nand2 VDD OUT A B VSS
X0 a_1640_n650 A.t0 OUT.t2 VSS.t3 nfet_03v3
**devattr s=17600,576 d=10400,304
X1 VDD.t1 B.t0 OUT.t3 VDD.t0 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X2 VSS.t1 B.t1 a_1640_n650 VSS.t0 nfet_03v3
**devattr s=10400,304 d=17600,576
X3 OUT.t0 A.t1 VDD.t3 VDD.t2 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X4 OUT.t1 A.t2 a_1640_n650 VSS.t2 nfet_03v3
**devattr s=10400,304 d=17600,576
X5 a_1640_n650 B.t2 VSS.t5 VSS.t4 nfet_03v3
**devattr s=17600,576 d=10400,304
R0 A.n1 A.t1 34.2529
R1 A.n0 A.t0 19.673
R2 A.n0 A.t2 19.4007
R3 A A.n1 6.43968
R4 A.n1 A.n0 0.106438
R5 OUT.n1 OUT.t2 18.7717
R6 OUT.n1 OUT.t1 9.2885
R7 OUT.n0 OUT.t3 4.23346
R8 OUT.n0 OUT.t0 3.85546
R9 OUT.n2 OUT.n1 0.4055
R10 OUT.n2 OUT.n0 0.352625
R11 OUT OUT.n2 0.254429
R12 VSS.n6 VSS.n5 61574.7
R13 VSS.t2 VSS.n3 849.126
R14 VSS.n5 VSS.t3 847.827
R15 VSS.n5 VSS.t0 847.827
R16 VSS.n6 VSS.t4 847.827
R17 VSS.t3 VSS.t2 720.653
R18 VSS.t0 VSS.t4 720.653
R19 VSS.n3 VSS.n1 87.3061
R20 VSS.n3 VSS.n2 87.3061
R21 VSS.n7 VSS.n1 87.3061
R22 VSS.n7 VSS.n2 87.3061
R23 VSS.n4 VSS.n1 20.8061
R24 VSS.n4 VSS.n2 20.8061
R25 VSS.n0 VSS.t1 4.7885
R26 VSS.n8 VSS.t5 4.7885
R27 VSS.n3 VSS 2.21437
R28 VSS.n4 VSS.n0 1.3005
R29 VSS.n5 VSS.n4 1.3005
R30 VSS.n8 VSS.n7 1.3005
R31 VSS.n7 VSS.n6 1.3005
R32 VSS.n9 VSS.n8 0.771017
R33 VSS.n9 VSS.n0 0.463217
R34 VSS.n9 VSS 0.00095
R35 B.n1 B.t0 34.1066
R36 B.n0 B.t1 19.673
R37 B.n0 B.t2 19.4007
R38 B B.n1 5.09932
R39 B.n1 B.n0 0.252687
R40 VDD.n1 VDD.t0 131.589
R41 VDD.n0 VDD.t2 131.589
R42 VDD.n1 VDD.t1 1.49467
R43 VDD.n0 VDD.t3 1.49467
R44 VDD VDD.n3 0.14689
R45 VDD.n2 VDD.n0 0.0313054
R46 VDD.n2 VDD.n1 0.0313054
R47 VDD VDD.n2 0.00224757
.ends

