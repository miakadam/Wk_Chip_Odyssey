magic
tech gf180mcuD
magscale 1 10
timestamp 1757409273
<< pwell >>
rect -958 -410 958 410
<< nmos >>
rect -708 -200 -508 200
rect -404 -200 -204 200
rect -100 -200 100 200
rect 204 -200 404 200
rect 508 -200 708 200
<< ndiff >>
rect -796 187 -708 200
rect -796 -187 -783 187
rect -737 -187 -708 187
rect -796 -200 -708 -187
rect -508 187 -404 200
rect -508 -187 -479 187
rect -433 -187 -404 187
rect -508 -200 -404 -187
rect -204 187 -100 200
rect -204 -187 -175 187
rect -129 -187 -100 187
rect -204 -200 -100 -187
rect 100 187 204 200
rect 100 -187 129 187
rect 175 -187 204 187
rect 100 -200 204 -187
rect 404 187 508 200
rect 404 -187 433 187
rect 479 -187 508 187
rect 404 -200 508 -187
rect 708 187 796 200
rect 708 -187 737 187
rect 783 -187 796 187
rect 708 -200 796 -187
<< ndiffc >>
rect -783 -187 -737 187
rect -479 -187 -433 187
rect -175 -187 -129 187
rect 129 -187 175 187
rect 433 -187 479 187
rect 737 -187 783 187
<< psubdiff >>
rect -934 314 934 386
rect -934 270 -862 314
rect -934 -270 -921 270
rect -875 -270 -862 270
rect 862 270 934 314
rect -934 -314 -862 -270
rect 862 -270 875 270
rect 921 -270 934 270
rect 862 -314 934 -270
rect -934 -386 934 -314
<< psubdiffcont >>
rect -921 -270 -875 270
rect 875 -270 921 270
<< polysilicon >>
rect -708 279 -508 292
rect -708 233 -695 279
rect -521 233 -508 279
rect -708 200 -508 233
rect -404 279 -204 292
rect -404 233 -391 279
rect -217 233 -204 279
rect -404 200 -204 233
rect -100 279 100 292
rect -100 233 -87 279
rect 87 233 100 279
rect -100 200 100 233
rect 204 279 404 292
rect 204 233 217 279
rect 391 233 404 279
rect 204 200 404 233
rect 508 279 708 292
rect 508 233 521 279
rect 695 233 708 279
rect 508 200 708 233
rect -708 -233 -508 -200
rect -708 -279 -695 -233
rect -521 -279 -508 -233
rect -708 -292 -508 -279
rect -404 -233 -204 -200
rect -404 -279 -391 -233
rect -217 -279 -204 -233
rect -404 -292 -204 -279
rect -100 -233 100 -200
rect -100 -279 -87 -233
rect 87 -279 100 -233
rect -100 -292 100 -279
rect 204 -233 404 -200
rect 204 -279 217 -233
rect 391 -279 404 -233
rect 204 -292 404 -279
rect 508 -233 708 -200
rect 508 -279 521 -233
rect 695 -279 708 -233
rect 508 -292 708 -279
<< polycontact >>
rect -695 233 -521 279
rect -391 233 -217 279
rect -87 233 87 279
rect 217 233 391 279
rect 521 233 695 279
rect -695 -279 -521 -233
rect -391 -279 -217 -233
rect -87 -279 87 -233
rect 217 -279 391 -233
rect 521 -279 695 -233
<< metal1 >>
rect -921 270 -875 281
rect -706 233 -695 279
rect -521 233 -510 279
rect -402 233 -391 279
rect -217 233 -206 279
rect -98 233 -87 279
rect 87 233 98 279
rect 206 233 217 279
rect 391 233 402 279
rect 510 233 521 279
rect 695 233 706 279
rect 875 270 921 281
rect -783 187 -737 198
rect -783 -198 -737 -187
rect -479 187 -433 198
rect -479 -198 -433 -187
rect -175 187 -129 198
rect -175 -198 -129 -187
rect 129 187 175 198
rect 129 -198 175 -187
rect 433 187 479 198
rect 433 -198 479 -187
rect 737 187 783 198
rect 737 -198 783 -187
rect -921 -281 -875 -270
rect -706 -279 -695 -233
rect -521 -279 -510 -233
rect -402 -279 -391 -233
rect -217 -279 -206 -233
rect -98 -279 -87 -233
rect 87 -279 98 -233
rect 206 -279 217 -233
rect 391 -279 402 -233
rect 510 -279 521 -233
rect 695 -279 706 -233
rect 875 -281 921 -270
<< properties >>
string FIXED_BBOX -898 -350 898 350
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
