** sch_path: /foss/designs/comparator/rslatch.sch
.subckt rslatch VDD Vout1 Vout2 Vin1 Vin2 VSS
*.PININFO VDD:B VSS:B Vin1:B Vin2:B Vout1:B Vout2:B
XM1 Vout1 Vin1 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM2 Vout2 Vin2 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM3 Vout1 Vout2 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
XM4 Vout2 Vout1 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
.ends
