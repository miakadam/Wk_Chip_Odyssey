magic
tech gf180mcuD
magscale 1 10
timestamp 1758099403
<< metal1 >>
rect 12038 19089 12108 19101
rect 19896 19089 19966 19091
rect 12038 19033 12050 19089
rect 12106 19033 19898 19089
rect 19954 19033 19966 19089
rect 12038 19031 12108 19033
rect 19896 19031 19966 19033
rect 16080 18913 16150 18925
rect 23938 18913 24008 18915
rect 16080 18857 16092 18913
rect 16148 18857 23940 18913
rect 23996 18857 24008 18913
rect 16080 18855 16150 18857
rect 23938 18855 24008 18857
rect 3900 18737 3970 18749
rect 11758 18737 11828 18739
rect 3900 18681 3912 18737
rect 3968 18681 11760 18737
rect 11816 18681 11828 18737
rect 3900 18679 3970 18681
rect 11758 18679 11828 18681
rect 20122 18737 20192 18749
rect 27980 18737 28050 18739
rect 20122 18681 20134 18737
rect 20190 18681 27982 18737
rect 28038 18681 28050 18737
rect 20122 18679 20192 18681
rect 27980 18679 28050 18681
rect 7996 18561 8066 18573
rect 15854 18561 15924 18563
rect 7996 18505 8008 18561
rect 8064 18505 15856 18561
rect 15912 18505 15924 18561
rect 7996 18503 8066 18505
rect 15854 18503 15924 18505
rect 24164 18561 24234 18573
rect 32022 18561 32092 18573
rect 24164 18505 24176 18561
rect 24232 18505 32024 18561
rect 32080 18505 32092 18561
rect 24164 18503 24234 18505
rect 32022 18503 32092 18505
rect 3546 17311 3616 17323
rect 3546 17255 3558 17311
rect 3614 17255 4088 17311
rect 7558 17308 7628 17320
rect 11600 17308 11670 17320
rect 15642 17308 15712 17320
rect 19684 17308 19754 17320
rect 23726 17308 23796 17320
rect 27768 17308 27848 17320
rect 3546 17253 3616 17255
rect 7558 17252 7570 17308
rect 7626 17252 8100 17308
rect 11600 17252 11612 17308
rect 11668 17252 12142 17308
rect 15642 17252 15654 17308
rect 15710 17252 16184 17308
rect 19684 17252 19696 17308
rect 19752 17252 20226 17308
rect 23726 17252 23738 17308
rect 23794 17252 24268 17308
rect 27768 17252 27780 17308
rect 27836 17252 28310 17308
rect 7558 17250 7628 17252
rect 11600 17250 11670 17252
rect 15642 17250 15712 17252
rect 19684 17250 19754 17252
rect 23726 17250 23796 17252
rect 27768 17250 27848 17252
rect 7704 14990 7774 14992
rect 7210 14934 7706 14990
rect 7762 14934 7774 14990
rect 11758 14987 11828 14999
rect 15854 14987 15924 14999
rect 19896 14987 19966 14999
rect 23938 14987 24008 14999
rect 27980 14987 28050 14999
rect 32022 14987 32092 14999
rect 7704 14922 7774 14934
rect 11210 14931 11760 14987
rect 11816 14931 11828 14987
rect 15306 14931 15856 14987
rect 15912 14931 15924 14987
rect 19348 14931 19898 14987
rect 19954 14931 19966 14987
rect 23390 14931 23940 14987
rect 23996 14931 24008 14987
rect 27432 14931 27982 14987
rect 28038 14931 28050 14987
rect 31474 14931 32024 14987
rect 32080 14931 32092 14987
rect 11758 14919 11828 14931
rect 15854 14919 15924 14931
rect 19896 14919 19966 14931
rect 23938 14919 24008 14931
rect 27980 14919 28050 14931
rect 32022 14919 32092 14931
rect 3900 14088 3970 14090
rect 3900 14032 3912 14088
rect 3968 14032 4024 14088
rect 7996 14085 8066 14087
rect 12038 14085 12108 14087
rect 16080 14085 16150 14087
rect 20122 14085 20192 14087
rect 24164 14085 24234 14087
rect 28162 14085 28240 14097
rect 3900 14020 3970 14032
rect 7996 14029 8008 14085
rect 8064 14029 8074 14085
rect 12038 14029 12050 14085
rect 12106 14029 12116 14085
rect 16080 14029 16092 14085
rect 16148 14029 16158 14085
rect 20122 14029 20134 14085
rect 20190 14029 20200 14085
rect 24164 14029 24176 14085
rect 24232 14029 24242 14085
rect 28162 14029 28173 14085
rect 28229 14029 28276 14085
rect 7996 14017 8066 14029
rect 12038 14017 12108 14029
rect 16080 14017 16150 14029
rect 20122 14017 20192 14029
rect 24164 14017 24234 14029
rect 28162 14017 28240 14029
rect 3274 10464 3344 10476
rect 3274 10408 3286 10464
rect 3342 10408 4078 10464
rect 7286 10461 7356 10473
rect 11328 10461 11398 10473
rect 15370 10461 15440 10473
rect 19412 10461 19482 10473
rect 23454 10461 23524 10473
rect 28162 10461 28240 10473
rect 3274 10396 3344 10408
rect 7286 10405 7298 10461
rect 7354 10405 8090 10461
rect 11328 10405 11340 10461
rect 11396 10405 12132 10461
rect 15370 10405 15382 10461
rect 15438 10405 16174 10461
rect 19412 10405 19424 10461
rect 19480 10405 20216 10461
rect 23454 10405 23466 10461
rect 23522 10405 24258 10461
rect 28162 10405 28173 10461
rect 28229 10405 28277 10461
rect 7286 10393 7356 10405
rect 11328 10393 11398 10405
rect 15370 10393 15440 10405
rect 19412 10393 19482 10405
rect 23454 10393 23524 10405
rect 28162 10393 28240 10405
rect 3818 9677 3888 9689
rect 3818 9621 3830 9677
rect 3886 9621 4098 9677
rect 7830 9674 7900 9686
rect 11872 9674 11942 9686
rect 15914 9674 15984 9686
rect 19956 9674 20026 9686
rect 23998 9674 24068 9686
rect 28040 9674 28110 9686
rect 3818 9619 3888 9621
rect 7830 9618 7842 9674
rect 7898 9618 8110 9674
rect 11872 9618 11884 9674
rect 11940 9618 12152 9674
rect 15914 9618 15926 9674
rect 15982 9618 16194 9674
rect 19956 9618 19968 9674
rect 20024 9618 20236 9674
rect 23998 9618 24010 9674
rect 24066 9618 24278 9674
rect 28040 9618 28052 9674
rect 28108 9618 28354 9674
rect 7830 9616 7900 9618
rect 11872 9616 11942 9618
rect 15914 9616 15984 9618
rect 19956 9616 20026 9618
rect 23998 9616 24068 9618
rect 28040 9606 28110 9618
rect -58 7732 12 7744
rect 4010 7732 4096 7744
rect -58 7676 -46 7732
rect 10 7676 20 7732
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect -58 7664 12 7676
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 3222 5355 4022 5411
rect 7222 5355 8034 5411
rect 11276 5355 12076 5411
rect 15318 5355 16118 5411
rect 19360 5355 20160 5411
rect 23402 5355 24202 5411
rect 3966 5233 4022 5355
rect 7978 5233 8034 5355
rect 12020 5233 12076 5355
rect 16062 5233 16118 5355
rect 20104 5233 20160 5355
rect 24146 5233 24202 5355
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect -330 4509 -260 4521
rect 3682 4509 3752 4521
rect 7694 4509 7764 4521
rect 11736 4509 11806 4521
rect 15778 4509 15848 4521
rect 19820 4509 19890 4521
rect 23862 4509 23932 4521
rect -330 4453 -318 4509
rect -262 4453 418 4509
rect 3682 4453 3694 4509
rect 3750 4453 4032 4509
rect 7694 4453 7706 4509
rect 7762 4453 8080 4509
rect 11736 4453 11748 4509
rect 11804 4453 12107 4509
rect 15778 4453 15790 4509
rect 15846 4453 16149 4509
rect 19820 4453 19832 4509
rect 19888 4453 20191 4509
rect 23862 4453 23874 4509
rect 23930 4453 24236 4509
rect -330 4441 -260 4453
rect 3682 4441 3752 4453
rect 7694 4441 7764 4453
rect 11736 4441 11806 4453
rect 15778 4441 15848 4453
rect 19820 4441 19890 4453
rect 23862 4441 23932 4453
rect -121 885 -41 897
rect 3954 885 4024 897
rect 7966 885 8046 897
rect 12008 885 12088 897
rect 16050 885 16130 897
rect 20092 885 20172 897
rect 24134 885 24214 897
rect -121 829 -109 885
rect -53 829 90 885
rect 3954 829 3966 885
rect 4022 829 4032 885
rect 7966 829 7978 885
rect 8034 829 8081 885
rect 12008 829 12020 885
rect 12076 829 12111 885
rect 16050 829 16062 885
rect 16118 829 16149 885
rect 20092 829 20104 885
rect 20160 829 20191 885
rect 24134 829 24146 885
rect 24202 829 24239 885
rect -121 817 -41 829
rect 3954 817 4024 829
rect 7966 817 8046 829
rect 12008 817 12088 829
rect 16050 817 16130 829
rect 20092 817 20172 829
rect 24134 817 24214 829
rect -121 98 -35 110
rect 3818 98 3888 110
rect 7830 98 7900 110
rect 11872 98 11942 110
rect 15914 98 15984 110
rect 19956 98 20026 110
rect 23998 98 24068 110
rect -121 42 -109 98
rect -53 42 27 98
rect 3818 42 3830 98
rect 3886 42 4039 98
rect 7830 42 7842 98
rect 7898 42 8081 98
rect 11872 42 11884 98
rect 11940 42 12123 98
rect 15914 42 15926 98
rect 15982 42 16165 98
rect 19956 42 19968 98
rect 20024 42 20207 98
rect 23998 42 24010 98
rect 24066 42 24249 98
rect -121 30 -35 42
rect 3818 30 3888 42
rect 7830 30 7900 42
rect 11872 30 11942 42
rect 15914 30 15984 42
rect 19956 30 20026 42
rect 23998 30 24068 42
<< via1 >>
rect 12050 19033 12106 19089
rect 19898 19033 19954 19089
rect 16092 18857 16148 18913
rect 23940 18857 23996 18913
rect 3912 18681 3968 18737
rect 11760 18681 11816 18737
rect 20134 18681 20190 18737
rect 27982 18681 28038 18737
rect 8008 18505 8064 18561
rect 15856 18505 15912 18561
rect 24176 18505 24232 18561
rect 32024 18505 32080 18561
rect 3558 17255 3614 17311
rect 7570 17252 7626 17308
rect 11612 17252 11668 17308
rect 15654 17252 15710 17308
rect 19696 17252 19752 17308
rect 23738 17252 23794 17308
rect 27780 17252 27836 17308
rect 7706 14934 7762 14990
rect 11760 14931 11816 14987
rect 15856 14931 15912 14987
rect 19898 14931 19954 14987
rect 23940 14931 23996 14987
rect 27982 14931 28038 14987
rect 32024 14931 32080 14987
rect 3912 14032 3968 14088
rect 8008 14029 8064 14085
rect 12050 14029 12106 14085
rect 16092 14029 16148 14085
rect 20134 14029 20190 14085
rect 24176 14029 24232 14085
rect 28173 14029 28229 14085
rect 3286 10408 3342 10464
rect 7298 10405 7354 10461
rect 11340 10405 11396 10461
rect 15382 10405 15438 10461
rect 19424 10405 19480 10461
rect 23466 10405 23522 10461
rect 28173 10405 28229 10461
rect 3830 9621 3886 9677
rect 7842 9618 7898 9674
rect 11884 9618 11940 9674
rect 15926 9618 15982 9674
rect 19968 9618 20024 9674
rect 24010 9618 24066 9674
rect 28052 9618 28108 9674
rect -46 7676 10 7732
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect 3966 5167 4022 5223
rect 7978 5167 8034 5223
rect 12020 5167 12076 5223
rect 16062 5167 16118 5223
rect 20104 5167 20160 5223
rect 24146 5167 24202 5223
rect -318 4453 -262 4509
rect 3694 4453 3750 4509
rect 7706 4453 7762 4509
rect 11748 4453 11804 4509
rect 15790 4453 15846 4509
rect 19832 4453 19888 4509
rect 23874 4453 23930 4509
rect -109 829 -53 885
rect 3966 829 4022 885
rect 7978 829 8034 885
rect 12020 829 12076 885
rect 16062 829 16118 885
rect 20104 829 20160 885
rect 24146 829 24202 885
rect -109 42 -53 98
rect 3830 42 3886 98
rect 7842 42 7898 98
rect 11884 42 11940 98
rect 15926 42 15982 98
rect 19968 42 20024 98
rect 24010 42 24066 98
<< metal2 >>
rect 3900 18737 3970 18749
rect 3900 18681 3912 18737
rect 3968 18681 3970 18737
rect 3900 18679 3970 18681
rect 3546 17311 3616 17323
rect 3546 17255 3558 17311
rect 3614 17255 3616 17311
rect 3546 17253 3616 17255
rect 3274 10464 3344 10476
rect 3274 10408 3286 10464
rect 3342 10408 3344 10464
rect 3274 10396 3344 10408
rect -201 9514 10 9524
rect -201 9414 -46 9514
rect -201 9404 10 9414
rect 3286 9514 3342 10396
rect 3286 9404 3342 9414
rect -201 9004 10 9014
rect -201 8904 -46 9004
rect -201 8894 10 8904
rect -46 7744 10 8894
rect -58 7732 12 7744
rect -58 7676 -46 7732
rect 10 7676 12 7732
rect -58 7664 12 7676
rect -330 4509 -260 4521
rect -330 4453 -318 4509
rect -262 4453 -260 4509
rect -330 4441 -260 4453
rect -318 -55 -262 4441
rect 3558 3207 3614 17253
rect 3912 14090 3968 18679
rect 7558 17308 7628 17320
rect 7558 17252 7570 17308
rect 7626 17252 7628 17308
rect 7558 17250 7628 17252
rect 3900 14088 3970 14090
rect 3900 14032 3912 14088
rect 3968 14032 3970 14088
rect 3900 14020 3970 14032
rect 7286 10461 7356 10473
rect 7286 10405 7298 10461
rect 7354 10405 7356 10461
rect 7286 10393 7356 10405
rect 3818 9677 3888 9689
rect 3818 9621 3830 9677
rect 3886 9621 3888 9677
rect 3818 9619 3888 9621
rect 3830 9007 3886 9619
rect 7298 9514 7354 10393
rect 7298 9404 7354 9414
rect 3682 4509 3752 4521
rect 3682 4453 3694 4509
rect 3750 4453 3752 4509
rect 3682 4441 3752 4453
rect 3478 3151 3614 3207
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect -473 -65 -262 -55
rect -473 -165 -318 -65
rect -473 -175 -262 -165
rect 3694 -65 3750 4441
rect 3830 110 3886 8907
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 3966 897 4022 5165
rect 7570 3207 7626 17250
rect 7706 14992 7762 19504
rect 11760 18739 11816 19501
rect 12038 19089 12108 19101
rect 12038 19033 12050 19089
rect 12106 19033 12108 19089
rect 12038 19031 12108 19033
rect 11758 18737 11828 18739
rect 11758 18681 11760 18737
rect 11816 18681 11828 18737
rect 11758 18679 11828 18681
rect 7996 18561 8066 18573
rect 7996 18505 8008 18561
rect 8064 18505 8066 18561
rect 7996 18503 8066 18505
rect 7704 14990 7774 14992
rect 7704 14934 7706 14990
rect 7762 14934 7774 14990
rect 7704 14922 7774 14934
rect 8008 14087 8064 18503
rect 11600 17308 11670 17320
rect 11600 17252 11612 17308
rect 11668 17252 11670 17308
rect 11600 17250 11670 17252
rect 7996 14085 8066 14087
rect 7996 14029 8008 14085
rect 8064 14029 8066 14085
rect 7996 14017 8066 14029
rect 11328 10461 11398 10473
rect 11328 10405 11340 10461
rect 11396 10405 11398 10461
rect 11328 10393 11398 10405
rect 7830 9674 7900 9686
rect 7830 9618 7842 9674
rect 7898 9618 7900 9674
rect 7830 9616 7900 9618
rect 7842 9004 7898 9616
rect 11340 9514 11396 10393
rect 11340 9404 11396 9414
rect 7694 4509 7764 4521
rect 7694 4453 7706 4509
rect 7762 4453 7764 4509
rect 7694 4441 7764 4453
rect 7490 3151 7626 3207
rect 3954 885 4024 897
rect 3954 829 3966 885
rect 4022 829 4024 885
rect 3954 817 4024 829
rect 3818 98 3888 110
rect 3818 42 3830 98
rect 3886 42 3888 98
rect 3818 30 3888 42
rect 3694 -175 3750 -165
rect 7706 -65 7762 4441
rect 7842 110 7898 8904
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 7978 897 8034 5165
rect 11612 3207 11668 17250
rect 11760 14999 11816 18679
rect 11758 14987 11828 14999
rect 11758 14931 11760 14987
rect 11816 14931 11828 14987
rect 11758 14919 11828 14931
rect 12050 14087 12106 19031
rect 15856 18563 15912 19501
rect 19898 19091 19954 19501
rect 19896 19089 19966 19091
rect 19896 19033 19898 19089
rect 19954 19033 19966 19089
rect 19896 19031 19966 19033
rect 16080 18913 16150 18925
rect 16080 18857 16092 18913
rect 16148 18857 16150 18913
rect 16080 18855 16150 18857
rect 15854 18561 15924 18563
rect 15854 18505 15856 18561
rect 15912 18505 15924 18561
rect 15854 18503 15924 18505
rect 15642 17308 15712 17320
rect 15642 17252 15654 17308
rect 15710 17252 15712 17308
rect 15642 17250 15712 17252
rect 12038 14085 12108 14087
rect 12038 14029 12050 14085
rect 12106 14029 12108 14085
rect 12038 14017 12108 14029
rect 15370 10461 15440 10473
rect 15370 10405 15382 10461
rect 15438 10405 15440 10461
rect 15370 10393 15440 10405
rect 11872 9674 11942 9686
rect 11872 9618 11884 9674
rect 11940 9618 11942 9674
rect 11872 9616 11942 9618
rect 11884 9004 11940 9616
rect 15382 9514 15438 10393
rect 15382 9404 15438 9414
rect 11736 4509 11806 4521
rect 11736 4453 11748 4509
rect 11804 4453 11806 4509
rect 11736 4441 11806 4453
rect 11532 3151 11668 3207
rect 7966 885 8046 897
rect 7966 829 7978 885
rect 8034 829 8046 885
rect 7966 817 8046 829
rect 7830 98 7900 110
rect 7830 42 7842 98
rect 7898 42 7900 98
rect 7830 30 7900 42
rect 7706 -175 7762 -165
rect 11748 -65 11804 4441
rect 11884 110 11940 8904
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 12020 897 12076 5165
rect 15654 3207 15710 17250
rect 15856 14999 15912 18503
rect 15854 14987 15924 14999
rect 15854 14931 15856 14987
rect 15912 14931 15924 14987
rect 15854 14919 15924 14931
rect 16092 14087 16148 18855
rect 19684 17308 19754 17320
rect 19684 17252 19696 17308
rect 19752 17252 19754 17308
rect 19684 17250 19754 17252
rect 16080 14085 16150 14087
rect 16080 14029 16092 14085
rect 16148 14029 16150 14085
rect 16080 14017 16150 14029
rect 19412 10461 19482 10473
rect 19412 10405 19424 10461
rect 19480 10405 19482 10461
rect 19412 10393 19482 10405
rect 15914 9674 15984 9686
rect 15914 9618 15926 9674
rect 15982 9618 15984 9674
rect 15914 9616 15984 9618
rect 15926 9004 15982 9616
rect 19424 9514 19480 10393
rect 19424 9404 19480 9414
rect 15778 4509 15848 4521
rect 15778 4453 15790 4509
rect 15846 4453 15848 4509
rect 15778 4441 15848 4453
rect 15574 3151 15710 3207
rect 12008 885 12088 897
rect 12008 829 12020 885
rect 12076 829 12088 885
rect 12008 817 12088 829
rect 11872 98 11942 110
rect 11872 42 11884 98
rect 11940 42 11942 98
rect 11872 30 11942 42
rect 11748 -175 11804 -165
rect 15790 -65 15846 4441
rect 15926 110 15982 8904
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 16062 897 16118 5165
rect 19696 3207 19752 17250
rect 19898 14999 19954 19031
rect 23940 18915 23996 19504
rect 23938 18913 24008 18915
rect 23938 18857 23940 18913
rect 23996 18857 24008 18913
rect 23938 18855 24008 18857
rect 20122 18737 20192 18749
rect 20122 18681 20134 18737
rect 20190 18681 20192 18737
rect 20122 18679 20192 18681
rect 19896 14987 19966 14999
rect 19896 14931 19898 14987
rect 19954 14931 19966 14987
rect 19896 14919 19966 14931
rect 20134 14087 20190 18679
rect 23726 17308 23796 17320
rect 23726 17252 23738 17308
rect 23794 17252 23796 17308
rect 23726 17250 23796 17252
rect 20122 14085 20192 14087
rect 20122 14029 20134 14085
rect 20190 14029 20192 14085
rect 20122 14017 20192 14029
rect 23454 10461 23524 10473
rect 23454 10405 23466 10461
rect 23522 10405 23524 10461
rect 23454 10393 23524 10405
rect 19956 9674 20026 9686
rect 19956 9618 19968 9674
rect 20024 9618 20026 9674
rect 19956 9616 20026 9618
rect 19968 9004 20024 9616
rect 23466 9514 23522 10393
rect 23466 9404 23522 9414
rect 19820 4509 19890 4521
rect 19820 4453 19832 4509
rect 19888 4453 19890 4509
rect 19820 4441 19890 4453
rect 19616 3151 19752 3207
rect 16050 885 16130 897
rect 16050 829 16062 885
rect 16118 829 16130 885
rect 16050 817 16130 829
rect 15914 98 15984 110
rect 15914 42 15926 98
rect 15982 42 15984 98
rect 15914 30 15984 42
rect 15790 -175 15846 -165
rect 19832 -65 19888 4441
rect 19968 110 20024 8904
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 20104 897 20160 5165
rect 23738 3207 23794 17250
rect 23940 14999 23996 18855
rect 27982 18739 28038 19501
rect 27980 18737 28050 18739
rect 27980 18681 27982 18737
rect 28038 18681 28050 18737
rect 27980 18679 28050 18681
rect 24164 18561 24234 18573
rect 24164 18505 24176 18561
rect 24232 18505 24234 18561
rect 24164 18503 24234 18505
rect 23938 14987 24008 14999
rect 23938 14931 23940 14987
rect 23996 14931 24008 14987
rect 23938 14919 24008 14931
rect 24176 14087 24232 18503
rect 27768 17308 27848 17320
rect 27768 17252 27780 17308
rect 27836 17252 27848 17308
rect 27768 17250 27848 17252
rect 24164 14085 24234 14087
rect 24164 14029 24176 14085
rect 24232 14029 24234 14085
rect 24164 14017 24234 14029
rect 23998 9674 24068 9686
rect 23998 9618 24010 9674
rect 24066 9618 24068 9674
rect 23998 9616 24068 9618
rect 24010 9004 24066 9616
rect 23862 4509 23932 4521
rect 23862 4453 23874 4509
rect 23930 4453 23932 4509
rect 23862 4441 23932 4453
rect 23658 3151 23794 3207
rect 20092 885 20172 897
rect 20092 829 20104 885
rect 20160 829 20172 885
rect 20092 817 20172 829
rect 19956 98 20026 110
rect 19956 42 19968 98
rect 20024 42 20026 98
rect 19956 30 20026 42
rect 19832 -175 19888 -165
rect 23874 -65 23930 4441
rect 24010 110 24066 8904
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect 24146 897 24202 5165
rect 27780 3207 27836 17250
rect 27982 14999 28038 18679
rect 32022 18561 32092 18573
rect 32022 18505 32024 18561
rect 32080 18505 32092 18561
rect 32022 18503 32092 18505
rect 32024 14999 32080 18503
rect 27980 14987 28050 14999
rect 27980 14931 27982 14987
rect 28038 14931 28050 14987
rect 27980 14919 28050 14931
rect 32022 14987 32092 14999
rect 32022 14931 32024 14987
rect 32080 14931 32092 14987
rect 32022 14919 32092 14931
rect 28162 14085 28240 14097
rect 28162 14029 28173 14085
rect 28229 14029 28240 14085
rect 28162 14017 28240 14029
rect 28162 10461 28240 10473
rect 28162 10405 28173 10461
rect 28229 10405 28240 10461
rect 28162 10393 28240 10405
rect 28040 9674 28110 9686
rect 28040 9618 28052 9674
rect 28108 9618 28110 9674
rect 28040 9606 28110 9618
rect 28052 9004 28108 9606
rect 28052 8894 28108 8904
rect 27608 3151 27836 3207
rect 24134 885 24214 897
rect 24134 829 24146 885
rect 24202 829 24214 885
rect 24134 817 24214 829
rect 23998 98 24068 110
rect 23998 42 24010 98
rect 24066 42 24068 98
rect 23998 30 24068 42
rect 23874 -175 23930 -165
<< via2 >>
rect -46 9414 10 9514
rect 3286 9414 3342 9514
rect -46 8904 10 9004
rect 7298 9414 7354 9514
rect 3830 8907 3886 9007
rect -109 829 -53 885
rect -109 42 -53 98
rect -318 -165 -262 -65
rect 4022 7676 4078 7732
rect 11340 9414 11396 9514
rect 7842 8904 7898 9004
rect 3694 -165 3750 -65
rect 8064 7676 8120 7732
rect 15382 9414 15438 9514
rect 11884 8904 11940 9004
rect 7706 -165 7762 -65
rect 12106 7676 12162 7732
rect 19424 9414 19480 9514
rect 15926 8904 15982 9004
rect 11748 -165 11804 -65
rect 16148 7676 16204 7732
rect 23466 9414 23522 9514
rect 19968 8904 20024 9004
rect 15790 -165 15846 -65
rect 20190 7676 20246 7732
rect 24010 8904 24066 9004
rect 19832 -165 19888 -65
rect 24232 7676 24288 7732
rect 28173 14029 28229 14085
rect 28173 10405 28229 10461
rect 28052 8904 28108 9004
rect 23874 -165 23930 -65
<< metal3 >>
rect 28162 14085 28240 14097
rect 28162 14029 28173 14085
rect 28229 14029 28240 14085
rect 28162 14017 28240 14029
rect 28162 10461 28240 10473
rect 28162 10405 28173 10461
rect 28229 10405 28240 10461
rect 28162 10393 28240 10405
rect -56 9414 -46 9514
rect 10 9414 3286 9514
rect 3342 9414 7298 9514
rect 7354 9414 11340 9514
rect 11396 9414 15382 9514
rect 15438 9414 19424 9514
rect 19480 9414 23466 9514
rect 23522 9414 23532 9514
rect 3820 9004 3830 9007
rect -56 8904 -46 9004
rect 10 8907 3830 9004
rect 3886 9004 3896 9007
rect 3886 8907 7842 9004
rect 10 8904 7842 8907
rect 7898 8904 11884 9004
rect 11940 8904 15926 9004
rect 15982 8904 19968 9004
rect 20024 8904 24010 9004
rect 24066 8904 28052 9004
rect 28108 8904 28118 9004
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect -328 -165 -318 -65
rect -262 -165 3694 -65
rect 3750 -165 7706 -65
rect 7762 -165 11748 -65
rect 11804 -165 15790 -65
rect 15846 -165 19832 -65
rect 19888 -165 23874 -65
rect 23930 -165 23940 -65
<< via3 >>
rect 28173 14029 28229 14085
rect 28173 10405 28229 10461
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect -109 829 -53 885
rect -109 42 -53 98
<< metal4 >>
rect 7460 9609 8202 18385
rect 4100 9606 8202 9609
rect 11502 9606 12244 18385
rect 15544 9606 16286 18385
rect 19586 9606 20328 18385
rect 23628 9606 24370 18385
rect 27670 14177 28412 18385
rect 27670 14085 28419 14177
rect 27670 14029 28173 14085
rect 28229 14029 28419 14085
rect 27670 14017 28419 14029
rect 27670 10473 28412 14017
rect 27670 10461 28417 10473
rect 27670 10405 28173 10461
rect 28229 10405 28417 10461
rect 27670 10313 28417 10405
rect 27670 9606 28412 10313
rect 4100 8809 27730 9606
rect 3448 7824 4160 8809
rect 7460 7824 8202 8809
rect 11502 7824 12244 8809
rect 15544 7824 16286 8809
rect 19586 7824 20328 8809
rect 23628 7824 24370 8809
rect 3448 7584 3930 7824
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 7460 7584 7972 7824
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 11502 7584 12014 7824
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 15544 7584 16056 7824
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 19586 7584 20098 7824
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 23628 7584 24140 7824
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect -121 885 156 897
rect -121 829 -109 885
rect -53 829 156 885
rect -121 737 156 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect 3448 30 4160 7584
rect 7460 30 8202 7584
rect 11502 30 12244 7584
rect 15544 30 16286 7584
rect 19586 30 20328 7584
rect 23628 30 24370 7584
<< via4 >>
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect -109 42 -53 98
<< metal5 >>
rect 7460 9609 8202 18385
rect 4100 9606 8202 9609
rect 11502 9606 12244 18385
rect 15544 9606 16286 18385
rect 19586 9606 20328 18385
rect 23628 9606 24370 18385
rect 27670 14177 28412 18385
rect 27670 13937 28082 14177
rect 28320 13937 28412 14177
rect 27670 10553 28412 13937
rect 27670 10313 28080 10553
rect 28322 10313 28412 10553
rect 27670 9606 28412 10313
rect 4100 8809 27730 9606
rect 3448 7732 4160 8809
rect 3448 7676 4022 7732
rect 4078 7676 4160 7732
rect -121 98 167 190
rect -121 42 -109 98
rect -53 42 167 98
rect -121 30 167 42
rect 3448 30 4160 7676
rect 7460 7732 8202 8809
rect 7460 7676 8064 7732
rect 8120 7676 8202 7732
rect 7460 30 8202 7676
rect 11502 7732 12244 8809
rect 11502 7676 12106 7732
rect 12162 7676 12244 7732
rect 11502 30 12244 7676
rect 15544 7732 16286 8809
rect 15544 7676 16148 7732
rect 16204 7676 16286 7732
rect 15544 30 16286 7676
rect 19586 7732 20328 8809
rect 19586 7676 20190 7732
rect 20246 7676 20328 7732
rect 19586 30 20328 7676
rect 20344 7664 20350 7744
rect 23628 7732 24370 8809
rect 23628 7676 24232 7732
rect 24288 7676 24370 7732
rect 23628 30 24370 7676
use dffrs  dffrs_0
timestamp 1758085300
transform 1 0 4870 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_1
timestamp 1758085300
transform 1 0 8912 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_2
timestamp 1758085300
transform 1 0 12954 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_3
timestamp 1758085300
transform 1 0 16996 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_4
timestamp 1758085300
transform 1 0 21038 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_5
timestamp 1758085300
transform 1 0 25080 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_7
timestamp 1758085300
transform 1 0 8912 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_8
timestamp 1758085300
transform 1 0 12954 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_9
timestamp 1758085300
transform 1 0 16996 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_10
timestamp 1758085300
transform 1 0 21038 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_11
timestamp 1758085300
transform 1 0 25080 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_12
timestamp 1758085300
transform 1 0 29122 0 1 15504
box -848 -5898 2620 2881
use dffrs  dffrs_13
timestamp 1758085300
transform 1 0 858 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_14
timestamp 1758085300
transform 1 0 4870 0 1 15507
box -848 -5898 2620 2881
<< labels >>
rlabel metal2 -473 -113 -473 -113 7 clk
port 2 w
rlabel metal2 -201 8954 -201 8954 7 reset
port 3 w
rlabel metal2 -201 9462 -201 9462 7 comp_in
port 4 w
rlabel metal2 7734 19504 7734 19504 1 d5
port 5 n
rlabel metal2 11789 19501 11789 19501 1 d4
port 6 n
rlabel metal2 15885 19501 15885 19501 1 d3
port 7 n
rlabel metal2 19926 19501 19926 19501 1 d2
port 8 n
rlabel metal2 23968 19504 23968 19504 1 d1
port 9 n
rlabel metal2 28012 19501 28012 19501 1 d0
port 10 n
rlabel metal5 19630 18385 19630 18385 1 vdd
port 0 n
rlabel metal4 15578 30 15578 30 5 vss
port 1 s
<< end >>
