magic
tech gf180mcuD
magscale 1 10
timestamp 1758262485
<< nwell >>
rect 16712 1249 16724 1269
rect 17860 1249 17870 1269
rect 16644 1189 16724 1193
<< pwell >>
rect 17579 558 17679 563
rect 18468 -524 18548 -402
rect 14770 -2740 19206 -524
rect 14770 -2764 16514 -2740
rect 14770 -2836 16538 -2764
rect 14770 -3320 16514 -2836
rect 17052 -3004 17108 -2740
rect 17462 -2764 19206 -2740
rect 17438 -2836 19206 -2764
rect 16847 -3199 17127 -3163
rect 16847 -3200 17134 -3199
rect 16842 -3219 17134 -3200
rect 17462 -3320 19206 -2836
<< nmos >>
rect 15216 -2324 15416 -2024
rect 15520 -2324 15720 -2024
rect 15824 -2324 16024 -2024
rect 16128 -2324 16328 -2024
rect 16432 -2324 16632 -2024
rect 16736 -2324 16936 -2024
rect 17040 -2324 17240 -2024
rect 17344 -2324 17544 -2024
rect 17648 -2324 17848 -2024
rect 17952 -2324 18152 -2024
rect 18256 -2324 18456 -2024
rect 18560 -2324 18760 -2024
<< ndiff >>
rect 15128 -2037 15216 -2024
rect 15128 -2311 15141 -2037
rect 15187 -2311 15216 -2037
rect 15128 -2324 15216 -2311
rect 15416 -2037 15520 -2024
rect 15416 -2311 15445 -2037
rect 15491 -2311 15520 -2037
rect 15416 -2324 15520 -2311
rect 15720 -2037 15824 -2024
rect 15720 -2311 15749 -2037
rect 15795 -2311 15824 -2037
rect 15720 -2324 15824 -2311
rect 16024 -2037 16128 -2024
rect 16024 -2311 16053 -2037
rect 16099 -2311 16128 -2037
rect 16024 -2324 16128 -2311
rect 16328 -2037 16432 -2024
rect 16328 -2311 16357 -2037
rect 16403 -2311 16432 -2037
rect 16328 -2324 16432 -2311
rect 16632 -2037 16736 -2024
rect 16632 -2311 16661 -2037
rect 16707 -2311 16736 -2037
rect 16632 -2324 16736 -2311
rect 16936 -2037 17040 -2024
rect 16936 -2311 16965 -2037
rect 17011 -2311 17040 -2037
rect 16936 -2324 17040 -2311
rect 17240 -2037 17344 -2024
rect 17240 -2311 17269 -2037
rect 17315 -2311 17344 -2037
rect 17240 -2324 17344 -2311
rect 17544 -2037 17648 -2024
rect 17544 -2311 17573 -2037
rect 17619 -2311 17648 -2037
rect 17544 -2324 17648 -2311
rect 17848 -2037 17952 -2024
rect 17848 -2311 17877 -2037
rect 17923 -2311 17952 -2037
rect 17848 -2324 17952 -2311
rect 18152 -2037 18256 -2024
rect 18152 -2311 18181 -2037
rect 18227 -2311 18256 -2037
rect 18152 -2324 18256 -2311
rect 18456 -2037 18560 -2024
rect 18456 -2311 18485 -2037
rect 18531 -2311 18560 -2037
rect 18456 -2324 18560 -2311
rect 18760 -2037 18848 -2024
rect 18760 -2311 18789 -2037
rect 18835 -2311 18848 -2037
rect 18760 -2324 18848 -2311
<< pdiff >>
rect 16712 1249 16724 1269
rect 17860 1249 17870 1269
<< ndiffc >>
rect 15141 -2311 15187 -2037
rect 15445 -2311 15491 -2037
rect 15749 -2311 15795 -2037
rect 16053 -2311 16099 -2037
rect 16357 -2311 16403 -2037
rect 16661 -2311 16707 -2037
rect 16965 -2311 17011 -2037
rect 17269 -2311 17315 -2037
rect 17573 -2311 17619 -2037
rect 17877 -2311 17923 -2037
rect 18181 -2311 18227 -2037
rect 18485 -2311 18531 -2037
rect 18789 -2311 18835 -2037
<< psubdiff >>
rect 17579 558 17679 563
rect 14795 -621 19181 -549
rect 14795 -720 14995 -621
rect 14795 -1220 14845 -720
rect 14945 -1220 14995 -720
rect 14795 -2165 14995 -1220
rect 18981 -720 19181 -621
rect 18981 -1220 19031 -720
rect 19131 -1220 19181 -720
rect 14795 -2665 14845 -2165
rect 14945 -2665 14995 -2165
rect 18981 -2165 19181 -1220
rect 14795 -2764 14995 -2665
rect 18981 -2665 19031 -2165
rect 19131 -2665 19181 -2165
rect 18981 -2764 19181 -2665
rect 14795 -2836 16538 -2764
rect 17438 -2836 19181 -2764
<< psubdiffcont >>
rect 14845 -1220 14945 -720
rect 19031 -1220 19131 -720
rect 14845 -2665 14945 -2165
rect 19031 -2665 19131 -2165
<< polysilicon >>
rect 15878 -1445 15968 -1375
rect 15878 -1455 15968 -1450
rect 15216 -1945 15416 -1932
rect 15216 -1991 15229 -1945
rect 15403 -1991 15416 -1945
rect 15216 -2024 15416 -1991
rect 15520 -1945 15720 -1932
rect 15520 -1991 15533 -1945
rect 15707 -1991 15720 -1945
rect 15520 -2024 15720 -1991
rect 15824 -1945 16024 -1932
rect 15824 -1991 15837 -1945
rect 16011 -1991 16024 -1945
rect 15824 -2024 16024 -1991
rect 16128 -1945 16328 -1932
rect 16128 -1991 16141 -1945
rect 16315 -1991 16328 -1945
rect 16128 -2024 16328 -1991
rect 16432 -1945 16632 -1932
rect 16432 -1991 16445 -1945
rect 16619 -1991 16632 -1945
rect 16432 -2024 16632 -1991
rect 16736 -1945 16936 -1932
rect 16736 -1991 16749 -1945
rect 16923 -1991 16936 -1945
rect 16736 -2024 16936 -1991
rect 17040 -1945 17240 -1932
rect 17040 -1991 17053 -1945
rect 17227 -1991 17240 -1945
rect 17040 -2024 17240 -1991
rect 17344 -1945 17544 -1932
rect 17344 -1991 17357 -1945
rect 17531 -1991 17544 -1945
rect 17344 -2024 17544 -1991
rect 17648 -1945 17848 -1932
rect 17648 -1991 17661 -1945
rect 17835 -1991 17848 -1945
rect 17648 -2024 17848 -1991
rect 17952 -1945 18152 -1932
rect 17952 -1991 17965 -1945
rect 18139 -1991 18152 -1945
rect 17952 -2024 18152 -1991
rect 18256 -1945 18456 -1932
rect 18256 -1991 18269 -1945
rect 18443 -1991 18456 -1945
rect 18256 -2024 18456 -1991
rect 18560 -1945 18760 -1932
rect 18560 -1991 18573 -1945
rect 18747 -1991 18760 -1945
rect 18560 -2024 18760 -1991
rect 15216 -2357 15416 -2324
rect 15216 -2403 15229 -2357
rect 15403 -2403 15416 -2357
rect 15216 -2416 15416 -2403
rect 15520 -2357 15720 -2324
rect 15520 -2403 15533 -2357
rect 15707 -2403 15720 -2357
rect 15520 -2416 15720 -2403
rect 15824 -2357 16024 -2324
rect 15824 -2403 15837 -2357
rect 16011 -2403 16024 -2357
rect 15824 -2416 16024 -2403
rect 16128 -2357 16328 -2324
rect 16128 -2403 16141 -2357
rect 16315 -2403 16328 -2357
rect 16128 -2416 16328 -2403
rect 16432 -2357 16632 -2324
rect 16432 -2403 16445 -2357
rect 16619 -2403 16632 -2357
rect 16432 -2416 16632 -2403
rect 16736 -2357 16936 -2324
rect 16736 -2403 16749 -2357
rect 16923 -2403 16936 -2357
rect 16736 -2416 16936 -2403
rect 17040 -2357 17240 -2324
rect 17040 -2403 17053 -2357
rect 17227 -2403 17240 -2357
rect 17040 -2416 17240 -2403
rect 17344 -2357 17544 -2324
rect 17344 -2403 17357 -2357
rect 17531 -2403 17544 -2357
rect 17344 -2416 17544 -2403
rect 17648 -2357 17848 -2324
rect 17648 -2403 17661 -2357
rect 17835 -2403 17848 -2357
rect 17648 -2416 17848 -2403
rect 17952 -2357 18152 -2324
rect 17952 -2403 17965 -2357
rect 18139 -2403 18152 -2357
rect 17952 -2416 18152 -2403
rect 18256 -2357 18456 -2324
rect 18256 -2403 18269 -2357
rect 18443 -2403 18456 -2357
rect 18256 -2416 18456 -2403
rect 18560 -2357 18760 -2324
rect 18560 -2403 18573 -2357
rect 18747 -2403 18760 -2357
rect 18560 -2416 18760 -2403
<< polycontact >>
rect 15229 -1991 15403 -1945
rect 15533 -1991 15707 -1945
rect 15837 -1991 16011 -1945
rect 16141 -1991 16315 -1945
rect 16445 -1991 16619 -1945
rect 16749 -1991 16923 -1945
rect 17053 -1991 17227 -1945
rect 17357 -1991 17531 -1945
rect 17661 -1991 17835 -1945
rect 17965 -1991 18139 -1945
rect 18269 -1991 18443 -1945
rect 18573 -1991 18747 -1945
rect 15229 -2403 15403 -2357
rect 15533 -2403 15707 -2357
rect 15837 -2403 16011 -2357
rect 16141 -2403 16315 -2357
rect 16445 -2403 16619 -2357
rect 16749 -2403 16923 -2357
rect 17053 -2403 17227 -2357
rect 17357 -2403 17531 -2357
rect 17661 -2403 17835 -2357
rect 17965 -2403 18139 -2357
rect 18269 -2403 18443 -2357
rect 18573 -2403 18747 -2357
<< metal1 >>
rect 13758 2115 13862 2129
rect 20114 2115 20218 2127
rect 13758 2039 13770 2115
rect 13850 2039 20126 2115
rect 20206 2039 20218 2115
rect 13758 2029 13862 2039
rect 14202 1439 14278 2039
rect 15062 1439 15138 2039
rect 15826 1459 16326 1515
rect 16434 1459 16934 1515
rect 17042 1459 17542 1515
rect 17650 1459 18150 1515
rect 18838 1439 18914 2039
rect 19698 1439 19774 2039
rect 20114 2027 20218 2039
rect 15732 1360 15812 1362
rect 14032 1347 14188 1349
rect 14032 1213 14120 1347
rect 14176 1213 14188 1347
rect 14032 1211 14188 1213
rect 14292 1347 14372 1349
rect 14292 1213 14304 1347
rect 14360 1213 14372 1347
rect 14292 1211 14372 1213
rect 14430 1347 14510 1349
rect 14430 1213 14442 1347
rect 14498 1213 14510 1347
rect 14430 1211 14510 1213
rect 14891 1347 15048 1349
rect 14891 1213 14980 1347
rect 15036 1213 15048 1347
rect 14891 1211 15048 1213
rect 15152 1347 15232 1349
rect 15152 1213 15164 1347
rect 15220 1213 15232 1347
rect 15152 1211 15232 1213
rect 15290 1347 15370 1349
rect 15290 1213 15302 1347
rect 15358 1213 15370 1347
rect 15732 1216 15744 1360
rect 15800 1216 15812 1360
rect 16340 1360 16420 1362
rect 15732 1214 15812 1216
rect 16036 1259 16116 1269
rect 15290 1211 15370 1213
rect 16036 1203 16048 1259
rect 16104 1203 16116 1259
rect 16340 1216 16352 1360
rect 16408 1216 16420 1360
rect 16948 1360 17028 1362
rect 16340 1214 16420 1216
rect 16644 1259 16724 1269
rect 16036 1193 16116 1203
rect 16644 1203 16656 1259
rect 16712 1203 16724 1259
rect 16948 1216 16960 1360
rect 17016 1216 17028 1360
rect 17556 1360 17636 1362
rect 16948 1214 17028 1216
rect 17252 1259 17332 1269
rect 16644 1193 16724 1203
rect 17252 1203 17264 1259
rect 17320 1203 17332 1259
rect 17556 1216 17568 1360
rect 17624 1216 17636 1360
rect 18164 1360 18244 1362
rect 17556 1214 17636 1216
rect 17860 1259 17940 1269
rect 17252 1193 17332 1203
rect 17860 1203 17872 1259
rect 17928 1203 17940 1259
rect 18164 1216 18176 1360
rect 18232 1216 18244 1360
rect 18164 1214 18244 1216
rect 18606 1347 18686 1349
rect 18606 1213 18618 1347
rect 18674 1213 18686 1347
rect 18606 1211 18686 1213
rect 18744 1347 18824 1349
rect 18744 1213 18756 1347
rect 18812 1213 18824 1347
rect 18744 1211 18824 1213
rect 18928 1347 19084 1349
rect 18928 1213 18940 1347
rect 18996 1213 19084 1347
rect 18928 1211 19084 1213
rect 19466 1347 19546 1349
rect 19466 1213 19478 1347
rect 19534 1213 19546 1347
rect 19466 1211 19546 1213
rect 19604 1347 19684 1349
rect 19604 1213 19616 1347
rect 19672 1213 19684 1347
rect 19604 1211 19684 1213
rect 19788 1347 19944 1349
rect 19788 1213 19800 1347
rect 19856 1213 19944 1347
rect 19788 1211 19944 1213
rect 17860 1193 17940 1203
rect 16839 1152 16919 1162
rect 14202 1091 14278 1121
rect 15062 1091 15138 1121
rect 16022 1101 16130 1136
rect 15886 1090 16326 1101
rect 16839 1096 16851 1152
rect 16907 1096 16919 1152
rect 14618 844 14722 856
rect 15140 844 15244 854
rect 15886 844 15990 1090
rect 16839 1086 16919 1096
rect 17057 1152 17137 1162
rect 17057 1096 17069 1152
rect 17125 1096 17137 1152
rect 17846 1101 17954 1136
rect 17986 1101 18090 1102
rect 17057 1086 17137 1096
rect 17650 1090 18090 1101
rect 18838 1091 18914 1121
rect 19698 1091 19774 1121
rect 16494 844 16734 852
rect 14618 760 14630 844
rect 14710 760 15152 844
rect 15232 842 16734 844
rect 15232 762 15898 842
rect 15978 762 16506 842
rect 16586 762 16644 842
rect 16724 762 16734 842
rect 15232 760 16734 762
rect 14618 750 14722 760
rect 15140 750 15244 760
rect 15886 748 15990 760
rect 16494 748 16734 760
rect 17240 844 17482 852
rect 17986 844 18090 1090
rect 18732 844 18836 854
rect 19254 844 19358 854
rect 17240 842 18744 844
rect 17240 762 17252 842
rect 17332 762 17390 842
rect 17470 762 17998 842
rect 18078 762 18744 842
rect 17240 760 18744 762
rect 18824 760 19266 844
rect 19346 760 19358 844
rect 17240 748 17482 760
rect 17986 749 18090 760
rect 18732 750 18836 760
rect 19254 750 19358 760
rect 15688 548 16492 563
rect 15688 503 16307 548
rect 16297 468 16307 503
rect 16387 503 16492 548
rect 17484 548 18288 563
rect 17484 503 17589 548
rect 16387 468 16397 503
rect 17579 468 17589 503
rect 17669 503 18288 548
rect 17669 468 17679 503
rect 17711 411 17757 422
rect 18319 411 18365 422
rect 15898 404 15978 406
rect 15898 260 15910 404
rect 15966 260 15978 404
rect 15898 258 15978 260
rect 16506 404 16586 406
rect 16506 260 16518 404
rect 16574 260 16586 404
rect 16506 258 16586 260
rect 17390 404 17470 406
rect 17390 260 17402 404
rect 17458 260 17470 404
rect 17390 258 17470 260
rect 17998 404 18078 406
rect 17998 260 18010 404
rect 18066 260 18078 404
rect 17998 258 18078 260
rect 15594 188 15674 190
rect 15152 98 15232 108
rect 15152 -46 15164 98
rect 15220 -46 15232 98
rect 15594 44 15606 188
rect 15662 44 15674 188
rect 15594 42 15674 44
rect 16202 188 16282 190
rect 16202 44 16214 188
rect 16270 44 16282 188
rect 16202 42 16282 44
rect 17694 188 17711 190
rect 17757 188 17774 190
rect 17694 44 17706 188
rect 17762 44 17774 188
rect 17694 42 17711 44
rect 17757 42 17774 44
rect 18302 188 18319 190
rect 18365 188 18382 190
rect 18302 44 18314 188
rect 18370 44 18382 188
rect 18302 42 18319 44
rect 18365 42 18382 44
rect 18744 98 18824 108
rect 17711 26 17757 37
rect 18319 26 18365 37
rect 15152 -57 15232 -46
rect 18744 -46 18756 98
rect 18812 -46 18824 98
rect 18744 -57 18824 -46
rect 14280 -322 14384 -312
rect 15416 -322 15520 -310
rect 15582 -322 15686 -310
rect 16190 -322 16294 -310
rect 14280 -402 14292 -322
rect 14372 -402 15428 -322
rect 15508 -402 15594 -322
rect 15674 -402 16202 -322
rect 16282 -402 16294 -322
rect 14280 -412 14384 -402
rect 15416 -414 15520 -402
rect 15582 -414 15686 -402
rect 16190 -414 16294 -402
rect 17682 -322 17786 -310
rect 18290 -322 18394 -310
rect 18456 -322 18560 -310
rect 19592 -322 19696 -312
rect 17682 -402 17694 -322
rect 17774 -402 18302 -322
rect 18382 -402 18468 -322
rect 18548 -402 19604 -322
rect 19684 -402 19696 -322
rect 17682 -414 17786 -402
rect 18290 -414 18394 -402
rect 18456 -414 18560 -402
rect 19592 -412 19696 -402
rect 14834 -720 14956 -709
rect 14834 -1220 14845 -720
rect 14945 -1220 14956 -720
rect 19020 -720 19142 -709
rect 16036 -1094 16116 -1084
rect 14834 -1231 14956 -1220
rect 15428 -1130 15508 -1120
rect 15428 -1291 15440 -1130
rect 15496 -1291 15508 -1130
rect 15428 -1301 15508 -1291
rect 15732 -1178 15812 -1168
rect 15732 -1339 15744 -1178
rect 15800 -1339 15812 -1178
rect 16036 -1311 16048 -1094
rect 16104 -1311 16116 -1094
rect 16644 -1094 16724 -1084
rect 16644 -1150 16656 -1094
rect 16712 -1150 16724 -1094
rect 16644 -1160 16724 -1150
rect 17252 -1094 17332 -1084
rect 17252 -1150 17264 -1094
rect 17320 -1150 17332 -1094
rect 17252 -1160 17332 -1150
rect 17860 -1094 17940 -1084
rect 16036 -1319 16116 -1311
rect 16340 -1178 16420 -1168
rect 15732 -1349 15812 -1339
rect 16340 -1339 16352 -1178
rect 16408 -1339 16420 -1178
rect 16340 -1349 16420 -1339
rect 16948 -1178 17028 -1168
rect 16948 -1339 16960 -1178
rect 17016 -1339 17028 -1178
rect 16948 -1349 17028 -1339
rect 17556 -1178 17636 -1168
rect 17556 -1339 17568 -1178
rect 17624 -1339 17636 -1178
rect 17556 -1349 17636 -1339
rect 17860 -1339 17872 -1094
rect 17928 -1339 17940 -1094
rect 18468 -1130 18548 -1120
rect 17860 -1349 17940 -1339
rect 18164 -1178 18244 -1168
rect 18164 -1339 18176 -1178
rect 18232 -1339 18244 -1178
rect 18468 -1291 18480 -1130
rect 18536 -1291 18548 -1130
rect 19020 -1220 19031 -720
rect 19131 -1220 19142 -720
rect 19020 -1231 19142 -1220
rect 18468 -1301 18548 -1291
rect 18164 -1349 18244 -1339
rect 15873 -1440 15888 -1385
rect 15523 -1495 15718 -1440
rect 15828 -1445 15888 -1440
rect 15958 -1440 15973 -1385
rect 15958 -1445 16013 -1440
rect 16178 -1445 16193 -1385
rect 16263 -1445 16278 -1385
rect 16433 -1495 16628 -1440
rect 16738 -1495 16933 -1440
rect 17088 -1445 17103 -1385
rect 17173 -1445 17188 -1385
rect 17393 -1445 17408 -1385
rect 17478 -1445 17493 -1385
rect 17653 -1495 17848 -1440
rect 17953 -1495 18148 -1440
rect 18308 -1445 18323 -1385
rect 18393 -1445 18408 -1385
rect 15523 -1510 19118 -1495
rect 15523 -1543 18638 -1510
rect 15523 -1570 15895 -1543
rect 15883 -1599 15895 -1570
rect 15951 -1570 17110 -1543
rect 15951 -1599 15963 -1570
rect 15883 -1609 15963 -1599
rect 17098 -1599 17110 -1570
rect 17166 -1570 18638 -1543
rect 18698 -1570 19118 -1510
rect 17166 -1599 17178 -1570
rect 17098 -1609 17178 -1599
rect 16188 -1791 16268 -1781
rect 16188 -1820 16200 -1791
rect 15523 -1847 16200 -1820
rect 16256 -1820 16268 -1791
rect 17403 -1791 17483 -1781
rect 17403 -1820 17415 -1791
rect 16256 -1847 17415 -1820
rect 17471 -1820 17483 -1791
rect 17471 -1847 18898 -1820
rect 15523 -1880 18898 -1847
rect 18958 -1880 19118 -1820
rect 15523 -1895 19118 -1880
rect 15523 -1945 15718 -1895
rect 16433 -1945 16628 -1895
rect 16738 -1945 16933 -1895
rect 17648 -1945 17843 -1895
rect 17953 -1945 18148 -1895
rect 15218 -1991 15229 -1945
rect 15403 -1991 15414 -1945
rect 15522 -1991 15533 -1945
rect 15707 -1991 15718 -1945
rect 15826 -1991 15837 -1945
rect 16011 -1991 16022 -1945
rect 16130 -1991 16141 -1945
rect 16315 -1991 16326 -1945
rect 16434 -1991 16445 -1945
rect 16619 -1991 16630 -1945
rect 16738 -1991 16749 -1945
rect 16923 -1991 16934 -1945
rect 17042 -1991 17053 -1945
rect 17227 -1991 17238 -1945
rect 17346 -1991 17357 -1945
rect 17531 -1991 17542 -1945
rect 17650 -1991 17661 -1945
rect 17835 -1991 17846 -1945
rect 17954 -1991 17965 -1945
rect 18139 -1991 18150 -1945
rect 18258 -1991 18269 -1945
rect 18443 -1991 18454 -1945
rect 18562 -1991 18573 -1945
rect 18747 -1991 18758 -1945
rect 15873 -2005 15888 -1991
rect 15958 -2005 15973 -1991
rect 16178 -2005 16193 -1991
rect 16263 -2005 16278 -1991
rect 17088 -2005 17103 -1991
rect 17173 -2005 17188 -1991
rect 17393 -2005 17408 -1991
rect 17478 -2005 17493 -1991
rect 18308 -2005 18323 -1991
rect 18393 -2005 18408 -1991
rect 15141 -2037 15187 -2026
rect 14834 -2165 14956 -2154
rect 14834 -2665 14845 -2165
rect 14945 -2665 14956 -2165
rect 15445 -2037 15491 -2026
rect 15428 -2238 15445 -2228
rect 15749 -2037 15795 -2026
rect 15732 -2049 15749 -2039
rect 16053 -2037 16099 -2026
rect 15795 -2049 15812 -2039
rect 15732 -2210 15744 -2049
rect 15800 -2210 15812 -2049
rect 15732 -2220 15749 -2210
rect 15491 -2238 15508 -2228
rect 15428 -2294 15440 -2238
rect 15496 -2294 15508 -2238
rect 15428 -2304 15445 -2294
rect 15141 -2322 15187 -2311
rect 15491 -2304 15508 -2294
rect 15445 -2322 15491 -2311
rect 15795 -2220 15812 -2210
rect 16036 -2083 16053 -2073
rect 16357 -2037 16403 -2026
rect 16340 -2049 16357 -2039
rect 16661 -2037 16707 -2026
rect 16403 -2049 16420 -2039
rect 16099 -2083 16116 -2073
rect 16036 -2294 16048 -2083
rect 16104 -2294 16116 -2083
rect 16340 -2210 16352 -2049
rect 16408 -2210 16420 -2049
rect 16340 -2220 16357 -2210
rect 16036 -2304 16053 -2294
rect 15749 -2322 15795 -2311
rect 16099 -2304 16116 -2294
rect 16053 -2322 16099 -2311
rect 16403 -2220 16420 -2210
rect 16644 -2049 16661 -2039
rect 16965 -2037 17011 -2026
rect 16707 -2049 16724 -2039
rect 16644 -2294 16656 -2049
rect 16712 -2294 16724 -2049
rect 16948 -2049 16965 -2039
rect 17269 -2037 17315 -2026
rect 17011 -2049 17028 -2039
rect 16948 -2210 16960 -2049
rect 17016 -2210 17028 -2049
rect 16948 -2220 16965 -2210
rect 16644 -2304 16661 -2294
rect 16357 -2322 16403 -2311
rect 16707 -2304 16724 -2294
rect 16661 -2322 16707 -2311
rect 17011 -2220 17028 -2210
rect 17252 -2083 17269 -2073
rect 17573 -2037 17619 -2026
rect 17556 -2049 17573 -2039
rect 17877 -2037 17923 -2026
rect 17619 -2049 17636 -2039
rect 17315 -2083 17332 -2073
rect 17252 -2294 17264 -2083
rect 17320 -2294 17332 -2083
rect 17556 -2210 17568 -2049
rect 17624 -2210 17636 -2049
rect 17556 -2220 17573 -2210
rect 17252 -2304 17269 -2294
rect 16965 -2322 17011 -2311
rect 17315 -2304 17332 -2294
rect 17269 -2322 17315 -2311
rect 17619 -2220 17636 -2210
rect 17860 -2049 17877 -2039
rect 18181 -2037 18227 -2026
rect 17923 -2049 17940 -2039
rect 17860 -2294 17872 -2049
rect 17928 -2294 17940 -2049
rect 17860 -2304 17877 -2294
rect 17573 -2322 17619 -2311
rect 17923 -2304 17940 -2294
rect 18164 -2049 18181 -2039
rect 18485 -2037 18531 -2026
rect 18227 -2049 18244 -2039
rect 18164 -2294 18176 -2049
rect 18232 -2294 18244 -2049
rect 18164 -2304 18181 -2294
rect 17877 -2322 17923 -2311
rect 18227 -2304 18244 -2294
rect 18468 -2237 18485 -2227
rect 18789 -2037 18835 -2026
rect 18531 -2237 18548 -2227
rect 18468 -2294 18480 -2237
rect 18536 -2294 18548 -2237
rect 18468 -2304 18485 -2294
rect 18181 -2322 18227 -2311
rect 18531 -2304 18548 -2294
rect 18485 -2322 18531 -2311
rect 18789 -2322 18835 -2311
rect 19020 -2165 19142 -2154
rect 15218 -2403 15229 -2357
rect 15403 -2403 15414 -2357
rect 15522 -2403 15533 -2357
rect 15707 -2403 15718 -2357
rect 15826 -2403 15837 -2357
rect 16011 -2403 16022 -2357
rect 16130 -2403 16141 -2357
rect 16315 -2403 16326 -2357
rect 16434 -2403 16445 -2357
rect 16619 -2403 16630 -2357
rect 16738 -2403 16749 -2357
rect 16923 -2403 16934 -2357
rect 17042 -2403 17053 -2357
rect 17227 -2403 17238 -2357
rect 17346 -2403 17357 -2357
rect 17531 -2403 17542 -2357
rect 17650 -2403 17661 -2357
rect 17835 -2403 17846 -2357
rect 17954 -2403 17965 -2357
rect 18139 -2403 18150 -2357
rect 18258 -2403 18269 -2357
rect 18443 -2403 18454 -2357
rect 18562 -2403 18573 -2357
rect 18747 -2403 18758 -2357
rect 14834 -2676 14956 -2665
rect 19020 -2665 19031 -2165
rect 19131 -2665 19142 -2165
rect 19020 -2676 19142 -2665
rect 16766 -2871 16842 -2841
rect 16950 -2871 17026 -2841
rect 17134 -2871 17210 -2841
rect 16534 -2969 16614 -2967
rect 16534 -3091 16546 -2969
rect 16602 -3091 16614 -2969
rect 16534 -3093 16614 -3091
rect 16856 -2969 16936 -2967
rect 16856 -3091 16868 -2969
rect 16924 -3091 16936 -2969
rect 16856 -3093 16936 -3091
rect 17040 -2969 17120 -2967
rect 17040 -3091 17052 -2969
rect 17108 -3091 17120 -2969
rect 17040 -3093 17120 -3091
rect 16766 -3219 16842 -3189
rect 13758 -3320 13862 -3310
rect 16950 -3320 17026 -3189
rect 17134 -3219 17210 -3189
rect 20114 -3320 20218 -3310
rect 13758 -3400 13770 -3320
rect 13850 -3400 20126 -3320
rect 20206 -3400 20218 -3320
rect 13758 -3410 13862 -3400
rect 20114 -3410 20218 -3400
<< via1 >>
rect 13770 2039 13850 2115
rect 20126 2039 20206 2115
rect 14120 1213 14176 1347
rect 14304 1213 14360 1347
rect 14442 1213 14498 1347
rect 14980 1213 15036 1347
rect 15164 1213 15220 1347
rect 15302 1213 15358 1347
rect 15744 1216 15800 1360
rect 16048 1203 16104 1259
rect 16352 1216 16408 1360
rect 16656 1203 16712 1259
rect 16960 1216 17016 1360
rect 17264 1203 17320 1259
rect 17568 1216 17624 1360
rect 17872 1203 17928 1259
rect 18176 1216 18232 1360
rect 18618 1213 18674 1347
rect 18756 1213 18812 1347
rect 18940 1213 18996 1347
rect 19478 1213 19534 1347
rect 19616 1213 19672 1347
rect 19800 1213 19856 1347
rect 16851 1096 16907 1152
rect 17069 1096 17125 1152
rect 14630 760 14710 844
rect 15152 760 15232 844
rect 15898 762 15978 842
rect 16506 762 16586 842
rect 16644 762 16724 842
rect 17252 762 17332 842
rect 17390 762 17470 842
rect 17998 762 18078 842
rect 18744 760 18824 844
rect 19266 760 19346 844
rect 16307 468 16387 548
rect 17589 468 17669 548
rect 15910 260 15966 404
rect 16518 260 16574 404
rect 17402 260 17458 404
rect 18010 260 18066 404
rect 15164 -46 15220 98
rect 15606 44 15662 188
rect 16214 44 16270 188
rect 17706 44 17762 188
rect 18314 44 18370 188
rect 18756 -46 18812 98
rect 14292 -402 14372 -322
rect 15428 -402 15508 -322
rect 15594 -402 15674 -322
rect 16202 -402 16282 -322
rect 17694 -402 17774 -322
rect 18302 -402 18382 -322
rect 18468 -402 18548 -322
rect 19604 -402 19684 -322
rect 14845 -881 14945 -720
rect 15440 -1291 15496 -1130
rect 15744 -1339 15800 -1178
rect 16048 -1311 16104 -1094
rect 16656 -1150 16712 -1094
rect 17264 -1150 17320 -1094
rect 16352 -1339 16408 -1178
rect 16960 -1339 17016 -1178
rect 17568 -1339 17624 -1178
rect 17872 -1339 17928 -1094
rect 18176 -1339 18232 -1178
rect 18480 -1291 18536 -1130
rect 19031 -881 19131 -720
rect 15888 -1445 15958 -1385
rect 16193 -1445 16263 -1385
rect 17103 -1445 17173 -1385
rect 17408 -1445 17478 -1385
rect 18323 -1445 18393 -1385
rect 15895 -1599 15951 -1543
rect 17110 -1599 17166 -1543
rect 18638 -1570 18698 -1510
rect 16200 -1847 16256 -1791
rect 17415 -1847 17471 -1791
rect 18898 -1880 18958 -1820
rect 15888 -1991 15958 -1945
rect 16193 -1991 16263 -1945
rect 17103 -1991 17173 -1945
rect 17408 -1991 17478 -1945
rect 18323 -1991 18393 -1945
rect 15888 -2005 15958 -1991
rect 16193 -2005 16263 -1991
rect 17103 -2005 17173 -1991
rect 17408 -2005 17478 -1991
rect 18323 -2005 18393 -1991
rect 14845 -2665 14945 -2504
rect 15744 -2210 15749 -2049
rect 15749 -2210 15795 -2049
rect 15795 -2210 15800 -2049
rect 15440 -2294 15445 -2238
rect 15445 -2294 15491 -2238
rect 15491 -2294 15496 -2238
rect 16048 -2294 16053 -2083
rect 16053 -2294 16099 -2083
rect 16099 -2294 16104 -2083
rect 16352 -2210 16357 -2049
rect 16357 -2210 16403 -2049
rect 16403 -2210 16408 -2049
rect 16656 -2294 16661 -2049
rect 16661 -2294 16707 -2049
rect 16707 -2294 16712 -2049
rect 16960 -2210 16965 -2049
rect 16965 -2210 17011 -2049
rect 17011 -2210 17016 -2049
rect 17264 -2294 17269 -2083
rect 17269 -2294 17315 -2083
rect 17315 -2294 17320 -2083
rect 17568 -2210 17573 -2049
rect 17573 -2210 17619 -2049
rect 17619 -2210 17624 -2049
rect 17872 -2294 17877 -2049
rect 17877 -2294 17923 -2049
rect 17923 -2294 17928 -2049
rect 18176 -2294 18181 -2049
rect 18181 -2294 18227 -2049
rect 18227 -2294 18232 -2049
rect 18480 -2294 18485 -2237
rect 18485 -2294 18531 -2237
rect 18531 -2294 18536 -2237
rect 16546 -3091 16602 -2969
rect 16868 -3091 16924 -2969
rect 17052 -3091 17108 -2969
rect 13770 -3400 13850 -3320
rect 20126 -3400 20206 -3320
<< metal2 >>
rect 13758 2115 13862 2129
rect 13758 2039 13770 2115
rect 13850 2039 13862 2115
rect 13758 2029 13862 2039
rect 20114 2115 20218 2127
rect 20114 2039 20126 2115
rect 20206 2039 20218 2115
rect 13770 -3310 13850 2029
rect 20114 2027 20218 2039
rect 14098 1806 14198 1816
rect 14098 1726 14108 1806
rect 14188 1726 14198 1806
rect 14098 1716 14198 1726
rect 14420 1806 14520 1816
rect 14420 1726 14430 1806
rect 14510 1726 14520 1806
rect 14420 1716 14520 1726
rect 14108 1347 14188 1716
rect 14304 1349 14360 1357
rect 14108 1213 14120 1347
rect 14176 1213 14188 1347
rect 14108 1211 14188 1213
rect 14292 1347 14372 1349
rect 14292 1213 14304 1347
rect 14360 1213 14372 1347
rect 14120 1203 14176 1211
rect 14292 -312 14372 1213
rect 14430 1347 14510 1716
rect 14430 1213 14442 1347
rect 14498 1213 14510 1347
rect 14430 1211 14510 1213
rect 14442 1203 14498 1211
rect 14630 856 14710 1960
rect 14958 1806 15058 1816
rect 14958 1726 14968 1806
rect 15048 1726 15058 1806
rect 14958 1716 15058 1726
rect 15280 1806 15380 1816
rect 15280 1726 15290 1806
rect 15370 1726 15380 1806
rect 15280 1716 15380 1726
rect 15722 1806 15822 1816
rect 15722 1726 15732 1806
rect 15812 1726 15822 1806
rect 15722 1716 15822 1726
rect 16330 1806 16430 1816
rect 16330 1726 16340 1806
rect 16420 1726 16430 1806
rect 16330 1716 16430 1726
rect 16938 1806 17038 1816
rect 16938 1726 16948 1806
rect 17028 1726 17038 1806
rect 16938 1716 17038 1726
rect 17546 1806 17646 1816
rect 17546 1726 17556 1806
rect 17636 1726 17646 1806
rect 17546 1716 17646 1726
rect 18154 1806 18254 1816
rect 18154 1726 18164 1806
rect 18244 1726 18254 1806
rect 18154 1716 18254 1726
rect 18596 1806 18696 1816
rect 18596 1726 18606 1806
rect 18686 1726 18696 1806
rect 18596 1716 18696 1726
rect 18918 1806 19018 1816
rect 18918 1726 18928 1806
rect 19008 1726 19018 1806
rect 18918 1716 19018 1726
rect 14968 1347 15048 1716
rect 15164 1349 15220 1357
rect 14968 1213 14980 1347
rect 15036 1213 15048 1347
rect 14968 1211 15048 1213
rect 15152 1347 15232 1349
rect 15152 1213 15164 1347
rect 15220 1213 15232 1347
rect 14980 1203 15036 1211
rect 14618 844 14722 856
rect 15152 854 15232 1213
rect 15290 1347 15370 1716
rect 15290 1213 15302 1347
rect 15358 1213 15370 1347
rect 15732 1360 15812 1716
rect 15732 1216 15744 1360
rect 15800 1216 15812 1360
rect 16340 1360 16420 1716
rect 15732 1214 15812 1216
rect 16036 1259 16116 1269
rect 15290 1211 15370 1213
rect 15302 1203 15358 1211
rect 15744 1206 15800 1214
rect 16036 1203 16048 1259
rect 16104 1203 16116 1259
rect 16340 1216 16352 1360
rect 16408 1216 16420 1360
rect 16948 1360 17028 1716
rect 16340 1214 16420 1216
rect 16644 1259 16724 1269
rect 16352 1206 16408 1214
rect 16036 1193 16116 1203
rect 16644 1203 16656 1259
rect 16712 1203 16724 1259
rect 16948 1216 16960 1360
rect 17016 1216 17028 1360
rect 17556 1360 17636 1716
rect 16948 1214 17028 1216
rect 17252 1259 17332 1269
rect 16960 1206 17016 1214
rect 14618 760 14630 844
rect 14710 760 14722 844
rect 14618 750 14722 760
rect 15140 844 15244 854
rect 16644 852 16724 1203
rect 17252 1203 17264 1259
rect 17320 1203 17332 1259
rect 17556 1216 17568 1360
rect 17624 1216 17636 1360
rect 18164 1360 18244 1716
rect 17556 1214 17636 1216
rect 17860 1259 17940 1269
rect 17568 1206 17624 1214
rect 16839 1152 16919 1162
rect 16839 1096 16851 1152
rect 16907 1096 16919 1152
rect 16839 1022 16919 1096
rect 17057 1152 17137 1162
rect 17057 1096 17069 1152
rect 17125 1096 17137 1152
rect 16829 1012 16929 1022
rect 16829 932 16839 1012
rect 16919 932 16929 1012
rect 16829 922 16929 932
rect 17057 852 17137 1096
rect 17252 1022 17332 1203
rect 17860 1203 17872 1259
rect 17928 1203 17940 1259
rect 18164 1216 18176 1360
rect 18232 1216 18244 1360
rect 18164 1214 18244 1216
rect 18606 1347 18686 1716
rect 18756 1349 18812 1357
rect 18176 1206 18232 1214
rect 18606 1213 18618 1347
rect 18674 1213 18686 1347
rect 18606 1211 18686 1213
rect 18744 1347 18824 1349
rect 18744 1213 18756 1347
rect 18812 1213 18824 1347
rect 18618 1203 18674 1211
rect 17860 1193 17940 1203
rect 17242 1012 17342 1022
rect 17242 932 17252 1012
rect 17332 932 17342 1012
rect 17242 922 17342 932
rect 17252 852 17332 922
rect 18744 854 18824 1213
rect 18928 1347 19008 1716
rect 18928 1213 18940 1347
rect 18996 1213 19008 1347
rect 18928 1211 19008 1213
rect 18940 1203 18996 1211
rect 19266 854 19346 1960
rect 19456 1806 19556 1816
rect 19456 1726 19466 1806
rect 19546 1726 19556 1806
rect 19456 1716 19556 1726
rect 19778 1806 19878 1816
rect 19778 1726 19788 1806
rect 19868 1726 19878 1806
rect 19778 1716 19878 1726
rect 19466 1347 19546 1716
rect 19616 1349 19672 1357
rect 19466 1213 19478 1347
rect 19534 1213 19546 1347
rect 19466 1211 19546 1213
rect 19604 1347 19684 1349
rect 19604 1213 19616 1347
rect 19672 1213 19684 1347
rect 19478 1203 19534 1211
rect 15140 760 15152 844
rect 15232 760 15244 844
rect 15140 750 15244 760
rect 15886 842 15990 852
rect 15886 762 15898 842
rect 15978 762 15990 842
rect 15886 748 15990 762
rect 16494 842 16734 852
rect 17047 842 17147 852
rect 16494 762 16506 842
rect 16586 762 16644 842
rect 16724 762 17057 842
rect 17137 762 17147 842
rect 16494 748 16734 762
rect 17047 752 17147 762
rect 17240 842 17482 852
rect 17240 762 17252 842
rect 17332 762 17390 842
rect 17470 762 17482 842
rect 17240 748 17482 762
rect 17986 842 18090 853
rect 17986 762 17998 842
rect 18078 762 18090 842
rect 17986 749 18090 762
rect 18732 844 18836 854
rect 18732 760 18744 844
rect 18824 760 18836 844
rect 18732 750 18836 760
rect 19254 844 19358 854
rect 19254 760 19266 844
rect 19346 760 19358 844
rect 19254 750 19358 760
rect 15898 404 15978 748
rect 16297 548 16397 558
rect 16297 468 16307 548
rect 16387 468 16397 548
rect 16297 458 16397 468
rect 15898 260 15910 404
rect 15966 260 15978 404
rect 15898 258 15978 260
rect 16506 404 16586 748
rect 16506 260 16518 404
rect 16574 260 16586 404
rect 16506 258 16586 260
rect 17390 404 17470 748
rect 17579 548 17679 558
rect 17579 468 17589 548
rect 17669 468 17679 548
rect 17579 458 17679 468
rect 17390 260 17402 404
rect 17458 260 17470 404
rect 17390 258 17470 260
rect 17998 404 18078 749
rect 17998 260 18010 404
rect 18066 260 18078 404
rect 17998 258 18078 260
rect 15910 250 15966 258
rect 16518 250 16574 258
rect 17402 250 17458 258
rect 18010 250 18066 258
rect 15606 190 15662 198
rect 16214 190 16270 198
rect 17706 190 17762 198
rect 18314 190 18370 198
rect 15594 188 15674 190
rect 15152 98 15232 108
rect 14843 -46 15164 98
rect 15220 -46 15232 98
rect 14280 -322 14384 -312
rect 14280 -402 14292 -322
rect 14372 -402 14384 -322
rect 14280 -412 14384 -402
rect 14843 -720 14947 -46
rect 15152 -57 15232 -46
rect 15594 44 15606 188
rect 15662 44 15674 188
rect 15594 -310 15674 44
rect 16202 188 16282 190
rect 16202 44 16214 188
rect 16270 44 16282 188
rect 16202 -310 16282 44
rect 17694 188 17774 190
rect 17694 44 17706 188
rect 17762 44 17774 188
rect 17694 -310 17774 44
rect 18302 188 18382 190
rect 18302 44 18314 188
rect 18370 44 18382 188
rect 18302 -310 18382 44
rect 18744 98 18824 108
rect 18744 -46 18756 98
rect 18812 -46 19133 98
rect 18744 -57 18824 -46
rect 15416 -322 15520 -310
rect 15416 -402 15428 -322
rect 15508 -402 15520 -322
rect 15416 -414 15520 -402
rect 15582 -322 15686 -310
rect 15582 -402 15594 -322
rect 15674 -402 15686 -322
rect 15582 -414 15686 -402
rect 16190 -322 16294 -310
rect 16190 -402 16202 -322
rect 16282 -402 16294 -322
rect 16190 -414 16294 -402
rect 17682 -322 17786 -310
rect 17682 -402 17694 -322
rect 17774 -402 17786 -322
rect 17682 -414 17786 -402
rect 18290 -322 18394 -310
rect 18290 -402 18302 -322
rect 18382 -402 18394 -322
rect 18290 -414 18394 -402
rect 18456 -322 18560 -310
rect 18456 -402 18468 -322
rect 18548 -402 18560 -322
rect 18456 -414 18560 -402
rect 14843 -881 14845 -720
rect 14945 -881 14947 -720
rect 14843 -893 14947 -881
rect 15428 -1130 15508 -414
rect 18468 -892 18548 -414
rect 15428 -1291 15440 -1130
rect 15496 -1291 15508 -1130
rect 16036 -948 18548 -892
rect 19029 -720 19133 -46
rect 19604 -312 19684 1213
rect 19788 1347 19868 1716
rect 19788 1213 19800 1347
rect 19856 1213 19868 1347
rect 19788 1211 19868 1213
rect 19800 1203 19856 1211
rect 19592 -322 19696 -312
rect 19592 -402 19604 -322
rect 19684 -402 19696 -322
rect 19592 -412 19696 -402
rect 19029 -881 19031 -720
rect 19131 -881 19133 -720
rect 19029 -893 19133 -881
rect 16036 -1094 16116 -948
rect 15428 -1301 15508 -1291
rect 15732 -1178 15812 -1168
rect 15732 -1339 15744 -1178
rect 15800 -1339 15812 -1178
rect 16036 -1311 16048 -1094
rect 16104 -1311 16116 -1094
rect 16644 -1094 16724 -1084
rect 16644 -1150 16656 -1094
rect 16712 -1150 16724 -1094
rect 16644 -1160 16724 -1150
rect 17252 -1094 17332 -948
rect 17252 -1150 17264 -1094
rect 17320 -1150 17332 -1094
rect 17252 -1160 17332 -1150
rect 17860 -1094 17940 -1084
rect 16036 -1319 16116 -1311
rect 16340 -1178 16420 -1168
rect 15732 -1669 15812 -1339
rect 16340 -1339 16352 -1178
rect 16408 -1339 16420 -1178
rect 15873 -1385 16278 -1375
rect 15873 -1445 15888 -1385
rect 15958 -1445 16193 -1385
rect 16263 -1445 16278 -1385
rect 15873 -1455 16278 -1445
rect 15883 -1543 15963 -1533
rect 15883 -1599 15895 -1543
rect 15951 -1599 15963 -1543
rect 15883 -1609 15963 -1599
rect 16340 -1669 16420 -1339
rect 16948 -1178 17028 -1168
rect 16948 -1339 16960 -1178
rect 17016 -1339 17028 -1178
rect 16948 -1669 17028 -1339
rect 17556 -1178 17636 -1168
rect 17556 -1339 17568 -1178
rect 17624 -1339 17636 -1178
rect 17088 -1385 17493 -1375
rect 17088 -1445 17103 -1385
rect 17173 -1445 17408 -1385
rect 17478 -1445 17493 -1385
rect 17088 -1455 17493 -1445
rect 17098 -1543 17178 -1533
rect 17098 -1599 17110 -1543
rect 17166 -1599 17178 -1543
rect 17098 -1609 17178 -1599
rect 17556 -1669 17636 -1339
rect 17860 -1339 17872 -1094
rect 17928 -1339 17940 -1094
rect 18468 -1130 18548 -948
rect 17860 -1349 17940 -1339
rect 18164 -1178 18244 -1168
rect 18164 -1339 18176 -1178
rect 18232 -1339 18244 -1178
rect 18468 -1291 18480 -1130
rect 18536 -1291 18548 -1130
rect 18468 -1301 18548 -1291
rect 18164 -1669 18244 -1339
rect 18308 -1385 18408 -1375
rect 18602 -1385 18828 -1384
rect 18308 -1445 18323 -1385
rect 18393 -1444 18828 -1385
rect 18393 -1445 18567 -1444
rect 18308 -1455 18408 -1445
rect 18623 -1510 18708 -1500
rect 18623 -1570 18638 -1510
rect 18698 -1570 18708 -1510
rect 18623 -1585 18708 -1570
rect 15732 -1725 18244 -1669
rect 15732 -2049 15812 -1725
rect 16188 -1791 16268 -1781
rect 16188 -1847 16200 -1791
rect 16256 -1847 16268 -1791
rect 16188 -1857 16268 -1847
rect 15873 -1945 16278 -1935
rect 15873 -2005 15888 -1945
rect 15958 -2005 16193 -1945
rect 16263 -2005 16278 -1945
rect 15873 -2015 16278 -2005
rect 15732 -2210 15744 -2049
rect 15800 -2210 15812 -2049
rect 16340 -2049 16420 -1725
rect 15428 -2238 15508 -2228
rect 15428 -2294 15440 -2238
rect 15496 -2294 15508 -2238
rect 15428 -2304 15508 -2294
rect 14843 -2504 14947 -2492
rect 14843 -2665 14845 -2504
rect 14945 -2665 14947 -2504
rect 15732 -2556 15812 -2210
rect 16036 -2083 16116 -2073
rect 16036 -2294 16048 -2083
rect 16104 -2294 16116 -2083
rect 16340 -2210 16352 -2049
rect 16408 -2210 16420 -2049
rect 16340 -2220 16420 -2210
rect 16644 -2049 16724 -2039
rect 16036 -2440 16116 -2294
rect 16644 -2294 16656 -2049
rect 16712 -2294 16724 -2049
rect 16948 -2049 17028 -1725
rect 17403 -1791 17483 -1781
rect 17403 -1847 17415 -1791
rect 17471 -1847 17483 -1791
rect 17403 -1857 17483 -1847
rect 17088 -1945 17493 -1935
rect 17088 -2005 17103 -1945
rect 17173 -2005 17408 -1945
rect 17478 -2005 17493 -1945
rect 17088 -2015 17493 -2005
rect 16948 -2210 16960 -2049
rect 17016 -2210 17028 -2049
rect 17556 -2049 17636 -1725
rect 16948 -2220 17028 -2210
rect 17252 -2083 17332 -2073
rect 16644 -2304 16724 -2294
rect 17252 -2294 17264 -2083
rect 17320 -2294 17332 -2083
rect 17556 -2210 17568 -2049
rect 17624 -2210 17636 -2049
rect 17556 -2220 17636 -2210
rect 17860 -2049 17940 -2039
rect 17252 -2440 17332 -2294
rect 17860 -2294 17872 -2049
rect 17928 -2294 17940 -2049
rect 17860 -2304 17940 -2294
rect 18164 -2049 18244 -1725
rect 18638 -1725 18698 -1585
rect 18768 -1605 18828 -1444
rect 18768 -1665 18958 -1605
rect 18638 -1785 18828 -1725
rect 18308 -1945 18408 -1935
rect 18768 -1945 18828 -1785
rect 18898 -1810 18958 -1665
rect 18888 -1820 18968 -1810
rect 18888 -1880 18898 -1820
rect 18958 -1880 18968 -1820
rect 18888 -1890 18968 -1880
rect 18308 -2005 18323 -1945
rect 18393 -2005 18828 -1945
rect 18308 -2015 18408 -2005
rect 18164 -2294 18176 -2049
rect 18232 -2294 18244 -2049
rect 18164 -2304 18244 -2294
rect 18468 -2237 18548 -2227
rect 18468 -2294 18480 -2237
rect 18536 -2294 18548 -2237
rect 18468 -2440 18548 -2294
rect 16036 -2496 18548 -2440
rect 15732 -2567 18254 -2556
rect 15732 -2623 18164 -2567
rect 18244 -2623 18254 -2567
rect 15732 -2633 18254 -2623
rect 14843 -2967 14947 -2665
rect 14843 -2969 16936 -2967
rect 14843 -3091 16546 -2969
rect 16602 -3091 16868 -2969
rect 16924 -3091 16936 -2969
rect 14843 -3093 16936 -3091
rect 17040 -2969 17120 -2633
rect 17040 -3091 17052 -2969
rect 17108 -3091 17120 -2969
rect 17040 -3093 17120 -3091
rect 20126 -3310 20206 2027
rect 13758 -3320 13862 -3310
rect 13615 -3400 13770 -3320
rect 13850 -3400 13862 -3320
rect 13758 -3410 13862 -3400
rect 20114 -3320 20218 -3310
rect 20114 -3400 20126 -3320
rect 20206 -3400 20218 -3320
rect 20114 -3410 20218 -3400
<< via2 >>
rect 14108 1726 14188 1806
rect 14430 1726 14510 1806
rect 14968 1726 15048 1806
rect 15290 1726 15370 1806
rect 15732 1726 15812 1806
rect 16340 1726 16420 1806
rect 16948 1726 17028 1806
rect 17556 1726 17636 1806
rect 18164 1726 18244 1806
rect 18606 1726 18686 1806
rect 18928 1726 19008 1806
rect 16048 1203 16104 1259
rect 16656 1203 16712 1259
rect 16839 932 16919 1012
rect 17872 1203 17928 1259
rect 17252 932 17332 1012
rect 19466 1726 19546 1806
rect 19788 1726 19868 1806
rect 17057 762 17137 842
rect 16307 468 16387 548
rect 17589 468 17669 548
rect 15440 -1291 15496 -1130
rect 16048 -1311 16104 -1255
rect 16656 -1150 16712 -1094
rect 16200 -1443 16256 -1387
rect 15895 -1599 15951 -1543
rect 17415 -1443 17471 -1387
rect 17110 -1599 17166 -1543
rect 17872 -1339 17928 -1094
rect 18480 -1291 18536 -1130
rect 16200 -1847 16256 -1791
rect 15895 -2003 15951 -1947
rect 15440 -2294 15496 -2238
rect 16048 -2139 16104 -2083
rect 16656 -2294 16712 -2049
rect 17415 -1847 17471 -1791
rect 17110 -2003 17166 -1947
rect 17264 -2139 17320 -2083
rect 17872 -2294 17928 -2049
rect 18176 -2294 18232 -2049
rect 18164 -2623 18244 -2567
<< metal3 >>
rect 14098 1806 14198 1816
rect 14420 1806 14520 1816
rect 14958 1806 15058 1816
rect 15280 1806 15380 1816
rect 15722 1806 15822 1816
rect 16938 1806 17038 1926
rect 17546 1806 17646 1816
rect 18154 1806 18254 1816
rect 18596 1806 18696 1816
rect 18918 1806 19018 1816
rect 19456 1806 19556 1816
rect 19778 1806 19878 1816
rect 14098 1726 14108 1806
rect 14188 1726 14430 1806
rect 14510 1726 14968 1806
rect 15048 1726 15290 1806
rect 15370 1726 15732 1806
rect 15812 1726 16340 1806
rect 16420 1726 16948 1806
rect 17028 1726 17556 1806
rect 17636 1726 18164 1806
rect 18244 1726 18606 1806
rect 18686 1726 18928 1806
rect 19008 1726 19466 1806
rect 19546 1726 19788 1806
rect 19868 1726 19878 1806
rect 14098 1716 14198 1726
rect 14420 1716 14520 1726
rect 14958 1716 15058 1726
rect 15280 1716 15380 1726
rect 15722 1716 15822 1726
rect 16330 1716 16430 1726
rect 16938 1716 17038 1726
rect 17546 1716 17646 1726
rect 18154 1716 18254 1726
rect 18596 1716 18696 1726
rect 18918 1716 19018 1726
rect 19456 1716 19556 1726
rect 19778 1716 19878 1726
rect 16036 1259 16116 1269
rect 16036 1203 16048 1259
rect 16104 1203 16116 1259
rect 16036 1193 16116 1203
rect 16644 1259 16724 1269
rect 17860 1259 17940 1269
rect 16644 1203 16656 1259
rect 16712 1203 17872 1259
rect 17928 1203 17940 1259
rect 16644 1193 16724 1203
rect 17860 1193 17940 1203
rect 16048 1012 16104 1193
rect 16829 1012 16929 1022
rect 17242 1012 17342 1022
rect 16048 932 16839 1012
rect 16919 932 17252 1012
rect 17332 932 17342 1012
rect 16297 548 16397 932
rect 16829 922 16929 932
rect 17242 922 17342 932
rect 17047 842 17147 852
rect 17047 762 17057 842
rect 17137 762 17147 842
rect 17047 714 17147 762
rect 17047 634 17669 714
rect 17589 558 17669 634
rect 16297 468 16307 548
rect 16387 468 16397 548
rect 16297 458 16397 468
rect 17579 548 17679 558
rect 17579 468 17589 548
rect 17669 468 17679 548
rect 17579 458 17679 468
rect 15428 -1094 17940 -1084
rect 15428 -1130 16656 -1094
rect 15428 -1291 15440 -1130
rect 15496 -1150 16656 -1130
rect 16712 -1150 17872 -1094
rect 15496 -1160 17872 -1150
rect 15496 -1291 15508 -1160
rect 15428 -1301 15508 -1291
rect 16036 -1255 16116 -1245
rect 15435 -1725 15500 -1301
rect 16036 -1311 16048 -1255
rect 16104 -1311 16116 -1255
rect 15883 -1543 15963 -1533
rect 15883 -1599 15895 -1543
rect 15951 -1599 15963 -1543
rect 15883 -1609 15963 -1599
rect 16036 -1609 16116 -1311
rect 17860 -1339 17872 -1160
rect 17928 -1339 17940 -1094
rect 18468 -1130 18548 -1120
rect 18468 -1291 18480 -1130
rect 18536 -1291 18548 -1130
rect 18468 -1301 18548 -1291
rect 16178 -1387 16278 -1375
rect 16178 -1443 16200 -1387
rect 16256 -1443 16278 -1387
rect 16178 -1455 16278 -1443
rect 17393 -1387 17493 -1375
rect 17393 -1443 17415 -1387
rect 17471 -1443 17493 -1387
rect 17393 -1455 17493 -1443
rect 17098 -1543 17178 -1533
rect 17098 -1599 17110 -1543
rect 17166 -1599 17178 -1543
rect 17098 -1609 17178 -1599
rect 17860 -1609 17940 -1339
rect 16036 -1669 16724 -1609
rect 15435 -1785 16116 -1725
rect 15873 -1947 15973 -1935
rect 15873 -2003 15895 -1947
rect 15951 -2003 15973 -1947
rect 15873 -2015 15973 -2003
rect 16036 -2083 16116 -1785
rect 16188 -1791 16268 -1781
rect 16188 -1847 16200 -1791
rect 16256 -1847 16268 -1791
rect 16188 -1857 16268 -1847
rect 16036 -2139 16048 -2083
rect 16104 -2139 16116 -2083
rect 16036 -2149 16116 -2139
rect 16644 -2049 16724 -1669
rect 17252 -1669 17940 -1609
rect 17088 -1947 17188 -1935
rect 17088 -2003 17110 -1947
rect 17166 -2003 17188 -1947
rect 17088 -2015 17188 -2003
rect 16644 -2228 16656 -2049
rect 15428 -2238 16656 -2228
rect 15428 -2294 15440 -2238
rect 15496 -2294 16656 -2238
rect 16712 -2228 16724 -2049
rect 17252 -2083 17332 -1669
rect 18475 -1725 18540 -1301
rect 17403 -1791 17483 -1781
rect 17403 -1847 17415 -1791
rect 17471 -1847 17483 -1791
rect 17403 -1857 17483 -1847
rect 17860 -1785 18540 -1725
rect 17252 -2139 17264 -2083
rect 17320 -2139 17332 -2083
rect 17252 -2149 17332 -2139
rect 17860 -2049 17940 -1785
rect 17860 -2228 17872 -2049
rect 16712 -2294 17872 -2228
rect 17928 -2294 17940 -2049
rect 15428 -2304 17940 -2294
rect 18164 -2049 18244 -2039
rect 18164 -2294 18176 -2049
rect 18232 -2294 18244 -2049
rect 18164 -2556 18244 -2294
rect 18154 -2567 18254 -2556
rect 18154 -2623 18164 -2567
rect 18244 -2623 18254 -2567
rect 18154 -2633 18254 -2623
<< via3 >>
rect 15895 -1599 15951 -1543
rect 16200 -1443 16256 -1387
rect 17415 -1443 17471 -1387
rect 17110 -1599 17166 -1543
rect 15895 -2003 15951 -1947
rect 16200 -1847 16256 -1791
rect 17110 -2003 17166 -1947
rect 17415 -1847 17471 -1791
<< metal4 >>
rect 16178 -1387 16278 -1375
rect 16178 -1443 16200 -1387
rect 16256 -1443 16278 -1387
rect 16178 -1455 16278 -1443
rect 17393 -1387 17493 -1375
rect 17393 -1443 17415 -1387
rect 17471 -1443 17493 -1387
rect 17393 -1455 17493 -1443
rect 15883 -1543 15963 -1533
rect 15883 -1599 15895 -1543
rect 15951 -1599 15963 -1543
rect 15883 -1609 15963 -1599
rect 15895 -1935 15951 -1609
rect 16200 -1781 16256 -1455
rect 17098 -1543 17178 -1533
rect 17098 -1599 17110 -1543
rect 17166 -1599 17178 -1543
rect 17098 -1609 17178 -1599
rect 16188 -1791 16268 -1781
rect 16188 -1847 16200 -1791
rect 16256 -1847 16268 -1791
rect 16188 -1857 16268 -1847
rect 17110 -1935 17166 -1609
rect 17415 -1781 17471 -1455
rect 17403 -1791 17483 -1781
rect 17403 -1847 17415 -1791
rect 17471 -1847 17483 -1791
rect 17403 -1857 17483 -1847
rect 15873 -1947 15973 -1935
rect 15873 -2003 15895 -1947
rect 15951 -2003 15973 -1947
rect 15873 -2015 15973 -2003
rect 17088 -1947 17188 -1935
rect 17088 -2003 17110 -1947
rect 17166 -2003 17188 -1947
rect 17088 -2015 17188 -2003
use nfet_03v3_6BEH2F  nfet_03v3_6BEH2F_0 comparator/final_magic/lvsclean_SAlatch
timestamp 1757405367
transform 1 0 16988 0 1 -2174
box -1884 -266 1884 266
use nfet_03v3_MJTYYT  nfet_03v3_MJTYYT_0 comparator/final_magic/lvsclean_SAlatch
timestamp 1757409273
transform 1 0 17886 0 1 224
box -958 -410 958 410
use nfet_03v3_MJTYYT  nfet_03v3_MJTYYT_1
timestamp 1757409273
transform 1 0 16090 0 1 224
box -958 -410 958 410
use pfet_03v3_CRJA84  pfet_03v3_CRJA84_0 comparator/final_magic/lvsclean_SAlatch
timestamp 1757500055
transform 1 0 15100 0 1 1280
box -290 -290 290 290
use pfet_03v3_USLA84  XM1 comparator/final_magic/lvsclean_SAlatch
timestamp 1757500055
transform 1 0 14240 0 1 1280
box -290 -290 290 290
use pfet_03v3_GABL2T  XM3 comparator/final_magic/lvsclean_SAlatch
timestamp 1757500055
transform 1 0 16988 0 1 1280
box -1718 -310 1718 310
use pfet_03v3_U2FB84  XM5 comparator/final_magic/lvsclean_SAlatch
timestamp 1757500055
transform 1 0 18876 0 1 1280
box -290 -290 290 290
use pfet_03v3_USLA84  XM6
timestamp 1757500055
transform 1 0 19736 0 1 1280
box -290 -290 290 290
use nfet_03v3_6BEH2F  XM9
timestamp 1757405367
transform 1 0 16988 0 1 -1211
box -1884 -266 1884 266
use nfet_03v3_W5F4U7  XM11 comparator/final_magic/lvsclean_SAlatch
timestamp 1757405367
transform 1 0 16988 0 1 -3030
box -474 -290 474 290
<< labels >>
rlabel metal2 16350 -3037 16350 -3037 7 VSS
port 4 w
rlabel metal2 14671 1960 14671 1960 1 Vout1
port 5 n
rlabel metal2 19307 1960 19307 1960 1 Vout2
port 6 n
rlabel metal1 16986 2115 16986 2115 1 Clk
port 0 n
rlabel metal1 19118 -1856 19118 -1856 3 Vin2
port 2 e
rlabel metal1 19118 -1535 19118 -1535 3 Vin1
port 1 e
rlabel metal1 15212 -322 15212 -322 1 Vp
rlabel metal1 18811 -322 18811 -322 1 Vq
rlabel metal3 16987 1926 16987 1926 1 VDD
port 3 n
<< end >>
