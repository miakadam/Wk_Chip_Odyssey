magic
tech gf180mcuD
magscale 1 10
timestamp 1757815838
<< metal1 >>
rect -365 2825 1182 2881
rect -365 1804 -309 2825
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -848 1748 -309 1804
rect -644 1688 -574 1700
rect 808 1688 878 1700
rect -644 1632 -632 1688
rect -576 1632 -360 1688
rect 669 1632 810 1688
rect 866 1632 878 1688
rect -644 1620 -574 1632
rect 808 1622 878 1632
rect -360 785 -304 1572
rect 621 835 701 915
rect 974 785 1054 795
rect -360 729 986 785
rect 1042 729 1054 785
rect 974 727 1054 729
rect 808 676 878 678
rect -360 675 878 676
rect -360 621 810 675
rect 866 621 878 675
rect -360 620 878 621
rect -360 -457 -304 620
rect 808 612 878 620
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 1126 -457 1182 2825
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect -780 -517 -710 -503
rect 984 -517 1044 -507
rect 2294 -517 2364 -505
rect -780 -573 -768 -517
rect -712 -573 -360 -517
rect 726 -573 986 -517
rect 1042 -573 1126 -517
rect 2095 -573 2296 -517
rect 2352 -573 2620 -517
rect -780 -585 -710 -573
rect 984 -585 1044 -573
rect 2294 -583 2364 -573
rect -496 -689 -360 -633
rect -496 -1419 -440 -689
rect -848 -1475 -440 -1419
rect 1126 -1419 1182 -671
rect 2460 -1419 2540 -1409
rect 1126 -1475 2472 -1419
rect 2528 -1475 2540 -1419
rect -496 -2722 -440 -1475
rect 2460 -1477 2540 -1475
rect 984 -1530 1054 -1528
rect 2284 -1529 2364 -1527
rect -360 -1586 986 -1530
rect 1042 -1586 1054 -1530
rect -360 -2662 -304 -1586
rect 984 -1598 1054 -1586
rect 1126 -1585 2296 -1529
rect 2352 -1585 2364 -1529
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 1126 -2661 1182 -1585
rect 2284 -1597 2364 -1585
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect 808 -2721 878 -2710
rect 2470 -2721 2540 -2711
rect 808 -2722 1126 -2721
rect -496 -2778 -360 -2722
rect 708 -2778 810 -2722
rect 866 -2778 1126 -2722
rect 2095 -2777 2472 -2721
rect 2528 -2777 2620 -2721
rect 808 -2788 878 -2778
rect 2470 -2789 2540 -2777
rect -644 -2838 -574 -2826
rect -644 -2894 -632 -2838
rect -576 -2883 -360 -2838
rect -576 -2894 -255 -2883
rect -644 -2906 -574 -2894
rect -360 -3625 -304 -2894
rect 974 -3625 1054 -3615
rect -360 -3681 986 -3625
rect 1042 -3681 1054 -3625
rect 974 -3683 1054 -3681
rect 808 -3734 878 -3732
rect -360 -3735 878 -3734
rect -360 -3789 810 -3735
rect 866 -3789 878 -3735
rect -360 -3790 878 -3789
rect -360 -4811 -304 -3790
rect 808 -3798 878 -3790
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect -360 -4822 -261 -4811
rect -349 -4867 -261 -4822
rect -780 -4927 -710 -4913
rect 984 -4927 1044 -4915
rect -780 -4983 -768 -4927
rect -712 -4981 -360 -4927
rect -322 -4979 -260 -4927
rect -351 -4981 -260 -4979
rect -712 -4983 -260 -4981
rect 714 -4983 986 -4927
rect 1042 -4983 1044 -4927
rect -780 -4995 -710 -4983
rect 984 -4995 1044 -4983
rect -848 -5099 -360 -5043
rect -354 -5099 -291 -5043
rect 621 -5780 701 -5700
rect -770 -5830 -710 -5826
rect 1126 -5830 1182 -2893
rect -831 -5886 -768 -5830
rect -712 -5886 1182 -5830
rect -770 -5898 -710 -5886
<< via1 >>
rect 316 2717 372 2773
rect -632 1632 -576 1688
rect 810 1632 866 1688
rect 986 729 1042 785
rect 810 621 866 675
rect 316 512 372 568
rect 1802 512 1858 568
rect -768 -573 -712 -517
rect 986 -573 1042 -517
rect 2296 -573 2352 -517
rect 2472 -1475 2528 -1419
rect 986 -1586 1042 -1530
rect 2296 -1585 2352 -1529
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect 810 -2778 866 -2722
rect 2472 -2777 2528 -2721
rect -632 -2894 -576 -2838
rect 986 -3681 1042 -3625
rect 810 -3789 866 -3735
rect 316 -3898 372 -3842
rect -768 -4983 -712 -4927
rect 986 -4983 1042 -4927
rect -768 -5886 -712 -5830
<< metal2 >>
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -644 1688 -574 1700
rect -644 1632 -632 1688
rect -576 1632 -574 1688
rect -644 1620 -574 1632
rect 808 1688 878 1700
rect 808 1632 810 1688
rect 866 1632 878 1688
rect 808 1622 878 1632
rect -780 -517 -710 -503
rect -780 -573 -768 -517
rect -712 -573 -710 -517
rect -780 -585 -710 -573
rect -768 -4913 -712 -585
rect -632 -2826 -576 1620
rect -185 903 -129 913
rect -185 837 -129 847
rect 621 903 701 915
rect 621 847 633 903
rect 689 847 701 903
rect 621 835 701 847
rect 810 678 866 1622
rect 974 785 1054 795
rect 974 729 986 785
rect 1042 729 1054 785
rect 974 727 1054 729
rect 808 675 878 678
rect 808 621 810 675
rect 866 621 878 675
rect 808 609 878 621
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 986 -507 1042 727
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect 984 -517 1044 -507
rect 984 -573 986 -517
rect 1042 -573 1044 -517
rect 984 -585 1044 -573
rect 2294 -517 2364 -505
rect 2294 -573 2296 -517
rect 2352 -573 2620 -517
rect 2294 -583 2364 -573
rect -185 -1302 -129 -1292
rect -185 -1368 -129 -1358
rect 633 -1302 689 -1292
rect 633 -1368 689 -1358
rect 986 -1528 1042 -585
rect 1301 -1302 1357 -1292
rect 1301 -1368 1357 -1358
rect 2119 -1302 2175 -1292
rect 2119 -1368 2175 -1358
rect 2296 -1527 2352 -583
rect 2460 -1419 2540 -1409
rect 2460 -1475 2472 -1419
rect 2528 -1475 2540 -1419
rect 2460 -1477 2540 -1475
rect 984 -1530 1054 -1528
rect 984 -1586 986 -1530
rect 1042 -1586 1054 -1530
rect 984 -1598 1054 -1586
rect 2284 -1529 2364 -1527
rect 2284 -1585 2296 -1529
rect 2352 -1585 2364 -1529
rect 2284 -1597 2364 -1585
rect 316 -1633 372 -1627
rect 1802 -1632 1858 -1626
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect 808 -2722 878 -2710
rect 2472 -2711 2528 -1477
rect 808 -2778 810 -2722
rect 866 -2778 878 -2722
rect 808 -2788 878 -2778
rect 2470 -2721 2540 -2711
rect 2470 -2777 2472 -2721
rect 2528 -2777 2620 -2721
rect -644 -2838 -574 -2826
rect -644 -2894 -632 -2838
rect -576 -2894 -574 -2838
rect -644 -2906 -574 -2894
rect -197 -3507 -117 -3495
rect -197 -3563 -185 -3507
rect -129 -3563 -117 -3507
rect -197 -3575 -117 -3563
rect 633 -3507 689 -3497
rect 633 -3573 689 -3563
rect 810 -3732 866 -2788
rect 2470 -2789 2540 -2777
rect 1301 -3506 1357 -3496
rect 1301 -3572 1357 -3562
rect 2119 -3506 2175 -3496
rect 2119 -3572 2175 -3562
rect 974 -3625 1054 -3615
rect 974 -3681 986 -3625
rect 1042 -3681 1054 -3625
rect 974 -3683 1054 -3681
rect 808 -3735 878 -3732
rect 808 -3789 810 -3735
rect 866 -3789 878 -3735
rect 808 -3801 878 -3789
rect 316 -3838 372 -3832
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect -780 -4927 -710 -4913
rect 986 -4915 1042 -3683
rect -780 -4983 -768 -4927
rect -712 -4983 -710 -4927
rect -780 -4995 -710 -4983
rect 984 -4927 1044 -4915
rect 984 -4983 986 -4927
rect 1042 -4983 1044 -4927
rect 984 -4995 1044 -4983
rect -768 -5826 -712 -4995
rect -197 -5712 -117 -5700
rect -197 -5768 -185 -5712
rect -129 -5768 -117 -5712
rect -197 -5780 -117 -5768
rect 621 -5712 701 -5700
rect 621 -5768 633 -5712
rect 689 -5768 701 -5712
rect 621 -5780 701 -5768
rect -770 -5830 -710 -5826
rect -770 -5886 -768 -5830
rect -712 -5886 -710 -5830
rect -770 -5898 -710 -5886
<< via2 >>
rect 316 2717 372 2773
rect -185 847 -129 903
rect 633 847 689 903
rect 316 512 372 568
rect 1802 512 1858 568
rect -185 -1358 -129 -1302
rect 633 -1358 689 -1302
rect 1301 -1358 1357 -1302
rect 2119 -1358 2175 -1302
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect -185 -3563 -129 -3507
rect 633 -3563 689 -3507
rect 1301 -3562 1357 -3506
rect 2119 -3562 2175 -3506
rect 316 -3898 372 -3842
rect -185 -5768 -129 -5712
rect 633 -5768 689 -5712
<< metal3 >>
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -197 903 -117 915
rect -197 847 -185 903
rect -129 847 -117 903
rect -197 835 -117 847
rect 621 903 701 915
rect 621 847 633 903
rect 689 847 701 903
rect 621 835 701 847
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect -197 -1302 -117 -1290
rect -197 -1358 -185 -1302
rect -129 -1358 -117 -1302
rect -197 -1370 -117 -1358
rect 621 -1302 701 -1290
rect 621 -1358 633 -1302
rect 689 -1358 701 -1302
rect 621 -1370 701 -1358
rect 1289 -1302 1369 -1290
rect 1289 -1358 1301 -1302
rect 1357 -1358 1369 -1302
rect 1289 -1370 1369 -1358
rect 2107 -1302 2187 -1290
rect 2107 -1358 2119 -1302
rect 2175 -1358 2187 -1302
rect 2107 -1370 2187 -1358
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect -197 -3507 -117 -3495
rect -197 -3563 -185 -3507
rect -129 -3563 -117 -3507
rect -197 -3575 -117 -3563
rect 621 -3507 701 -3495
rect 621 -3563 633 -3507
rect 689 -3563 701 -3507
rect 621 -3575 701 -3563
rect 1289 -3506 1369 -3494
rect 1289 -3562 1301 -3506
rect 1357 -3562 1369 -3506
rect 1289 -3574 1369 -3562
rect 2107 -3506 2187 -3494
rect 2107 -3562 2119 -3506
rect 2175 -3562 2187 -3506
rect 2107 -3574 2187 -3562
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect -197 -5712 -117 -5700
rect -197 -5768 -185 -5712
rect -129 -5768 -117 -5712
rect -197 -5780 -117 -5768
rect 621 -5712 701 -5700
rect 621 -5768 633 -5712
rect 689 -5768 701 -5712
rect 621 -5780 701 -5768
<< via3 >>
rect 316 2717 372 2773
rect -185 847 -129 903
rect 633 847 689 903
rect 316 512 372 568
rect 1802 512 1858 568
rect -185 -1358 -129 -1302
rect 633 -1358 689 -1302
rect 1301 -1358 1357 -1302
rect 2119 -1358 2175 -1302
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect -185 -3563 -129 -3507
rect 633 -3563 689 -3507
rect 1301 -3562 1357 -3506
rect 2119 -3562 2175 -3506
rect 316 -3898 372 -3842
rect -185 -5768 -129 -5712
rect 633 -5768 689 -5712
<< metal4 >>
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -710 903 2590 2569
rect -710 847 -185 903
rect -129 847 633 903
rect 689 847 2590 903
rect -710 729 2590 847
rect -710 364 122 729
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 572 364 1608 729
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect 2058 364 2590 729
rect -710 -1302 2590 364
rect -710 -1358 -185 -1302
rect -129 -1358 633 -1302
rect 689 -1358 1301 -1302
rect 1357 -1358 2119 -1302
rect 2175 -1358 2590 -1302
rect -710 -1476 2590 -1358
rect -710 -1841 122 -1476
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 572 -1841 1608 -1476
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect 2058 -1841 2590 -1476
rect -710 -3506 2590 -1841
rect -710 -3507 1301 -3506
rect -710 -3563 -185 -3507
rect -129 -3563 633 -3507
rect 689 -3562 1301 -3507
rect 1357 -3562 2119 -3506
rect 2175 -3562 2590 -3506
rect 689 -3563 2590 -3562
rect -710 -3681 2590 -3563
rect -710 -4046 122 -3681
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect 572 -4046 2590 -3681
rect -710 -5712 2590 -4046
rect -710 -5768 -185 -5712
rect -129 -5768 633 -5712
rect 689 -5768 2590 -5712
rect -710 -5898 2590 -5768
<< via4 >>
rect 316 2717 372 2773
rect 316 512 372 568
rect 1802 512 1858 568
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect 316 -3898 372 -3842
<< metal5 >>
rect -710 2773 2590 2881
rect -710 2717 316 2773
rect 372 2717 2590 2773
rect -710 568 2590 2717
rect -710 512 316 568
rect 372 512 1802 568
rect 1858 512 2590 568
rect -710 -1636 2590 512
rect -710 -1637 1802 -1636
rect -710 -1693 316 -1637
rect 372 -1692 1802 -1637
rect 1858 -1692 2590 -1636
rect 372 -1693 2590 -1692
rect -710 -3842 2590 -1693
rect -710 -3898 316 -3842
rect 372 -3898 2590 -3842
rect -710 -5898 2590 -3898
use nand3  nand3_0 nand3
timestamp 1757649945
transform 1 0 -2072 0 1 2640
box 1712 -1805 2798 145
use nand3  nand3_1
timestamp 1757649945
transform 1 0 -2072 0 1 435
box 1712 -1805 2798 145
use nand3  nand3_2
timestamp 1757649945
transform 1 0 -586 0 1 435
box 1712 -1805 2798 145
use nand3  nand3_3
timestamp 1757649945
transform 1 0 -2072 0 1 -1770
box 1712 -1805 2798 145
use nand3  nand3_4
timestamp 1757649945
transform 1 0 -586 0 1 -1769
box 1712 -1805 2798 145
use nand3  nand3_5
timestamp 1757649945
transform 1 0 -2072 0 1 -3975
box 1712 -1805 2798 145
<< labels >>
rlabel metal1 -848 1776 -848 1776 7 setb
port 4 w
rlabel metal1 -848 -1447 -848 -1447 7 clk
port 3 w
rlabel metal1 -848 -5072 -848 -5072 7 d
port 2 w
rlabel metal1 -831 -5859 -831 -5859 7 resetb
port 5 w
rlabel metal2 2620 -545 2620 -545 3 Q
port 6 e
rlabel metal2 2620 -2750 2620 -2750 3 Qb
port 7 e
rlabel metal5 1260 2881 1260 2881 1 vdd
port 0 n
<< end >>
