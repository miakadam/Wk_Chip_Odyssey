magic
tech gf180mcuD
magscale 1 10
timestamp 1757551291
<< error_s >>
rect 1675 -397 1686 -351
rect 1169 -643 1226 -633
rect 1286 -643 1337 -633
rect 1423 -643 1543 -548
rect 1193 -656 1313 -646
rect 1185 -691 1215 -679
rect 1009 -770 1059 -714
rect 1155 -725 1220 -714
rect 1226 -725 1268 -679
rect 1400 -702 1543 -643
rect 1155 -737 1230 -725
rect 1153 -758 1184 -742
rect 1133 -770 1213 -758
rect 1065 -1168 1115 -770
rect 1133 -778 1184 -770
rect 1138 -1145 1184 -778
rect 1233 -783 1293 -754
rect 1338 -760 1354 -726
rect 1262 -1150 1293 -783
rect 1322 -771 1354 -760
rect 1322 -1145 1356 -771
rect 1262 -1157 1313 -1150
rect 1322 -1156 1354 -1145
rect 1293 -1158 1313 -1157
rect 1387 -1158 1543 -702
rect 1233 -1168 1313 -1158
rect 1065 -1170 1153 -1168
rect 1233 -1170 1321 -1168
rect 1400 -1194 1543 -1158
rect 1153 -1224 1166 -1208
rect 1220 -1224 1231 -1208
rect 1093 -1236 1253 -1224
rect 1133 -1237 1253 -1236
rect 1357 -1237 1543 -1194
rect 1133 -1240 1543 -1237
rect 1133 -1244 1403 -1240
rect 1153 -1251 1403 -1244
rect 1092 -1262 1403 -1251
rect 1092 -1283 1400 -1262
rect 1423 -1320 1543 -1240
rect 1675 -1309 1686 -1263
rect 1423 -1343 1492 -1320
rect 1423 -1380 1483 -1343
<< metal1 >>
rect 1129 325 1187 593
rect 1226 -711 1286 -396
rect 1338 -961 1395 -183
rect 1116 -1249 1174 -981
use nfet_03v3_WAQWUP  M3
timestamp 0
transform 1 0 1193 0 1 -970
box -290 -410 290 410
use pfet_03v3_LSTY94  M4
timestamp 0
transform 1 0 1713 0 1 -830
box -290 -610 290 610
use nfet_03v3_Q7US5R  XM3
timestamp 1757549261
transform 1 0 1253 0 1 -934
box -290 -386 290 386
use pfet_03v3_YXHA8C  XM4
timestamp 1757549261
transform 1 0 1253 0 1 47
box -290 -586 290 586
<< labels >>
rlabel metal1 1130 -1220 1140 -1210 7 avss
port 3 w
rlabel metal1 1140 530 1150 540 7 avdd
port 0 w
rlabel metal1 1240 -550 1250 -540 7 in
port 1 w
rlabel metal1 1350 -540 1360 -530 7 out
port 2 w
<< end >>
