magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< pwell >>
rect -958 -310 958 310
<< nmos >>
rect -708 -100 -508 100
rect -404 -100 -204 100
rect -100 -100 100 100
rect 204 -100 404 100
rect 508 -100 708 100
<< ndiff >>
rect -796 87 -708 100
rect -796 -87 -783 87
rect -737 -87 -708 87
rect -796 -100 -708 -87
rect -508 87 -404 100
rect -508 -87 -479 87
rect -433 -87 -404 87
rect -508 -100 -404 -87
rect -204 87 -100 100
rect -204 -87 -175 87
rect -129 -87 -100 87
rect -204 -100 -100 -87
rect 100 87 204 100
rect 100 -87 129 87
rect 175 -87 204 87
rect 100 -100 204 -87
rect 404 87 508 100
rect 404 -87 433 87
rect 479 -87 508 87
rect 404 -100 508 -87
rect 708 87 796 100
rect 708 -87 737 87
rect 783 -87 796 87
rect 708 -100 796 -87
<< ndiffc >>
rect -783 -87 -737 87
rect -479 -87 -433 87
rect -175 -87 -129 87
rect 129 -87 175 87
rect 433 -87 479 87
rect 737 -87 783 87
<< psubdiff >>
rect -934 214 934 286
rect -934 170 -862 214
rect -934 -170 -921 170
rect -875 -170 -862 170
rect 862 170 934 214
rect -934 -214 -862 -170
rect 862 -170 875 170
rect 921 -170 934 170
rect 862 -214 934 -170
rect -934 -286 934 -214
<< psubdiffcont >>
rect -921 -170 -875 170
rect 875 -170 921 170
<< polysilicon >>
rect -708 179 -508 192
rect -708 133 -695 179
rect -521 133 -508 179
rect -708 100 -508 133
rect -404 179 -204 192
rect -404 133 -391 179
rect -217 133 -204 179
rect -404 100 -204 133
rect -100 179 100 192
rect -100 133 -87 179
rect 87 133 100 179
rect -100 100 100 133
rect 204 179 404 192
rect 204 133 217 179
rect 391 133 404 179
rect 204 100 404 133
rect 508 179 708 192
rect 508 133 521 179
rect 695 133 708 179
rect 508 100 708 133
rect -708 -133 -508 -100
rect -708 -179 -695 -133
rect -521 -179 -508 -133
rect -708 -192 -508 -179
rect -404 -133 -204 -100
rect -404 -179 -391 -133
rect -217 -179 -204 -133
rect -404 -192 -204 -179
rect -100 -133 100 -100
rect -100 -179 -87 -133
rect 87 -179 100 -133
rect -100 -192 100 -179
rect 204 -133 404 -100
rect 204 -179 217 -133
rect 391 -179 404 -133
rect 204 -192 404 -179
rect 508 -133 708 -100
rect 508 -179 521 -133
rect 695 -179 708 -133
rect 508 -192 708 -179
<< polycontact >>
rect -695 133 -521 179
rect -391 133 -217 179
rect -87 133 87 179
rect 217 133 391 179
rect 521 133 695 179
rect -695 -179 -521 -133
rect -391 -179 -217 -133
rect -87 -179 87 -133
rect 217 -179 391 -133
rect 521 -179 695 -133
<< metal1 >>
rect -921 227 921 273
rect -921 170 -875 227
rect -706 133 -695 179
rect -521 133 -510 179
rect -402 133 -391 179
rect -217 133 -206 179
rect -98 133 -87 179
rect 87 133 98 179
rect 206 133 217 179
rect 391 133 402 179
rect 510 133 521 179
rect 695 133 706 179
rect 875 170 921 227
rect -783 87 -737 98
rect -783 -98 -737 -87
rect -479 87 -433 98
rect -479 -98 -433 -87
rect -175 87 -129 98
rect -175 -98 -129 -87
rect 129 87 175 98
rect 129 -98 175 -87
rect 433 87 479 98
rect 433 -98 479 -87
rect 737 87 783 98
rect 737 -98 783 -87
rect -921 -227 -875 -170
rect -706 -179 -695 -133
rect -521 -179 -510 -133
rect -402 -179 -391 -133
rect -217 -179 -206 -133
rect -98 -179 -87 -133
rect 87 -179 98 -133
rect 206 -179 217 -133
rect 391 -179 402 -133
rect 510 -179 521 -133
rect 695 -179 706 -133
rect 875 -227 921 -170
rect -921 -273 921 -227
<< properties >>
string FIXED_BBOX -898 -250 898 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
