** sch_path: /foss/designs/FinalBlocksLayout/comparator/comparator_no_offsetcal.sch
.subckt comparator_no_offsetcal VDD VSS CLK Vin1 Vin2 Vout
*.PININFO VDD:B VSS:B CLK:B Vin1:B Vin2:B Vout:B
* noconn #net1
x2 VDD latch net1 inv1 inv2 VSS rslatch
x4 VDD latch Vout VSS osu_sc_buf_4
x1 CLK Vin1 Vin2 VDD VSS out1 out2 no_offsetLatch
x3 VDD out1 inv1 VSS inv_mia
x5 VDD out2 inv2 VSS inv_mia
.ends

* expanding   symbol:  comparator/final_magic/RSlatch/rslatch.sym # of pins=6
** sym_path: /foss/designs/comparator/final_magic/RSlatch/rslatch.sym
** sch_path: /foss/designs/comparator/final_magic/RSlatch/rslatch.sch
.subckt rslatch VDD Vout1 Vout2 Vin1 Vin2 VSS
*.PININFO VDD:B VSS:B Vin1:B Vin2:B Vout1:B Vout2:B
XM1 Vout1 Vin1 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM2 Vout2 Vin2 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM3 Vout1 Vout2 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
XM4 Vout2 Vout1 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
.ends


* expanding   symbol:  comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sym # of pins=4
** sym_path: /foss/designs/comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sym
** sch_path: /foss/designs/comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sch
.subckt osu_sc_buf_4 VDD A Y VSS
*.PININFO A:I Y:O VDD:I VSS:I
XM1 net1 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 net1 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM3 Y net1 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=4
XM4 Y net1 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=4
.ends


* expanding   symbol:  FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sym # of pins=7
** sym_path: /foss/designs/FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sym
** sch_path: /foss/designs/FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sch
.subckt no_offsetLatch Clk Vin1 Vin2 VDD VSS Vout1 Vout2
*.PININFO Clk:I Vin1:I Vin2:I VDD:B VSS:B Vout1:O Vout2:O
XM1 Vp Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM2 Vout1 Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM3 Vout1 Vout2 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=4
XM4 Vout2 Vout1 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=4
XM5 Vout2 Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM6 Vq Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM7 Vout1 Vout2 Vp VSS nfet_03v3 L=1u W=2u nf=1 m=3
XM8 Vout2 Vout1 Vq VSS nfet_03v3 L=1u W=2u nf=1 m=3
XM9 Vp Vin1 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM10 Vq Vin2 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM11 net1 Clk VSS VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM20 Vp Vin1 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM21 Vq Vin2 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM24 Vp net2 net3 VSS nfet_03v3 L=1u W=1.5u nf=1 m=2
* noconn #net3
* noconn #net2
XM25 Vq net4 net5 VSS nfet_03v3 L=1u W=1.5u nf=1 m=2
* noconn #net5
* noconn #net4
XM26 Vout1 net6 net7 VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net7
* noconn #net6
XM27 Vout2 net8 net9 VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net9
* noconn #net8
* noconn #net10
* noconn #net11
* noconn #net12
* noconn #net13
XM30 net1 net14 net15 VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM31 net16 net17 VSS VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
* noconn #net15
* noconn #net16
* noconn #net17
* noconn #net14
XM32 net18 net19 Vq VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net18
* noconn #net19
XM33 net20 net21 Vp VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net20
* noconn #net21
XM28 net10 net11 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=1
XM29 net12 net13 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=1
.ends


* expanding   symbol:  FinalBlocksLayout/inverter/inv_mia.sym # of pins=4
** sym_path: /foss/designs/FinalBlocksLayout/inverter/inv_mia.sym
** sch_path: /foss/designs/FinalBlocksLayout/inverter/inv_mia.sch
.subckt inv_mia avdd in out avss
*.PININFO avdd:B avss:B in:B out:B
XM3 out in avss avss nfet_03v3 L=0.4u W=2u nf=1 m=1
XM4 out in avdd avdd pfet_03v3 L=0.4u W=4u nf=1 m=1
.ends

