magic
tech gf180mcuD
magscale 1 10
timestamp 1755271904
<< error_p >>
rect -34 233 -23 279
rect 23 233 34 244
rect -80 -198 -57 -187
rect 57 -198 80 -187
rect -34 -279 -23 -233
<< nwell >>
rect -278 -410 278 410
<< pmos >>
rect -28 -200 28 200
<< pdiff >>
rect -116 187 -28 200
rect -116 -187 -103 187
rect -57 -187 -28 187
rect -116 -200 -28 -187
rect 28 187 116 200
rect 28 -187 57 187
rect 103 -187 116 187
rect 28 -200 116 -187
<< pdiffc >>
rect -103 -187 -57 187
rect 57 -187 103 187
<< nsubdiff >>
rect -254 314 254 386
rect -254 270 -182 314
rect -254 -270 -241 270
rect -195 -270 -182 270
rect 182 270 254 314
rect -254 -314 -182 -270
rect 182 -270 195 270
rect 241 -270 254 270
rect 182 -314 254 -270
rect -254 -386 254 -314
<< nsubdiffcont >>
rect -241 -270 -195 270
rect 195 -270 241 270
<< polysilicon >>
rect -36 279 36 292
rect -36 233 -23 279
rect 23 233 36 279
rect -36 220 36 233
rect -28 200 28 220
rect -28 -220 28 -200
rect -36 -233 36 -220
rect -36 -279 -23 -233
rect 23 -279 36 -233
rect -36 -292 36 -279
<< polycontact >>
rect -23 233 23 279
rect -23 -279 23 -233
<< metal1 >>
rect -241 327 241 373
rect -241 270 -195 327
rect -34 233 -23 279
rect 23 233 34 279
rect 195 270 241 327
rect -103 187 -57 198
rect -103 -198 -57 -187
rect 57 187 103 198
rect 57 -198 103 -187
rect -241 -327 -195 -270
rect -34 -279 -23 -233
rect 23 -279 34 -233
rect 195 -327 241 -270
rect -241 -373 241 -327
<< properties >>
string FIXED_BBOX -218 -350 218 350
string gencell pfet_03v3
string library gf180mcu
string parameters w 2.0 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
