magic
tech gf180mcuD
magscale 1 10
timestamp 1757998313
<< pwell >>
rect 1502 -539 1588 -459
<< metal1 >>
rect 1250 570 1850 770
rect 1287 441 1333 570
rect 1502 439 1598 470
rect 1767 441 1813 570
rect 1327 -238 1429 358
rect 1612 63 1692 73
rect 1612 -177 1624 63
rect 1680 -177 1692 63
rect 1612 -187 1692 -177
rect 1502 -460 1598 -319
rect 1434 -472 1598 -460
rect 1434 -528 1446 -472
rect 1502 -528 1598 -472
rect 1434 -540 1598 -528
rect 1502 -681 1598 -540
rect 1330 -958 1426 -762
rect 1612 -832 1692 -822
rect 1612 -888 1624 -832
rect 1680 -888 1692 -832
rect 1612 -898 1692 -888
rect 1287 -1170 1333 -1041
rect 1502 -1070 1598 -1039
rect 1767 -1170 1813 -1041
rect 1250 -1370 1850 -1170
<< via1 >>
rect 1624 -177 1680 63
rect 1446 -528 1502 -472
rect 1624 -888 1680 -832
<< metal2 >>
rect 1612 63 1692 73
rect 1612 -177 1624 63
rect 1680 -177 1692 63
rect 1434 -472 1504 -460
rect 1250 -528 1446 -472
rect 1502 -528 1504 -472
rect 1434 -540 1504 -528
rect 1612 -472 1692 -177
rect 1612 -528 1850 -472
rect 1612 -832 1692 -528
rect 1612 -888 1624 -832
rect 1680 -888 1692 -832
rect 1612 -898 1692 -888
use pfet_03v3_LJVJK4  M1
timestamp 1757998004
transform 1 0 1550 0 1 60
box -300 -510 300 510
use nfet_03v3_EKBWUP  M2
timestamp 1757998004
transform 1 0 1550 0 1 -860
box -300 -310 300 310
<< labels >>
rlabel metal2 1250 -499 1250 -499 7 in
port 0 w
rlabel metal1 1545 770 1545 770 1 vdd
port 1 n
rlabel metal2 1850 -499 1850 -499 3 out
port 2 e
rlabel metal1 1555 -1370 1555 -1370 5 vss
port 3 s
<< end >>
