** sch_path: /foss/designs/FinalBlocksLayout/comp_SAR_final/comp_SAR_final.sch
.subckt comp_SAR_final Clk_piso Vdd Vss Load Clk Piso_out Vin1 Vin2 Comp_out Reset SAR_in
*.PININFO Vdd:B Vss:B Clk:B Vin1:B Vin2:B Comp_out:B Reset:B SAR_in:B Clk_piso:B Load:B Piso_out:B
x1 Vdd Vss Clk Vin1 Vin2 Comp_out comparator_no_offsetcal
x2 Vdd Vss Clk Reset SAR_in d5 d4 d3 d2 d1 d0 SARlogic
x4 loadb d5 d4 d3 Piso_out Vdd d2 Vss d1 d0 Clk_piso adc_PISO
x3 Load Vdd loadb Vss inv2
.ends

* expanding   symbol:  FinalBlocksLayout/comparator/comparator_no_offsetcal.sym # of pins=6
** sym_path: /foss/designs/FinalBlocksLayout/comparator/comparator_no_offsetcal.sym
** sch_path: /foss/designs/FinalBlocksLayout/comparator/comparator_no_offsetcal.sch
.subckt comparator_no_offsetcal VDD VSS CLK Vin1 Vin2 Vout
*.PININFO VDD:B VSS:B CLK:B Vin1:B Vin2:B Vout:B
* noconn #net1
x2 VDD latch net1 inv1 inv2 VSS rslatch
x4 VDD latch Vout VSS osu_sc_buf_4
x1 CLK Vin1 Vin2 VDD VSS out1 out2 no_offsetLatch
x3 VDD out1 inv1 VSS inv_mia
x5 VDD out2 inv2 VSS inv_mia
.ends


* expanding   symbol:  FinalBlocksLayout/SARlogic/SARlogic.sym # of pins=11
** sym_path: /foss/designs/FinalBlocksLayout/SARlogic/SARlogic.sym
** sch_path: /foss/designs/FinalBlocksLayout/SARlogic/SARlogic.sch
.subckt SARlogic vdd vss clk reset comp_in d5 d4 d3 d2 d1 d0
*.PININFO comp_in:I vdd:B vss:B clk:I reset:I d5:B d4:B d3:B d2:B d1:B d0:B
* noconn #net15
* noconn #net16
* noconn #net17
* noconn #net18
* noconn #net19
* noconn #net20
* noconn #net21
x1 vdd vss vss clk reset vdd net1 net7 dffrs
x2 vdd vss net1 clk vdd reset net2 net8 dffrs
x3 vdd vss net2 clk vdd reset net3 net9 dffrs
x4 vdd vss net3 clk vdd reset net4 net10 dffrs
x5 vdd vss net4 clk vdd reset net5 net11 dffrs
x6 vdd vss net5 clk vdd reset net6 net12 dffrs
x7 vdd vss net6 clk vdd reset net22 net13 dffrs
x8 vdd vss vss vss net13 reset net14 net21 dffrs
x9 vdd vss comp_in net14 net12 reset d0 net20 dffrs
x10 vdd vss comp_in d0 net11 reset d1 net19 dffrs
x11 vdd vss comp_in d1 net10 reset d2 net18 dffrs
x12 vdd vss comp_in d2 net9 reset d3 net17 dffrs
x13 vdd vss comp_in d3 net8 reset d4 net16 dffrs
x14 vdd vss comp_in d4 net7 reset d5 net15 dffrs
.ends


* expanding   symbol:  FinalBlocksLayout/piso/adc_PISO.sym # of pins=11
** sym_path: /foss/designs/FinalBlocksLayout/piso/adc_PISO.sym
** sch_path: /foss/designs/FinalBlocksLayout/piso/adc_PISO.sch
.subckt adc_PISO load B6 B5 B4 serial_out avdd B3 avss B2 B1 clk
*.PININFO avdd:B avss:B clk:B B6:B B5:B B4:B B3:B B2:B B1:B load:B serial_out:B
x7 avss load avdd D6 avss B6 2inmux
x8 Q6 load avdd D5 avss B5 2inmux
x27 Q5 load avdd D4 avss B4 2inmux
x28 Q4 load avdd D3 avss B3 2inmux
x29 Q3 load avdd D2 avss B2 2inmux
x30 Q2 load avdd D1 avss B1 2inmux
x1 avdd avss D6 clk avdd avdd Q6 net1 dffrs
x2 avdd avss D5 clk avdd avdd Q5 net2 dffrs
x3 avdd avss D4 clk avdd avdd Q4 net3 dffrs
x4 avdd avss D3 clk avdd avdd Q3 net4 dffrs
x5 avdd avss D2 clk avdd avdd Q2 net5 dffrs
x6 avdd avss D1 clk avdd avdd serial_out net6 dffrs
.ends


* expanding   symbol:  FinalBlocksLayout/inv2/inv2.sym # of pins=4
** sym_path: /foss/designs/FinalBlocksLayout/inv2/inv2.sym
** sch_path: /foss/designs/FinalBlocksLayout/inv2/inv2.sch
.subckt inv2 in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
XM1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
XM2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends


* expanding   symbol:  comparator/final_magic/RSlatch/rslatch.sym # of pins=6
** sym_path: /foss/designs/comparator/final_magic/RSlatch/rslatch.sym
** sch_path: /foss/designs/comparator/final_magic/RSlatch/rslatch.sch
.subckt rslatch VDD Vout1 Vout2 Vin1 Vin2 VSS
*.PININFO VDD:B VSS:B Vin1:B Vin2:B Vout1:B Vout2:B
XM1 Vout1 Vin1 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM2 Vout2 Vin2 VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM3 Vout1 Vout2 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
XM4 Vout2 Vout1 VDD VDD pfet_03v3 L=0.4u W=1u nf=1 m=1
.ends


* expanding   symbol:  comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sym # of pins=4
** sym_path: /foss/designs/comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sym
** sch_path: /foss/designs/comparator/final_magic/osu_sc/buff4x/osu_sc_buf_4.sch
.subckt osu_sc_buf_4 VDD A Y VSS
*.PININFO A:I Y:O VDD:I VSS:I
XM1 net1 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 net1 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM3 Y net1 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=4
XM4 Y net1 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=4
.ends


* expanding   symbol:  FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sym # of pins=7
** sym_path: /foss/designs/FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sym
** sch_path: /foss/designs/FinalBlocksLayout/no_offsetLatch/no_offsetLatch.sch
.subckt no_offsetLatch Clk Vin1 Vin2 VDD VSS Vout1 Vout2
*.PININFO Clk:I Vin1:I Vin2:I VDD:B VSS:B Vout1:O Vout2:O
XM1 Vp Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM2 Vout1 Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM3 Vout1 Vout2 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=4
XM4 Vout2 Vout1 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=4
XM5 Vout2 Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM6 Vq Clk VDD VDD pfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM7 Vout1 Vout2 Vp VSS nfet_03v3 L=1u W=2u nf=1 m=3
XM8 Vout2 Vout1 Vq VSS nfet_03v3 L=1u W=2u nf=1 m=3
XM9 Vp Vin1 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM10 Vq Vin2 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM11 net1 Clk VSS VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM20 Vp Vin1 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM21 Vq Vin2 net1 VSS nfet_03v3 L=1u W=1.5u nf=1 m=5
XM24 Vp net2 net3 VSS nfet_03v3 L=1u W=1.5u nf=1 m=2
* noconn #net3
* noconn #net2
XM25 Vq net4 net5 VSS nfet_03v3 L=1u W=1.5u nf=1 m=2
* noconn #net5
* noconn #net4
XM26 Vout1 net6 net7 VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net7
* noconn #net6
XM27 Vout2 net8 net9 VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net9
* noconn #net8
* noconn #net10
* noconn #net11
* noconn #net12
* noconn #net13
XM30 net1 net14 net15 VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
XM31 net16 net17 VSS VSS nfet_03v3 L=0.40u W=0.80u nf=1 m=1
* noconn #net15
* noconn #net16
* noconn #net17
* noconn #net14
XM32 net18 net19 Vq VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net18
* noconn #net19
XM33 net20 net21 Vp VSS nfet_03v3 L=1u W=2u nf=1 m=1
* noconn #net20
* noconn #net21
XM28 net10 net11 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=1
XM29 net12 net13 VDD VDD pfet_03v3 L=1u W=1u nf=1 m=1
.ends


* expanding   symbol:  FinalBlocksLayout/inverter/inv_mia.sym # of pins=4
** sym_path: /foss/designs/FinalBlocksLayout/inverter/inv_mia.sym
** sch_path: /foss/designs/FinalBlocksLayout/inverter/inv_mia.sch
.subckt inv_mia avdd in out avss
*.PININFO avdd:B avss:B in:B out:B
XM3 out in avss avss nfet_03v3 L=0.4u W=2u nf=1 m=1
XM4 out in avdd avdd pfet_03v3 L=0.4u W=4u nf=1 m=1
.ends


* expanding   symbol:  FinalBlocksLayout/dffrs/dffrs.sym # of pins=8
** sym_path: /foss/designs/FinalBlocksLayout/dffrs/dffrs.sym
** sch_path: /foss/designs/FinalBlocksLayout/dffrs/dffrs.sch
.subckt dffrs vdd vss d clk setb resetb Q Qb
*.PININFO vdd:B vss:B Q:B Qb:B d:B clk:B resetb:B setb:B
x1 vdd net2 net1 net3 setb vss nand3
x2 vdd net1 clk resetb net2 vss nand3
x3 vdd Q Qb net1 setb vss nand3
x4 vdd Qb resetb net4 Q vss nand3
x5 vdd net4 net3 clk net1 vss nand3
x6 vdd net3 d resetb net4 vss nand3
.ends


* expanding   symbol:  FinalBlocksLayout/2inmux/2inmux.sym # of pins=6
** sym_path: /foss/designs/FinalBlocksLayout/2inmux/2inmux.sym
** sch_path: /foss/designs/FinalBlocksLayout/2inmux/2inmux.sch
.subckt 2inmux Bit Load VDD OUT VSS In
*.PININFO VDD:B Bit:B In:B VSS:B Load:B OUT:B
x1 VDD net3 Bit Load VSS and2
x2 VDD net2 net1 In VSS and2
x3 VDD VSS OUT net3 net2 or2
x4 Load VDD net1 VSS inv2
.ends


* expanding   symbol:  comparator/final_magic/nand3/nand3.sym # of pins=6
** sym_path: /foss/designs/comparator/final_magic/nand3/nand3.sym
** sch_path: /foss/designs/comparator/final_magic/nand3/nand3.sch
.subckt nand3 VDD Z A B C VSS
*.PININFO VDD:B VSS:B Z:B A:B B:B C:B
XM1 Z A net1 VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM2 net1 B net2 VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM3 Z B VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM4 Z A VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM5 Z C VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM6 net2 C VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
.ends


* expanding   symbol:  FinalBlocksLayout/and2/and2.sym # of pins=5
** sym_path: /foss/designs/FinalBlocksLayout/and2/and2.sym
** sch_path: /foss/designs/FinalBlocksLayout/and2/and2.sch
.subckt and2 VDD OUT A B VSS
*.PININFO VDD:B A:B B:B VSS:B OUT:B
x1 VDD net1 B A VSS nand2
x2 net1 VDD OUT VSS inv2
.ends


* expanding   symbol:  FinalBlocksLayout/or2/or2.sym # of pins=5
** sym_path: /foss/designs/FinalBlocksLayout/or2/or2.sym
** sch_path: /foss/designs/FinalBlocksLayout/or2/or2.sch
.subckt or2 VDD VSS OUT A B
*.PININFO VDD:B A:B B:B VSS:B OUT:B
x1 VDD VSS net1 A B nor2
x2 net1 VDD OUT VSS inv2
.ends


* expanding   symbol:  FinalBlocksLayout/nand2/nand2.sym # of pins=5
** sym_path: /foss/designs/FinalBlocksLayout/nand2/nand2.sym
** sch_path: /foss/designs/FinalBlocksLayout/nand2/nand2.sch
.subckt nand2 VDD OUT A B VSS
*.PININFO VDD:B VSS:B B:B A:B OUT:B
XM1 OUT A net1 VSS nfet_03v3 L=0.5u W=1u nf=1 m=2
XM2 OUT A VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=1
XM3 net1 B VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=2
XM4 OUT B VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=1
.ends


* expanding   symbol:  FinalBlocksLayout/nor2/nor2.sym # of pins=5
** sym_path: /foss/designs/FinalBlocksLayout/nor2/nor2.sym
** sch_path: /foss/designs/FinalBlocksLayout/nor2/nor2.sch
.subckt nor2 VDD VSS OUT A B
*.PININFO VDD:B VSS:B B:B A:B OUT:B
XM1 OUT A VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=1
XM2 OUT B VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=1
XM3 OUT B net1 VDD pfet_03v3 L=0.5u W=3u nf=1 m=2
XM4 net1 A VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=2
.ends

