magic
tech gf180mcuD
magscale 1 10
timestamp 1758265644
<< metal1 >>
rect -12288 31314 -10879 31362
rect -12288 31114 -10769 31314
rect -12288 28819 -12030 31114
rect -12288 28619 -12088 28819
rect -10803 27724 -10603 27815
rect -10921 27689 -10603 27724
rect -10921 26879 -10568 27689
rect -12030 26679 -10568 26879
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -13680 4940 -13603 4954
rect -12380 4940 -12294 4954
rect -13680 4939 -12366 4940
rect -13680 4881 -13665 4939
rect -13607 4881 -12366 4939
rect -13680 4880 -12366 4881
rect -12306 4880 -12294 4940
rect -13680 4867 -13603 4880
rect -12380 4866 -12294 4880
rect -13722 -1178 -13632 -1166
rect -13722 -1179 -12440 -1178
rect -13722 -1252 -13707 -1179
rect -13634 -1252 -12440 -1179
rect -13722 -1253 -12440 -1252
rect -13722 -1266 -13632 -1253
rect -13717 -1503 -13627 -1491
rect -13717 -1504 -12438 -1503
rect -13717 -1577 -13704 -1504
rect -13631 -1577 -12438 -1504
rect -13717 -1578 -12438 -1577
rect -13717 -1591 -13627 -1578
rect -13382 -3003 -13286 -3000
rect -13382 -3004 -12446 -3003
rect -13382 -3082 -13368 -3004
rect -13290 -3082 -12446 -3004
rect -13382 -3083 -12446 -3082
rect -13382 -3096 -13286 -3083
rect -4464 -3363 -2407 -3321
rect -4464 -3663 -4454 -3363
rect -2454 -3663 -2407 -3363
rect -4464 -3701 -2407 -3663
<< via1 >>
rect -4454 6134 -2454 6434
rect -13665 4881 -13607 4939
rect -12366 4880 -12306 4940
rect -13707 -1252 -13634 -1179
rect -13704 -1577 -13631 -1504
rect -13368 -3082 -13290 -3004
rect -4454 -3663 -2454 -3363
<< metal2 >>
rect -8093 33382 -8037 38726
rect 4049 38341 4105 38603
rect 4045 38285 45751 38341
rect 45695 37436 45751 38285
rect -8103 33372 -8027 33382
rect -8103 33316 -8093 33372
rect -8037 33316 -8027 33372
rect -8103 33306 -8027 33316
rect -11840 27577 -11764 27587
rect -13170 27521 -12630 27577
rect -12030 27521 -11830 27577
rect -11774 27521 -11764 27577
rect -11840 27511 -11764 27521
rect -11141 26474 -11085 27345
rect -1669 26484 -1613 27350
rect 3069 27289 7859 27345
rect -11141 26418 -5025 26474
rect -1669 26428 -971 26484
rect 3069 26417 3125 27289
rect 17275 27078 17331 27346
rect 7111 27022 17331 27078
rect 7111 26391 7167 27022
rect 26747 26814 26803 27350
rect 11153 26758 26803 26814
rect 11153 26397 11209 26758
rect 36219 26445 36275 27346
rect 15195 26389 36275 26445
rect -13224 16389 -12868 16509
rect -13233 15879 -12868 15999
rect -13369 6810 -13259 6930
rect -13680 4940 -13603 4954
rect -13894 4939 -13603 4940
rect -13894 4881 -13665 4939
rect -13607 4881 -13603 4939
rect -13894 4880 -13603 4881
rect -13680 4867 -13603 4880
rect -13722 -1177 -13632 -1166
rect -13880 -1179 -13632 -1177
rect -13880 -1252 -13707 -1179
rect -13634 -1252 -13632 -1179
rect -13722 -1266 -13632 -1252
rect -13717 -1502 -13627 -1491
rect -13878 -1504 -13627 -1502
rect -13878 -1577 -13704 -1504
rect -13631 -1577 -13627 -1504
rect -13717 -1591 -13627 -1577
rect -13369 -3000 -13289 6810
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -12380 4940 -12294 4954
rect -12380 4880 -12366 4940
rect -12306 4880 -12294 4940
rect -12380 4866 -12294 4880
rect -13382 -3004 -13286 -3000
rect -13784 -3082 -13368 -3004
rect -13290 -3082 -13286 -3004
rect -13382 -3096 -13286 -3082
rect -4464 -3363 -2407 -3321
rect -4464 -3663 -4454 -3363
rect -2454 -3663 -2407 -3363
rect -4464 -3701 -2407 -3663
<< via2 >>
rect -8093 33316 -8037 33372
rect -11830 27521 -11774 27577
rect -4454 6134 -2454 6434
rect -4454 -3663 -2454 -3363
<< metal3 >>
rect -8103 33372 -8027 33382
rect -8103 33316 -8093 33372
rect -8037 33316 -8027 33372
rect -8103 33306 -8027 33316
rect -11840 27577 -11764 27587
rect -11840 27521 -11830 27577
rect -11774 27521 -11764 27577
rect -11840 27511 -11764 27521
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -4464 -3363 -2407 -3321
rect -4464 -3663 -4454 -3363
rect -2454 -3663 -2407 -3363
rect -4464 -3701 -2407 -3663
<< via3 >>
rect -4454 6134 -2454 6434
rect -4454 -3663 -2454 -3363
<< metal4 >>
rect -8627 25373 24343 27880
rect 32519 26106 35819 28897
rect 41533 26106 43287 27880
rect -5327 25370 18925 25373
rect 32519 22673 43287 26106
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -4464 -3322 30646 -3321
rect 32519 -3322 35819 22673
rect -4464 -3363 35819 -3322
rect -4464 -3663 -4454 -3363
rect -2454 -3663 35819 -3363
rect -4464 -3701 35819 -3663
rect 30646 -3702 35819 -3701
<< via4 >>
rect -4454 6134 -2454 6434
<< metal5 >>
rect -5369 25370 -2069 28896
rect 4103 25370 7403 28896
rect 13575 25370 16875 28897
rect 23047 25370 26347 28897
rect 18925 21844 26347 25370
rect 22821 6477 26347 21844
rect -4464 6434 26347 6477
rect -4464 6134 -4454 6434
rect -2454 6134 26347 6434
rect -4464 6097 26347 6134
rect 22821 -3206 26347 6097
use adc_PISO  adc_PISO_0
timestamp 1758101161
transform 1 0 -11151 0 1 27659
box -689 -370 56902 10017
use comparator_no_offsetcal  comparator_no_offsetcal_0
timestamp 1758264283
transform 1 0 -16096 0 1 2097
box 2794 -5798 12429 4380
use inv2  inv2_0
timestamp 1757998295
transform 1 0 -13880 0 1 28049
box 1250 -1370 1850 770
use SARlogic  SARlogic_0
timestamp 1757846223
transform 1 0 -12787 0 1 6985
box -473 -175 32092 19504
<< labels >>
rlabel metal2 -13784 -3047 -13784 -3047 7 Clk
port 2 w
rlabel metal2 -13233 15938 -13233 15938 7 Reset
port 6 w
rlabel metal2 -13224 16448 -13224 16448 7 SAR_in
port 7 w
rlabel metal2 -13170 27549 -13170 27549 7 Load
port 8 w
rlabel metal2 4077 38603 4077 38603 1 Piso_out
port 10 n
rlabel metal2 -8063 38726 -8063 38726 1 Clk_piso
port 9 n
rlabel metal5 24711 -3206 24711 -3206 5 Vdd
port 0 s
rlabel metal4 34239 -3702 34239 -3702 5 Vss
port 1 s
rlabel metal2 -13880 -1213 -13880 -1213 7 Vin1
port 3 w
rlabel metal2 -13878 -1540 -13878 -1540 7 Vin2
port 4 w
rlabel metal2 -13894 4909 -13894 4909 7 Comp_out
port 5 w
<< end >>
