* NGSPICE file created from comp_SAR_final.ext - technology: (null)

.subckt comp_SAR_final Clk_piso Vdd Vss Load Clk Piso_out Vin1 Vin2 Comp_out Reset SAR_in
X0 Vdd.t103 SARlogic_0.d3.t4 SARlogic_0.dffrs_7.nand3_8.C.t0 Vdd.t102 pfet_03v3
**devattr s=26000,604 d=26000,604
X1 a_5803_9634 SARlogic_0.dffrs_4.d.t4 Vss.t656 Vss.t655 nfet_03v3
**devattr s=17600,576 d=10400,304
X2 adc_PISO_0.dffrs_4.Qb Vdd.t738 Vdd.t740 Vdd.t739 pfet_03v3
**devattr s=26000,604 d=44000,1176
X3 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t4 Vdd.t343 Vdd.t342 pfet_03v3
**devattr s=26000,604 d=44000,1176
X4 a_37687_30440 inv2_0.out.t2 a_37499_31160.t2 Vss.t548 nfet_03v3
**devattr s=17600,576 d=10400,304
X5 a_n7937_n2793 a_n8017_n2885 a_n9429_n2007.t17 Vss.t450 nfet_03v3
**devattr s=8320,264 d=14080,496
X6 a_28027_28820.t3 SARlogic_0.d1.t4 Vdd.t585 Vdd.t584 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X7 Vss.t109 a_8377_29020 a_9271_28100 Vss.t108 nfet_03v3
**devattr s=10400,304 d=17600,576
X8 Vdd.t507 Reset.t0 SARlogic_0.dffrs_14.nand3_6.C.t1 Vdd.t506 pfet_03v3
**devattr s=26000,604 d=26000,604
X9 a_n7809_21417 SARlogic_0.dffrs_14.nand3_1.C Vss.t358 Vss.t357 nfet_03v3
**devattr s=17600,576 d=10400,304
X10 SARlogic_0.dffrs_2.nand3_1.C.t1 SARlogic_0.dffrs_2.nand3_6.C.t4 a_459_14043 Vss.t373 nfet_03v3
**devattr s=10400,304 d=17600,576
X11 SARlogic_0.d3.t3 SARlogic_0.dffrs_1.Qb.t4 Vdd.t369 Vdd.t368 pfet_03v3
**devattr s=44000,1176 d=26000,604
X12 SARlogic_0.dffrs_4.nand3_8.C.t2 SARlogic_0.dffrs_4.nand3_8.Z.t4 a_8543_9633 Vss.t367 nfet_03v3
**devattr s=10400,304 d=17600,576
X13 Vdd.t531 SARlogic_0.dffrs_1.nand3_8.C.t4 SARlogic_0.dffrs_1.Qb.t3 Vdd.t530 pfet_03v3
**devattr s=26000,604 d=26000,604
X14 adc_PISO_0.dffrs_0.Qb Vdd.t735 Vdd.t737 Vdd.t736 pfet_03v3
**devattr s=26000,604 d=44000,1176
X15 a_12401_7428 SARlogic_0.dffrs_5.nand3_8.C.t4 Vss.t531 Vss.t530 nfet_03v3
**devattr s=17600,576 d=10400,304
X16 SARlogic_0.dffrs_3.nand3_8.C.t2 SARlogic_0.dffrs_3.nand3_8.Z.t4 Vdd.t535 Vdd.t534 pfet_03v3
**devattr s=26000,604 d=44000,1176
X17 Vdd.t734 Vdd.t732 a_33257_31423.t1 Vdd.t733 pfet_03v3
**devattr s=26000,604 d=26000,604
X18 SARlogic_0.dffrs_5.nand3_8.C.t3 SARlogic_0.dffrs_5.nand3_6.C.t4 Vdd.t742 Vdd.t741 pfet_03v3
**devattr s=44000,1176 d=26000,604
X19 a_14071_9634 SARlogic_0.dffrs_5.nand3_8.C.t5 a_13887_9634 Vss.t353 nfet_03v3
**devattr s=10400,304 d=10400,304
X20 SARlogic_0.dffrs_1.Qb.t2 Reset.t1 Vdd.t417 Vdd.t416 pfet_03v3
**devattr s=26000,604 d=44000,1176
X21 a_18113_19210 SARlogic_0.dffrs_12.nand3_8.C.t4 a_17929_19210 Vss.t383 nfet_03v3
**devattr s=10400,304 d=10400,304
X22 Vdd.t567 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t8 Vdd.t566 pfet_03v3
**devattr s=10400,304 d=10400,304
X23 a_10029_9634 SARlogic_0.dffrs_4.nand3_8.C.t4 a_9845_9634 Vss.t350 nfet_03v3
**devattr s=10400,304 d=10400,304
X24 SARlogic_0.dffrs_1.nand3_6.C.t2 Clk.t0 a_n3583_11838 Vss.t23 nfet_03v3
**devattr s=10400,304 d=17600,576
X25 a_n4367_29309 Vdd.t955 a_n4551_29309 Vss.t529 nfet_03v3
**devattr s=10400,304 d=10400,304
X26 SARlogic_0.dffrs_9.Qb SARlogic_0.d2.t4 Vdd.t305 Vdd.t304 pfet_03v3
**devattr s=44000,1176 d=26000,604
X27 a_4841_33627.t2 a_4841_31422.t4 Vdd.t471 Vdd.t470 pfet_03v3
**devattr s=26000,604 d=44000,1176
X28 Vdd.t451 adc_PISO_0.2inmux_1.Bit.t4 a_37499_31160.t3 Vdd.t450 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X29 SARlogic_0.dffrs_5.nand3_6.C.t3 SARlogic_0.dffrs_5.nand3_1.C.t4 Vdd.t830 Vdd.t829 pfet_03v3
**devattr s=44000,1176 d=26000,604
X30 SARlogic_0.dffrs_4.d.t3 Vdd.t729 Vdd.t731 Vdd.t730 pfet_03v3
**devattr s=44000,1176 d=26000,604
X31 SARlogic_0.dffrs_3.nand3_6.C.t3 Clk.t1 Vdd.t43 Vdd.t42 pfet_03v3
**devattr s=26000,604 d=44000,1176
X32 Vdd.t419 Reset.t2 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t418 pfet_03v3
**devattr s=26000,604 d=26000,604
X33 Vdd.t509 a_33337_30170.t4 a_33257_33628.t2 Vdd.t508 pfet_03v3
**devattr s=26000,604 d=26000,604
X34 SARlogic_0.dffrs_13.Qb.t3 SARlogic_0.dffrs_0.d.t4 Vdd.t824 Vdd.t823 pfet_03v3
**devattr s=44000,1176 d=26000,604
X35 Vdd.t754 a_n10831_4320 Comp_out.t7 Vdd.t753 pfet_03v3
**devattr s=18700,450 d=18700,450
X36 a_10639_28100 a_9083_28820.t4 Vdd.t912 Vdd.t911 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X37 a_5987_21414 SARlogic_0.dffrs_9.nand3_6.C.t4 a_5803_21414 Vss.t647 nfet_03v3
**devattr s=10400,304 d=10400,304
X38 a_275_7428 SARlogic_0.dffrs_2.nand3_8.C.t4 Vss.t659 Vss.t658 nfet_03v3
**devattr s=17600,576 d=10400,304
X39 adc_PISO_0.2inmux_5.OUT.t0 a_30255_29264.t4 Vss.t258 Vss.t257 nfet_03v3
**devattr s=17600,576 d=17600,576
X40 SARlogic_0.dffrs_10.nand3_6.C.t3 SARlogic_0.d0.t4 Vdd.t944 Vdd.t943 pfet_03v3
**devattr s=26000,604 d=44000,1176
X41 SARlogic_0.d1.t2 SARlogic_0.dffrs_3.Qb.t4 Vdd.t167 Vdd.t166 pfet_03v3
**devattr s=44000,1176 d=26000,604
X42 a_12585_21414 Reset.t3 a_12401_21414 Vss.t318 nfet_03v3
**devattr s=10400,304 d=10400,304
X43 SARlogic_0.dffrs_3.Qb.t2 Reset.t4 a_5987_9634 Vss.t319 nfet_03v3
**devattr s=10400,304 d=17600,576
X44 SARlogic_0.dffrs_12.nand3_6.C.t3 SARlogic_0.dffrs_12.nand3_1.C Vdd.t884 Vdd.t883 pfet_03v3
**devattr s=44000,1176 d=26000,604
X45 SARlogic_0.dffrs_1.Qb.t1 Reset.t5 a_n2097_9634 Vss.t320 nfet_03v3
**devattr s=10400,304 d=17600,576
X46 a_n11637_11838 Vdd.t956 a_n11821_11838 Vss.t528 nfet_03v3
**devattr s=10400,304 d=10400,304
X47 a_n4551_35924 Vdd.t957 Vss.t527 Vss.t526 nfet_03v3
**devattr s=17600,576 d=10400,304
X48 SARlogic_0.dffrs_4.nand3_8.Z.t1 SARlogic_0.dffrs_4.nand3_8.C.t5 Vdd.t457 Vdd.t456 pfet_03v3
**devattr s=44000,1176 d=26000,604
X49 a_1761_19210 SARlogic_0.d3.t5 Vss.t59 Vss.t58 nfet_03v3
**devattr s=17600,576 d=10400,304
X50 a_14393_33720 a_14313_33628.t4 Vss.t372 Vss.t371 nfet_03v3
**devattr s=17600,576 d=10400,304
X51 a_9271_28100 SARlogic_0.d3.t6 a_9083_28820.t1 Vss.t57 nfet_03v3
**devattr s=17600,576 d=10400,304
X52 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t4 Vdd.t287 Vdd.t286 pfet_03v3
**devattr s=26000,604 d=44000,1176
X53 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_5.Qb.t4 Vdd.t846 Vdd.t845 pfet_03v3
**devattr s=44000,1176 d=26000,604
X54 a_12585_23619 SARlogic_0.dffrs_11.nand3_8.Z a_12401_23619 Vss.t118 nfet_03v3
**devattr s=10400,304 d=10400,304
X55 adc_PISO_0.dffrs_1.Qb adc_PISO_0.dffrs_1.Q.t4 Vdd.t844 Vdd.t843 pfet_03v3
**devattr s=44000,1176 d=26000,604
X56 Vdd.t377 SARlogic_0.dffrs_14.nand3_6.C.t4 SARlogic_0.d5.t0 Vdd.t376 pfet_03v3
**devattr s=26000,604 d=26000,604
X57 a_275_14043 Vdd.t958 Vss.t525 Vss.t524 nfet_03v3
**devattr s=17600,576 d=10400,304
X58 a_33257_29218.t1 a_33337_30170.t5 a_33521_31515 Vss.t384 nfet_03v3
**devattr s=10400,304 d=17600,576
X59 SARlogic_0.dffrs_0.Qb.t3 Reset.t6 a_n6139_9634 Vss.t321 nfet_03v3
**devattr s=10400,304 d=17600,576
X60 a_14393_35925 Vdd.t959 Vss.t523 Vss.t522 nfet_03v3
**devattr s=17600,576 d=10400,304
X61 SARlogic_0.dffrs_3.nand3_8.C.t1 SARlogic_0.dffrs_3.nand3_6.C.t4 Vdd.t383 Vdd.t382 pfet_03v3
**devattr s=44000,1176 d=26000,604
X62 a_9083_31160.t1 inv2_0.out.t3 a_9271_30440 Vss.t549 nfet_03v3
**devattr s=10400,304 d=17600,576
X63 a_23865_30170.t1 a_23785_29218.t4 Vdd.t217 Vdd.t216 pfet_03v3
**devattr s=44000,1176 d=26000,604
X64 a_18743_28100 a_17849_29020 Vss.t456 Vss.t455 nfet_03v3
**devattr s=17600,576 d=10400,304
X65 Vdd.t549 a_40051_37983 Piso_out.t7 Vdd.t548 pfet_03v3
**devattr s=18700,450 d=18700,450
X66 a_9845_19210 SARlogic_0.d1.t5 Vss.t428 Vss.t427 nfet_03v3
**devattr s=17600,576 d=10400,304
X67 SARlogic_0.dffrs_3.nand3_6.C.t0 SARlogic_0.dffrs_3.nand3_1.C.t4 Vdd.t223 Vdd.t222 pfet_03v3
**devattr s=44000,1176 d=26000,604
X68 a_42729_31423.t0 a_42729_33628.t4 Vdd.t193 Vdd.t192 pfet_03v3
**devattr s=44000,1176 d=26000,604
X69 a_29583_30440 a_28027_31160.t4 Vdd.t812 Vdd.t811 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X70 SARlogic_0.dffrs_13.Qb.t2 Vdd.t726 Vdd.t728 Vdd.t727 pfet_03v3
**devattr s=26000,604 d=44000,1176
X71 a_23785_29218.t0 a_23785_31423.t4 Vdd.t237 Vdd.t236 pfet_03v3
**devattr s=44000,1176 d=26000,604
X72 Vdd.t121 a_20111_30440 a_20971_29984 Vdd.t120 pfet_03v3
**devattr s=31200,704 d=52800,1376
X73 a_n9429_n2007.t7 Vin1.t0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t9 Vss.t260 nfet_03v3
**devattr s=15600,404 d=15600,404
X74 a_28027_31160.t1 inv2_0.out.t4 a_28215_30440 Vss.t550 nfet_03v3
**devattr s=10400,304 d=17600,576
X75 SARlogic_0.dffrs_10.nand3_6.C.t0 SARlogic_0.dffrs_10.nand3_1.C Vdd.t123 Vdd.t122 pfet_03v3
**devattr s=44000,1176 d=26000,604
X76 a_42729_33628.t2 Vdd.t723 Vdd.t725 Vdd.t724 pfet_03v3
**devattr s=44000,1176 d=26000,604
X77 a_n4631_33627.t0 a_n4631_31422.t4 a_n4367_35924 Vss.t670 nfet_03v3
**devattr s=10400,304 d=17600,576
X78 a_12401_17004 SARlogic_0.dffrs_11.nand3_8.C.t4 Vss.t184 Vss.t183 nfet_03v3
**devattr s=17600,576 d=10400,304
X79 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t0 a_4501_17004 Vss.t77 nfet_03v3
**devattr s=10400,304 d=17600,576
X80 a_n8305_30439 a_n9861_31159.t4 Vdd.t191 Vdd.t190 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X81 a_n6139_19213 SARlogic_0.dffrs_14.nand3_8.C.t4 a_n6323_19213 Vss.t272 nfet_03v3
**devattr s=10400,304 d=10400,304
X82 a_n201_28099 a_n1095_29019 Vss.t547 Vss.t546 nfet_03v3
**devattr s=17600,576 d=10400,304
X83 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_3.Qb.t5 Vdd.t169 Vdd.t168 pfet_03v3
**devattr s=44000,1176 d=26000,604
X84 SARlogic_0.d1.t0 SARlogic_0.dffrs_10.Qb Vdd.t127 Vdd.t126 pfet_03v3
**devattr s=26000,604 d=44000,1176
X85 Vdd.t722 Vdd.t720 SARlogic_0.dffrs_13.nand3_8.Z.t3 Vdd.t721 pfet_03v3
**devattr s=26000,604 d=26000,604
X86 SARlogic_0.dffrs_5.Qb.t1 Reset.t7 Vdd.t421 Vdd.t420 pfet_03v3
**devattr s=26000,604 d=44000,1176
X87 a_1167_30439 a_n389_31159.t4 Vdd.t107 Vdd.t106 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X88 SARlogic_0.dffrs_9.nand3_8.C.t1 SARlogic_0.dffrs_9.nand3_8.Z a_4501_19209 Vss.t112 nfet_03v3
**devattr s=10400,304 d=17600,576
X89 SARlogic_0.dffrs_0.nand3_8.C.t2 SARlogic_0.dffrs_0.nand3_6.C.t4 Vdd.t33 Vdd.t32 pfet_03v3
**devattr s=44000,1176 d=26000,604
X90 a_12401_19209 SARlogic_0.dffrs_11.nand3_6.C.t4 Vss.t40 Vss.t39 nfet_03v3
**devattr s=17600,576 d=10400,304
X91 a_33337_31515 a_33257_31423.t4 Vss.t405 Vss.t404 nfet_03v3
**devattr s=17600,576 d=10400,304
X92 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_13.Qb.t4 Vdd.t814 Vdd.t813 pfet_03v3
**devattr s=44000,1176 d=26000,604
X93 SARlogic_0.dffrs_3.nand3_8.C.t3 SARlogic_0.dffrs_3.nand3_8.Z.t5 a_4501_9633 Vss.t411 nfet_03v3
**devattr s=10400,304 d=17600,576
X94 a_10639_30440 a_9083_31160.t4 Vss.t580 Vss.t579 nfet_03v3
**devattr s=17600,576 d=17600,576
X95 Vdd.t461 SARlogic_0.dffrs_5.nand3_8.C.t6 SARlogic_0.dffrs_5.Qb.t3 Vdd.t460 pfet_03v3
**devattr s=26000,604 d=26000,604
X96 Piso_out.t3 a_40051_37983 Vss.t420 Vss.t419 nfet_03v3
**devattr s=9350,280 d=9350,280
X97 Vss.t87 a_29583_30440 a_30255_29264.t0 Vss.t86 nfet_03v3
**devattr s=17600,576 d=17600,576
X98 Vss.t341 adc_PISO_0.2inmux_1.Bit.t5 a_37687_30440 Vss.t340 nfet_03v3
**devattr s=10400,304 d=17600,576
X99 SARlogic_0.dffrs_8.nand3_6.C.t3 SARlogic_0.d2.t5 Vdd.t307 Vdd.t306 pfet_03v3
**devattr s=26000,604 d=44000,1176
X100 Vdd.t756 a_n1095_29019 a_n389_28819.t2 Vdd.t755 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X101 Vss.t83 a_1167_30439 a_1839_29263.t0 Vss.t82 nfet_03v3
**devattr s=17600,576 d=17600,576
X102 a_5987_9634 SARlogic_0.dffrs_3.nand3_8.C.t4 a_5803_9634 Vss.t401 nfet_03v3
**devattr s=10400,304 d=10400,304
X103 SARlogic_0.dffrs_0.nand3_6.C.t1 SARlogic_0.dffrs_0.nand3_1.C.t4 Vdd.t367 Vdd.t366 pfet_03v3
**devattr s=44000,1176 d=26000,604
X104 SARlogic_0.dffrs_5.nand3_1.C.t2 Vdd.t717 Vdd.t719 Vdd.t718 pfet_03v3
**devattr s=44000,1176 d=26000,604
X105 SARlogic_0.dffrs_3.nand3_1.C.t2 SARlogic_0.dffrs_3.nand3_6.C.t5 Vdd.t385 Vdd.t384 pfet_03v3
**devattr s=26000,604 d=44000,1176
X106 a_20971_29984 a_20111_28100 a_20783_29264.t1 Vdd.t29 pfet_03v3
**devattr s=52800,1376 d=31200,704
X107 a_n3065_31515 adc_PISO_0.2inmux_2.Bit.t4 Vss.t34 Vss.t33 nfet_03v3
**devattr s=17600,576 d=10400,304
X108 SARlogic_0.dffrs_12.Q.t3 SARlogic_0.dffrs_12.Qb Vdd.t153 Vdd.t152 pfet_03v3
**devattr s=26000,604 d=44000,1176
X109 SARlogic_0.dffrs_12.nand3_8.Z Vss.t687 Vdd.t11 Vdd.t10 pfet_03v3
**devattr s=26000,604 d=44000,1176
X110 a_4921_30169.t1 adc_PISO_0.2inmux_2.OUT.t2 a_5105_29309 Vss.t148 nfet_03v3
**devattr s=10400,304 d=17600,576
X111 Vdd.t197 a_27321_29020 a_28027_28820.t0 Vdd.t196 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X112 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t4 Vdd.t87 Vdd.t86 pfet_03v3
**devattr s=26000,604 d=44000,1176
X113 a_n2881_31515 a_n4631_29217.t4 a_n3065_31515 Vss.t421 nfet_03v3
**devattr s=10400,304 d=10400,304
X114 a_12585_7428 Reset.t8 a_12401_7428 Vss.t322 nfet_03v3
**devattr s=10400,304 d=10400,304
X115 SARlogic_0.dffrs_10.Qb Reset.t9 a_10029_19210 Vss.t323 nfet_03v3
**devattr s=10400,304 d=17600,576
X116 a_17849_29020 inv2_0.out.t5 Vdd.t758 Vdd.t757 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X117 SARlogic_0.dffrs_3.nand3_8.Z.t3 SARlogic_0.dffrs_3.nand3_8.C.t5 Vdd.t521 Vdd.t520 pfet_03v3
**devattr s=44000,1176 d=26000,604
X118 a_4317_17004 SARlogic_0.dffrs_9.nand3_8.C.t4 Vss.t442 Vss.t441 nfet_03v3
**devattr s=17600,576 d=10400,304
X119 Vdd.t423 Reset.t10 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t422 pfet_03v3
**devattr s=26000,604 d=26000,604
X120 SARlogic_0.dffrs_7.nand3_8.C.t3 SARlogic_0.dffrs_7.nand3_6.C.t4 Vdd.t579 Vdd.t578 pfet_03v3
**devattr s=44000,1176 d=26000,604
X121 SARlogic_0.d3.t1 SARlogic_0.dffrs_8.Qb Vdd.t131 Vdd.t130 pfet_03v3
**devattr s=26000,604 d=44000,1176
X122 Vdd.t445 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t1 Vdd.t444 pfet_03v3
**devattr s=10400,304 d=10400,304
X123 a_14393_30170.t1 adc_PISO_0.2inmux_3.OUT.t2 Vdd.t267 Vdd.t266 pfet_03v3
**devattr s=26000,604 d=44000,1176
X124 Vdd.t89 SARlogic_0.dffrs_8.nand3_6.C.t5 SARlogic_0.d3.t0 Vdd.t88 pfet_03v3
**devattr s=26000,604 d=26000,604
X125 a_4317_19209 SARlogic_0.dffrs_9.nand3_6.C.t5 Vss.t649 Vss.t648 nfet_03v3
**devattr s=17600,576 d=10400,304
X126 a_459_7428 Reset.t11 a_275_7428 Vss.t324 nfet_03v3
**devattr s=10400,304 d=10400,304
X127 a_n9429_n2007.t18 Vin2.t0 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t263 nfet_03v3
**devattr s=15600,404 d=15600,404
X128 Vdd.t45 Clk.t2 SARlogic_0.dffrs_5.nand3_8.C.t0 Vdd.t44 pfet_03v3
**devattr s=26000,604 d=26000,604
X129 a_33257_31423.t3 Clk_piso.t0 Vdd.t876 Vdd.t875 pfet_03v3
**devattr s=26000,604 d=44000,1176
X130 adc_PISO_0.2inmux_1.Bit.t3 Vdd.t714 Vdd.t716 Vdd.t715 pfet_03v3
**devattr s=44000,1176 d=26000,604
X131 SARlogic_0.dffrs_8.nand3_6.C.t0 SARlogic_0.dffrs_8.nand3_1.C Vdd.t129 Vdd.t128 pfet_03v3
**devattr s=44000,1176 d=26000,604
X132 SARlogic_0.dffrs_12.Qb Reset.t12 a_18113_19210 Vss.t325 nfet_03v3
**devattr s=10400,304 d=17600,576
X133 a_14313_29218.t1 a_14393_30170.t4 Vdd.t329 Vdd.t328 pfet_03v3
**devattr s=26000,604 d=44000,1176
X134 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t1 a_n7971_249 a_n8059_341 Vss.t134 nfet_03v3
**devattr s=35200,976 d=20800,504
X135 SARlogic_0.dffrs_3.nand3_1.C.t3 Vdd.t711 Vdd.t713 Vdd.t712 pfet_03v3
**devattr s=44000,1176 d=26000,604
X136 Vdd.t587 SARlogic_0.dffrs_9.nand3_8.C.t5 SARlogic_0.dffrs_9.Qb Vdd.t586 pfet_03v3
**devattr s=26000,604 d=26000,604
X137 SARlogic_0.dffrs_5.nand3_6.C.t1 Clk.t3 a_12585_11838 Vss.t24 nfet_03v3
**devattr s=10400,304 d=17600,576
X138 Vdd.t425 Reset.t13 SARlogic_0.dffrs_5.nand3_6.C.t2 Vdd.t424 pfet_03v3
**devattr s=26000,604 d=26000,604
X139 Vdd.t387 SARlogic_0.dffrs_3.nand3_6.C.t6 SARlogic_0.dffrs_4.d.t2 Vdd.t386 pfet_03v3
**devattr s=26000,604 d=26000,604
X140 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_8.C.t5 Vdd.t491 Vdd.t490 pfet_03v3
**devattr s=44000,1176 d=26000,604
X141 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t1 Vdd.t259 Vdd.t258 pfet_03v3
**devattr s=26000,604 d=44000,1176
X142 a_33257_33628.t1 a_33257_31423.t5 Vdd.t525 Vdd.t524 pfet_03v3
**devattr s=26000,604 d=44000,1176
X143 a_6591_31515 a_4841_29217.t4 a_6407_31515 Vss.t629 nfet_03v3
**devattr s=10400,304 d=10400,304
X144 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_1.Qb.t5 Vdd.t371 Vdd.t370 pfet_03v3
**devattr s=44000,1176 d=26000,604
X145 SARlogic_0.dffrs_14.nand3_6.C.t3 SARlogic_0.d4.t4 a_n7625_21417 Vss.t634 nfet_03v3
**devattr s=10400,304 d=17600,576
X146 a_n6323_21417 SARlogic_0.dffrs_13.Qb.t5 Vss.t587 Vss.t586 nfet_03v3
**devattr s=17600,576 d=10400,304
X147 a_13887_21414 SARlogic_0.dffrs_4.Qb.t4 Vss.t681 Vss.t680 nfet_03v3
**devattr s=17600,576 d=10400,304
X148 Vdd.t289 SARlogic_0.dffrs_10.nand3_6.C.t5 SARlogic_0.d1.t3 Vdd.t288 pfet_03v3
**devattr s=26000,604 d=26000,604
X149 Vdd.t427 Reset.t14 SARlogic_0.dffrs_12.nand3_6.C.t2 Vdd.t426 pfet_03v3
**devattr s=26000,604 d=26000,604
X150 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t1 a_n9429_n2007.t19 Vss.t261 nfet_03v3
**devattr s=15600,404 d=15600,404
X151 a_n3583_9633 Clk.t4 a_n3767_9633 Vss.t25 nfet_03v3
**devattr s=10400,304 d=10400,304
X152 a_n6139_9634 SARlogic_0.dffrs_0.nand3_8.C.t4 a_n6323_9634 Vss.t60 nfet_03v3
**devattr s=10400,304 d=10400,304
X153 SARlogic_0.dffrs_8.Qb Reset.t15 a_1945_19210 Vss.t326 nfet_03v3
**devattr s=10400,304 d=17600,576
X154 a_44295_33720 Vdd.t960 Vss.t521 Vss.t520 nfet_03v3
**devattr s=17600,576 d=10400,304
X155 a_n7445_29983 a_n8305_30439 Vdd.t139 Vdd.t138 pfet_03v3
**devattr s=52800,1376 d=31200,704
X156 a_23785_29218.t1 a_23865_30170.t4 a_24049_31515 Vss.t604 nfet_03v3
**devattr s=10400,304 d=17600,576
X157 a_1945_19210 SARlogic_0.dffrs_8.nand3_8.C.t4 a_1761_19210 Vss.t127 nfet_03v3
**devattr s=10400,304 d=10400,304
X158 a_5105_35924 a_4921_30169.t4 a_4921_35924 Vss.t657 nfet_03v3
**devattr s=10400,304 d=10400,304
X159 a_n201_30439 adc_PISO_0.2inmux_2.Bit.t5 Vss.t36 Vss.t35 nfet_03v3
**devattr s=17600,576 d=10400,304
X160 Vdd.t23 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_1.C Vdd.t22 pfet_03v3
**devattr s=26000,604 d=26000,604
X161 SARlogic_0.dffrs_7.nand3_8.C.t1 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t279 Vdd.t278 pfet_03v3
**devattr s=26000,604 d=44000,1176
X162 a_4501_11838 Reset.t16 a_4317_11838 Vss.t327 nfet_03v3
**devattr s=10400,304 d=10400,304
X163 a_42993_33720 Vdd.t961 a_42809_33720 Vss.t519 nfet_03v3
**devattr s=10400,304 d=10400,304
X164 a_4921_35924 Vdd.t962 Vss.t518 Vss.t517 nfet_03v3
**devattr s=17600,576 d=10400,304
X165 adc_PISO_0.dffrs_4.Qb adc_PISO_0.2inmux_1.Bit.t6 Vdd.t453 Vdd.t452 pfet_03v3
**devattr s=44000,1176 d=26000,604
X166 a_459_14043 SARlogic_0.dffrs_2.nand3_8.Z.t4 a_275_14043 Vss.t200 nfet_03v3
**devattr s=10400,304 d=10400,304
X167 a_28215_30440 adc_PISO_0.dffrs_3.Q.t4 Vss.t445 Vss.t444 nfet_03v3
**devattr s=17600,576 d=10400,304
X168 a_39727_29264.t2 a_39055_28100 a_39915_29984 Vdd.t281 pfet_03v3
**devattr s=31200,704 d=52800,1376
X169 a_8543_21414 Reset.t17 a_8359_21414 Vss.t328 nfet_03v3
**devattr s=10400,304 d=10400,304
X170 a_n7809_9633 SARlogic_0.dffrs_0.nand3_6.C.t5 Vss.t15 Vss.t14 nfet_03v3
**devattr s=17600,576 d=10400,304
X171 comparator_no_offsetcal_0.no_offsetLatch_0.Vq a_n9933_n2099 a_n10021_n2007 Vss.t217 nfet_03v3
**devattr s=26400,776 d=15600,404
X172 SARlogic_0.dffrs_0.nand3_1.C.t3 Vdd.t708 Vdd.t710 Vdd.t709 pfet_03v3
**devattr s=44000,1176 d=26000,604
X173 a_n7809_17007 SARlogic_0.dffrs_14.nand3_8.C.t5 Vss.t274 Vss.t273 nfet_03v3
**devattr s=17600,576 d=10400,304
X174 a_42993_35925 a_42809_30170.t4 a_42809_35925 Vss.t639 nfet_03v3
**devattr s=10400,304 d=10400,304
X175 a_33257_31423.t2 a_33257_33628.t4 Vdd.t820 Vdd.t819 pfet_03v3
**devattr s=44000,1176 d=26000,604
X176 a_28215_28100 SARlogic_0.d1.t6 a_28027_28820.t2 Vss.t429 nfet_03v3
**devattr s=17600,576 d=10400,304
X177 Vdd.t707 Vdd.t705 a_23865_30170.t2 Vdd.t706 pfet_03v3
**devattr s=26000,604 d=26000,604
X178 a_8543_23619 SARlogic_0.dffrs_10.nand3_8.Z a_8359_23619 Vss.t276 nfet_03v3
**devattr s=10400,304 d=10400,304
X179 a_10029_19210 SARlogic_0.dffrs_10.nand3_8.C.t4 a_9845_19210 Vss.t244 nfet_03v3
**devattr s=10400,304 d=10400,304
X180 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_8.C.t5 Vdd.t319 Vdd.t318 pfet_03v3
**devattr s=44000,1176 d=26000,604
X181 a_33257_33628.t3 Vdd.t702 Vdd.t704 Vdd.t703 pfet_03v3
**devattr s=44000,1176 d=26000,604
X182 Vdd.t878 Clk_piso.t1 a_23785_29218.t3 Vdd.t877 pfet_03v3
**devattr s=26000,604 d=26000,604
X183 SARlogic_0.d5.t2 SARlogic_0.dffrs_14.Qb a_n6139_21417 Vss.t265 nfet_03v3
**devattr s=10400,304 d=17600,576
X184 a_44295_31516 adc_PISO_0.serial_out.t4 Vss.t641 Vss.t640 nfet_03v3
**devattr s=17600,576 d=10400,304
X185 a_n4367_35924 a_n4551_30169.t4 a_n4551_35924 Vss.t226 nfet_03v3
**devattr s=10400,304 d=10400,304
X186 a_n4551_30169.t3 a_n4631_29217.t5 Vdd.t551 Vdd.t550 pfet_03v3
**devattr s=44000,1176 d=26000,604
X187 a_12585_17004 Reset.t18 a_12401_17004 Vss.t329 nfet_03v3
**devattr s=10400,304 d=10400,304
X188 a_40051_37983 adc_PISO_0.serial_out.t5 Vss.t643 Vss.t642 nfet_03v3
**devattr s=9350,280 d=17000,540
X189 a_8377_29020 inv2_0.out.t6 Vss.t552 Vss.t551 nfet_03v3
**devattr s=17600,576 d=17600,576
X190 SARlogic_0.dffrs_0.nand3_8.Z.t3 SARlogic_0.dffrs_0.d.t5 Vdd.t826 Vdd.t825 pfet_03v3
**devattr s=26000,604 d=44000,1176
X191 a_14393_29310 a_14313_29218.t4 Vss.t252 Vss.t251 nfet_03v3
**devattr s=17600,576 d=10400,304
X192 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t2 Vdd.t261 Vdd.t260 pfet_03v3
**devattr s=26000,604 d=44000,1176
X193 a_12585_19209 SARlogic_0.dffrs_12.Q.t4 a_12401_19209 Vss.t53 nfet_03v3
**devattr s=10400,304 d=10400,304
X194 a_39727_29264.t0 a_39055_28100 Vss.t216 Vss.t215 nfet_03v3
**devattr s=17600,576 d=17600,576
X195 a_11499_29984 a_10639_28100 a_11311_29264.t2 Vdd.t599 pfet_03v3
**devattr s=52800,1376 d=31200,704
X196 a_n6555_341 a_n6755_249 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t175 nfet_03v3
**devattr s=20800,504 d=35200,976
X197 Vdd.t804 SARlogic_0.dffrs_5.nand3_8.Z.t4 SARlogic_0.dffrs_5.nand3_1.C.t3 Vdd.t803 pfet_03v3
**devattr s=26000,604 d=26000,604
X198 a_n10151_9634 SARlogic_0.dffrs_13.nand3_8.C.t4 a_n10335_9634 Vss.t13 nfet_03v3
**devattr s=10400,304 d=10400,304
X199 SARlogic_0.d2.t2 SARlogic_0.dffrs_9.Qb Vdd.t822 Vdd.t821 pfet_03v3
**devattr s=26000,604 d=44000,1176
X200 adc_PISO_0.2inmux_1.Bit.t1 adc_PISO_0.dffrs_4.Qb a_35007_33720 Vss.t460 nfet_03v3
**devattr s=10400,304 d=17600,576
X201 adc_PISO_0.2inmux_0.OUT.t1 a_n7633_29263.t4 Vdd.t776 Vdd.t775 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X202 SARlogic_0.d4.t2 SARlogic_0.dffrs_0.Qb.t4 Vdd.t229 Vdd.t228 pfet_03v3
**devattr s=44000,1176 d=26000,604
X203 SARlogic_0.dffrs_0.nand3_8.C.t1 SARlogic_0.dffrs_0.nand3_8.Z.t4 Vdd.t125 Vdd.t124 pfet_03v3
**devattr s=26000,604 d=44000,1176
X204 a_36793_29020 inv2_0.out.t7 Vdd.t760 Vdd.t759 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X205 Vdd.t569 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t7 Vdd.t568 pfet_03v3
**devattr s=10400,304 d=10400,304
X206 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t5 Vdd.t379 Vdd.t378 pfet_03v3
**devattr s=26000,604 d=44000,1176
X207 SARlogic_0.dffrs_5.nand3_8.Z.t0 SARlogic_0.dffrs_4.Q.t4 Vdd.t225 Vdd.t224 pfet_03v3
**devattr s=26000,604 d=44000,1176
X208 a_n9429_n2007.t20 Vin2.t2 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t262 nfet_03v3
**devattr s=15600,404 d=15600,404
X209 SARlogic_0.dffrs_0.nand3_6.C.t2 Clk.t5 Vdd.t47 Vdd.t46 pfet_03v3
**devattr s=26000,604 d=44000,1176
X210 a_n4551_30169.t0 adc_PISO_0.2inmux_0.OUT.t2 Vdd.t199 Vdd.t198 pfet_03v3
**devattr s=26000,604 d=44000,1176
X211 SARlogic_0.dffrs_0.Q.t1 Vdd.t699 Vdd.t701 Vdd.t700 pfet_03v3
**devattr s=44000,1176 d=26000,604
X212 adc_PISO_0.dffrs_3.Q.t3 Vdd.t696 Vdd.t698 Vdd.t697 pfet_03v3
**devattr s=44000,1176 d=26000,604
X213 a_18555_28820.t3 SARlogic_0.d2.t6 Vdd.t309 Vdd.t308 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X214 a_18113_21414 SARlogic_0.dffrs_12.nand3_6.C.t5 a_17929_21414 Vss.t266 nfet_03v3
**devattr s=10400,304 d=10400,304
X215 a_23785_31423.t3 Clk_piso.t2 Vdd.t880 Vdd.t879 pfet_03v3
**devattr s=26000,604 d=44000,1176
X216 SARlogic_0.dffrs_13.nand3_8.Z.t1 Vss.t100 a_n11637_7428 Vss.t101 nfet_03v3
**devattr s=10400,304 d=17600,576
X217 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t331 Vdd.t330 pfet_03v3
**devattr s=17600,576 d=17600,576
X218 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_8.C.t5 Vdd.t187 Vdd.t186 pfet_03v3
**devattr s=44000,1176 d=26000,604
X219 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x3.out Vss.t287 Vss.t286 nfet_03v3
**devattr s=17600,576 d=17600,576
X220 SARlogic_0.dffrs_12.nand3_6.C.t0 Vss.t98 a_16627_21414 Vss.t99 nfet_03v3
**devattr s=10400,304 d=17600,576
X221 a_n3767_9633 SARlogic_0.dffrs_1.nand3_6.C.t4 Vss.t103 Vss.t102 nfet_03v3
**devattr s=17600,576 d=10400,304
X222 Vdd.t527 a_33257_31423.t6 adc_PISO_0.2inmux_1.Bit.t0 Vdd.t526 pfet_03v3
**devattr s=26000,604 d=26000,604
X223 SARlogic_0.dffrs_9.Qb Reset.t19 a_5987_19210 Vss.t330 nfet_03v3
**devattr s=10400,304 d=17600,576
X224 a_23785_33628.t0 a_23785_31423.t5 Vdd.t239 Vdd.t238 pfet_03v3
**devattr s=26000,604 d=44000,1176
X225 Vdd.t429 Reset.t20 SARlogic_0.dffrs_8.nand3_6.C.t1 Vdd.t428 pfet_03v3
**devattr s=26000,604 d=26000,604
X226 SARlogic_0.dffrs_14.Qb SARlogic_0.d5.t4 Vdd.t299 Vdd.t298 pfet_03v3
**devattr s=44000,1176 d=26000,604
X227 a_n2281_19210 SARlogic_0.d4.t5 Vss.t636 Vss.t635 nfet_03v3
**devattr s=17600,576 d=10400,304
X228 a_n3583_14043 SARlogic_0.dffrs_1.nand3_8.Z.t4 a_n3767_14043 Vss.t147 nfet_03v3
**devattr s=10400,304 d=10400,304
X229 a_n7633_29263.t3 a_n8305_28099 a_n7445_29983 Vdd.t323 pfet_03v3
**devattr s=31200,704 d=52800,1376
X230 SARlogic_0.dffrs_2.nand3_8.Z.t0 SARlogic_0.dffrs_2.d.t4 Vdd.t39 Vdd.t38 pfet_03v3
**devattr s=26000,604 d=44000,1176
X231 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t6 a_16627_23619 Vss.t267 nfet_03v3
**devattr s=10400,304 d=17600,576
X232 SARlogic_0.dffrs_11.Qb SARlogic_0.d0.t5 Vdd.t946 Vdd.t945 pfet_03v3
**devattr s=44000,1176 d=26000,604
X233 adc_PISO_0.dffrs_4.Qb Vdd.t963 a_35007_31516 Vss.t516 nfet_03v3
**devattr s=10400,304 d=17600,576
X234 SARlogic_0.dffrs_5.Q.t3 Vdd.t693 Vdd.t695 Vdd.t694 pfet_03v3
**devattr s=44000,1176 d=26000,604
X235 Vdd.t431 Reset.t21 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t430 pfet_03v3
**devattr s=26000,604 d=26000,604
X236 a_n389_31159.t1 inv2_0.out.t8 Vdd.t762 Vdd.t761 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X237 a_n7625_21417 Reset.t22 a_n7809_21417 Vss.t331 nfet_03v3
**devattr s=10400,304 d=10400,304
X238 Vdd.t327 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_1.C Vdd.t326 pfet_03v3
**devattr s=26000,604 d=26000,604
X239 adc_PISO_0.dffrs_0.Qb Vdd.t964 a_n2881_31515 Vss.t515 nfet_03v3
**devattr s=10400,304 d=17600,576
X240 a_1761_21414 SARlogic_0.dffrs_1.Qb.t6 Vss.t289 Vss.t288 nfet_03v3
**devattr s=17600,576 d=10400,304
X241 a_n10567_29019 inv2_0.out.t9 Vss.t554 Vss.t553 nfet_03v3
**devattr s=17600,576 d=17600,576
X242 a_n201_28099 SARlogic_0.d4.t6 a_n389_28819.t3 Vss.t637 nfet_03v3
**devattr s=17600,576 d=10400,304
X243 SARlogic_0.dffrs_12.Q.t1 SARlogic_0.dffrs_5.Qb.t5 Vdd.t848 Vdd.t847 pfet_03v3
**devattr s=44000,1176 d=26000,604
X244 a_n11821_14043 Reset.t23 Vss.t333 Vss.t332 nfet_03v3
**devattr s=17600,576 d=10400,304
X245 a_33521_33720 Vdd.t965 a_33337_33720 Vss.t514 nfet_03v3
**devattr s=10400,304 d=10400,304
X246 Vdd.t49 Clk.t6 SARlogic_0.dffrs_4.nand3_8.C.t0 Vdd.t48 pfet_03v3
**devattr s=26000,604 d=26000,604
X247 SARlogic_0.dffrs_1.nand3_8.Z.t2 SARlogic_0.dffrs_0.Q.t4 Vdd.t774 Vdd.t773 pfet_03v3
**devattr s=26000,604 d=44000,1176
X248 SARlogic_0.dffrs_0.Q.t3 SARlogic_0.dffrs_0.Qb.t5 Vdd.t231 Vdd.t230 pfet_03v3
**devattr s=26000,604 d=44000,1176
X249 adc_PISO_0.dffrs_3.Qb adc_PISO_0.dffrs_3.Q.t5 Vdd.t591 Vdd.t590 pfet_03v3
**devattr s=44000,1176 d=26000,604
X250 a_30255_29264.t3 a_29583_28100 a_30443_29984 Vdd.t249 pfet_03v3
**devattr s=31200,704 d=52800,1376
X251 a_5803_11838 Vdd.t966 Vss.t513 Vss.t512 nfet_03v3
**devattr s=17600,576 d=10400,304
X252 a_4841_33627.t1 a_4841_31422.t5 a_5105_35924 Vss.t359 nfet_03v3
**devattr s=10400,304 d=17600,576
X253 a_1839_29263.t3 a_1167_28099 a_2027_29983 Vdd.t283 pfet_03v3
**devattr s=31200,704 d=52800,1376
X254 a_12401_11838 SARlogic_0.dffrs_5.nand3_1.C.t5 Vss.t300 Vss.t299 nfet_03v3
**devattr s=17600,576 d=10400,304
X255 SARlogic_0.dffrs_3.nand3_6.C.t2 Clk.t7 a_4501_11838 Vss.t26 nfet_03v3
**devattr s=10400,304 d=17600,576
X256 Vdd.t433 Reset.t24 SARlogic_0.dffrs_4.nand3_6.C.t0 Vdd.t432 pfet_03v3
**devattr s=26000,604 d=26000,604
X257 a_33521_35925 a_33337_30170.t6 a_33337_35925 Vss.t385 nfet_03v3
**devattr s=10400,304 d=10400,304
X258 a_42809_30170.t2 adc_PISO_0.2inmux_1.OUT.t2 Vdd.t834 Vdd.t833 pfet_03v3
**devattr s=26000,604 d=44000,1176
X259 inv2_0.out.t0 Load.t0 Vss.t116 Vss.t115 nfet_03v3
**devattr s=17600,576 d=17600,576
X260 Vdd.t692 Vdd.t690 a_14393_30170.t3 Vdd.t691 pfet_03v3
**devattr s=26000,604 d=26000,604
X261 Comp_out.t3 a_n10831_4320 Vss.t543 Vss.t542 nfet_03v3
**devattr s=17000,540 d=9350,280
X262 Vdd.t808 a_33257_29218.t4 adc_PISO_0.dffrs_4.Qb Vdd.t807 pfet_03v3
**devattr s=26000,604 d=26000,604
X263 SARlogic_0.dffrs_11.nand3_8.C.t2 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t173 Vdd.t172 pfet_03v3
**devattr s=26000,604 d=44000,1176
X264 SARlogic_0.dffrs_10.nand3_6.C.t2 SARlogic_0.d0.t6 a_8543_21414 Vss.t682 nfet_03v3
**devattr s=10400,304 d=17600,576
X265 a_9845_21414 SARlogic_0.dffrs_3.Qb.t6 Vss.t120 Vss.t119 nfet_03v3
**devattr s=17600,576 d=10400,304
X266 a_16443_21414 SARlogic_0.dffrs_12.nand3_1.C Vss.t631 Vss.t630 nfet_03v3
**devattr s=17600,576 d=10400,304
X267 a_42729_29218.t1 a_42809_30170.t5 Vdd.t896 Vdd.t895 pfet_03v3
**devattr s=26000,604 d=44000,1176
X268 Piso_out.t6 a_40051_37983 Vdd.t547 Vdd.t546 pfet_03v3
**devattr s=18700,450 d=18700,450
X269 a_8359_7428 SARlogic_0.dffrs_4.nand3_8.C.t6 Vss.t352 Vss.t351 nfet_03v3
**devattr s=17600,576 d=10400,304
X270 Vdd.t882 Clk_piso.t3 a_14313_29218.t3 Vdd.t881 pfet_03v3
**devattr s=26000,604 d=26000,604
X271 SARlogic_0.dffrs_14.Qb Reset.t25 Vdd.t435 Vdd.t434 pfet_03v3
**devattr s=26000,604 d=44000,1176
X272 inv2_0.out.t1 Load.t1 Vdd.t375 Vdd.t374 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X273 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t6 a_8543_23619 Vss.t222 nfet_03v3
**devattr s=10400,304 d=17600,576
X274 a_16443_23619 SARlogic_0.dffrs_5.Qb.t6 Vss.t616 Vss.t615 nfet_03v3
**devattr s=17600,576 d=10400,304
X275 a_17929_19210 SARlogic_0.dffrs_12.Q.t5 Vss.t425 Vss.t424 nfet_03v3
**devattr s=17600,576 d=10400,304
X276 a_n9429_n2007.t21 Vin2.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t260 nfet_03v3
**devattr s=15600,404 d=15600,404
X277 a_6407_31515 adc_PISO_0.dffrs_1.Q.t5 Vss.t612 Vss.t611 nfet_03v3
**devattr s=17600,576 d=10400,304
X278 a_18555_31160.t1 inv2_0.out.t10 a_18743_30440 Vss.t555 nfet_03v3
**devattr s=10400,304 d=17600,576
X279 Vdd.t561 SARlogic_0.d1.t7 SARlogic_0.dffrs_9.nand3_8.C.t2 Vdd.t560 pfet_03v3
**devattr s=26000,604 d=26000,604
X280 Vdd.t437 Reset.t26 SARlogic_0.dffrs_0.nand3_8.Z.t1 Vdd.t436 pfet_03v3
**devattr s=26000,604 d=26000,604
X281 a_n6139_21417 SARlogic_0.dffrs_14.nand3_6.C.t6 a_n6323_21417 Vss.t293 nfet_03v3
**devattr s=10400,304 d=10400,304
X282 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t11 Vss.t434 Vss.t433 nfet_03v3
**devattr s=35200,976 d=35200,976
X283 SARlogic_0.dffrs_13.nand3_1.C.t1 SARlogic_0.dffrs_13.nand3_6.C.t4 a_n11637_14043 Vss.t625 nfet_03v3
**devattr s=10400,304 d=17600,576
X284 SARlogic_0.dffrs_0.nand3_1.C.t2 SARlogic_0.dffrs_0.nand3_6.C.t6 Vdd.t35 Vdd.t34 pfet_03v3
**devattr s=26000,604 d=44000,1176
X285 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t3 a_n7625_17007 Vss.t192 nfet_03v3
**devattr s=10400,304 d=17600,576
X286 adc_PISO_0.2inmux_5.OUT.t1 a_30255_29264.t5 Vdd.t339 Vdd.t338 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X287 a_n10335_9634 SARlogic_0.dffrs_0.d.t6 Vss.t596 Vss.t595 nfet_03v3
**devattr s=17600,576 d=10400,304
X288 a_42809_33720 a_42729_33628.t5 Vss.t607 Vss.t606 nfet_03v3
**devattr s=17600,576 d=10400,304
X289 Vdd.t689 Vdd.t687 a_4921_30169.t3 Vdd.t688 pfet_03v3
**devattr s=26000,604 d=26000,604
X290 a_4317_11838 SARlogic_0.dffrs_3.nand3_1.C.t5 Vss.t155 Vss.t154 nfet_03v3
**devattr s=17600,576 d=10400,304
X291 a_23865_31515 a_23785_31423.t6 Vss.t170 Vss.t169 nfet_03v3
**devattr s=17600,576 d=10400,304
X292 a_4921_30169.t2 a_4841_29217.t5 Vdd.t315 Vdd.t314 pfet_03v3
**devattr s=44000,1176 d=26000,604
X293 a_42993_29310 Vdd.t967 a_42809_29310 Vss.t511 nfet_03v3
**devattr s=10400,304 d=10400,304
X294 Vss.t74 a_20111_30440 a_20783_29264.t3 Vss.t73 nfet_03v3
**devattr s=17600,576 d=17600,576
X295 a_8359_21414 SARlogic_0.dffrs_10.nand3_1.C Vss.t76 Vss.t75 nfet_03v3
**devattr s=17600,576 d=10400,304
X296 a_42809_35925 Vdd.t968 Vss.t510 Vss.t509 nfet_03v3
**devattr s=17600,576 d=10400,304
X297 a_n9673_28099 a_n10567_29019 Vss.t283 Vss.t282 nfet_03v3
**devattr s=17600,576 d=10400,304
X298 a_8543_17004 Reset.t27 a_8359_17004 Vss.t334 nfet_03v3
**devattr s=10400,304 d=10400,304
X299 SARlogic_0.d1.t1 SARlogic_0.dffrs_10.Qb a_10029_21414 Vss.t78 nfet_03v3
**devattr s=10400,304 d=17600,576
X300 a_8359_23619 SARlogic_0.dffrs_3.Qb.t7 Vss.t122 Vss.t121 nfet_03v3
**devattr s=17600,576 d=10400,304
X301 a_n11637_7428 Vdd.t969 a_n11821_7428 Vss.t508 nfet_03v3
**devattr s=10400,304 d=10400,304
X302 Vdd.t601 a_17849_29020 a_18555_28820.t0 Vdd.t600 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X303 Vdd.t439 Reset.t28 SARlogic_0.dffrs_7.nand3_6.C.t2 Vdd.t438 pfet_03v3
**devattr s=26000,604 d=26000,604
X304 Vdd.t51 Clk.t8 SARlogic_0.dffrs_0.nand3_8.C.t3 Vdd.t50 pfet_03v3
**devattr s=26000,604 d=26000,604
X305 a_n201_30439 inv2_0.out.t11 a_n389_31159.t3 Vss.t556 nfet_03v3
**devattr s=17600,576 d=10400,304
X306 a_20111_28100 a_18555_28820.t4 Vss.t144 Vss.t143 nfet_03v3
**devattr s=17600,576 d=17600,576
X307 a_8543_19209 SARlogic_0.d0.t7 a_8359_19209 Vss.t683 nfet_03v3
**devattr s=10400,304 d=10400,304
X308 Vdd.t365 a_n10567_29019 a_n9861_28819.t0 Vdd.t364 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X309 Vdd.t27 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_1.C Vdd.t26 pfet_03v3
**devattr s=26000,604 d=26000,604
X310 a_n7809_23622 SARlogic_0.dffrs_13.Qb.t6 Vss.t589 Vss.t588 nfet_03v3
**devattr s=17600,576 d=10400,304
X311 Vss.t614 adc_PISO_0.dffrs_1.Q.t6 a_9271_30440 Vss.t613 nfet_03v3
**devattr s=10400,304 d=17600,576
X312 a_37499_28820.t2 SARlogic_0.d0.t8 a_37687_28100 Vss.t684 nfet_03v3
**devattr s=10400,304 d=17600,576
X313 Vdd.t277 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_1.C Vdd.t276 pfet_03v3
**devattr s=26000,604 d=26000,604
X314 SARlogic_0.dffrs_8.nand3_6.C.t2 SARlogic_0.d2.t7 a_459_21414 Vss.t236 nfet_03v3
**devattr s=10400,304 d=17600,576
X315 Vdd.t940 SARlogic_0.dffrs_12.nand3_8.C.t6 SARlogic_0.dffrs_12.Qb Vdd.t939 pfet_03v3
**devattr s=26000,604 d=26000,604
X316 Vdd.t686 Vdd.t684 a_n4551_30169.t2 Vdd.t685 pfet_03v3
**devattr s=26000,604 d=26000,604
X317 a_12401_9633 SARlogic_0.dffrs_5.nand3_6.C.t5 Vss.t533 Vss.t532 nfet_03v3
**devattr s=17600,576 d=10400,304
X318 a_n7809_11838 SARlogic_0.dffrs_0.nand3_1.C.t5 Vss.t285 Vss.t284 nfet_03v3
**devattr s=17600,576 d=10400,304
X319 Vdd.t441 Reset.t29 SARlogic_0.dffrs_0.nand3_6.C.t0 Vdd.t440 pfet_03v3
**devattr s=26000,604 d=26000,604
X320 Vdd.t483 SARlogic_0.dffrs_4.nand3_8.Z.t5 SARlogic_0.dffrs_4.nand3_1.C.t1 Vdd.t482 pfet_03v3
**devattr s=26000,604 d=26000,604
X321 a_1761_9634 SARlogic_0.dffrs_2.Q.t4 Vss.t365 Vss.t364 nfet_03v3
**devattr s=17600,576 d=10400,304
X322 Vdd.t241 a_23785_31423.t7 adc_PISO_0.dffrs_3.Q.t0 Vdd.t240 pfet_03v3
**devattr s=26000,604 d=26000,604
X323 SARlogic_0.dffrs_12.Q.t2 SARlogic_0.dffrs_12.Qb a_18113_21414 Vss.t110 nfet_03v3
**devattr s=10400,304 d=17600,576
X324 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t6 a_459_23619 Vss.t49 nfet_03v3
**devattr s=10400,304 d=17600,576
X325 Vdd.t443 Reset.t30 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t442 pfet_03v3
**devattr s=26000,604 d=26000,604
X326 Piso_out.t2 a_40051_37983 Vss.t418 Vss.t417 nfet_03v3
**devattr s=17000,540 d=9350,280
X327 Vdd.t53 Clk.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vdd.t52 pfet_03v3
**devattr s=14080,496 d=14080,496
X328 a_275_9633 SARlogic_0.dffrs_2.nand3_6.C.t5 Vss.t375 Vss.t374 nfet_03v3
**devattr s=17600,576 d=10400,304
X329 adc_PISO_0.dffrs_1.Q.t1 adc_PISO_0.dffrs_1.Qb Vdd.t159 Vdd.t158 pfet_03v3
**devattr s=26000,604 d=44000,1176
X330 a_4317_7428 SARlogic_0.dffrs_3.nand3_8.C.t6 Vss.t403 Vss.t402 nfet_03v3
**devattr s=17600,576 d=10400,304
X331 a_n3767_14043 Vdd.t970 Vss.t507 Vss.t506 nfet_03v3
**devattr s=17600,576 d=10400,304
X332 SARlogic_0.dffrs_8.Qb SARlogic_0.d3.t7 Vdd.t101 Vdd.t100 pfet_03v3
**devattr s=44000,1176 d=26000,604
X333 a_30443_29984 a_29583_30440 Vdd.t143 Vdd.t142 pfet_03v3
**devattr s=52800,1376 d=31200,704
X334 SARlogic_0.dffrs_2.Q.t1 Vdd.t681 Vdd.t683 Vdd.t682 pfet_03v3
**devattr s=44000,1176 d=26000,604
X335 SARlogic_0.d3.t2 SARlogic_0.dffrs_8.Qb a_1945_21414 Vss.t81 nfet_03v3
**devattr s=10400,304 d=17600,576
X336 a_2027_29983 a_1167_30439 Vdd.t135 Vdd.t134 pfet_03v3
**devattr s=52800,1376 d=31200,704
X337 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t8 Vin1.t1 a_n9429_n2007.t8 Vss.t261 nfet_03v3
**devattr s=15600,404 d=15600,404
X338 a_9271_30440 inv2_0.out.t12 a_9083_31160.t0 Vss.t557 nfet_03v3
**devattr s=17600,576 d=10400,304
X339 a_39055_28100 a_37499_28820.t4 Vss.t379 Vss.t378 nfet_03v3
**devattr s=17600,576 d=17600,576
X340 Vdd.t581 SARlogic_0.dffrs_7.nand3_6.C.t5 SARlogic_0.d4.t3 Vdd.t580 pfet_03v3
**devattr s=26000,604 d=26000,604
X341 comparator_no_offsetcal_0.no_offsetLatch_0.Vq comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t4 Vss.t435 nfet_03v3
**devattr s=20800,504 d=20800,504
X342 a_n7633_29263.t1 a_n8305_28099 Vss.t248 Vss.t247 nfet_03v3
**devattr s=17600,576 d=17600,576
X343 a_1945_21414 SARlogic_0.dffrs_8.nand3_6.C.t7 a_1761_21414 Vss.t50 nfet_03v3
**devattr s=10400,304 d=10400,304
X344 SARlogic_0.dffrs_3.Qb.t3 SARlogic_0.dffrs_4.d.t5 Vdd.t541 Vdd.t540 pfet_03v3
**devattr s=44000,1176 d=26000,604
X345 a_33257_31423.t0 Clk_piso.t4 a_33521_33720 Vss.t202 nfet_03v3
**devattr s=10400,304 d=17600,576
X346 a_34823_33720 Vdd.t971 Vss.t505 Vss.t504 nfet_03v3
**devattr s=17600,576 d=10400,304
X347 SARlogic_0.d4.t1 SARlogic_0.dffrs_7.Qb Vdd.t265 Vdd.t264 pfet_03v3
**devattr s=26000,604 d=44000,1176
X348 SARlogic_0.dffrs_4.nand3_8.C.t3 SARlogic_0.dffrs_4.nand3_8.Z.t6 Vdd.t485 Vdd.t484 pfet_03v3
**devattr s=26000,604 d=44000,1176
X349 a_14313_29218.t0 a_14393_30170.t5 a_14577_31515 Vss.t206 nfet_03v3
**devattr s=10400,304 d=17600,576
X350 a_275_21414 SARlogic_0.dffrs_8.nand3_1.C Vss.t80 Vss.t79 nfet_03v3
**devattr s=17600,576 d=10400,304
X351 a_9083_31160.t2 inv2_0.out.t13 Vdd.t764 Vdd.t763 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X352 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t10 Vdd.t447 Vdd.t446 pfet_03v3
**devattr s=10400,304 d=10400,304
X353 Vdd.t37 SARlogic_0.dffrs_0.nand3_6.C.t7 SARlogic_0.dffrs_0.Q.t0 Vdd.t36 pfet_03v3
**devattr s=26000,604 d=26000,604
X354 a_40051_37983 adc_PISO_0.serial_out.t6 Vdd.t892 Vdd.t891 pfet_03v3
**devattr s=18700,450 d=34000,880
X355 Vdd.t219 a_23785_29218.t5 adc_PISO_0.dffrs_3.Qb Vdd.t218 pfet_03v3
**devattr s=26000,604 d=26000,604
X356 SARlogic_0.dffrs_10.Qb SARlogic_0.d1.t8 Vdd.t563 Vdd.t562 pfet_03v3
**devattr s=44000,1176 d=26000,604
X357 a_5987_11838 SARlogic_0.dffrs_3.nand3_6.C.t7 a_5803_11838 Vss.t301 nfet_03v3
**devattr s=10400,304 d=10400,304
X358 a_n1095_29019 inv2_0.out.t14 Vss.t559 Vss.t558 nfet_03v3
**devattr s=17600,576 d=17600,576
X359 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vss.t449 Vss.t448 nfet_03v3
**devattr s=9350,280 d=17000,540
X360 a_12585_11838 Reset.t31 a_12401_11838 Vss.t335 nfet_03v3
**devattr s=10400,304 d=10400,304
X361 SARlogic_0.dffrs_4.Q.t3 Vdd.t678 Vdd.t680 Vdd.t679 pfet_03v3
**devattr s=44000,1176 d=26000,604
X362 SARlogic_0.dffrs_4.nand3_6.C.t3 Clk.t10 Vdd.t55 Vdd.t54 pfet_03v3
**devattr s=26000,604 d=44000,1176
X363 a_33257_33628.t0 a_33257_31423.t7 a_33521_35925 Vss.t406 nfet_03v3
**devattr s=10400,304 d=17600,576
X364 a_18743_30440 adc_PISO_0.dffrs_2.Q.t4 Vss.t628 Vss.t627 nfet_03v3
**devattr s=17600,576 d=10400,304
X365 a_275_23619 SARlogic_0.dffrs_1.Qb.t7 Vss.t291 Vss.t290 nfet_03v3
**devattr s=17600,576 d=10400,304
X366 a_n6389_n1044 a_n6589_n1136 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t382 nfet_03v3
**devattr s=15600,404 d=26400,776
X367 a_23785_31423.t0 a_23785_33628.t4 Vdd.t221 Vdd.t220 pfet_03v3
**devattr s=44000,1176 d=26000,604
X368 a_28027_31160.t2 inv2_0.out.t15 Vdd.t766 Vdd.t765 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X369 a_10029_21414 SARlogic_0.dffrs_10.nand3_6.C.t7 a_9845_21414 Vss.t223 nfet_03v3
**devattr s=10400,304 d=10400,304
X370 a_16627_21414 Reset.t32 a_16443_21414 Vss.t303 nfet_03v3
**devattr s=10400,304 d=10400,304
X371 a_n9673_30439 Vss.t95 Vss.t97 Vss.t96 nfet_03v3
**devattr s=17600,576 d=10400,304
X372 Vdd.t349 SARlogic_0.dffrs_14.nand3_8.C.t6 SARlogic_0.dffrs_14.Qb Vdd.t348 pfet_03v3
**devattr s=26000,604 d=26000,604
X373 a_n2097_19210 SARlogic_0.dffrs_7.nand3_8.C.t4 a_n2281_19210 Vss.t126 nfet_03v3
**devattr s=10400,304 d=10400,304
X374 SARlogic_0.dffrs_1.nand3_1.C.t2 SARlogic_0.dffrs_1.nand3_6.C.t5 a_n3583_14043 Vss.t104 nfet_03v3
**devattr s=10400,304 d=17600,576
X375 SARlogic_0.dffrs_12.nand3_8.Z Vss.t93 a_16627_17004 Vss.t94 nfet_03v3
**devattr s=10400,304 d=17600,576
X376 a_23785_33628.t2 Vdd.t675 Vdd.t677 Vdd.t676 pfet_03v3
**devattr s=44000,1176 d=26000,604
X377 a_1839_29263.t1 a_1167_28099 Vss.t219 Vss.t218 nfet_03v3
**devattr s=17600,576 d=17600,576
X378 adc_PISO_0.2inmux_4.OUT.t0 a_20783_29264.t4 Vss.t438 Vss.t437 nfet_03v3
**devattr s=17600,576 d=17600,576
X379 a_16627_23619 SARlogic_0.dffrs_12.nand3_8.Z a_16443_23619 Vss.t8 nfet_03v3
**devattr s=10400,304 d=10400,304
X380 SARlogic_0.dffrs_7.Qb Reset.t33 a_n2097_19210 Vss.t304 nfet_03v3
**devattr s=10400,304 d=17600,576
X381 SARlogic_0.dffrs_9.nand3_8.C.t0 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t157 Vdd.t156 pfet_03v3
**devattr s=26000,604 d=44000,1176
X382 SARlogic_0.dffrs_11.nand3_8.C.t0 SARlogic_0.dffrs_11.nand3_6.C.t5 Vdd.t77 Vdd.t76 pfet_03v3
**devattr s=44000,1176 d=26000,604
X383 Vdd.t389 Reset.t34 SARlogic_0.dffrs_4.nand3_8.Z.t0 Vdd.t388 pfet_03v3
**devattr s=26000,604 d=26000,604
X384 a_34823_31516 adc_PISO_0.2inmux_1.Bit.t7 Vss.t343 Vss.t342 nfet_03v3
**devattr s=17600,576 d=10400,304
X385 a_9271_28100 a_8377_29020 Vss.t107 Vss.t106 nfet_03v3
**devattr s=17600,576 d=10400,304
X386 SARlogic_0.dffrs_12.nand3_8.C.t0 SARlogic_0.dffrs_12.nand3_8.Z a_16627_19209 Vss.t7 nfet_03v3
**devattr s=10400,304 d=17600,576
X387 Vdd.t117 SARlogic_0.dffrs_0.nand3_8.Z.t5 SARlogic_0.dffrs_0.nand3_1.C.t0 Vdd.t116 pfet_03v3
**devattr s=26000,604 d=26000,604
X388 a_10639_30440 a_9083_31160.t5 Vdd.t806 Vdd.t805 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X389 a_27321_29020 inv2_0.out.t16 Vss.t561 Vss.t560 nfet_03v3
**devattr s=17600,576 d=17600,576
X390 SARlogic_0.dffrs_4.nand3_8.C.t1 SARlogic_0.dffrs_4.nand3_6.C.t4 Vdd.t109 Vdd.t108 pfet_03v3
**devattr s=44000,1176 d=26000,604
X391 a_n11637_14043 SARlogic_0.dffrs_13.nand3_8.Z.t4 a_n11821_14043 Vss.t71 nfet_03v3
**devattr s=10400,304 d=10400,304
X392 a_n7625_17007 Reset.t35 a_n7809_17007 Vss.t305 nfet_03v3
**devattr s=10400,304 d=10400,304
X393 a_33337_33720 a_33257_33628.t5 Vss.t591 Vss.t590 nfet_03v3
**devattr s=17600,576 d=10400,304
X394 a_n9861_28819.t2 SARlogic_0.d5.t5 a_n9673_28099 Vss.t228 nfet_03v3
**devattr s=10400,304 d=17600,576
X395 a_33521_29310 Vdd.t972 a_33337_29310 Vss.t503 nfet_03v3
**devattr s=10400,304 d=10400,304
X396 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t0 Clk.t11 Vdd.t57 Vdd.t56 pfet_03v3
**devattr s=14080,496 d=14080,496
X397 a_4921_30169.t0 adc_PISO_0.2inmux_2.OUT.t3 Vdd.t215 Vdd.t214 pfet_03v3
**devattr s=26000,604 d=44000,1176
X398 SARlogic_0.dffrs_4.nand3_6.C.t1 SARlogic_0.dffrs_4.nand3_1.C.t4 Vdd.t487 Vdd.t486 pfet_03v3
**devattr s=44000,1176 d=26000,604
X399 a_33337_35925 Vdd.t973 Vss.t502 Vss.t501 nfet_03v3
**devattr s=17600,576 d=10400,304
X400 a_24049_31515 Clk_piso.t5 a_23865_31515 Vss.t203 nfet_03v3
**devattr s=10400,304 d=10400,304
X401 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t15 Clk.t12 Vdd.t59 Vdd.t58 pfet_03v3
**devattr s=14080,496 d=14080,496
X402 a_n9861_28819.t3 SARlogic_0.d5.t6 Vdd.t301 Vdd.t300 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X403 a_37687_28100 a_36793_29020 Vss.t197 Vss.t196 nfet_03v3
**devattr s=17600,576 d=10400,304
X404 SARlogic_0.dffrs_10.Qb Reset.t36 Vdd.t391 Vdd.t390 pfet_03v3
**devattr s=26000,604 d=44000,1176
X405 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t14 Vss.t336 nfet_03v3
**devattr s=20800,504 d=20800,504
X406 a_12585_9633 Clk.t13 a_12401_9633 Vss.t27 nfet_03v3
**devattr s=10400,304 d=10400,304
X407 SARlogic_0.dffrs_4.Q.t2 SARlogic_0.dffrs_4.Qb.t5 Vdd.t942 Vdd.t941 pfet_03v3
**devattr s=26000,604 d=44000,1176
X408 Vdd.t393 Reset.t37 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t392 pfet_03v3
**devattr s=26000,604 d=26000,604
X409 SARlogic_0.dffrs_2.nand3_8.C.t0 SARlogic_0.dffrs_2.nand3_8.Z.t5 Vdd.t269 Vdd.t268 pfet_03v3
**devattr s=26000,604 d=44000,1176
X410 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t4 a_8543_17004 Vss.t193 nfet_03v3
**devattr s=10400,304 d=17600,576
X411 a_16443_17004 SARlogic_0.dffrs_12.nand3_8.C.t7 Vss.t679 Vss.t678 nfet_03v3
**devattr s=17600,576 d=10400,304
X412 a_1945_9634 SARlogic_0.dffrs_2.nand3_8.C.t5 a_1761_9634 Vss.t660 nfet_03v3
**devattr s=10400,304 d=10400,304
X413 SARlogic_0.d0.t2 SARlogic_0.dffrs_11.Qb Vdd.t245 Vdd.t244 pfet_03v3
**devattr s=26000,604 d=44000,1176
X414 a_13887_9634 SARlogic_0.dffrs_5.Q.t4 Vss.t355 Vss.t354 nfet_03v3
**devattr s=17600,576 d=10400,304
X415 SARlogic_0.dffrs_7.nand3_6.C.t3 SARlogic_0.dffrs_7.nand3_1.C Vdd.t455 Vdd.t454 pfet_03v3
**devattr s=44000,1176 d=26000,604
X416 SARlogic_0.dffrs_0.nand3_8.Z.t2 SARlogic_0.dffrs_0.d.t7 a_n7625_7428 Vss.t597 nfet_03v3
**devattr s=10400,304 d=17600,576
X417 SARlogic_0.dffrs_9.nand3_8.C.t3 SARlogic_0.dffrs_9.nand3_6.C.t6 Vdd.t904 Vdd.t903 pfet_03v3
**devattr s=44000,1176 d=26000,604
X418 SARlogic_0.dffrs_2.nand3_6.C.t0 Clk.t14 Vdd.t61 Vdd.t60 pfet_03v3
**devattr s=26000,604 d=44000,1176
X419 a_16443_19209 SARlogic_0.dffrs_12.nand3_6.C.t7 Vss.t269 Vss.t268 nfet_03v3
**devattr s=17600,576 d=10400,304
X420 SARlogic_0.dffrs_10.nand3_8.C.t0 SARlogic_0.dffrs_10.nand3_8.Z a_8543_19209 Vss.t275 nfet_03v3
**devattr s=10400,304 d=17600,576
X421 Vdd.t79 SARlogic_0.dffrs_11.nand3_6.C.t6 SARlogic_0.d0.t0 Vdd.t78 pfet_03v3
**devattr s=26000,604 d=26000,604
X422 a_n9429_n2007.t9 Vin1.t2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t7 Vss.t262 nfet_03v3
**devattr s=15600,404 d=15600,404
X423 SARlogic_0.dffrs_12.Qb Reset.t38 Vdd.t395 Vdd.t394 pfet_03v3
**devattr s=26000,604 d=44000,1176
X424 a_459_9633 Clk.t15 a_275_9633 Vss.t28 nfet_03v3
**devattr s=10400,304 d=10400,304
X425 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_0.Qb.t6 Vdd.t233 Vdd.t232 pfet_03v3
**devattr s=44000,1176 d=26000,604
X426 SARlogic_0.dffrs_13.nand3_8.Z.t0 SARlogic_0.dffrs_13.nand3_8.C.t5 Vdd.t31 Vdd.t30 pfet_03v3
**devattr s=44000,1176 d=26000,604
X427 SARlogic_0.dffrs_4.nand3_1.C.t3 SARlogic_0.dffrs_4.nand3_6.C.t5 Vdd.t111 Vdd.t110 pfet_03v3
**devattr s=26000,604 d=44000,1176
X428 a_14313_31423.t3 Clk_piso.t6 Vdd.t273 Vdd.t272 pfet_03v3
**devattr s=26000,604 d=44000,1176
X429 Vss.t338 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t12 comparator_no_offsetcal_0.x5.out Vss.t337 nfet_03v3
**devattr s=35200,976 d=35200,976
X430 adc_PISO_0.dffrs_3.Q.t2 adc_PISO_0.dffrs_3.Qb Vdd.t337 Vdd.t336 pfet_03v3
**devattr s=26000,604 d=44000,1176
X431 SARlogic_0.d2.t1 SARlogic_0.dffrs_9.Qb a_5987_21414 Vss.t594 nfet_03v3
**devattr s=10400,304 d=17600,576
X432 a_8377_29020 inv2_0.out.t17 Vdd.t768 Vdd.t767 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X433 a_n2281_21414 SARlogic_0.dffrs_0.Qb.t7 Vss.t162 Vss.t161 nfet_03v3
**devattr s=17600,576 d=10400,304
X434 Comp_out.t2 a_n10831_4320 Vss.t541 Vss.t540 nfet_03v3
**devattr s=9350,280 d=9350,280
X435 Comp_out.t6 a_n10831_4320 Vdd.t752 Vdd.t751 pfet_03v3
**devattr s=34000,880 d=18700,450
X436 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t7 a_n7625_23622 Vss.t294 nfet_03v3
**devattr s=10400,304 d=17600,576
X437 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t6 Vin1.t3 a_n9429_n2007.t10 Vss.t212 nfet_03v3
**devattr s=15600,404 d=15600,404
X438 a_14313_33628.t2 a_14313_31423.t4 Vdd.t856 Vdd.t855 pfet_03v3
**devattr s=26000,604 d=44000,1176
X439 a_42809_29310 a_42729_29218.t4 Vss.t600 Vss.t599 nfet_03v3
**devattr s=17600,576 d=10400,304
X440 SARlogic_0.dffrs_8.Qb Reset.t39 Vdd.t397 Vdd.t396 pfet_03v3
**devattr s=26000,604 d=44000,1176
X441 SARlogic_0.dffrs_5.nand3_8.Z.t1 SARlogic_0.dffrs_4.Q.t5 a_12585_7428 Vss.t156 nfet_03v3
**devattr s=10400,304 d=17600,576
X442 SARlogic_0.dffrs_5.Qb.t0 Reset.t40 a_14071_9634 Vss.t306 nfet_03v3
**devattr s=10400,304 d=17600,576
X443 SARlogic_0.dffrs_2.Q.t2 SARlogic_0.dffrs_2.Qb.t4 Vdd.t840 Vdd.t839 pfet_03v3
**devattr s=26000,604 d=44000,1176
X444 SARlogic_0.dffrs_11.Qb Reset.t41 a_14071_19210 Vss.t307 nfet_03v3
**devattr s=10400,304 d=17600,576
X445 a_39915_29984 a_39055_28100 a_39727_29264.t1 Vdd.t280 pfet_03v3
**devattr s=52800,1376 d=31200,704
X446 a_n6323_11838 Vdd.t974 Vss.t500 Vss.t499 nfet_03v3
**devattr s=17600,576 d=10400,304
X447 SARlogic_0.dffrs_0.nand3_6.C.t3 Clk.t16 a_n7625_11838 Vss.t29 nfet_03v3
**devattr s=10400,304 d=17600,576
X448 a_29583_28100 a_28027_28820.t4 Vss.t578 Vss.t577 nfet_03v3
**devattr s=17600,576 d=17600,576
X449 Vdd.t189 SARlogic_0.dffrs_8.nand3_8.C.t6 SARlogic_0.dffrs_8.Qb Vdd.t188 pfet_03v3
**devattr s=26000,604 d=26000,604
X450 SARlogic_0.dffrs_2.nand3_8.C.t2 SARlogic_0.dffrs_2.nand3_6.C.t6 Vdd.t495 Vdd.t494 pfet_03v3
**devattr s=44000,1176 d=26000,604
X451 a_8359_17004 SARlogic_0.dffrs_10.nand3_8.C.t6 Vss.t246 Vss.t245 nfet_03v3
**devattr s=17600,576 d=10400,304
X452 Vdd.t73 adc_PISO_0.2inmux_2.Bit.t6 a_n389_31159.t0 Vdd.t72 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X453 Vdd.t497 SARlogic_0.dffrs_2.nand3_6.C.t7 SARlogic_0.dffrs_2.Q.t0 Vdd.t496 pfet_03v3
**devattr s=26000,604 d=26000,604
X454 a_14071_19210 SARlogic_0.dffrs_11.nand3_8.C.t5 a_13887_19210 Vss.t185 nfet_03v3
**devattr s=10400,304 d=10400,304
X455 a_23785_31423.t1 Clk_piso.t7 a_24049_33720 Vss.t204 nfet_03v3
**devattr s=10400,304 d=17600,576
X456 a_25351_33720 Vdd.t975 Vss.t498 Vss.t497 nfet_03v3
**devattr s=17600,576 d=10400,304
X457 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t13 Vdd.t571 Vdd.t570 pfet_03v3
**devattr s=10400,304 d=10400,304
X458 SARlogic_0.dffrs_7.nand3_6.C.t1 SARlogic_0.d3.t8 Vdd.t99 Vdd.t98 pfet_03v3
**devattr s=26000,604 d=44000,1176
X459 Vdd.t399 Reset.t42 SARlogic_0.dffrs_3.nand3_8.Z.t0 Vdd.t398 pfet_03v3
**devattr s=26000,604 d=26000,604
X460 SARlogic_0.dffrs_2.nand3_6.C.t2 SARlogic_0.dffrs_2.nand3_1.C.t4 Vdd.t71 Vdd.t70 pfet_03v3
**devattr s=44000,1176 d=26000,604
X461 a_8359_19209 SARlogic_0.dffrs_10.nand3_6.C.t8 Vss.t225 Vss.t224 nfet_03v3
**devattr s=17600,576 d=10400,304
X462 a_35007_33720 a_33257_31423.t8 a_34823_33720 Vss.t407 nfet_03v3
**devattr s=10400,304 d=10400,304
X463 Vdd.t247 adc_PISO_0.dffrs_3.Q.t6 a_28027_31160.t3 Vdd.t246 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X464 a_n2097_9634 SARlogic_0.dffrs_1.nand3_8.C.t5 a_n2281_9634 Vss.t408 nfet_03v3
**devattr s=10400,304 d=10400,304
X465 Vdd.t523 SARlogic_0.dffrs_3.nand3_8.C.t7 SARlogic_0.dffrs_3.Qb.t0 Vdd.t522 pfet_03v3
**devattr s=26000,604 d=26000,604
X466 a_23785_33628.t1 a_23785_31423.t8 a_24049_35925 Vss.t171 nfet_03v3
**devattr s=10400,304 d=17600,576
X467 a_n9861_31159.t1 inv2_0.out.t18 a_n9673_30439 Vss.t562 nfet_03v3
**devattr s=10400,304 d=17600,576
X468 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t6 Vdd.t303 Vdd.t302 pfet_03v3
**devattr s=26000,604 d=44000,1176
X469 a_459_21414 Reset.t43 a_275_21414 Vss.t308 nfet_03v3
**devattr s=10400,304 d=10400,304
X470 a_n7809_19212 SARlogic_0.dffrs_14.nand3_6.C.t8 Vss.t296 Vss.t295 nfet_03v3
**devattr s=17600,576 d=10400,304
X471 Vss.t138 a_27321_29020 a_28215_28100 Vss.t137 nfet_03v3
**devattr s=10400,304 d=17600,576
X472 SARlogic_0.dffrs_2.nand3_8.Z.t1 SARlogic_0.dffrs_2.d.t5 a_459_7428 Vss.t17 nfet_03v3
**devattr s=10400,304 d=17600,576
X473 SARlogic_0.dffrs_4.nand3_1.C.t0 Vdd.t672 Vdd.t674 Vdd.t673 pfet_03v3
**devattr s=44000,1176 d=26000,604
X474 adc_PISO_0.dffrs_3.Qb Vdd.t669 Vdd.t671 Vdd.t670 pfet_03v3
**devattr s=26000,604 d=44000,1176
X475 Vdd.t321 SARlogic_0.dffrs_10.nand3_8.C.t7 SARlogic_0.dffrs_10.Qb Vdd.t320 pfet_03v3
**devattr s=26000,604 d=26000,604
X476 a_13887_11838 Vdd.t976 Vss.t496 Vss.t495 nfet_03v3
**devattr s=17600,576 d=10400,304
X477 a_28215_30440 inv2_0.out.t19 a_28027_31160.t0 Vss.t563 nfet_03v3
**devattr s=17600,576 d=10400,304
X478 Vdd.t113 SARlogic_0.dffrs_4.nand3_6.C.t6 SARlogic_0.dffrs_4.Q.t0 Vdd.t112 pfet_03v3
**devattr s=26000,604 d=26000,604
X479 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t5 a_459_17004 Vss.t277 nfet_03v3
**devattr s=10400,304 d=17600,576
X480 SARlogic_0.dffrs_4.nand3_8.Z.t3 SARlogic_0.dffrs_4.d.t6 Vdd.t539 Vdd.t538 pfet_03v3
**devattr s=26000,604 d=44000,1176
X481 a_459_23619 SARlogic_0.dffrs_8.nand3_8.Z a_275_23619 Vss.t250 nfet_03v3
**devattr s=10400,304 d=10400,304
X482 Vdd.t668 Vdd.t666 a_23785_31423.t2 Vdd.t667 pfet_03v3
**devattr s=26000,604 d=26000,604
X483 a_17929_21414 SARlogic_0.dffrs_5.Qb.t7 Vss.t618 Vss.t617 nfet_03v3
**devattr s=17600,576 d=10400,304
X484 adc_PISO_0.2inmux_1.OUT.t0 a_39727_29264.t4 Vss.t610 Vss.t609 nfet_03v3
**devattr s=17600,576 d=17600,576
X485 SARlogic_0.dffrs_8.nand3_8.C.t1 SARlogic_0.dffrs_8.nand3_8.Z a_459_19209 Vss.t249 nfet_03v3
**devattr s=10400,304 d=17600,576
X486 SARlogic_0.dffrs_1.nand3_8.Z.t1 SARlogic_0.dffrs_0.Q.t5 a_n3583_7428 Vss.t564 nfet_03v3
**devattr s=10400,304 d=17600,576
X487 a_25351_31516 adc_PISO_0.dffrs_3.Q.t7 Vss.t178 Vss.t177 nfet_03v3
**devattr s=17600,576 d=10400,304
X488 SARlogic_0.dffrs_0.Q.t2 SARlogic_0.dffrs_0.Qb.t8 a_n6139_11838 Vss.t622 nfet_03v3
**devattr s=10400,304 d=17600,576
X489 a_n4631_29217.t0 a_n4631_31422.t5 Vdd.t932 Vdd.t931 pfet_03v3
**devattr s=44000,1176 d=26000,604
X490 a_n6323_9634 SARlogic_0.dffrs_0.Q.t6 Vss.t133 Vss.t132 nfet_03v3
**devattr s=17600,576 d=10400,304
X491 Vdd.t836 a_23865_30170.t5 a_23785_33628.t3 Vdd.t835 pfet_03v3
**devattr s=26000,604 d=26000,604
X492 a_8543_11838 Reset.t44 a_8359_11838 Vss.t309 nfet_03v3
**devattr s=10400,304 d=10400,304
X493 SARlogic_0.dffrs_5.nand3_1.C.t0 SARlogic_0.dffrs_5.nand3_6.C.t6 a_12585_14043 Vss.t534 nfet_03v3
**devattr s=10400,304 d=17600,576
X494 SARlogic_0.dffrs_2.nand3_1.C.t2 SARlogic_0.dffrs_2.nand3_6.C.t8 Vdd.t499 Vdd.t498 pfet_03v3
**devattr s=26000,604 d=44000,1176
X495 a_14393_30170.t2 a_14313_29218.t5 Vdd.t333 Vdd.t332 pfet_03v3
**devattr s=44000,1176 d=26000,604
X496 Vdd.t555 SARlogic_0.dffrs_12.Q.t6 SARlogic_0.dffrs_11.nand3_8.C.t3 Vdd.t554 pfet_03v3
**devattr s=26000,604 d=26000,604
X497 a_35007_31516 a_33257_29218.t5 a_34823_31516 Vss.t581 nfet_03v3
**devattr s=10400,304 d=10400,304
X498 a_n4631_31422.t1 a_n4631_33627.t4 Vdd.t583 Vdd.t582 pfet_03v3
**devattr s=44000,1176 d=26000,604
X499 a_42729_29218.t0 a_42809_30170.t6 a_42993_31515 Vss.t644 nfet_03v3
**devattr s=10400,304 d=17600,576
X500 a_14313_29218.t2 a_14313_31423.t5 Vdd.t858 Vdd.t857 pfet_03v3
**devattr s=44000,1176 d=26000,604
X501 a_14577_31515 Clk_piso.t8 a_14393_31515 Vss.t205 nfet_03v3
**devattr s=10400,304 d=10400,304
X502 a_n10567_29019 inv2_0.out.t20 Vdd.t770 Vdd.t769 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X503 a_33337_30170.t0 adc_PISO_0.2inmux_5.OUT.t2 a_33521_29310 Vss.t264 nfet_03v3
**devattr s=10400,304 d=17600,576
X504 a_4501_14043 SARlogic_0.dffrs_3.nand3_8.Z.t6 a_4317_14043 Vss.t412 nfet_03v3
**devattr s=10400,304 d=10400,304
X505 a_275_17004 SARlogic_0.dffrs_8.nand3_8.C.t7 Vss.t129 Vss.t128 nfet_03v3
**devattr s=17600,576 d=10400,304
X506 a_n7625_7428 Reset.t45 a_n7809_7428 Vss.t310 nfet_03v3
**devattr s=10400,304 d=10400,304
X507 Piso_out.t5 a_40051_37983 Vdd.t545 Vdd.t544 pfet_03v3
**devattr s=34000,880 d=18700,450
X508 a_275_19209 SARlogic_0.dffrs_8.nand3_6.C.t8 Vss.t52 Vss.t51 nfet_03v3
**devattr s=17600,576 d=10400,304
X509 Vdd.t449 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t4 Vdd.t448 pfet_03v3
**devattr s=10400,304 d=10400,304
X510 SARlogic_0.dffrs_4.Qb.t1 Reset.t46 a_10029_9634 Vss.t311 nfet_03v3
**devattr s=10400,304 d=17600,576
X511 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_8.C.t5 Vdd.t185 Vdd.t184 pfet_03v3
**devattr s=44000,1176 d=26000,604
X512 a_16627_17004 Reset.t47 a_16443_17004 Vss.t312 nfet_03v3
**devattr s=10400,304 d=10400,304
X513 a_n4631_29217.t1 a_n4551_30169.t5 Vdd.t293 Vdd.t292 pfet_03v3
**devattr s=26000,604 d=44000,1176
X514 Vdd.t137 a_n8305_30439 a_n7445_29983 Vdd.t136 pfet_03v3
**devattr s=31200,704 d=52800,1376
X515 SARlogic_0.dffrs_2.nand3_1.C.t3 Vdd.t663 Vdd.t665 Vdd.t664 pfet_03v3
**devattr s=44000,1176 d=26000,604
X516 SARlogic_0.dffrs_13.nand3_8.C.t1 SARlogic_0.dffrs_13.nand3_8.Z.t5 a_n11637_9633 Vss.t72 nfet_03v3
**devattr s=10400,304 d=17600,576
X517 a_16627_19209 Vss.t91 a_16443_19209 Vss.t92 nfet_03v3
**devattr s=10400,304 d=10400,304
X518 a_n4631_31422.t0 Clk_piso.t9 Vdd.t275 Vdd.t274 pfet_03v3
**devattr s=26000,604 d=44000,1176
X519 adc_PISO_0.2inmux_2.Bit.t3 Vdd.t660 Vdd.t662 Vdd.t661 pfet_03v3
**devattr s=44000,1176 d=26000,604
X520 adc_PISO_0.dffrs_2.Q.t1 adc_PISO_0.dffrs_2.Qb Vdd.t481 Vdd.t480 pfet_03v3
**devattr s=26000,604 d=44000,1176
X521 SARlogic_0.dffrs_9.Qb Reset.t48 Vdd.t401 Vdd.t400 pfet_03v3
**devattr s=26000,604 d=44000,1176
X522 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t14 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t436 nfet_03v3
**devattr s=20800,504 d=20800,504
X523 SARlogic_0.dffrs_7.Qb SARlogic_0.d4.t7 Vdd.t890 Vdd.t889 pfet_03v3
**devattr s=44000,1176 d=26000,604
X524 SARlogic_0.dffrs_4.d.t0 SARlogic_0.dffrs_3.Qb.t8 Vdd.t181 Vdd.t180 pfet_03v3
**devattr s=26000,604 d=44000,1176
X525 adc_PISO_0.serial_out.t1 adc_PISO_0.dffrs_5.Qb Vdd.t513 Vdd.t512 pfet_03v3
**devattr s=26000,604 d=44000,1176
X526 SARlogic_0.dffrs_2.d.t0 Vdd.t657 Vdd.t659 Vdd.t658 pfet_03v3
**devattr s=44000,1176 d=26000,604
X527 Vdd.t934 a_n4631_31422.t6 adc_PISO_0.2inmux_2.Bit.t2 Vdd.t933 pfet_03v3
**devattr s=26000,604 d=26000,604
X528 Vdd.t860 a_14313_31423.t6 adc_PISO_0.dffrs_2.Q.t3 Vdd.t859 pfet_03v3
**devattr s=26000,604 d=26000,604
X529 a_33337_29310 a_33257_29218.t6 Vss.t583 Vss.t582 nfet_03v3
**devattr s=17600,576 d=10400,304
X530 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vdd.t597 Vdd.t596 pfet_03v3
**devattr s=18700,450 d=34000,880
X531 a_n3583_21414 Reset.t49 a_n3767_21414 Vss.t313 nfet_03v3
**devattr s=10400,304 d=10400,304
X532 SARlogic_0.dffrs_3.nand3_8.Z.t2 SARlogic_0.dffrs_2.Q.t5 Vdd.t479 Vdd.t478 pfet_03v3
**devattr s=26000,604 d=44000,1176
X533 SARlogic_0.dffrs_0.Qb.t1 SARlogic_0.dffrs_0.Q.t7 Vdd.t195 Vdd.t194 pfet_03v3
**devattr s=44000,1176 d=26000,604
X534 a_n7625_23622 SARlogic_0.dffrs_14.nand3_8.Z a_n7809_23622 Vss.t10 nfet_03v3
**devattr s=10400,304 d=10400,304
X535 a_n3583_23619 SARlogic_0.dffrs_7.nand3_8.Z a_n3767_23619 Vss.t208 nfet_03v3
**devattr s=10400,304 d=10400,304
X536 a_20971_29984 a_20111_30440 Vdd.t119 Vdd.t118 pfet_03v3
**devattr s=52800,1376 d=31200,704
X537 Vdd.t63 Clk.t17 SARlogic_0.dffrs_2.nand3_8.C.t3 Vdd.t62 pfet_03v3
**devattr s=26000,604 d=26000,604
X538 a_n7625_11838 Reset.t50 a_n7809_11838 Vss.t314 nfet_03v3
**devattr s=10400,304 d=10400,304
X539 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t6 Vdd.t357 Vdd.t356 pfet_03v3
**devattr s=26000,604 d=44000,1176
X540 a_25535_33720 a_23785_31423.t9 a_25351_33720 Vss.t172 nfet_03v3
**devattr s=10400,304 d=10400,304
X541 Vss.t646 a_39055_30440 a_39727_29264.t3 Vss.t645 nfet_03v3
**devattr s=17600,576 d=17600,576
X542 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t16 a_n9767_249 a_n9855_341 Vss.t685 nfet_03v3
**devattr s=35200,976 d=20800,504
X543 Vdd.t403 Reset.t51 SARlogic_0.dffrs_2.nand3_6.C.t3 Vdd.t402 pfet_03v3
**devattr s=26000,604 d=26000,604
X544 adc_PISO_0.dffrs_2.Qb Vdd.t654 Vdd.t656 Vdd.t655 pfet_03v3
**devattr s=26000,604 d=44000,1176
X545 adc_PISO_0.dffrs_5.Qb Vdd.t651 Vdd.t653 Vdd.t652 pfet_03v3
**devattr s=26000,604 d=44000,1176
X546 a_20111_28100 a_18555_28820.t5 Vdd.t205 Vdd.t204 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X547 SARlogic_0.dffrs_11.nand3_6.C.t2 SARlogic_0.dffrs_12.Q.t7 Vdd.t557 Vdd.t556 pfet_03v3
**devattr s=26000,604 d=44000,1176
X548 SARlogic_0.dffrs_5.Qb.t2 SARlogic_0.dffrs_5.Q.t5 Vdd.t465 Vdd.t464 pfet_03v3
**devattr s=44000,1176 d=26000,604
X549 Vdd.t473 a_4841_31422.t6 adc_PISO_0.dffrs_1.Q.t2 Vdd.t472 pfet_03v3
**devattr s=26000,604 d=26000,604
X550 adc_PISO_0.dffrs_1.Q.t0 adc_PISO_0.dffrs_1.Qb a_6591_33719 Vss.t113 nfet_03v3
**devattr s=10400,304 d=17600,576
X551 Vdd.t335 a_14313_29218.t6 adc_PISO_0.dffrs_2.Qb Vdd.t334 pfet_03v3
**devattr s=26000,604 d=26000,604
X552 a_37499_28820.t3 SARlogic_0.d0.t9 Vdd.t948 Vdd.t947 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X553 a_42729_31423.t2 Clk_piso.t10 Vdd.t862 Vdd.t861 pfet_03v3
**devattr s=26000,604 d=44000,1176
X554 a_8359_9633 SARlogic_0.dffrs_4.nand3_6.C.t7 Vss.t64 Vss.t63 nfet_03v3
**devattr s=17600,576 d=10400,304
X555 Vdd.t650 Vdd.t648 a_14313_31423.t1 Vdd.t649 pfet_03v3
**devattr s=26000,604 d=26000,604
X556 SARlogic_0.dffrs_12.Qb SARlogic_0.dffrs_12.Q.t8 Vdd.t559 Vdd.t558 pfet_03v3
**devattr s=44000,1176 d=26000,604
X557 a_1761_11838 Vdd.t977 Vss.t494 Vss.t493 nfet_03v3
**devattr s=17600,576 d=10400,304
X558 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t7 Vdd.t81 Vdd.t80 pfet_03v3
**devattr s=26000,604 d=44000,1176
X559 a_n6389_n2007 a_n6589_n2099 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t11 Vss.t382 nfet_03v3
**devattr s=15600,404 d=26400,776
X560 a_18555_31160.t2 inv2_0.out.t21 Vdd.t772 Vdd.t771 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X561 adc_PISO_0.2inmux_2.OUT.t0 a_1839_29263.t4 Vss.t168 Vss.t167 nfet_03v3
**devattr s=17600,576 d=17600,576
X562 a_n2097_21414 SARlogic_0.dffrs_7.nand3_6.C.t7 a_n2281_21414 Vss.t232 nfet_03v3
**devattr s=10400,304 d=10400,304
X563 SARlogic_0.dffrs_0.Qb.t2 Reset.t52 Vdd.t405 Vdd.t404 pfet_03v3
**devattr s=26000,604 d=44000,1176
X564 a_42729_33628.t0 a_42729_31423.t4 Vdd.t175 Vdd.t174 pfet_03v3
**devattr s=26000,604 d=44000,1176
X565 Vdd.t407 Reset.t53 SARlogic_0.dffrs_9.nand3_6.C.t0 Vdd.t406 pfet_03v3
**devattr s=26000,604 d=26000,604
X566 Vdd.t910 a_14393_30170.t6 a_14313_33628.t3 Vdd.t909 pfet_03v3
**devattr s=26000,604 d=26000,604
X567 SARlogic_0.d4.t0 SARlogic_0.dffrs_7.Qb a_n2097_21414 Vss.t198 nfet_03v3
**devattr s=10400,304 d=17600,576
X568 Vdd.t854 SARlogic_0.dffrs_13.nand3_6.C.t5 SARlogic_0.dffrs_0.d.t3 Vdd.t853 pfet_03v3
**devattr s=26000,604 d=26000,604
X569 SARlogic_0.dffrs_14.nand3_8.C.t0 SARlogic_0.dffrs_14.nand3_8.Z a_n7625_19212 Vss.t9 nfet_03v3
**devattr s=10400,304 d=17600,576
X570 a_25535_31516 a_23785_29218.t6 a_25351_31516 Vss.t149 nfet_03v3
**devattr s=10400,304 d=10400,304
X571 adc_PISO_0.2inmux_3.OUT.t1 a_11311_29264.t4 Vss.t160 Vss.t159 nfet_03v3
**devattr s=17600,576 d=17600,576
X572 a_n8351_341 a_n8551_249 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t6 Vss.t356 nfet_03v3
**devattr s=20800,504 d=35200,976
X573 a_n6139_11838 SARlogic_0.dffrs_0.nand3_6.C.t8 a_n6323_11838 Vss.t16 nfet_03v3
**devattr s=10400,304 d=10400,304
X574 Vdd.t155 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_1.C Vdd.t154 pfet_03v3
**devattr s=26000,604 d=26000,604
X575 SARlogic_0.dffrs_4.nand3_6.C.t2 Clk.t18 a_8543_11838 Vss.t30 nfet_03v3
**devattr s=10400,304 d=17600,576
X576 a_9845_11838 Vdd.t978 Vss.t492 Vss.t491 nfet_03v3
**devattr s=17600,576 d=10400,304
X577 a_18743_28100 SARlogic_0.d2.t8 a_18555_28820.t2 Vss.t237 nfet_03v3
**devattr s=17600,576 d=10400,304
X578 Vdd.t409 Reset.t54 SARlogic_0.dffrs_1.nand3_8.Z.t0 Vdd.t408 pfet_03v3
**devattr s=26000,604 d=26000,604
X579 Vdd.t864 Clk_piso.t11 a_4841_29217.t3 Vdd.t863 pfet_03v3
**devattr s=26000,604 d=26000,604
X580 Vdd.t647 Vdd.t645 a_42809_30170.t1 Vdd.t646 pfet_03v3
**devattr s=26000,604 d=26000,604
X581 a_39055_28100 a_37499_28820.t5 Vdd.t503 Vdd.t502 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X582 a_23865_30170.t0 adc_PISO_0.2inmux_4.OUT.t2 a_24049_29310 Vss.t70 nfet_03v3
**devattr s=10400,304 d=17600,576
X583 Vdd.t133 a_1167_30439 a_2027_29983 Vdd.t132 pfet_03v3
**devattr s=31200,704 d=52800,1376
X584 a_23865_33720 a_23785_33628.t5 Vss.t153 Vss.t152 nfet_03v3
**devattr s=17600,576 d=10400,304
X585 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 Vdd.t573 Vdd.t572 pfet_03v3
**devattr s=10400,304 d=10400,304
X586 a_n7445_29983 a_n8305_28099 a_n7633_29263.t2 Vdd.t322 pfet_03v3
**devattr s=52800,1376 d=31200,704
X587 a_4841_29217.t2 a_4841_31422.t7 Vdd.t475 Vdd.t474 pfet_03v3
**devattr s=44000,1176 d=26000,604
X588 a_n9429_n2007.t1 Vin2.t4 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t209 nfet_03v3
**devattr s=15600,404 d=15600,404
X589 Vdd.t644 Vdd.t642 a_4841_31422.t2 Vdd.t643 pfet_03v3
**devattr s=26000,604 d=26000,604
X590 Vdd.t866 Clk_piso.t12 a_42729_29218.t3 Vdd.t865 pfet_03v3
**devattr s=26000,604 d=26000,604
X591 a_459_17004 Reset.t55 a_275_17004 Vss.t315 nfet_03v3
**devattr s=10400,304 d=10400,304
X592 SARlogic_0.dffrs_3.nand3_1.C.t1 SARlogic_0.dffrs_3.nand3_6.C.t8 a_4501_14043 Vss.t302 nfet_03v3
**devattr s=10400,304 d=17600,576
X593 a_12401_14043 Vdd.t980 Vss.t488 Vss.t487 nfet_03v3
**devattr s=17600,576 d=10400,304
X594 Vdd.t888 a_10639_30440 a_11499_29984 Vdd.t887 pfet_03v3
**devattr s=31200,704 d=52800,1376
X595 a_23865_35925 Vdd.t979 Vss.t490 Vss.t489 nfet_03v3
**devattr s=17600,576 d=10400,304
X596 Comp_out.t5 a_n10831_4320 Vdd.t750 Vdd.t749 pfet_03v3
**devattr s=18700,450 d=18700,450
X597 a_8543_7428 Reset.t56 a_8359_7428 Vss.t316 nfet_03v3
**devattr s=10400,304 d=10400,304
X598 a_4841_31422.t1 a_4841_33627.t4 Vdd.t505 Vdd.t504 pfet_03v3
**devattr s=44000,1176 d=26000,604
X599 SARlogic_0.dffrs_0.nand3_8.Z.t0 SARlogic_0.dffrs_0.nand3_8.C.t5 Vdd.t105 Vdd.t104 pfet_03v3
**devattr s=44000,1176 d=26000,604
X600 Vdd.t950 SARlogic_0.d0.t10 SARlogic_0.dffrs_10.nand3_8.C.t3 Vdd.t949 pfet_03v3
**devattr s=26000,604 d=26000,604
X601 a_n1095_29019 inv2_0.out.t22 Vdd.t920 Vdd.t919 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X602 a_n11637_9633 Clk.t19 a_n11821_9633 Vss.t31 nfet_03v3
**devattr s=10400,304 d=10400,304
X603 a_459_19209 SARlogic_0.d2.t9 a_275_19209 Vss.t238 nfet_03v3
**devattr s=10400,304 d=10400,304
X604 a_20111_30440 a_18555_31160.t4 Vss.t21 Vss.t20 nfet_03v3
**devattr s=17600,576 d=17600,576
X605 a_37499_31160.t1 inv2_0.out.t23 a_37687_30440 Vss.t661 nfet_03v3
**devattr s=10400,304 d=17600,576
X606 a_30255_29264.t1 a_29583_28100 Vss.t182 Vss.t181 nfet_03v3
**devattr s=17600,576 d=17600,576
X607 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t5 a_n9429_n2007.t2 Vss.t210 nfet_03v3
**devattr s=15600,404 d=15600,404
X608 Vdd.t868 Clk_piso.t13 a_n4631_29217.t3 Vdd.t867 pfet_03v3
**devattr s=26000,604 d=26000,604
X609 Vdd.t271 SARlogic_0.dffrs_2.nand3_8.Z.t6 SARlogic_0.dffrs_2.nand3_1.C.t0 Vdd.t270 pfet_03v3
**devattr s=26000,604 d=26000,604
X610 a_8359_11838 SARlogic_0.dffrs_4.nand3_1.C.t5 Vss.t370 Vss.t369 nfet_03v3
**devattr s=17600,576 d=10400,304
X611 Vss.t387 a_n8385_n2885 a_n8473_n2793 Vss.t386 nfet_03v3
**devattr s=14080,496 d=8320,264
X612 Vdd.t65 Clk.t20 SARlogic_0.dffrs_1.nand3_8.C.t1 Vdd.t64 pfet_03v3
**devattr s=26000,604 d=26000,604
X613 adc_PISO_0.2inmux_4.OUT.t1 a_20783_29264.t5 Vdd.t577 Vdd.t576 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X614 a_2027_29983 a_1167_28099 a_1839_29263.t2 Vdd.t282 pfet_03v3
**devattr s=52800,1376 d=31200,704
X615 Vss.t416 a_40051_37983 Piso_out.t1 Vss.t415 nfet_03v3
**devattr s=9350,280 d=9350,280
X616 SARlogic_0.dffrs_4.Q.t1 SARlogic_0.dffrs_4.Qb.t6 a_10029_11838 Vss.t189 nfet_03v3
**devattr s=10400,304 d=17600,576
X617 Vdd.t641 Vdd.t639 a_n4631_31422.t2 Vdd.t640 pfet_03v3
**devattr s=26000,604 d=26000,604
X618 Vdd.t151 a_8377_29020 a_9083_28820.t3 Vdd.t150 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X619 Vdd.t411 Reset.t57 SARlogic_0.dffrs_1.nand3_6.C.t0 Vdd.t410 pfet_03v3
**devattr s=26000,604 d=26000,604
X620 a_27321_29020 inv2_0.out.t24 Vdd.t922 Vdd.t921 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X621 a_4317_9633 SARlogic_0.dffrs_3.nand3_6.C.t9 Vss.t298 Vss.t297 nfet_03v3
**devattr s=17600,576 d=10400,304
X622 a_4317_14043 Vdd.t981 Vss.t486 Vss.t485 nfet_03v3
**devattr s=17600,576 d=10400,304
X623 SARlogic_0.dffrs_13.nand3_8.C.t3 SARlogic_0.dffrs_13.nand3_6.C.t6 Vdd.t952 Vdd.t951 pfet_03v3
**devattr s=44000,1176 d=26000,604
X624 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t6 a_n9429_n2007.t3 Vss.t211 nfet_03v3
**devattr s=15600,404 d=15600,404
X625 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t7 a_n9429_n2007.t4 Vss.t212 nfet_03v3
**devattr s=15600,404 d=15600,404
X626 SARlogic_0.d0.t1 SARlogic_0.dffrs_11.Qb a_14071_21414 Vss.t176 nfet_03v3
**devattr s=10400,304 d=17600,576
X627 a_n3767_21414 SARlogic_0.dffrs_7.nand3_1.C Vss.t347 Vss.t346 nfet_03v3
**devattr s=17600,576 d=10400,304
X628 Vss.t545 a_n1095_29019 a_n201_28099 Vss.t544 nfet_03v3
**devattr s=10400,304 d=17600,576
X629 Vss.t633 a_10639_30440 a_11311_29264.t3 Vss.t632 nfet_03v3
**devattr s=17600,576 d=17600,576
X630 SARlogic_0.dffrs_2.nand3_6.C.t1 Clk.t21 a_459_11838 Vss.t32 nfet_03v3
**devattr s=10400,304 d=17600,576
X631 a_14071_21414 SARlogic_0.dffrs_11.nand3_6.C.t8 a_13887_21414 Vss.t41 nfet_03v3
**devattr s=10400,304 d=10400,304
X632 SARlogic_0.dffrs_13.nand3_6.C.t0 SARlogic_0.dffrs_13.nand3_1.C.t4 Vdd.t603 Vdd.t602 pfet_03v3
**devattr s=44000,1176 d=26000,604
X633 a_n11821_7428 SARlogic_0.dffrs_13.nand3_8.C.t6 Vss.t142 Vss.t141 nfet_03v3
**devattr s=17600,576 d=10400,304
X634 a_n3767_23619 SARlogic_0.dffrs_0.Qb.t9 Vss.t624 Vss.t623 nfet_03v3
**devattr s=17600,576 d=10400,304
X635 a_39055_30440 a_37499_31160.t4 Vss.t271 Vss.t270 nfet_03v3
**devattr s=17600,576 d=17600,576
X636 Vdd.t263 a_36793_29020 a_37499_28820.t0 Vdd.t262 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X637 a_14313_31423.t2 Clk_piso.t14 a_14577_33720 Vss.t626 nfet_03v3
**devattr s=10400,304 d=17600,576
X638 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t7 Vdd.t359 Vdd.t358 pfet_03v3
**devattr s=26000,604 d=44000,1176
X639 a_n9429_n2007.t11 Vin1.t4 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t5 Vss.t213 nfet_03v3
**devattr s=15600,404 d=15600,404
X640 adc_PISO_0.dffrs_3.Q.t1 adc_PISO_0.dffrs_3.Qb a_25535_33720 Vss.t259 nfet_03v3
**devattr s=10400,304 d=17600,576
X641 adc_PISO_0.dffrs_1.Qb Vdd.t636 Vdd.t638 Vdd.t637 pfet_03v3
**devattr s=26000,604 d=44000,1176
X642 Vdd.t874 adc_PISO_0.dffrs_2.Q.t5 a_18555_31160.t3 Vdd.t873 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X643 SARlogic_0.dffrs_2.Qb.t3 SARlogic_0.dffrs_2.Q.t6 Vdd.t477 Vdd.t476 pfet_03v3
**devattr s=44000,1176 d=26000,604
X644 a_14313_33628.t0 a_14313_31423.t7 a_14577_35925 Vss.t391 nfet_03v3
**devattr s=10400,304 d=17600,576
X645 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t16 Vdd.t575 Vdd.t574 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X646 SARlogic_0.dffrs_2.Q.t3 SARlogic_0.dffrs_2.Qb.t5 a_1945_11838 Vss.t608 nfet_03v3
**devattr s=10400,304 d=17600,576
X647 Vdd.t13 Vss.t688 a_n9861_31159.t3 Vdd.t12 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X648 a_n7809_14043 Vdd.t982 Vss.t484 Vss.t483 nfet_03v3
**devattr s=17600,576 d=10400,304
X649 Vdd.t183 SARlogic_0.dffrs_7.nand3_8.C.t6 SARlogic_0.dffrs_7.Qb Vdd.t182 pfet_03v3
**devattr s=26000,604 d=26000,604
X650 Vss.t454 a_17849_29020 a_18743_28100 Vss.t453 nfet_03v3
**devattr s=10400,304 d=17600,576
X651 Vdd.t177 a_42729_31423.t5 adc_PISO_0.serial_out.t2 Vdd.t176 pfet_03v3
**devattr s=26000,604 d=26000,604
X652 Vdd.t145 SARlogic_0.dffrs_1.nand3_6.C.t6 SARlogic_0.dffrs_2.d.t1 Vdd.t144 pfet_03v3
**devattr s=26000,604 d=26000,604
X653 Vdd.t413 Reset.t58 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t412 pfet_03v3
**devattr s=26000,604 d=26000,604
X654 a_1945_11838 SARlogic_0.dffrs_2.nand3_6.C.t9 a_1761_11838 Vss.t376 nfet_03v3
**devattr s=10400,304 d=10400,304
X655 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t4 Vin1.t5 a_n9429_n2007.t12 Vss.t214 nfet_03v3
**devattr s=15600,404 d=15600,404
X656 Vdd.t67 Clk.t22 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t0 Vdd.t66 pfet_03v3
**devattr s=14080,496 d=14080,496
X657 adc_PISO_0.dffrs_2.Q.t2 Vdd.t633 Vdd.t635 Vdd.t634 pfet_03v3
**devattr s=44000,1176 d=26000,604
X658 adc_PISO_0.2inmux_2.Bit.t1 adc_PISO_0.dffrs_0.Qb Vdd.t1 Vdd.t0 pfet_03v3
**devattr s=26000,604 d=44000,1176
X659 SARlogic_0.dffrs_13.nand3_8.C.t2 SARlogic_0.dffrs_13.nand3_8.Z.t6 Vdd.t93 Vdd.t92 pfet_03v3
**devattr s=26000,604 d=44000,1176
X660 SARlogic_0.dffrs_7.Qb Reset.t59 Vdd.t415 Vdd.t414 pfet_03v3
**devattr s=26000,604 d=44000,1176
X661 SARlogic_0.dffrs_2.d.t3 SARlogic_0.dffrs_1.Qb.t8 Vdd.t373 Vdd.t372 pfet_03v3
**devattr s=26000,604 d=44000,1176
X662 a_4501_7428 Reset.t60 a_4317_7428 Vss.t317 nfet_03v3
**devattr s=10400,304 d=10400,304
X663 SARlogic_0.dffrs_7.nand3_6.C.t0 SARlogic_0.d3.t9 a_n3583_21414 Vss.t56 nfet_03v3
**devattr s=10400,304 d=17600,576
X664 a_275_11838 SARlogic_0.dffrs_2.nand3_1.C.t5 Vss.t396 Vss.t395 nfet_03v3
**devattr s=17600,576 d=10400,304
X665 Vdd.t83 SARlogic_0.dffrs_0.nand3_8.C.t6 SARlogic_0.dffrs_0.Qb.t0 Vdd.t82 pfet_03v3
**devattr s=26000,604 d=26000,604
X666 SARlogic_0.dffrs_1.nand3_8.Z.t3 SARlogic_0.dffrs_1.nand3_8.C.t6 Vdd.t533 Vdd.t532 pfet_03v3
**devattr s=44000,1176 d=26000,604
X667 SARlogic_0.dffrs_12.nand3_8.C.t1 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t21 Vdd.t20 pfet_03v3
**devattr s=26000,604 d=44000,1176
X668 SARlogic_0.dffrs_11.nand3_6.C.t1 SARlogic_0.dffrs_11.nand3_1.C Vdd.t243 Vdd.t242 pfet_03v3
**devattr s=44000,1176 d=26000,604
X669 SARlogic_0.d2.t0 SARlogic_0.dffrs_2.Qb.t6 Vdd.t517 Vdd.t516 pfet_03v3
**devattr s=44000,1176 d=26000,604
X670 SARlogic_0.dffrs_9.nand3_6.C.t3 SARlogic_0.d1.t9 Vdd.t565 Vdd.t564 pfet_03v3
**devattr s=26000,604 d=44000,1176
X671 a_n3583_17004 Reset.t61 a_n3767_17004 Vss.t567 nfet_03v3
**devattr s=10400,304 d=10400,304
X672 SARlogic_0.dffrs_13.nand3_6.C.t3 Clk.t23 Vdd.t69 Vdd.t68 pfet_03v3
**devattr s=26000,604 d=44000,1176
X673 SARlogic_0.dffrs_4.Qb.t0 SARlogic_0.dffrs_4.Q.t6 Vdd.t227 Vdd.t226 pfet_03v3
**devattr s=44000,1176 d=26000,604
X674 SARlogic_0.dffrs_0.d.t0 Reset.t62 Vdd.t778 Vdd.t777 pfet_03v3
**devattr s=44000,1176 d=26000,604
X675 a_n7625_19212 SARlogic_0.d4.t8 a_n7809_19212 Vss.t638 nfet_03v3
**devattr s=10400,304 d=10400,304
X676 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t8 a_n3583_23619 Vss.t233 nfet_03v3
**devattr s=10400,304 d=17600,576
X677 a_37687_28100 SARlogic_0.d0.t11 a_37499_28820.t1 Vss.t254 nfet_03v3
**devattr s=17600,576 d=10400,304
X678 a_9271_30440 adc_PISO_0.dffrs_1.Q.t7 Vss.t621 Vss.t620 nfet_03v3
**devattr s=17600,576 d=10400,304
X679 Vdd.t632 Vdd.t630 a_33337_30170.t2 Vdd.t631 pfet_03v3
**devattr s=26000,604 d=26000,604
X680 adc_PISO_0.dffrs_3.Qb Vdd.t983 a_25535_31516 Vss.t482 nfet_03v3
**devattr s=10400,304 d=17600,576
X681 a_10029_11838 SARlogic_0.dffrs_4.nand3_6.C.t8 a_9845_11838 Vss.t65 nfet_03v3
**devattr s=10400,304 d=10400,304
X682 Vdd.t313 a_n9629_1405 a_n9717_1497 Vdd.t312 pfet_03v3
**devattr s=17600,576 d=10400,304
X683 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_4.Qb.t7 Vdd.t255 Vdd.t254 pfet_03v3
**devattr s=44000,1176 d=26000,604
X684 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t7 Vdd.t906 Vdd.t905 pfet_03v3
**devattr s=26000,604 d=44000,1176
X685 a_n8305_28099 a_n9861_28819.t4 Vss.t390 Vss.t389 nfet_03v3
**devattr s=17600,576 d=17600,576
X686 a_n3583_19209 SARlogic_0.d3.t10 a_n3767_19209 Vss.t55 nfet_03v3
**devattr s=10400,304 d=10400,304
X687 a_29583_28100 a_28027_28820.t5 Vdd.t467 Vdd.t466 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X688 SARlogic_0.dffrs_4.nand3_8.Z.t2 SARlogic_0.dffrs_4.d.t7 a_8543_7428 Vss.t654 nfet_03v3
**devattr s=10400,304 d=17600,576
X689 a_4841_29217.t1 a_4921_30169.t5 Vdd.t914 Vdd.t913 pfet_03v3
**devattr s=26000,604 d=44000,1176
X690 a_1167_28099 a_n389_28819.t4 Vss.t447 Vss.t446 nfet_03v3
**devattr s=17600,576 d=17600,576
X691 Vdd.t870 Clk_piso.t15 a_33257_29218.t3 Vdd.t869 pfet_03v3
**devattr s=26000,604 d=26000,604
X692 Vdd.t211 SARlogic_0.dffrs_1.nand3_8.Z.t5 SARlogic_0.dffrs_1.nand3_1.C.t0 Vdd.t210 pfet_03v3
**devattr s=26000,604 d=26000,604
X693 a_24049_33720 Vdd.t984 a_23865_33720 Vss.t481 nfet_03v3
**devattr s=10400,304 d=10400,304
X694 Vdd.t832 a_42729_29218.t5 adc_PISO_0.dffrs_5.Qb Vdd.t831 pfet_03v3
**devattr s=26000,604 d=26000,604
X695 a_n8305_28099 a_n9861_28819.t5 Vdd.t515 Vdd.t514 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X696 adc_PISO_0.dffrs_2.Qb adc_PISO_0.dffrs_2.Q.t6 Vdd.t85 Vdd.t84 pfet_03v3
**devattr s=44000,1176 d=26000,604
X697 adc_PISO_0.dffrs_1.Q.t3 Vdd.t627 Vdd.t629 Vdd.t628 pfet_03v3
**devattr s=44000,1176 d=26000,604
X698 a_20783_29264.t0 a_20111_28100 a_20971_29984 Vdd.t28 pfet_03v3
**devattr s=31200,704 d=52800,1376
X699 a_4841_31422.t3 Clk_piso.t16 Vdd.t938 Vdd.t937 pfet_03v3
**devattr s=26000,604 d=44000,1176
X700 a_5803_19210 SARlogic_0.d2.t10 Vss.t240 Vss.t239 nfet_03v3
**devattr s=17600,576 d=10400,304
X701 a_37687_30440 adc_PISO_0.2inmux_1.Bit.t8 Vss.t345 Vss.t344 nfet_03v3
**devattr s=17600,576 d=10400,304
X702 a_n4551_31514 a_n4631_31422.t7 Vss.t672 Vss.t671 nfet_03v3
**devattr s=17600,576 d=10400,304
X703 a_12585_14043 SARlogic_0.dffrs_5.nand3_8.Z.t5 a_12401_14043 Vss.t145 nfet_03v3
**devattr s=10400,304 d=10400,304
X704 Vss.t38 adc_PISO_0.2inmux_2.Bit.t7 a_n201_30439 Vss.t37 nfet_03v3
**devattr s=10400,304 d=17600,576
X705 a_24049_35925 a_23865_30170.t6 a_23865_35925 Vss.t605 nfet_03v3
**devattr s=10400,304 d=10400,304
X706 a_1167_28099 a_n389_28819.t5 Vdd.t593 Vdd.t592 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X707 SARlogic_0.dffrs_13.nand3_1.C.t0 Reset.t63 Vdd.t780 Vdd.t779 pfet_03v3
**devattr s=44000,1176 d=26000,604
X708 SARlogic_0.dffrs_12.nand3_8.C.t2 SARlogic_0.dffrs_12.nand3_6.C.t8 Vdd.t345 Vdd.t344 pfet_03v3
**devattr s=44000,1176 d=26000,604
X709 SARlogic_0.dffrs_10.nand3_8.C.t1 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t355 Vdd.t354 pfet_03v3
**devattr s=26000,604 d=44000,1176
X710 SARlogic_0.dffrs_0.nand3_8.C.t0 SARlogic_0.dffrs_0.nand3_8.Z.t6 a_n7625_9633 Vss.t68 nfet_03v3
**devattr s=10400,304 d=17600,576
X711 SARlogic_0.dffrs_9.nand3_6.C.t1 SARlogic_0.dffrs_9.nand3_1.C Vdd.t285 Vdd.t284 pfet_03v3
**devattr s=44000,1176 d=26000,604
X712 a_n4551_33719 a_n4631_33627.t5 Vss.t440 Vss.t439 nfet_03v3
**devattr s=17600,576 d=10400,304
X713 SARlogic_0.dffrs_0.d.t1 SARlogic_0.dffrs_13.Qb.t7 Vdd.t816 Vdd.t815 pfet_03v3
**devattr s=26000,604 d=44000,1176
X714 a_14393_31515 a_14313_31423.t8 Vss.t393 Vss.t392 nfet_03v3
**devattr s=17600,576 d=10400,304
X715 adc_PISO_0.2inmux_1.OUT.t1 a_39727_29264.t5 Vdd.t842 Vdd.t841 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X716 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_2.Qb.t7 Vdd.t519 Vdd.t518 pfet_03v3
**devattr s=44000,1176 d=26000,604
X717 SARlogic_0.dffrs_4.Qb.t2 Reset.t64 Vdd.t782 Vdd.t781 pfet_03v3
**devattr s=26000,604 d=44000,1176
X718 SARlogic_0.dffrs_1.nand3_8.C.t2 SARlogic_0.dffrs_1.nand3_6.C.t7 Vdd.t147 Vdd.t146 pfet_03v3
**devattr s=44000,1176 d=26000,604
X719 a_9083_28820.t0 SARlogic_0.d3.t11 a_9271_28100 Vss.t54 nfet_03v3
**devattr s=10400,304 d=17600,576
X720 a_42809_30170.t0 a_42729_29218.t6 Vdd.t115 Vdd.t114 pfet_03v3
**devattr s=44000,1176 d=26000,604
X721 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t13 Vss.t339 nfet_03v3
**devattr s=20800,504 d=20800,504
X722 SARlogic_0.dffrs_11.Qb Reset.t65 Vdd.t784 Vdd.t783 pfet_03v3
**devattr s=26000,604 d=44000,1176
X723 SARlogic_0.dffrs_5.Q.t1 SARlogic_0.dffrs_5.Qb.t8 Vdd.t850 Vdd.t849 pfet_03v3
**devattr s=26000,604 d=44000,1176
X724 SARlogic_0.dffrs_5.nand3_8.C.t1 SARlogic_0.dffrs_5.nand3_8.Z.t6 a_12585_9633 Vss.t146 nfet_03v3
**devattr s=10400,304 d=17600,576
X725 SARlogic_0.dffrs_1.nand3_6.C.t3 SARlogic_0.dffrs_1.nand3_1.C.t4 Vdd.t872 Vdd.t871 pfet_03v3
**devattr s=44000,1176 d=26000,604
X726 a_23865_29310 a_23785_29218.t7 Vss.t151 Vss.t150 nfet_03v3
**devattr s=17600,576 d=10400,304
X727 Vdd.t251 SARlogic_0.dffrs_11.nand3_8.C.t6 SARlogic_0.dffrs_11.Qb Vdd.t250 pfet_03v3
**devattr s=26000,604 d=26000,604
X728 Vdd.t902 a_39055_30440 a_39915_29984 Vdd.t901 pfet_03v3
**devattr s=31200,704 d=52800,1376
X729 a_42729_29218.t2 a_42729_31423.t6 Vdd.t179 Vdd.t178 pfet_03v3
**devattr s=44000,1176 d=26000,604
X730 Vdd.t744 SARlogic_0.dffrs_5.nand3_6.C.t7 SARlogic_0.dffrs_5.Q.t2 Vdd.t743 pfet_03v3
**devattr s=26000,604 d=26000,604
X731 a_28027_28820.t1 SARlogic_0.d1.t10 a_28215_28100 Vss.t430 nfet_03v3
**devattr s=10400,304 d=17600,576
X732 a_n4631_29217.t2 a_n4551_30169.t6 a_n4367_31514 Vss.t227 nfet_03v3
**devattr s=10400,304 d=17600,576
X733 comparator_no_offsetcal_0.no_offsetLatch_0.Vq comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t17 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t2 Vss.t459 nfet_03v3
**devattr s=20800,504 d=20800,504
X734 a_29583_30440 a_28027_31160.t5 Vss.t585 Vss.t584 nfet_03v3
**devattr s=17600,576 d=17600,576
X735 SARlogic_0.dffrs_13.nand3_1.C.t2 SARlogic_0.dffrs_13.nand3_6.C.t7 Vdd.t954 Vdd.t953 pfet_03v3
**devattr s=26000,604 d=44000,1176
X736 SARlogic_0.dffrs_10.nand3_8.C.t2 SARlogic_0.dffrs_10.nand3_6.C.t9 Vdd.t291 Vdd.t290 pfet_03v3
**devattr s=44000,1176 d=26000,604
X737 a_n4631_31422.t3 Clk_piso.t17 a_n4367_33719 Vss.t674 nfet_03v3
**devattr s=10400,304 d=17600,576
X738 SARlogic_0.dffrs_4.d.t1 SARlogic_0.dffrs_3.Qb.t9 a_5987_11838 Vss.t123 nfet_03v3
**devattr s=10400,304 d=17600,576
X739 adc_PISO_0.dffrs_2.Q.t0 adc_PISO_0.dffrs_2.Qb a_16063_33720 Vss.t366 nfet_03v3
**devattr s=10400,304 d=17600,576
X740 a_n3065_33719 Vdd.t985 Vss.t480 Vss.t479 nfet_03v3
**devattr s=17600,576 d=10400,304
X741 SARlogic_0.dffrs_14.nand3_8.C.t3 SARlogic_0.dffrs_14.nand3_6.C.t9 Vdd.t381 Vdd.t380 pfet_03v3
**devattr s=44000,1176 d=26000,604
X742 a_n9861_31159.t2 inv2_0.out.t25 Vdd.t924 Vdd.t923 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X743 adc_PISO_0.serial_out.t0 adc_PISO_0.dffrs_5.Qb a_44479_33720 Vss.t388 nfet_03v3
**devattr s=10400,304 d=17600,576
X744 a_n2281_11838 Vdd.t986 Vss.t478 Vss.t477 nfet_03v3
**devattr s=17600,576 d=10400,304
X745 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t15 Vdd.t928 Vdd.t927 pfet_03v3
**devattr s=10400,304 d=10400,304
X746 a_n8305_30439 a_n9861_31159.t5 Vss.t131 Vss.t130 nfet_03v3
**devattr s=17600,576 d=17600,576
X747 a_16063_33720 a_14313_31423.t9 a_15879_33720 Vss.t394 nfet_03v3
**devattr s=10400,304 d=10400,304
X748 a_n2881_33719 a_n4631_31422.t8 a_n3065_33719 Vss.t673 nfet_03v3
**devattr s=10400,304 d=10400,304
X749 SARlogic_0.dffrs_2.nand3_8.C.t1 SARlogic_0.dffrs_2.nand3_8.Z.t7 a_459_9633 Vss.t201 nfet_03v3
**devattr s=10400,304 d=17600,576
X750 SARlogic_0.dffrs_2.Qb.t1 Reset.t66 Vdd.t786 Vdd.t785 pfet_03v3
**devattr s=26000,604 d=44000,1176
X751 Vss.t539 a_n10831_4320 Comp_out.t1 Vss.t538 nfet_03v3
**devattr s=9350,280 d=9350,280
X752 a_10639_28100 a_9083_28820.t5 Vss.t653 Vss.t652 nfet_03v3
**devattr s=17600,576 d=17600,576
X753 SARlogic_0.dffrs_1.nand3_8.C.t3 SARlogic_0.dffrs_1.nand3_8.Z.t6 Vdd.t213 Vdd.t212 pfet_03v3
**devattr s=26000,604 d=44000,1176
X754 SARlogic_0.dffrs_3.nand3_8.Z.t1 SARlogic_0.dffrs_2.Q.t7 a_4501_7428 Vss.t363 nfet_03v3
**devattr s=10400,304 d=17600,576
X755 SARlogic_0.dffrs_14.nand3_6.C.t2 SARlogic_0.dffrs_14.nand3_1.C Vdd.t469 Vdd.t468 pfet_03v3
**devattr s=44000,1176 d=26000,604
X756 Vss.t180 adc_PISO_0.dffrs_3.Q.t8 a_28215_30440 Vss.t179 nfet_03v3
**devattr s=10400,304 d=17600,576
X757 Vss.t195 a_36793_29020 a_37687_28100 Vss.t194 nfet_03v3
**devattr s=10400,304 d=17600,576
X758 a_1167_30439 a_n389_31159.t5 Vss.t62 Vss.t61 nfet_03v3
**devattr s=17600,576 d=17600,576
X759 Vdd.t916 SARlogic_0.dffrs_2.nand3_8.C.t6 SARlogic_0.dffrs_2.Qb.t2 Vdd.t915 pfet_03v3
**devattr s=26000,604 d=26000,604
X760 SARlogic_0.dffrs_5.nand3_8.Z.t3 SARlogic_0.dffrs_5.nand3_8.C.t7 Vdd.t463 Vdd.t462 pfet_03v3
**devattr s=44000,1176 d=26000,604
X761 SARlogic_0.dffrs_8.nand3_8.C.t2 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t325 Vdd.t324 pfet_03v3
**devattr s=26000,604 d=44000,1176
X762 SARlogic_0.dffrs_1.nand3_6.C.t1 Clk.t24 Vdd.t3 Vdd.t2 pfet_03v3
**devattr s=26000,604 d=44000,1176
X763 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t8 Vdd.t361 Vdd.t360 pfet_03v3
**devattr s=26000,604 d=44000,1176
X764 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_8.C.t7 Vdd.t253 Vdd.t252 pfet_03v3
**devattr s=44000,1176 d=26000,604
X765 Vdd.t5 Clk.t25 SARlogic_0.dffrs_13.nand3_8.C.t0 Vdd.t4 pfet_03v3
**devattr s=26000,604 d=26000,604
X766 SARlogic_0.dffrs_1.nand3_8.C.t0 SARlogic_0.dffrs_1.nand3_8.Z.t7 a_n3583_9633 Vss.t22 nfet_03v3
**devattr s=10400,304 d=17600,576
X767 a_459_11838 Reset.t67 a_275_11838 Vss.t568 nfet_03v3
**devattr s=10400,304 d=10400,304
X768 SARlogic_0.dffrs_2.nand3_8.Z.t3 SARlogic_0.dffrs_2.nand3_8.C.t7 Vdd.t918 Vdd.t917 pfet_03v3
**devattr s=44000,1176 d=26000,604
X769 SARlogic_0.dffrs_11.nand3_6.C.t3 SARlogic_0.dffrs_12.Q.t9 a_12585_21414 Vss.t426 nfet_03v3
**devattr s=10400,304 d=17600,576
X770 Vdd.t788 Reset.t68 SARlogic_0.dffrs_11.nand3_6.C.t0 Vdd.t787 pfet_03v3
**devattr s=26000,604 d=26000,604
X771 Vdd.t908 SARlogic_0.dffrs_9.nand3_6.C.t8 SARlogic_0.d2.t3 Vdd.t907 pfet_03v3
**devattr s=26000,604 d=26000,604
X772 adc_PISO_0.dffrs_2.Qb Vdd.t987 a_16063_31516 Vss.t476 nfet_03v3
**devattr s=10400,304 d=17600,576
X773 a_n3767_17004 SARlogic_0.dffrs_7.nand3_8.C.t7 Vss.t125 Vss.t124 nfet_03v3
**devattr s=17600,576 d=10400,304
X774 Vdd.t626 Vdd.t624 SARlogic_0.dffrs_13.nand3_6.C.t1 Vdd.t625 pfet_03v3
**devattr s=26000,604 d=26000,604
X775 Vdd.t459 SARlogic_0.dffrs_4.nand3_8.C.t7 SARlogic_0.dffrs_4.Qb.t3 Vdd.t458 pfet_03v3
**devattr s=26000,604 d=26000,604
X776 adc_PISO_0.dffrs_5.Qb Vdd.t988 a_44479_31516 Vss.t475 nfet_03v3
**devattr s=10400,304 d=17600,576
X777 a_16063_31516 a_14313_29218.t7 a_15879_31516 Vss.t253 nfet_03v3
**devattr s=10400,304 d=10400,304
X778 a_6591_33719 a_4841_31422.t8 a_6407_33719 Vss.t360 nfet_03v3
**devattr s=10400,304 d=10400,304
X779 a_n4631_33627.t3 Vdd.t621 Vdd.t623 Vdd.t622 pfet_03v3
**devattr s=44000,1176 d=26000,604
X780 SARlogic_0.dffrs_0.nand3_1.C.t1 SARlogic_0.dffrs_0.nand3_6.C.t9 a_n7625_14043 Vss.t377 nfet_03v3
**devattr s=10400,304 d=17600,576
X781 a_42729_31423.t3 Clk_piso.t18 a_42993_33720 Vss.t675 nfet_03v3
**devattr s=10400,304 d=17600,576
X782 a_33337_30170.t1 adc_PISO_0.2inmux_5.OUT.t3 Vdd.t501 Vdd.t500 pfet_03v3
**devattr s=26000,604 d=44000,1176
X783 a_n3767_19209 SARlogic_0.dffrs_7.nand3_6.C.t9 Vss.t235 Vss.t234 nfet_03v3
**devattr s=17600,576 d=10400,304
X784 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t9 a_12585_23619 Vss.t42 nfet_03v3
**devattr s=10400,304 d=17600,576
X785 Vdd.t171 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_1.C Vdd.t170 pfet_03v3
**devattr s=26000,604 d=26000,604
X786 a_14577_33720 Vdd.t989 a_14393_33720 Vss.t474 nfet_03v3
**devattr s=10400,304 d=10400,304
X787 a_14313_31423.t0 a_14313_33628.t5 Vdd.t489 Vdd.t488 pfet_03v3
**devattr s=44000,1176 d=26000,604
X788 a_n2281_9634 SARlogic_0.dffrs_2.d.t6 Vss.t19 Vss.t18 nfet_03v3
**devattr s=17600,576 d=10400,304
X789 a_n7625_9633 Clk.t26 a_n7809_9633 Vss.t1 nfet_03v3
**devattr s=10400,304 d=10400,304
X790 a_14393_30170.t0 adc_PISO_0.2inmux_3.OUT.t3 a_14577_29310 Vss.t199 nfet_03v3
**devattr s=10400,304 d=17600,576
X791 a_11311_29264.t1 a_10639_28100 a_11499_29984 Vdd.t598 pfet_03v3
**devattr s=31200,704 d=52800,1376
X792 a_42729_33628.t1 a_42729_31423.t7 a_42993_35925 Vss.t163 nfet_03v3
**devattr s=10400,304 d=17600,576
X793 Vdd.t543 a_40051_37983 Piso_out.t4 Vdd.t542 pfet_03v3
**devattr s=18700,450 d=18700,450
X794 a_4501_21414 Reset.t69 a_4317_21414 Vss.t569 nfet_03v3
**devattr s=10400,304 d=10400,304
X795 a_33257_29218.t2 a_33337_30170.t7 Vdd.t511 Vdd.t510 pfet_03v3
**devattr s=26000,604 d=44000,1176
X796 SARlogic_0.dffrs_1.nand3_1.C.t1 Vdd.t615 Vdd.t617 Vdd.t616 pfet_03v3
**devattr s=44000,1176 d=26000,604
X797 a_n9429_n2007.t13 Vin1.t6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t3 Vss.t209 nfet_03v3
**devattr s=15600,404 d=15600,404
X798 SARlogic_0.dffrs_8.nand3_8.C.t0 SARlogic_0.dffrs_8.nand3_6.C.t9 Vdd.t91 Vdd.t90 pfet_03v3
**devattr s=44000,1176 d=26000,604
X799 a_39915_29984 a_39055_30440 Vdd.t900 Vdd.t899 pfet_03v3
**devattr s=52800,1376 d=31200,704
X800 a_14577_35925 a_14393_30170.t7 a_14393_35925 Vss.t651 nfet_03v3
**devattr s=10400,304 d=10400,304
X801 a_14313_33628.t1 Vdd.t618 Vdd.t620 Vdd.t619 pfet_03v3
**devattr s=44000,1176 d=26000,604
X802 a_n10151_11838 SARlogic_0.dffrs_13.nand3_6.C.t8 a_n10335_11838 Vss.t686 nfet_03v3
**devattr s=10400,304 d=10400,304
X803 a_5987_19210 SARlogic_0.dffrs_9.nand3_8.C.t6 a_5803_19210 Vss.t443 nfet_03v3
**devattr s=10400,304 d=10400,304
X804 a_4501_23619 SARlogic_0.dffrs_9.nand3_8.Z a_4317_23619 Vss.t111 nfet_03v3
**devattr s=10400,304 d=10400,304
X805 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_8.C.t7 Vdd.t589 Vdd.t588 pfet_03v3
**devattr s=44000,1176 d=26000,604
X806 Vdd.t930 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t16 comparator_no_offsetcal_0.x5.out Vdd.t929 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X807 a_n3583_7428 Reset.t70 a_n3767_7428 Vss.t570 nfet_03v3
**devattr s=10400,304 d=10400,304
X808 Vdd.t15 Vss.t689 SARlogic_0.dffrs_12.nand3_8.C.t3 Vdd.t14 pfet_03v3
**devattr s=26000,604 d=26000,604
X809 a_5105_31514 Clk_piso.t19 a_4921_31514 Vss.t676 nfet_03v3
**devattr s=10400,304 d=10400,304
X810 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t9 a_n3583_17004 Vss.t278 nfet_03v3
**devattr s=10400,304 d=17600,576
X811 adc_PISO_0.2inmux_2.OUT.t1 a_1839_29263.t5 Vdd.t235 Vdd.t234 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X812 a_4921_31514 a_4841_31422.t9 Vss.t362 Vss.t361 nfet_03v3
**devattr s=17600,576 d=10400,304
X813 a_20783_29264.t2 a_20111_28100 Vss.t12 Vss.t11 nfet_03v3
**devattr s=17600,576 d=17600,576
X814 a_5105_33719 Vdd.t990 a_4921_33719 Vss.t473 nfet_03v3
**devattr s=10400,304 d=10400,304
X815 a_n4631_33627.t1 a_n4631_31422.t9 Vdd.t936 Vdd.t935 pfet_03v3
**devattr s=26000,604 d=44000,1176
X816 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t2 Vin1.t7 a_n9429_n2007.t14 Vss.t210 nfet_03v3
**devattr s=15600,404 d=15600,404
X817 SARlogic_0.dffrs_2.Qb.t0 Reset.t71 a_1945_9634 Vss.t571 nfet_03v3
**devattr s=10400,304 d=17600,576
X818 a_33337_30170.t3 a_33257_29218.t7 Vdd.t810 Vdd.t809 pfet_03v3
**devattr s=44000,1176 d=26000,604
X819 a_42993_31515 Clk_piso.t20 a_42809_31515 Vss.t677 nfet_03v3
**devattr s=10400,304 d=10400,304
X820 a_8543_14043 SARlogic_0.dffrs_4.nand3_8.Z.t7 a_8359_14043 Vss.t368 nfet_03v3
**devattr s=10400,304 d=10400,304
X821 SARlogic_0.dffrs_7.nand3_8.C.t2 SARlogic_0.dffrs_7.nand3_8.Z a_n3583_19209 Vss.t207 nfet_03v3
**devattr s=10400,304 d=17600,576
X822 a_28215_28100 a_27321_29020 Vss.t136 Vss.t135 nfet_03v3
**devattr s=17600,576 d=10400,304
X823 adc_PISO_0.2inmux_3.OUT.t0 a_11311_29264.t5 Vdd.t209 Vdd.t208 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X824 a_4921_33719 a_4841_33627.t5 Vss.t381 Vss.t380 nfet_03v3
**devattr s=17600,576 d=10400,304
X825 a_n7809_7428 SARlogic_0.dffrs_0.nand3_8.C.t7 Vss.t44 Vss.t43 nfet_03v3
**devattr s=17600,576 d=10400,304
X826 Vss.t537 a_n10831_4320 Comp_out.t0 Vss.t536 nfet_03v3
**devattr s=9350,280 d=9350,280
X827 SARlogic_0.dffrs_13.Qb.t1 Vdd.t991 a_n10151_9634 Vss.t472 nfet_03v3
**devattr s=10400,304 d=17600,576
X828 SARlogic_0.dffrs_1.nand3_1.C.t3 SARlogic_0.dffrs_1.nand3_6.C.t8 Vdd.t149 Vdd.t148 pfet_03v3
**devattr s=26000,604 d=44000,1176
X829 a_17849_29020 inv2_0.out.t26 Vss.t663 Vss.t662 nfet_03v3
**devattr s=17600,576 d=17600,576
X830 a_33257_29218.t0 a_33257_31423.t9 Vdd.t529 Vdd.t528 pfet_03v3
**devattr s=44000,1176 d=26000,604
X831 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t1 Vin1.t8 a_n9429_n2007.t15 Vss.t211 nfet_03v3
**devattr s=15600,404 d=15600,404
X832 a_24049_29310 Vdd.t992 a_23865_29310 Vss.t471 nfet_03v3
**devattr s=10400,304 d=10400,304
X833 a_n4367_31514 Clk_piso.t21 a_n4551_31514 Vss.t186 nfet_03v3
**devattr s=10400,304 d=10400,304
X834 adc_PISO_0.dffrs_0.Qb adc_PISO_0.2inmux_2.Bit.t8 Vdd.t75 Vdd.t74 pfet_03v3
**devattr s=44000,1176 d=26000,604
X835 SARlogic_0.dffrs_3.Qb.t1 Reset.t72 Vdd.t790 Vdd.t789 pfet_03v3
**devattr s=26000,604 d=44000,1176
X836 a_n9429_n2007.t0 Clk.t27 Vss.t3 Vss.t2 nfet_03v3
**devattr s=8320,264 d=8320,264
X837 SARlogic_0.dffrs_1.Qb.t0 SARlogic_0.dffrs_2.d.t7 Vdd.t41 Vdd.t40 pfet_03v3
**devattr s=44000,1176 d=26000,604
X838 a_n389_28819.t0 SARlogic_0.d4.t9 a_n201_28099 Vss.t114 nfet_03v3
**devattr s=10400,304 d=17600,576
X839 Vdd.t95 SARlogic_0.dffrs_13.nand3_8.Z.t7 SARlogic_0.dffrs_13.nand3_1.C.t3 Vdd.t94 pfet_03v3
**devattr s=26000,604 d=26000,604
X840 Vdd.t553 a_n4631_29217.t6 adc_PISO_0.dffrs_0.Qb Vdd.t552 pfet_03v3
**devattr s=26000,604 d=26000,604
X841 Vdd.t792 Reset.t73 SARlogic_0.dffrs_5.nand3_8.Z.t2 Vdd.t791 pfet_03v3
**devattr s=26000,604 d=26000,604
X842 a_n4367_33719 Vdd.t993 a_n4551_33719 Vss.t470 nfet_03v3
**devattr s=10400,304 d=10400,304
X843 a_n3583_11838 Reset.t74 a_n3767_11838 Vss.t572 nfet_03v3
**devattr s=10400,304 d=10400,304
X844 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_8.C.t7 Vdd.t351 Vdd.t350 pfet_03v3
**devattr s=44000,1176 d=26000,604
X845 a_n4551_29309 a_n4631_29217.t7 Vss.t423 Vss.t422 nfet_03v3
**devattr s=17600,576 d=10400,304
X846 a_n9429_n2007.t5 Vin2.t8 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t213 nfet_03v3
**devattr s=15600,404 d=15600,404
X847 a_n389_28819.t1 SARlogic_0.d4.t10 Vdd.t161 Vdd.t160 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X848 Vss.t414 a_40051_37983 Piso_out.t0 Vss.t413 nfet_03v3
**devattr s=9350,280 d=9350,280
X849 a_30443_29984 a_29583_28100 a_30255_29264.t2 Vdd.t248 pfet_03v3
**devattr s=52800,1376 d=31200,704
X850 Vdd.t794 Reset.t75 SARlogic_0.dffrs_2.nand3_8.Z.t2 Vdd.t793 pfet_03v3
**devattr s=26000,604 d=26000,604
X851 a_n11821_11838 SARlogic_0.dffrs_13.nand3_1.C.t5 Vss.t458 Vss.t457 nfet_03v3
**devattr s=17600,576 d=10400,304
X852 SARlogic_0.dffrs_5.nand3_8.C.t2 SARlogic_0.dffrs_5.nand3_8.Z.t7 Vdd.t207 Vdd.t206 pfet_03v3
**devattr s=26000,604 d=44000,1176
X853 Vss.t85 a_n8305_30439 a_n7633_29263.t0 Vss.t84 nfet_03v3
**devattr s=17600,576 d=17600,576
X854 SARlogic_0.dffrs_14.nand3_8.C.t1 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t25 Vdd.t24 pfet_03v3
**devattr s=26000,604 d=44000,1176
X855 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t9 a_n9429_n2007.t6 Vss.t214 nfet_03v3
**devattr s=15600,404 d=15600,404
X856 Vdd.t796 Reset.t76 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t795 pfet_03v3
**devattr s=26000,604 d=26000,604
X857 SARlogic_0.dffrs_5.nand3_6.C.t0 Clk.t28 Vdd.t7 Vdd.t6 pfet_03v3
**devattr s=26000,604 d=44000,1176
X858 SARlogic_0.dffrs_14.nand3_6.C.t0 SARlogic_0.d4.t11 Vdd.t163 Vdd.t162 pfet_03v3
**devattr s=26000,604 d=44000,1176
X859 SARlogic_0.d5.t3 SARlogic_0.dffrs_13.Qb.t8 Vdd.t818 Vdd.t817 pfet_03v3
**devattr s=44000,1176 d=26000,604
X860 Vdd.t595 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t594 pfet_03v3
**devattr s=17600,576 d=17600,576
X861 a_n9673_28099 SARlogic_0.d5.t7 a_n9861_28819.t1 Vss.t229 nfet_03v3
**devattr s=17600,576 d=10400,304
X862 adc_PISO_0.dffrs_1.Qb Vdd.t994 a_6591_31515 Vss.t469 nfet_03v3
**devattr s=10400,304 d=17600,576
X863 Vdd.t317 a_4841_29217.t6 adc_PISO_0.dffrs_1.Qb Vdd.t316 pfet_03v3
**devattr s=26000,604 d=26000,604
X864 a_11499_29984 a_10639_30440 Vdd.t886 Vdd.t885 pfet_03v3
**devattr s=52800,1376 d=31200,704
X865 a_23865_30170.t3 adc_PISO_0.2inmux_4.OUT.t3 Vdd.t828 Vdd.t827 pfet_03v3
**devattr s=26000,604 d=44000,1176
X866 SARlogic_0.d0.t3 SARlogic_0.dffrs_4.Qb.t8 Vdd.t257 Vdd.t256 pfet_03v3
**devattr s=44000,1176 d=26000,604
X867 Vss.t349 comparator_no_offsetcal_0.x5.out comparator_no_offsetcal_0.x2.Vout2 Vss.t348 nfet_03v3
**devattr s=17600,576 d=17600,576
X868 a_18743_30440 inv2_0.out.t27 a_18555_31160.t0 Vss.t664 nfet_03v3
**devattr s=17600,576 d=10400,304
X869 Vdd.t9 Clk.t29 SARlogic_0.dffrs_3.nand3_8.C.t0 Vdd.t8 pfet_03v3
**devattr s=26000,604 d=26000,604
X870 a_n9429_n2007.t16 Vin1.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t0 Vss.t263 nfet_03v3
**devattr s=15600,404 d=15600,404
X871 adc_PISO_0.serial_out.t3 Vdd.t612 Vdd.t614 Vdd.t613 pfet_03v3
**devattr s=44000,1176 d=26000,604
X872 a_44479_33720 a_42729_31423.t8 a_44295_33720 Vss.t164 nfet_03v3
**devattr s=10400,304 d=10400,304
X873 a_n2097_11838 SARlogic_0.dffrs_1.nand3_6.C.t9 a_n2281_11838 Vss.t105 nfet_03v3
**devattr s=10400,304 d=10400,304
X874 a_n7625_14043 SARlogic_0.dffrs_0.nand3_8.Z.t7 a_n7809_14043 Vss.t69 nfet_03v3
**devattr s=10400,304 d=10400,304
X875 adc_PISO_0.2inmux_2.Bit.t0 adc_PISO_0.dffrs_0.Qb a_n2881_33719 Vss.t0 nfet_03v3
**devattr s=10400,304 d=17600,576
X876 a_15879_33720 Vdd.t995 Vss.t468 Vss.t467 nfet_03v3
**devattr s=17600,576 d=10400,304
X877 a_23785_29218.t2 a_23865_30170.t7 Vdd.t838 Vdd.t837 pfet_03v3
**devattr s=26000,604 d=44000,1176
X878 a_n4551_30169.t1 adc_PISO_0.2inmux_0.OUT.t3 a_n4367_29309 Vss.t139 nfet_03v3
**devattr s=10400,304 d=17600,576
X879 Vdd.t201 a_4921_30169.t6 a_4841_33627.t0 Vdd.t200 pfet_03v3
**devattr s=26000,604 d=26000,604
X880 Vdd.t798 Reset.t77 SARlogic_0.dffrs_3.nand3_6.C.t1 Vdd.t797 pfet_03v3
**devattr s=26000,604 d=26000,604
X881 Vdd.t611 Vdd.t609 a_42729_31423.t1 Vdd.t610 pfet_03v3
**devattr s=26000,604 d=26000,604
X882 Vdd.t203 SARlogic_0.dffrs_13.nand3_8.C.t7 SARlogic_0.dffrs_13.Qb.t0 Vdd.t202 pfet_03v3
**devattr s=26000,604 d=26000,604
X883 SARlogic_0.dffrs_2.d.t2 SARlogic_0.dffrs_1.Qb.t9 a_n2097_11838 Vss.t292 nfet_03v3
**devattr s=10400,304 d=17600,576
X884 a_n3767_7428 SARlogic_0.dffrs_1.nand3_8.C.t7 Vss.t410 Vss.t409 nfet_03v3
**devattr s=17600,576 d=10400,304
X885 a_4841_33627.t3 Vdd.t606 Vdd.t608 Vdd.t607 pfet_03v3
**devattr s=44000,1176 d=26000,604
X886 SARlogic_0.dffrs_9.nand3_6.C.t2 SARlogic_0.d1.t11 a_4501_21414 Vss.t431 nfet_03v3
**devattr s=10400,304 d=17600,576
X887 a_5803_21414 SARlogic_0.dffrs_2.Qb.t8 Vss.t400 Vss.t399 nfet_03v3
**devattr s=17600,576 d=10400,304
X888 a_12401_21414 SARlogic_0.dffrs_11.nand3_1.C Vss.t174 Vss.t173 nfet_03v3
**devattr s=17600,576 d=10400,304
X889 a_8543_9633 Clk.t30 a_8359_9633 Vss.t4 nfet_03v3
**devattr s=10400,304 d=10400,304
X890 Vdd.t800 Reset.t78 SARlogic_0.dffrs_10.nand3_6.C.t1 Vdd.t799 pfet_03v3
**devattr s=26000,604 d=26000,604
X891 Vdd.t311 SARlogic_0.d2.t11 SARlogic_0.dffrs_8.nand3_8.C.t3 Vdd.t310 pfet_03v3
**devattr s=26000,604 d=26000,604
X892 SARlogic_0.dffrs_13.nand3_6.C.t2 Clk.t31 a_n11637_11838 Vss.t5 nfet_03v3
**devattr s=10400,304 d=17600,576
X893 Vdd.t898 a_42809_30170.t7 a_42729_33628.t3 Vdd.t897 pfet_03v3
**devattr s=26000,604 d=26000,604
X894 a_20111_30440 a_18555_31160.t5 Vdd.t802 Vdd.t801 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X895 a_n10335_11838 Reset.t79 Vss.t574 Vss.t573 nfet_03v3
**devattr s=17600,576 d=10400,304
X896 a_n6693_1497 a_n6893_1405 Vdd.t493 Vdd.t492 pfet_03v3
**devattr s=10400,304 d=17600,576
X897 a_n6323_19213 SARlogic_0.d5.t8 Vss.t231 Vss.t230 nfet_03v3
**devattr s=17600,576 d=10400,304
X898 a_9845_9634 SARlogic_0.dffrs_4.Q.t7 Vss.t158 Vss.t157 nfet_03v3
**devattr s=17600,576 d=10400,304
X899 a_37499_31160.t0 inv2_0.out.t28 Vdd.t926 Vdd.t925 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X900 Vss.t281 a_n10567_29019 a_n9673_28099 Vss.t280 nfet_03v3
**devattr s=10400,304 d=17600,576
X901 Vdd.t353 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_1.C Vdd.t352 pfet_03v3
**devattr s=26000,604 d=26000,604
X902 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t9 a_4501_23619 Vss.t650 nfet_03v3
**devattr s=10400,304 d=17600,576
X903 a_12401_23619 SARlogic_0.dffrs_4.Qb.t9 Vss.t191 Vss.t190 nfet_03v3
**devattr s=17600,576 d=10400,304
X904 a_13887_19210 SARlogic_0.d0.t12 Vss.t256 Vss.t255 nfet_03v3
**devattr s=17600,576 d=10400,304
X905 a_n389_31159.t2 inv2_0.out.t29 a_n201_30439 Vss.t665 nfet_03v3
**devattr s=10400,304 d=17600,576
X906 a_4841_29217.t0 a_4921_30169.t7 a_5105_31514 Vss.t140 nfet_03v3
**devattr s=10400,304 d=17600,576
X907 a_11311_29264.t0 a_10639_28100 Vss.t452 Vss.t451 nfet_03v3
**devattr s=17600,576 d=17600,576
X908 SARlogic_0.d5.t1 SARlogic_0.dffrs_14.Qb Vdd.t341 Vdd.t340 pfet_03v3
**devattr s=26000,604 d=44000,1176
X909 a_33521_31515 Clk_piso.t22 a_33337_31515 Vss.t187 nfet_03v3
**devattr s=10400,304 d=10400,304
X910 adc_PISO_0.dffrs_5.Qb adc_PISO_0.serial_out.t7 Vdd.t894 Vdd.t893 pfet_03v3
**devattr s=44000,1176 d=26000,604
X911 a_44479_31516 a_42729_29218.t7 a_44295_31516 Vss.t67 nfet_03v3
**devattr s=10400,304 d=10400,304
X912 Vdd.t295 a_n4551_30169.t7 a_n4631_33627.t2 Vdd.t294 pfet_03v3
**devattr s=26000,604 d=26000,604
X913 a_4841_31422.t0 Clk_piso.t23 a_5105_33719 Vss.t188 nfet_03v3
**devattr s=10400,304 d=17600,576
X914 a_6407_33719 Vdd.t996 Vss.t466 Vss.t465 nfet_03v3
**devattr s=17600,576 d=10400,304
X915 a_15879_31516 adc_PISO_0.dffrs_2.Q.t7 Vss.t46 Vss.t45 nfet_03v3
**devattr s=17600,576 d=10400,304
X916 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t10 a_n9933_n1136 a_n10021_n1044 Vss.t217 nfet_03v3
**devattr s=26400,776 d=15600,404
X917 adc_PISO_0.2inmux_0.OUT.t0 a_n7633_29263.t5 Vss.t566 Vss.t565 nfet_03v3
**devattr s=17600,576 d=17600,576
X918 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t10 a_12585_17004 Vss.t279 nfet_03v3
**devattr s=10400,304 d=17600,576
X919 a_36793_29020 inv2_0.out.t30 Vss.t667 Vss.t666 nfet_03v3
**devattr s=17600,576 d=17600,576
X920 Vdd.t748 a_n10831_4320 Comp_out.t4 Vdd.t747 pfet_03v3
**devattr s=18700,450 d=18700,450
X921 SARlogic_0.dffrs_4.nand3_1.C.t2 SARlogic_0.dffrs_4.nand3_6.C.t9 a_8543_14043 Vss.t66 nfet_03v3
**devattr s=10400,304 d=17600,576
X922 a_42809_30170.t3 adc_PISO_0.2inmux_1.OUT.t3 a_42993_29310 Vss.t603 nfet_03v3
**devattr s=10400,304 d=17600,576
X923 a_14577_29310 Vdd.t997 a_14393_29310 Vss.t464 nfet_03v3
**devattr s=10400,304 d=10400,304
X924 SARlogic_0.dffrs_11.nand3_8.C.t1 SARlogic_0.dffrs_11.nand3_8.Z a_12585_19209 Vss.t117 nfet_03v3
**devattr s=10400,304 d=17600,576
X925 a_4317_21414 SARlogic_0.dffrs_9.nand3_1.C Vss.t221 Vss.t220 nfet_03v3
**devattr s=17600,576 d=10400,304
X926 SARlogic_0.dffrs_0.d.t2 SARlogic_0.dffrs_13.Qb.t9 a_n10151_11838 Vss.t598 nfet_03v3
**devattr s=10400,304 d=17600,576
X927 a_39055_30440 a_37499_31160.t5 Vdd.t347 Vdd.t346 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X928 Vdd.t141 a_29583_30440 a_30443_29984 Vdd.t140 pfet_03v3
**devattr s=31200,704 d=52800,1376
X929 a_4501_17004 Reset.t80 a_4317_17004 Vss.t575 nfet_03v3
**devattr s=10400,304 d=10400,304
X930 a_18555_28820.t1 SARlogic_0.d2.t12 a_18743_28100 Vss.t241 nfet_03v3
**devattr s=10400,304 d=17600,576
X931 SARlogic_0.dffrs_14.Qb Reset.t81 a_n6139_19213 Vss.t576 nfet_03v3
**devattr s=10400,304 d=17600,576
X932 a_n11821_9633 SARlogic_0.dffrs_13.nand3_6.C.t9 Vss.t602 Vss.t601 nfet_03v3
**devattr s=17600,576 d=10400,304
X933 SARlogic_0.dffrs_5.nand3_1.C.t1 SARlogic_0.dffrs_5.nand3_6.C.t8 Vdd.t746 Vdd.t745 pfet_03v3
**devattr s=26000,604 d=44000,1176
X934 a_4317_23619 SARlogic_0.dffrs_2.Qb.t9 Vss.t593 Vss.t592 nfet_03v3
**devattr s=17600,576 d=10400,304
X935 adc_PISO_0.2inmux_1.Bit.t2 adc_PISO_0.dffrs_4.Qb Vdd.t605 Vdd.t604 pfet_03v3
**devattr s=26000,604 d=44000,1176
X936 a_n9673_30439 inv2_0.out.t31 a_n9861_31159.t0 Vss.t668 nfet_03v3
**devattr s=17600,576 d=10400,304
X937 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t17 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t8 Vss.t669 nfet_03v3
**devattr s=20800,504 d=20800,504
X938 a_4501_19209 SARlogic_0.d1.t12 a_4317_19209 Vss.t432 nfet_03v3
**devattr s=10400,304 d=10400,304
X939 SARlogic_0.dffrs_5.Q.t0 SARlogic_0.dffrs_5.Qb.t9 a_14071_11838 Vss.t619 nfet_03v3
**devattr s=10400,304 d=17600,576
X940 a_n3767_11838 SARlogic_0.dffrs_1.nand3_1.C.t5 Vss.t398 Vss.t397 nfet_03v3
**devattr s=17600,576 d=10400,304
X941 Vdd.t537 SARlogic_0.dffrs_3.nand3_8.Z.t7 SARlogic_0.dffrs_3.nand3_1.C.t0 Vdd.t536 pfet_03v3
**devattr s=26000,604 d=26000,604
X942 a_42809_31515 a_42729_31423.t9 Vss.t166 Vss.t165 nfet_03v3
**devattr s=17600,576 d=10400,304
X943 a_14071_11838 SARlogic_0.dffrs_5.nand3_6.C.t9 a_13887_11838 Vss.t535 nfet_03v3
**devattr s=10400,304 d=10400,304
X944 Vss.t48 adc_PISO_0.dffrs_2.Q.t8 a_18743_30440 Vss.t47 nfet_03v3
**devattr s=10400,304 d=17600,576
X945 a_5105_29309 Vdd.t998 a_4921_29309 Vss.t463 nfet_03v3
**devattr s=10400,304 d=10400,304
X946 Vdd.t297 SARlogic_0.dffrs_12.nand3_6.C.t9 SARlogic_0.dffrs_12.Q.t0 Vdd.t296 pfet_03v3
**devattr s=26000,604 d=26000,604
X947 SARlogic_0.dffrs_13.nand3_8.Z.t2 Vss.t690 Vdd.t17 Vdd.t16 pfet_03v3
**devattr s=26000,604 d=44000,1176
X948 a_8359_14043 Vdd.t999 Vss.t462 Vss.t461 nfet_03v3
**devattr s=17600,576 d=10400,304
X949 a_4921_29309 a_4841_29217.t7 Vss.t243 Vss.t242 nfet_03v3
**devattr s=17600,576 d=10400,304
X950 SARlogic_0.dffrs_12.nand3_6.C.t1 Vss.t691 Vdd.t19 Vdd.t18 pfet_03v3
**devattr s=26000,604 d=44000,1176
X951 a_4501_9633 Clk.t32 a_4317_9633 Vss.t6 nfet_03v3
**devattr s=10400,304 d=10400,304
X952 a_9083_28820.t2 SARlogic_0.d3.t12 Vdd.t97 Vdd.t96 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X953 Vdd.t165 SARlogic_0.d4.t12 SARlogic_0.dffrs_14.nand3_8.C.t2 Vdd.t164 pfet_03v3
**devattr s=26000,604 d=26000,604
X954 Vdd.t852 adc_PISO_0.dffrs_1.Q.t8 a_9083_31160.t3 Vdd.t851 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X955 Vss.t90 Vss.t88 a_n9673_30439 Vss.t89 nfet_03v3
**devattr s=10400,304 d=17600,576
X956 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t11 Vdd.t363 Vdd.t362 pfet_03v3
**devattr s=26000,604 d=44000,1176
R0 SARlogic_0.d3.n3 SARlogic_0.d3.t8 41.0041
R1 SARlogic_0.d3.n4 SARlogic_0.d3.t4 40.8177
R2 SARlogic_0.d3.n7 SARlogic_0.d3.t7 40.6313
R3 SARlogic_0.d3.n1 SARlogic_0.d3.t12 34.2529
R4 SARlogic_0.d3.n6 SARlogic_0.dffrs_7.clk 33.3108
R5 SARlogic_0.d3.n7 SARlogic_0.d3.t5 27.3166
R6 SARlogic_0.d3.n4 SARlogic_0.d3.t10 27.1302
R7 SARlogic_0.d3.n3 SARlogic_0.d3.t9 26.9438
R8 SARlogic_0.d3.n0 SARlogic_0.d3.t6 19.673
R9 SARlogic_0.d3.n0 SARlogic_0.d3.t11 19.4007
R10 SARlogic_0.d3.n9 SARlogic_0.d3.n8 14.0582
R11 SARlogic_0.d3.n9 SARlogic_0.d3.n6 11.1633
R12 SARlogic_0.d3 SARlogic_0.d3.n2 10.6816
R13 SARlogic_0.d3.n12 SARlogic_0.d3.t2 10.0473
R14 SARlogic_0.d3.n2 SARlogic_0.d3.n1 8.05164
R15 SARlogic_0.d3.n11 SARlogic_0.d3.t1 6.51042
R16 SARlogic_0.d3.n11 SARlogic_0.d3.n10 6.04952
R17 SARlogic_0.dffrs_7.nand3_1.A SARlogic_0.d3.n3 5.7755
R18 SARlogic_0.dffrs_7.nand3_6.B SARlogic_0.d3.n4 5.47979
R19 SARlogic_0.d3.n8 SARlogic_0.d3.n7 5.13907
R20 SARlogic_0.dffrs_8.nand3_2.Z SARlogic_0.d3.n12 4.72925
R21 SARlogic_0.d3.n5 SARlogic_0.dffrs_7.nand3_6.B 2.17818
R22 SARlogic_0.d3.n6 SARlogic_0.d3 1.54657
R23 SARlogic_0.d3.n5 SARlogic_0.dffrs_7.nand3_1.A 1.34729
R24 SARlogic_0.d3.n12 SARlogic_0.d3.n11 0.732092
R25 SARlogic_0.d3.n10 SARlogic_0.d3.t0 0.7285
R26 SARlogic_0.d3.n10 SARlogic_0.d3.t3 0.7285
R27 SARlogic_0.dffrs_7.clk SARlogic_0.d3.n5 0.610571
R28 SARlogic_0.dffrs_8.nand3_2.Z SARlogic_0.d3.n9 0.166901
R29 SARlogic_0.d3.n1 SARlogic_0.d3.n0 0.106438
R30 SARlogic_0.d3.n8 SARlogic_0.dffrs_8.nand3_7.C 0.0455
R31 SARlogic_0.d3.n2 adc_PISO_0.2inmux_3.In 0.0455
R32 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t6 40.8177
R33 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t5 40.6313
R34 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t7 27.3166
R35 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t4 27.1302
R36 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_8.C.n2 14.119
R37 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.t2 10.0473
R38 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.t1 6.51042
R39 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.n4 6.04952
R40 SARlogic_0.dffrs_7.nand3_7.B SARlogic_0.dffrs_7.nand3_8.C.n0 5.47979
R41 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C.n1 5.13907
R42 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n6 4.72925
R43 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.n5 0.732092
R44 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t0 0.7285
R45 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t3 0.7285
R46 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_7.B 0.438233
R47 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n3 0.166901
R48 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C 0.0455
R49 Vdd.n1033 Vdd.t574 869.717
R50 Vdd.n1022 Vdd.t929 869.717
R51 Vdd.t448 Vdd.t492 490.324
R52 Vdd.t927 Vdd.t448 490.324
R53 Vdd.t566 Vdd.t927 490.324
R54 Vdd.t572 Vdd.t566 490.324
R55 Vdd.t444 Vdd.t572 490.324
R56 Vdd.t446 Vdd.t444 490.324
R57 Vdd.t568 Vdd.t446 490.324
R58 Vdd.t570 Vdd.t568 490.324
R59 Vdd.t312 Vdd.t570 490.324
R60 Vdd.t492 Vdd.n1069 467.743
R61 Vdd.n1071 Vdd.t312 467.743
R62 Vdd.n1072 Vdd.t56 398.652
R63 Vdd.n1054 Vdd.t66 398.652
R64 Vdd.t56 Vdd.n1071 389.878
R65 Vdd.n1069 Vdd.t66 389.878
R66 Vdd.t594 Vdd.n1026 372.543
R67 Vdd.n1029 Vdd.t330 372.543
R68 Vdd.n1028 Vdd.t594 370.969
R69 Vdd.t330 Vdd.n1028 370.969
R70 Vdd.n1049 Vdd.n1047 287.351
R71 Vdd.n1050 Vdd.n1048 287.351
R72 Vdd.t749 Vdd.t747 265.625
R73 Vdd.t546 Vdd.t542 265.625
R74 Vdd.t238 Vdd.n4 250.9
R75 Vdd.n5 Vdd.t676 250.9
R76 Vdd.t879 Vdd.n1108 250.9
R77 Vdd.n1109 Vdd.t220 250.9
R78 Vdd.t336 Vdd.n9 250.9
R79 Vdd.n10 Vdd.t697 250.9
R80 Vdd.t837 Vdd.n1096 250.9
R81 Vdd.n1097 Vdd.t236 250.9
R82 Vdd.t670 Vdd.n1102 250.9
R83 Vdd.n1103 Vdd.t590 250.9
R84 Vdd.t827 Vdd.n1089 250.9
R85 Vdd.n1090 Vdd.t216 250.9
R86 Vdd.t174 Vdd.n63 250.9
R87 Vdd.n64 Vdd.t724 250.9
R88 Vdd.t861 Vdd.n75 250.9
R89 Vdd.n76 Vdd.t192 250.9
R90 Vdd.t512 Vdd.n70 250.9
R91 Vdd.n71 Vdd.t613 250.9
R92 Vdd.t895 Vdd.n87 250.9
R93 Vdd.n88 Vdd.t178 250.9
R94 Vdd.t652 Vdd.n81 250.9
R95 Vdd.n82 Vdd.t893 250.9
R96 Vdd.t833 Vdd.n98 250.9
R97 Vdd.n99 Vdd.t114 250.9
R98 Vdd.t524 Vdd.n137 250.9
R99 Vdd.n138 Vdd.t703 250.9
R100 Vdd.t875 Vdd.n148 250.9
R101 Vdd.n149 Vdd.t819 250.9
R102 Vdd.t604 Vdd.n143 250.9
R103 Vdd.n144 Vdd.t715 250.9
R104 Vdd.t510 Vdd.n160 250.9
R105 Vdd.n161 Vdd.t528 250.9
R106 Vdd.t739 Vdd.n154 250.9
R107 Vdd.n155 Vdd.t452 250.9
R108 Vdd.t500 Vdd.n171 250.9
R109 Vdd.n172 Vdd.t809 250.9
R110 Vdd.t480 Vdd.n217 250.9
R111 Vdd.n218 Vdd.t634 250.9
R112 Vdd.t655 Vdd.n222 250.9
R113 Vdd.n223 Vdd.t84 250.9
R114 Vdd.t342 Vdd.n211 250.9
R115 Vdd.n212 Vdd.t845 250.9
R116 Vdd.t18 Vdd.n1014 250.9
R117 Vdd.n1015 Vdd.t883 250.9
R118 Vdd.t152 Vdd.n997 250.9
R119 Vdd.n998 Vdd.t847 250.9
R120 Vdd.t20 Vdd.n1002 250.9
R121 Vdd.n1003 Vdd.t344 250.9
R122 Vdd.t394 Vdd.n1008 250.9
R123 Vdd.n1009 Vdd.t558 250.9
R124 Vdd.t10 Vdd.n990 250.9
R125 Vdd.n991 Vdd.t490 250.9
R126 Vdd.t855 Vdd.n518 250.9
R127 Vdd.n519 Vdd.t619 250.9
R128 Vdd.t272 Vdd.n524 250.9
R129 Vdd.n525 Vdd.t488 250.9
R130 Vdd.t328 Vdd.n530 250.9
R131 Vdd.n531 Vdd.t857 250.9
R132 Vdd.t266 Vdd.n981 250.9
R133 Vdd.n982 Vdd.t332 250.9
R134 Vdd.t378 Vdd.n767 250.9
R135 Vdd.n768 Vdd.t813 250.9
R136 Vdd.t302 Vdd.n806 250.9
R137 Vdd.n807 Vdd.t232 250.9
R138 Vdd.t86 Vdd.n844 250.9
R139 Vdd.n845 Vdd.t370 250.9
R140 Vdd.t905 Vdd.n882 250.9
R141 Vdd.n883 Vdd.t518 250.9
R142 Vdd.t286 Vdd.n921 250.9
R143 Vdd.n922 Vdd.t168 250.9
R144 Vdd.t80 Vdd.n959 250.9
R145 Vdd.n960 Vdd.t254 250.9
R146 Vdd.t162 Vdd.n685 250.9
R147 Vdd.n686 Vdd.t468 250.9
R148 Vdd.t340 Vdd.n778 250.9
R149 Vdd.n779 Vdd.t817 250.9
R150 Vdd.t98 Vdd.n411 250.9
R151 Vdd.n412 Vdd.t454 250.9
R152 Vdd.t264 Vdd.n817 250.9
R153 Vdd.n818 Vdd.t228 250.9
R154 Vdd.t306 Vdd.n381 250.9
R155 Vdd.n382 Vdd.t128 250.9
R156 Vdd.t130 Vdd.n855 250.9
R157 Vdd.n856 Vdd.t368 250.9
R158 Vdd.t564 Vdd.n351 250.9
R159 Vdd.n352 Vdd.t284 250.9
R160 Vdd.t821 Vdd.n894 250.9
R161 Vdd.n895 Vdd.t516 250.9
R162 Vdd.t943 Vdd.n315 250.9
R163 Vdd.n316 Vdd.t122 250.9
R164 Vdd.t126 Vdd.n932 250.9
R165 Vdd.n933 Vdd.t166 250.9
R166 Vdd.t556 Vdd.n285 250.9
R167 Vdd.n286 Vdd.t242 250.9
R168 Vdd.t244 Vdd.n970 250.9
R169 Vdd.n971 Vdd.t256 250.9
R170 Vdd.t24 Vdd.n762 250.9
R171 Vdd.n763 Vdd.t380 250.9
R172 Vdd.t434 Vdd.n675 250.9
R173 Vdd.n676 Vdd.t298 250.9
R174 Vdd.t278 Vdd.n801 250.9
R175 Vdd.n802 Vdd.t578 250.9
R176 Vdd.t414 Vdd.n401 250.9
R177 Vdd.n402 Vdd.t889 250.9
R178 Vdd.t324 Vdd.n839 250.9
R179 Vdd.n840 Vdd.t90 250.9
R180 Vdd.t396 Vdd.n371 250.9
R181 Vdd.n372 Vdd.t100 250.9
R182 Vdd.t156 Vdd.n877 250.9
R183 Vdd.n878 Vdd.t903 250.9
R184 Vdd.t400 Vdd.n335 250.9
R185 Vdd.n336 Vdd.t304 250.9
R186 Vdd.t354 Vdd.n916 250.9
R187 Vdd.n917 Vdd.t290 250.9
R188 Vdd.t390 Vdd.n305 250.9
R189 Vdd.n306 Vdd.t562 250.9
R190 Vdd.t172 Vdd.n954 250.9
R191 Vdd.n955 Vdd.t76 250.9
R192 Vdd.t783 Vdd.n275 250.9
R193 Vdd.n276 Vdd.t945 250.9
R194 Vdd.t362 Vdd.n690 250.9
R195 Vdd.n691 Vdd.t350 250.9
R196 Vdd.t356 Vdd.n416 250.9
R197 Vdd.n417 Vdd.t184 250.9
R198 Vdd.t260 Vdd.n386 250.9
R199 Vdd.n387 Vdd.t186 250.9
R200 Vdd.t360 Vdd.n356 250.9
R201 Vdd.n357 Vdd.t588 250.9
R202 Vdd.t258 Vdd.n320 250.9
R203 Vdd.n321 Vdd.t318 250.9
R204 Vdd.t358 Vdd.n290 250.9
R205 Vdd.n291 Vdd.t252 250.9
R206 Vdd.t34 Vdd.n757 250.9
R207 Vdd.n758 Vdd.t709 250.9
R208 Vdd.t46 Vdd.n695 250.9
R209 Vdd.n696 Vdd.t366 250.9
R210 Vdd.t148 Vdd.n796 250.9
R211 Vdd.n797 Vdd.t616 250.9
R212 Vdd.t230 Vdd.n773 250.9
R213 Vdd.n774 Vdd.t700 250.9
R214 Vdd.t2 Vdd.n421 250.9
R215 Vdd.n422 Vdd.t871 250.9
R216 Vdd.t498 Vdd.n834 250.9
R217 Vdd.n835 Vdd.t664 250.9
R218 Vdd.t372 Vdd.n812 250.9
R219 Vdd.n813 Vdd.t658 250.9
R220 Vdd.t60 Vdd.n391 250.9
R221 Vdd.n392 Vdd.t70 250.9
R222 Vdd.t384 Vdd.n872 250.9
R223 Vdd.n873 Vdd.t712 250.9
R224 Vdd.t839 Vdd.n850 250.9
R225 Vdd.n851 Vdd.t682 250.9
R226 Vdd.t42 Vdd.n361 250.9
R227 Vdd.n362 Vdd.t222 250.9
R228 Vdd.t110 Vdd.n911 250.9
R229 Vdd.n912 Vdd.t673 250.9
R230 Vdd.t180 Vdd.n889 250.9
R231 Vdd.n890 Vdd.t730 250.9
R232 Vdd.t54 Vdd.n325 250.9
R233 Vdd.n326 Vdd.t486 250.9
R234 Vdd.t745 Vdd.n949 250.9
R235 Vdd.n950 Vdd.t718 250.9
R236 Vdd.t941 Vdd.n927 250.9
R237 Vdd.n928 Vdd.t679 250.9
R238 Vdd.t6 Vdd.n295 250.9
R239 Vdd.n296 Vdd.t829 250.9
R240 Vdd.t849 Vdd.n965 250.9
R241 Vdd.n966 Vdd.t694 250.9
R242 Vdd.t124 Vdd.n752 250.9
R243 Vdd.n753 Vdd.t32 250.9
R244 Vdd.t404 Vdd.n680 250.9
R245 Vdd.n681 Vdd.t194 250.9
R246 Vdd.t212 Vdd.n791 250.9
R247 Vdd.n792 Vdd.t146 250.9
R248 Vdd.t416 Vdd.n406 250.9
R249 Vdd.n407 Vdd.t40 250.9
R250 Vdd.t268 Vdd.n829 250.9
R251 Vdd.n830 Vdd.t494 250.9
R252 Vdd.t785 Vdd.n376 250.9
R253 Vdd.n377 Vdd.t476 250.9
R254 Vdd.t534 Vdd.n867 250.9
R255 Vdd.n868 Vdd.t382 250.9
R256 Vdd.t789 Vdd.n340 250.9
R257 Vdd.n341 Vdd.t540 250.9
R258 Vdd.t484 Vdd.n906 250.9
R259 Vdd.n907 Vdd.t108 250.9
R260 Vdd.t781 Vdd.n310 250.9
R261 Vdd.n311 Vdd.t226 250.9
R262 Vdd.t206 Vdd.n944 250.9
R263 Vdd.n945 Vdd.t741 250.9
R264 Vdd.t420 Vdd.n280 250.9
R265 Vdd.n281 Vdd.t464 250.9
R266 Vdd.t825 Vdd.n700 250.9
R267 Vdd.n701 Vdd.t104 250.9
R268 Vdd.t773 Vdd.n426 250.9
R269 Vdd.n427 Vdd.t532 250.9
R270 Vdd.t38 Vdd.n396 250.9
R271 Vdd.n397 Vdd.t917 250.9
R272 Vdd.t478 Vdd.n366 250.9
R273 Vdd.n367 Vdd.t520 250.9
R274 Vdd.t538 Vdd.n330 250.9
R275 Vdd.n331 Vdd.t456 250.9
R276 Vdd.t224 Vdd.n300 250.9
R277 Vdd.n301 Vdd.t462 250.9
R278 Vdd.t953 Vdd.n705 250.9
R279 Vdd.n706 Vdd.t779 250.9
R280 Vdd.t68 Vdd.n721 250.9
R281 Vdd.n722 Vdd.t602 250.9
R282 Vdd.t815 Vdd.n716 250.9
R283 Vdd.n717 Vdd.t777 250.9
R284 Vdd.t92 Vdd.n739 250.9
R285 Vdd.n740 Vdd.t951 250.9
R286 Vdd.t727 Vdd.n745 250.9
R287 Vdd.n746 Vdd.t823 250.9
R288 Vdd.t16 Vdd.n733 250.9
R289 Vdd.n734 Vdd.t30 250.9
R290 Vdd.t935 Vdd.n638 250.9
R291 Vdd.n639 Vdd.t622 250.9
R292 Vdd.t274 Vdd.n649 250.9
R293 Vdd.n650 Vdd.t582 250.9
R294 Vdd.t0 Vdd.n644 250.9
R295 Vdd.n645 Vdd.t661 250.9
R296 Vdd.t292 Vdd.n661 250.9
R297 Vdd.n662 Vdd.t931 250.9
R298 Vdd.t736 Vdd.n655 250.9
R299 Vdd.n656 Vdd.t74 250.9
R300 Vdd.t198 Vdd.n668 250.9
R301 Vdd.n669 Vdd.t550 250.9
R302 Vdd.t470 Vdd.n569 250.9
R303 Vdd.n570 Vdd.t607 250.9
R304 Vdd.t937 Vdd.n580 250.9
R305 Vdd.n581 Vdd.t504 250.9
R306 Vdd.t158 Vdd.n575 250.9
R307 Vdd.n576 Vdd.t628 250.9
R308 Vdd.t913 Vdd.n592 250.9
R309 Vdd.n593 Vdd.t474 250.9
R310 Vdd.t637 Vdd.n586 250.9
R311 Vdd.n587 Vdd.t843 250.9
R312 Vdd.t214 Vdd.n599 250.9
R313 Vdd.n600 Vdd.t314 250.9
R314 Vdd.n1040 Vdd.t596 242.189
R315 Vdd.t891 Vdd.n59 242.189
R316 Vdd.n199 Vdd.t811 236.083
R317 Vdd.t765 Vdd.n196 236.083
R318 Vdd.t466 Vdd.n179 236.083
R319 Vdd.n185 Vdd.t584 236.083
R320 Vdd.n126 Vdd.t346 236.083
R321 Vdd.t925 Vdd.n123 236.083
R322 Vdd.t502 Vdd.n106 236.083
R323 Vdd.n112 Vdd.t947 236.083
R324 Vdd.n45 Vdd.t841 236.083
R325 Vdd.n39 Vdd.t899 236.083
R326 Vdd.n29 Vdd.t338 236.083
R327 Vdd.n23 Vdd.t142 236.083
R328 Vdd.t204 Vdd.n244 236.083
R329 Vdd.n250 Vdd.t308 236.083
R330 Vdd.n627 Vdd.t106 236.083
R331 Vdd.t761 Vdd.n624 236.083
R332 Vdd.t592 Vdd.n607 236.083
R333 Vdd.n613 Vdd.t160 236.083
R334 Vdd.n558 Vdd.t805 236.083
R335 Vdd.t763 Vdd.n555 236.083
R336 Vdd.t911 Vdd.n538 236.083
R337 Vdd.n544 Vdd.t96 236.083
R338 Vdd.n512 Vdd.t208 236.083
R339 Vdd.n506 Vdd.t885 236.083
R340 Vdd.n496 Vdd.t234 236.083
R341 Vdd.n490 Vdd.t134 236.083
R342 Vdd.t514 Vdd.n466 236.083
R343 Vdd.n472 Vdd.t300 236.083
R344 Vdd.t190 Vdd.n448 236.083
R345 Vdd.n458 Vdd.t923 236.083
R346 Vdd.t775 Vdd.n435 236.083
R347 Vdd.n446 Vdd.t138 236.083
R348 Vdd.t801 Vdd.n260 236.083
R349 Vdd.n264 Vdd.t771 236.083
R350 Vdd.t576 Vdd.n234 236.083
R351 Vdd.n236 Vdd.t118 236.083
R352 Vdd.t811 Vdd.n198 235.294
R353 Vdd.n198 Vdd.t765 235.294
R354 Vdd.n184 Vdd.t466 235.294
R355 Vdd.t584 Vdd.n184 235.294
R356 Vdd.t346 Vdd.n125 235.294
R357 Vdd.n125 Vdd.t925 235.294
R358 Vdd.n111 Vdd.t502 235.294
R359 Vdd.t947 Vdd.n111 235.294
R360 Vdd.t841 Vdd.n44 235.294
R361 Vdd.n44 Vdd.t281 235.294
R362 Vdd.t280 Vdd.n42 235.294
R363 Vdd.n42 Vdd.t901 235.294
R364 Vdd.t338 Vdd.n28 235.294
R365 Vdd.n28 Vdd.t249 235.294
R366 Vdd.t248 Vdd.n26 235.294
R367 Vdd.n26 Vdd.t140 235.294
R368 Vdd.n249 Vdd.t204 235.294
R369 Vdd.t308 Vdd.n249 235.294
R370 Vdd.t106 Vdd.n626 235.294
R371 Vdd.n626 Vdd.t761 235.294
R372 Vdd.n612 Vdd.t592 235.294
R373 Vdd.t160 Vdd.n612 235.294
R374 Vdd.t805 Vdd.n557 235.294
R375 Vdd.n557 Vdd.t763 235.294
R376 Vdd.n543 Vdd.t911 235.294
R377 Vdd.t96 Vdd.n543 235.294
R378 Vdd.t208 Vdd.n511 235.294
R379 Vdd.n511 Vdd.t598 235.294
R380 Vdd.t599 Vdd.n509 235.294
R381 Vdd.n509 Vdd.t887 235.294
R382 Vdd.t234 Vdd.n495 235.294
R383 Vdd.n495 Vdd.t283 235.294
R384 Vdd.t282 Vdd.n493 235.294
R385 Vdd.n493 Vdd.t132 235.294
R386 Vdd.n471 Vdd.t514 235.294
R387 Vdd.t300 Vdd.n471 235.294
R388 Vdd.n457 Vdd.t190 235.294
R389 Vdd.t923 Vdd.n457 235.294
R390 Vdd.n443 Vdd.t775 235.294
R391 Vdd.t323 Vdd.n443 235.294
R392 Vdd.n445 Vdd.t322 235.294
R393 Vdd.t136 Vdd.n445 235.294
R394 Vdd.n263 Vdd.t801 235.294
R395 Vdd.t771 Vdd.n263 235.294
R396 Vdd.n240 Vdd.t576 235.294
R397 Vdd.n240 Vdd.t28 235.294
R398 Vdd.t29 Vdd.n239 235.294
R399 Vdd.n239 Vdd.t120 235.294
R400 Vdd.t835 Vdd.t238 200
R401 Vdd.t676 Vdd.t835 200
R402 Vdd.t667 Vdd.t879 200
R403 Vdd.t220 Vdd.t667 200
R404 Vdd.t240 Vdd.t336 200
R405 Vdd.t697 Vdd.t240 200
R406 Vdd.t877 Vdd.t837 200
R407 Vdd.t236 Vdd.t877 200
R408 Vdd.t218 Vdd.t670 200
R409 Vdd.t590 Vdd.t218 200
R410 Vdd.t706 Vdd.t827 200
R411 Vdd.t216 Vdd.t706 200
R412 Vdd.t897 Vdd.t174 200
R413 Vdd.t724 Vdd.t897 200
R414 Vdd.t610 Vdd.t861 200
R415 Vdd.t192 Vdd.t610 200
R416 Vdd.t176 Vdd.t512 200
R417 Vdd.t613 Vdd.t176 200
R418 Vdd.t865 Vdd.t895 200
R419 Vdd.t178 Vdd.t865 200
R420 Vdd.t831 Vdd.t652 200
R421 Vdd.t893 Vdd.t831 200
R422 Vdd.t646 Vdd.t833 200
R423 Vdd.t114 Vdd.t646 200
R424 Vdd.t281 Vdd.t280 200
R425 Vdd.t899 Vdd.t901 200
R426 Vdd.t508 Vdd.t524 200
R427 Vdd.t703 Vdd.t508 200
R428 Vdd.t733 Vdd.t875 200
R429 Vdd.t819 Vdd.t733 200
R430 Vdd.t526 Vdd.t604 200
R431 Vdd.t715 Vdd.t526 200
R432 Vdd.t869 Vdd.t510 200
R433 Vdd.t528 Vdd.t869 200
R434 Vdd.t807 Vdd.t739 200
R435 Vdd.t452 Vdd.t807 200
R436 Vdd.t631 Vdd.t500 200
R437 Vdd.t809 Vdd.t631 200
R438 Vdd.t249 Vdd.t248 200
R439 Vdd.t142 Vdd.t140 200
R440 Vdd.t859 Vdd.t480 200
R441 Vdd.t634 Vdd.t859 200
R442 Vdd.t334 Vdd.t655 200
R443 Vdd.t84 Vdd.t334 200
R444 Vdd.t22 Vdd.t342 200
R445 Vdd.t845 Vdd.t22 200
R446 Vdd.t426 Vdd.t18 200
R447 Vdd.t883 Vdd.t426 200
R448 Vdd.t296 Vdd.t152 200
R449 Vdd.t847 Vdd.t296 200
R450 Vdd.t14 Vdd.t20 200
R451 Vdd.t344 Vdd.t14 200
R452 Vdd.t939 Vdd.t394 200
R453 Vdd.t558 Vdd.t939 200
R454 Vdd.t430 Vdd.t10 200
R455 Vdd.t490 Vdd.t430 200
R456 Vdd.t909 Vdd.t855 200
R457 Vdd.t619 Vdd.t909 200
R458 Vdd.t649 Vdd.t272 200
R459 Vdd.t488 Vdd.t649 200
R460 Vdd.t881 Vdd.t328 200
R461 Vdd.t857 Vdd.t881 200
R462 Vdd.t691 Vdd.t266 200
R463 Vdd.t332 Vdd.t691 200
R464 Vdd.t26 Vdd.t378 200
R465 Vdd.t813 Vdd.t26 200
R466 Vdd.t276 Vdd.t302 200
R467 Vdd.t232 Vdd.t276 200
R468 Vdd.t326 Vdd.t86 200
R469 Vdd.t370 Vdd.t326 200
R470 Vdd.t154 Vdd.t905 200
R471 Vdd.t518 Vdd.t154 200
R472 Vdd.t352 Vdd.t286 200
R473 Vdd.t168 Vdd.t352 200
R474 Vdd.t170 Vdd.t80 200
R475 Vdd.t254 Vdd.t170 200
R476 Vdd.t506 Vdd.t162 200
R477 Vdd.t468 Vdd.t506 200
R478 Vdd.t376 Vdd.t340 200
R479 Vdd.t817 Vdd.t376 200
R480 Vdd.t438 Vdd.t98 200
R481 Vdd.t454 Vdd.t438 200
R482 Vdd.t580 Vdd.t264 200
R483 Vdd.t228 Vdd.t580 200
R484 Vdd.t428 Vdd.t306 200
R485 Vdd.t128 Vdd.t428 200
R486 Vdd.t88 Vdd.t130 200
R487 Vdd.t368 Vdd.t88 200
R488 Vdd.t406 Vdd.t564 200
R489 Vdd.t284 Vdd.t406 200
R490 Vdd.t907 Vdd.t821 200
R491 Vdd.t516 Vdd.t907 200
R492 Vdd.t799 Vdd.t943 200
R493 Vdd.t122 Vdd.t799 200
R494 Vdd.t288 Vdd.t126 200
R495 Vdd.t166 Vdd.t288 200
R496 Vdd.t787 Vdd.t556 200
R497 Vdd.t242 Vdd.t787 200
R498 Vdd.t78 Vdd.t244 200
R499 Vdd.t256 Vdd.t78 200
R500 Vdd.t164 Vdd.t24 200
R501 Vdd.t380 Vdd.t164 200
R502 Vdd.t348 Vdd.t434 200
R503 Vdd.t298 Vdd.t348 200
R504 Vdd.t102 Vdd.t278 200
R505 Vdd.t578 Vdd.t102 200
R506 Vdd.t182 Vdd.t414 200
R507 Vdd.t889 Vdd.t182 200
R508 Vdd.t310 Vdd.t324 200
R509 Vdd.t90 Vdd.t310 200
R510 Vdd.t188 Vdd.t396 200
R511 Vdd.t100 Vdd.t188 200
R512 Vdd.t560 Vdd.t156 200
R513 Vdd.t903 Vdd.t560 200
R514 Vdd.t586 Vdd.t400 200
R515 Vdd.t304 Vdd.t586 200
R516 Vdd.t949 Vdd.t354 200
R517 Vdd.t290 Vdd.t949 200
R518 Vdd.t320 Vdd.t390 200
R519 Vdd.t562 Vdd.t320 200
R520 Vdd.t554 Vdd.t172 200
R521 Vdd.t76 Vdd.t554 200
R522 Vdd.t250 Vdd.t783 200
R523 Vdd.t945 Vdd.t250 200
R524 Vdd.t422 Vdd.t362 200
R525 Vdd.t350 Vdd.t422 200
R526 Vdd.t392 Vdd.t356 200
R527 Vdd.t184 Vdd.t392 200
R528 Vdd.t442 Vdd.t260 200
R529 Vdd.t186 Vdd.t442 200
R530 Vdd.t412 Vdd.t360 200
R531 Vdd.t588 Vdd.t412 200
R532 Vdd.t418 Vdd.t258 200
R533 Vdd.t318 Vdd.t418 200
R534 Vdd.t795 Vdd.t358 200
R535 Vdd.t252 Vdd.t795 200
R536 Vdd.t116 Vdd.t34 200
R537 Vdd.t709 Vdd.t116 200
R538 Vdd.t440 Vdd.t46 200
R539 Vdd.t366 Vdd.t440 200
R540 Vdd.t210 Vdd.t148 200
R541 Vdd.t616 Vdd.t210 200
R542 Vdd.t36 Vdd.t230 200
R543 Vdd.t700 Vdd.t36 200
R544 Vdd.t410 Vdd.t2 200
R545 Vdd.t871 Vdd.t410 200
R546 Vdd.t270 Vdd.t498 200
R547 Vdd.t664 Vdd.t270 200
R548 Vdd.t144 Vdd.t372 200
R549 Vdd.t658 Vdd.t144 200
R550 Vdd.t402 Vdd.t60 200
R551 Vdd.t70 Vdd.t402 200
R552 Vdd.t536 Vdd.t384 200
R553 Vdd.t712 Vdd.t536 200
R554 Vdd.t496 Vdd.t839 200
R555 Vdd.t682 Vdd.t496 200
R556 Vdd.t797 Vdd.t42 200
R557 Vdd.t222 Vdd.t797 200
R558 Vdd.t482 Vdd.t110 200
R559 Vdd.t673 Vdd.t482 200
R560 Vdd.t386 Vdd.t180 200
R561 Vdd.t730 Vdd.t386 200
R562 Vdd.t432 Vdd.t54 200
R563 Vdd.t486 Vdd.t432 200
R564 Vdd.t803 Vdd.t745 200
R565 Vdd.t718 Vdd.t803 200
R566 Vdd.t112 Vdd.t941 200
R567 Vdd.t679 Vdd.t112 200
R568 Vdd.t424 Vdd.t6 200
R569 Vdd.t829 Vdd.t424 200
R570 Vdd.t743 Vdd.t849 200
R571 Vdd.t694 Vdd.t743 200
R572 Vdd.t50 Vdd.t124 200
R573 Vdd.t32 Vdd.t50 200
R574 Vdd.t82 Vdd.t404 200
R575 Vdd.t194 Vdd.t82 200
R576 Vdd.t64 Vdd.t212 200
R577 Vdd.t146 Vdd.t64 200
R578 Vdd.t530 Vdd.t416 200
R579 Vdd.t40 Vdd.t530 200
R580 Vdd.t62 Vdd.t268 200
R581 Vdd.t494 Vdd.t62 200
R582 Vdd.t915 Vdd.t785 200
R583 Vdd.t476 Vdd.t915 200
R584 Vdd.t8 Vdd.t534 200
R585 Vdd.t382 Vdd.t8 200
R586 Vdd.t522 Vdd.t789 200
R587 Vdd.t540 Vdd.t522 200
R588 Vdd.t48 Vdd.t484 200
R589 Vdd.t108 Vdd.t48 200
R590 Vdd.t458 Vdd.t781 200
R591 Vdd.t226 Vdd.t458 200
R592 Vdd.t44 Vdd.t206 200
R593 Vdd.t741 Vdd.t44 200
R594 Vdd.t460 Vdd.t420 200
R595 Vdd.t464 Vdd.t460 200
R596 Vdd.t436 Vdd.t825 200
R597 Vdd.t104 Vdd.t436 200
R598 Vdd.t408 Vdd.t773 200
R599 Vdd.t532 Vdd.t408 200
R600 Vdd.t793 Vdd.t38 200
R601 Vdd.t917 Vdd.t793 200
R602 Vdd.t398 Vdd.t478 200
R603 Vdd.t520 Vdd.t398 200
R604 Vdd.t388 Vdd.t538 200
R605 Vdd.t456 Vdd.t388 200
R606 Vdd.t791 Vdd.t224 200
R607 Vdd.t462 Vdd.t791 200
R608 Vdd.t94 Vdd.t953 200
R609 Vdd.t779 Vdd.t94 200
R610 Vdd.t625 Vdd.t68 200
R611 Vdd.t602 Vdd.t625 200
R612 Vdd.t853 Vdd.t815 200
R613 Vdd.t777 Vdd.t853 200
R614 Vdd.t4 Vdd.t92 200
R615 Vdd.t951 Vdd.t4 200
R616 Vdd.t202 Vdd.t727 200
R617 Vdd.t823 Vdd.t202 200
R618 Vdd.t721 Vdd.t16 200
R619 Vdd.t30 Vdd.t721 200
R620 Vdd.t294 Vdd.t935 200
R621 Vdd.t622 Vdd.t294 200
R622 Vdd.t640 Vdd.t274 200
R623 Vdd.t582 Vdd.t640 200
R624 Vdd.t933 Vdd.t0 200
R625 Vdd.t661 Vdd.t933 200
R626 Vdd.t867 Vdd.t292 200
R627 Vdd.t931 Vdd.t867 200
R628 Vdd.t552 Vdd.t736 200
R629 Vdd.t74 Vdd.t552 200
R630 Vdd.t685 Vdd.t198 200
R631 Vdd.t550 Vdd.t685 200
R632 Vdd.t200 Vdd.t470 200
R633 Vdd.t607 Vdd.t200 200
R634 Vdd.t643 Vdd.t937 200
R635 Vdd.t504 Vdd.t643 200
R636 Vdd.t472 Vdd.t158 200
R637 Vdd.t628 Vdd.t472 200
R638 Vdd.t863 Vdd.t913 200
R639 Vdd.t474 Vdd.t863 200
R640 Vdd.t316 Vdd.t637 200
R641 Vdd.t843 Vdd.t316 200
R642 Vdd.t688 Vdd.t214 200
R643 Vdd.t314 Vdd.t688 200
R644 Vdd.t598 Vdd.t599 200
R645 Vdd.t885 Vdd.t887 200
R646 Vdd.t283 Vdd.t282 200
R647 Vdd.t134 Vdd.t132 200
R648 Vdd.t322 Vdd.t323 200
R649 Vdd.t138 Vdd.t136 200
R650 Vdd.t28 Vdd.t29 200
R651 Vdd.t118 Vdd.t120 200
R652 Vdd.t753 Vdd.n1042 195.312
R653 Vdd.t548 Vdd.n55 195.312
R654 Vdd.n1076 Vdd.t58 190.464
R655 Vdd.n1052 Vdd.t52 190.464
R656 Vdd.n1043 Vdd.t753 179.689
R657 Vdd.n56 Vdd.t548 179.689
R658 Vdd.t596 Vdd.n1039 145.413
R659 Vdd.n60 Vdd.t891 145.413
R660 Vdd.n15 Vdd.t246 131.589
R661 Vdd.n187 Vdd.t196 131.589
R662 Vdd.n31 Vdd.t450 131.589
R663 Vdd.n114 Vdd.t262 131.589
R664 Vdd.n252 Vdd.t600 131.589
R665 Vdd.n266 Vdd.t873 131.589
R666 Vdd.n482 Vdd.t72 131.589
R667 Vdd.n615 Vdd.t755 131.589
R668 Vdd.n498 Vdd.t851 131.589
R669 Vdd.n546 Vdd.t150 131.589
R670 Vdd.n474 Vdd.t364 131.589
R671 Vdd.n460 Vdd.t12 131.589
R672 Vdd.n1019 Vdd.n272 130.231
R673 Vdd.n1019 Vdd.n995 121.085
R674 Vdd.n130 Vdd.t759 118.543
R675 Vdd.n203 Vdd.t921 118.543
R676 Vdd.n562 Vdd.t767 118.543
R677 Vdd.n631 Vdd.t919 118.543
R678 Vdd.n451 Vdd.t769 118.543
R679 Vdd.n268 Vdd.t757 118.543
R680 Vdd.n450 Vdd.t374 118.519
R681 Vdd.n272 Vdd.n271 117.481
R682 Vdd.n39 Vdd.n38 96.0755
R683 Vdd.n40 Vdd.n39 96.0755
R684 Vdd.n23 Vdd.n22 96.0755
R685 Vdd.n24 Vdd.n23 96.0755
R686 Vdd.n506 Vdd.n505 96.0755
R687 Vdd.n507 Vdd.n506 96.0755
R688 Vdd.n490 Vdd.n489 96.0755
R689 Vdd.n491 Vdd.n490 96.0755
R690 Vdd.n446 Vdd.n438 96.0755
R691 Vdd.n446 Vdd.n439 96.0755
R692 Vdd.n236 Vdd.n235 96.0755
R693 Vdd.n237 Vdd.n236 96.0755
R694 Vdd.n1043 Vdd.t749 85.938
R695 Vdd.n56 Vdd.t546 85.938
R696 Vdd.n181 Vdd.n179 78.2255
R697 Vdd.n185 Vdd.n181 78.2255
R698 Vdd.n185 Vdd.n182 78.2255
R699 Vdd.n182 Vdd.n179 78.2255
R700 Vdd.n108 Vdd.n106 78.2255
R701 Vdd.n112 Vdd.n108 78.2255
R702 Vdd.n112 Vdd.n109 78.2255
R703 Vdd.n109 Vdd.n106 78.2255
R704 Vdd.n45 Vdd.n36 78.2255
R705 Vdd.n45 Vdd.n37 78.2255
R706 Vdd.n126 Vdd.n121 78.2255
R707 Vdd.n126 Vdd.n122 78.2255
R708 Vdd.n123 Vdd.n121 78.2255
R709 Vdd.n123 Vdd.n122 78.2255
R710 Vdd.n29 Vdd.n20 78.2255
R711 Vdd.n29 Vdd.n21 78.2255
R712 Vdd.n199 Vdd.n194 78.2255
R713 Vdd.n199 Vdd.n195 78.2255
R714 Vdd.n196 Vdd.n194 78.2255
R715 Vdd.n196 Vdd.n195 78.2255
R716 Vdd.n246 Vdd.n244 78.2255
R717 Vdd.n250 Vdd.n246 78.2255
R718 Vdd.n250 Vdd.n247 78.2255
R719 Vdd.n247 Vdd.n244 78.2255
R720 Vdd.n609 Vdd.n607 78.2255
R721 Vdd.n613 Vdd.n609 78.2255
R722 Vdd.n613 Vdd.n610 78.2255
R723 Vdd.n610 Vdd.n607 78.2255
R724 Vdd.n540 Vdd.n538 78.2255
R725 Vdd.n544 Vdd.n540 78.2255
R726 Vdd.n544 Vdd.n541 78.2255
R727 Vdd.n541 Vdd.n538 78.2255
R728 Vdd.n512 Vdd.n503 78.2255
R729 Vdd.n512 Vdd.n504 78.2255
R730 Vdd.n558 Vdd.n553 78.2255
R731 Vdd.n558 Vdd.n554 78.2255
R732 Vdd.n555 Vdd.n553 78.2255
R733 Vdd.n555 Vdd.n554 78.2255
R734 Vdd.n496 Vdd.n487 78.2255
R735 Vdd.n496 Vdd.n488 78.2255
R736 Vdd.n627 Vdd.n622 78.2255
R737 Vdd.n627 Vdd.n623 78.2255
R738 Vdd.n624 Vdd.n622 78.2255
R739 Vdd.n624 Vdd.n623 78.2255
R740 Vdd.n468 Vdd.n466 78.2255
R741 Vdd.n472 Vdd.n468 78.2255
R742 Vdd.n472 Vdd.n469 78.2255
R743 Vdd.n469 Vdd.n466 78.2255
R744 Vdd.n454 Vdd.n448 78.2255
R745 Vdd.n458 Vdd.n454 78.2255
R746 Vdd.n458 Vdd.n455 78.2255
R747 Vdd.n455 Vdd.n448 78.2255
R748 Vdd.n440 Vdd.n435 78.2255
R749 Vdd.n441 Vdd.n435 78.2255
R750 Vdd.n260 Vdd.n228 78.2255
R751 Vdd.n264 Vdd.n228 78.2255
R752 Vdd.n264 Vdd.n229 78.2255
R753 Vdd.n260 Vdd.n229 78.2255
R754 Vdd.n234 Vdd.n232 78.2255
R755 Vdd.n234 Vdd.n233 78.2255
R756 Vdd.n1042 Vdd.t751 70.313
R757 Vdd.n55 Vdd.t544 70.313
R758 Vdd.n5 Vdd.n4 68.0765
R759 Vdd.n1109 Vdd.n1108 68.0765
R760 Vdd.n10 Vdd.n9 68.0765
R761 Vdd.n1097 Vdd.n1096 68.0765
R762 Vdd.n1103 Vdd.n1102 68.0765
R763 Vdd.n1090 Vdd.n1089 68.0765
R764 Vdd.n64 Vdd.n63 68.0765
R765 Vdd.n76 Vdd.n75 68.0765
R766 Vdd.n71 Vdd.n70 68.0765
R767 Vdd.n88 Vdd.n87 68.0765
R768 Vdd.n82 Vdd.n81 68.0765
R769 Vdd.n99 Vdd.n98 68.0765
R770 Vdd.n138 Vdd.n137 68.0765
R771 Vdd.n149 Vdd.n148 68.0765
R772 Vdd.n144 Vdd.n143 68.0765
R773 Vdd.n161 Vdd.n160 68.0765
R774 Vdd.n155 Vdd.n154 68.0765
R775 Vdd.n172 Vdd.n171 68.0765
R776 Vdd.n218 Vdd.n217 68.0765
R777 Vdd.n223 Vdd.n222 68.0765
R778 Vdd.n212 Vdd.n211 68.0765
R779 Vdd.n1015 Vdd.n1014 68.0765
R780 Vdd.n998 Vdd.n997 68.0765
R781 Vdd.n1003 Vdd.n1002 68.0765
R782 Vdd.n1009 Vdd.n1008 68.0765
R783 Vdd.n991 Vdd.n990 68.0765
R784 Vdd.n519 Vdd.n518 68.0765
R785 Vdd.n525 Vdd.n524 68.0765
R786 Vdd.n531 Vdd.n530 68.0765
R787 Vdd.n982 Vdd.n981 68.0765
R788 Vdd.n768 Vdd.n767 68.0765
R789 Vdd.n807 Vdd.n806 68.0765
R790 Vdd.n845 Vdd.n844 68.0765
R791 Vdd.n883 Vdd.n882 68.0765
R792 Vdd.n922 Vdd.n921 68.0765
R793 Vdd.n960 Vdd.n959 68.0765
R794 Vdd.n686 Vdd.n685 68.0765
R795 Vdd.n779 Vdd.n778 68.0765
R796 Vdd.n412 Vdd.n411 68.0765
R797 Vdd.n818 Vdd.n817 68.0765
R798 Vdd.n382 Vdd.n381 68.0765
R799 Vdd.n856 Vdd.n855 68.0765
R800 Vdd.n352 Vdd.n351 68.0765
R801 Vdd.n895 Vdd.n894 68.0765
R802 Vdd.n316 Vdd.n315 68.0765
R803 Vdd.n933 Vdd.n932 68.0765
R804 Vdd.n286 Vdd.n285 68.0765
R805 Vdd.n971 Vdd.n970 68.0765
R806 Vdd.n763 Vdd.n762 68.0765
R807 Vdd.n676 Vdd.n675 68.0765
R808 Vdd.n802 Vdd.n801 68.0765
R809 Vdd.n402 Vdd.n401 68.0765
R810 Vdd.n840 Vdd.n839 68.0765
R811 Vdd.n372 Vdd.n371 68.0765
R812 Vdd.n878 Vdd.n877 68.0765
R813 Vdd.n336 Vdd.n335 68.0765
R814 Vdd.n917 Vdd.n916 68.0765
R815 Vdd.n306 Vdd.n305 68.0765
R816 Vdd.n955 Vdd.n954 68.0765
R817 Vdd.n276 Vdd.n275 68.0765
R818 Vdd.n691 Vdd.n690 68.0765
R819 Vdd.n417 Vdd.n416 68.0765
R820 Vdd.n387 Vdd.n386 68.0765
R821 Vdd.n357 Vdd.n356 68.0765
R822 Vdd.n321 Vdd.n320 68.0765
R823 Vdd.n291 Vdd.n290 68.0765
R824 Vdd.n758 Vdd.n757 68.0765
R825 Vdd.n696 Vdd.n695 68.0765
R826 Vdd.n797 Vdd.n796 68.0765
R827 Vdd.n774 Vdd.n773 68.0765
R828 Vdd.n422 Vdd.n421 68.0765
R829 Vdd.n835 Vdd.n834 68.0765
R830 Vdd.n813 Vdd.n812 68.0765
R831 Vdd.n392 Vdd.n391 68.0765
R832 Vdd.n873 Vdd.n872 68.0765
R833 Vdd.n851 Vdd.n850 68.0765
R834 Vdd.n362 Vdd.n361 68.0765
R835 Vdd.n912 Vdd.n911 68.0765
R836 Vdd.n890 Vdd.n889 68.0765
R837 Vdd.n326 Vdd.n325 68.0765
R838 Vdd.n950 Vdd.n949 68.0765
R839 Vdd.n928 Vdd.n927 68.0765
R840 Vdd.n296 Vdd.n295 68.0765
R841 Vdd.n966 Vdd.n965 68.0765
R842 Vdd.n753 Vdd.n752 68.0765
R843 Vdd.n681 Vdd.n680 68.0765
R844 Vdd.n792 Vdd.n791 68.0765
R845 Vdd.n407 Vdd.n406 68.0765
R846 Vdd.n830 Vdd.n829 68.0765
R847 Vdd.n377 Vdd.n376 68.0765
R848 Vdd.n868 Vdd.n867 68.0765
R849 Vdd.n341 Vdd.n340 68.0765
R850 Vdd.n907 Vdd.n906 68.0765
R851 Vdd.n311 Vdd.n310 68.0765
R852 Vdd.n945 Vdd.n944 68.0765
R853 Vdd.n281 Vdd.n280 68.0765
R854 Vdd.n701 Vdd.n700 68.0765
R855 Vdd.n427 Vdd.n426 68.0765
R856 Vdd.n397 Vdd.n396 68.0765
R857 Vdd.n367 Vdd.n366 68.0765
R858 Vdd.n331 Vdd.n330 68.0765
R859 Vdd.n301 Vdd.n300 68.0765
R860 Vdd.n706 Vdd.n705 68.0765
R861 Vdd.n722 Vdd.n721 68.0765
R862 Vdd.n717 Vdd.n716 68.0765
R863 Vdd.n740 Vdd.n739 68.0765
R864 Vdd.n746 Vdd.n745 68.0765
R865 Vdd.n734 Vdd.n733 68.0765
R866 Vdd.n639 Vdd.n638 68.0765
R867 Vdd.n650 Vdd.n649 68.0765
R868 Vdd.n645 Vdd.n644 68.0765
R869 Vdd.n662 Vdd.n661 68.0765
R870 Vdd.n656 Vdd.n655 68.0765
R871 Vdd.n669 Vdd.n668 68.0765
R872 Vdd.n570 Vdd.n569 68.0765
R873 Vdd.n581 Vdd.n580 68.0765
R874 Vdd.n576 Vdd.n575 68.0765
R875 Vdd.n593 Vdd.n592 68.0765
R876 Vdd.n587 Vdd.n586 68.0765
R877 Vdd.n600 Vdd.n599 68.0765
R878 Vdd.n38 Vdd.n36 59.8505
R879 Vdd.n40 Vdd.n37 59.8505
R880 Vdd.n22 Vdd.n20 59.8505
R881 Vdd.n24 Vdd.n21 59.8505
R882 Vdd.n505 Vdd.n503 59.8505
R883 Vdd.n507 Vdd.n504 59.8505
R884 Vdd.n489 Vdd.n487 59.8505
R885 Vdd.n491 Vdd.n488 59.8505
R886 Vdd.n440 Vdd.n438 59.8505
R887 Vdd.n441 Vdd.n439 59.8505
R888 Vdd.n235 Vdd.n232 59.8505
R889 Vdd.n237 Vdd.n233 59.8505
R890 Vdd.n1026 Vdd.n1024 58.9755
R891 Vdd.n1029 Vdd.n1024 58.9755
R892 Vdd.n1029 Vdd.n1025 58.9755
R893 Vdd.n1026 Vdd.n1025 58.9755
R894 Vdd.n1072 Vdd.n1047 54.0755
R895 Vdd.n1054 Vdd.n1049 54.0755
R896 Vdd.n1054 Vdd.n1050 54.0755
R897 Vdd.n1072 Vdd.n1048 54.0755
R898 Vdd.n205 Vdd.t669 41.0041
R899 Vdd.n92 Vdd.t651 41.0041
R900 Vdd.n165 Vdd.t738 41.0041
R901 Vdd.n975 Vdd.t654 41.0041
R902 Vdd.n726 Vdd.t726 41.0041
R903 Vdd.n430 Vdd.t735 41.0041
R904 Vdd.n344 Vdd.t636 41.0041
R905 Vdd.n207 Vdd.t705 40.8177
R906 Vdd.n206 Vdd.t666 40.8177
R907 Vdd.n94 Vdd.t645 40.8177
R908 Vdd.n93 Vdd.t609 40.8177
R909 Vdd.n167 Vdd.t630 40.8177
R910 Vdd.n166 Vdd.t732 40.8177
R911 Vdd.n977 Vdd.t690 40.8177
R912 Vdd.n976 Vdd.t648 40.8177
R913 Vdd.n729 Vdd.t720 40.8177
R914 Vdd.n728 Vdd.t624 40.8177
R915 Vdd.n432 Vdd.t684 40.8177
R916 Vdd.n431 Vdd.t639 40.8177
R917 Vdd.n346 Vdd.t687 40.8177
R918 Vdd.n345 Vdd.t642 40.8177
R919 Vdd.n47 Vdd.t723 40.6313
R920 Vdd.n46 Vdd.t612 40.6313
R921 Vdd.n133 Vdd.t702 40.6313
R922 Vdd.n132 Vdd.t714 40.6313
R923 Vdd.n514 Vdd.t618 40.6313
R924 Vdd.n513 Vdd.t633 40.6313
R925 Vdd.n786 Vdd.t615 40.6313
R926 Vdd.n784 Vdd.t657 40.6313
R927 Vdd.n824 Vdd.t663 40.6313
R928 Vdd.n822 Vdd.t681 40.6313
R929 Vdd.n862 Vdd.t711 40.6313
R930 Vdd.n860 Vdd.t729 40.6313
R931 Vdd.n901 Vdd.t672 40.6313
R932 Vdd.n899 Vdd.t678 40.6313
R933 Vdd.n939 Vdd.t717 40.6313
R934 Vdd.n937 Vdd.t693 40.6313
R935 Vdd.n711 Vdd.t708 40.6313
R936 Vdd.n709 Vdd.t699 40.6313
R937 Vdd.n565 Vdd.t606 40.6313
R938 Vdd.n564 Vdd.t627 40.6313
R939 Vdd.n634 Vdd.t621 40.6313
R940 Vdd.n633 Vdd.t660 40.6313
R941 Vdd.n1 Vdd.t675 40.6313
R942 Vdd.n0 Vdd.t696 40.6313
R943 Vdd.n183 Vdd.n181 36.2255
R944 Vdd.n183 Vdd.n182 36.2255
R945 Vdd.n110 Vdd.n108 36.2255
R946 Vdd.n110 Vdd.n109 36.2255
R947 Vdd.n41 Vdd.n38 36.2255
R948 Vdd.n41 Vdd.n40 36.2255
R949 Vdd.n43 Vdd.n36 36.2255
R950 Vdd.n43 Vdd.n37 36.2255
R951 Vdd.n124 Vdd.n121 36.2255
R952 Vdd.n124 Vdd.n122 36.2255
R953 Vdd.n25 Vdd.n22 36.2255
R954 Vdd.n25 Vdd.n24 36.2255
R955 Vdd.n27 Vdd.n20 36.2255
R956 Vdd.n27 Vdd.n21 36.2255
R957 Vdd.n197 Vdd.n194 36.2255
R958 Vdd.n197 Vdd.n195 36.2255
R959 Vdd.n248 Vdd.n246 36.2255
R960 Vdd.n248 Vdd.n247 36.2255
R961 Vdd.n611 Vdd.n609 36.2255
R962 Vdd.n611 Vdd.n610 36.2255
R963 Vdd.n542 Vdd.n540 36.2255
R964 Vdd.n542 Vdd.n541 36.2255
R965 Vdd.n508 Vdd.n505 36.2255
R966 Vdd.n508 Vdd.n507 36.2255
R967 Vdd.n510 Vdd.n503 36.2255
R968 Vdd.n510 Vdd.n504 36.2255
R969 Vdd.n556 Vdd.n553 36.2255
R970 Vdd.n556 Vdd.n554 36.2255
R971 Vdd.n492 Vdd.n489 36.2255
R972 Vdd.n492 Vdd.n491 36.2255
R973 Vdd.n494 Vdd.n487 36.2255
R974 Vdd.n494 Vdd.n488 36.2255
R975 Vdd.n625 Vdd.n622 36.2255
R976 Vdd.n625 Vdd.n623 36.2255
R977 Vdd.n470 Vdd.n468 36.2255
R978 Vdd.n470 Vdd.n469 36.2255
R979 Vdd.n456 Vdd.n454 36.2255
R980 Vdd.n456 Vdd.n455 36.2255
R981 Vdd.n444 Vdd.n438 36.2255
R982 Vdd.n444 Vdd.n439 36.2255
R983 Vdd.n442 Vdd.n440 36.2255
R984 Vdd.n442 Vdd.n441 36.2255
R985 Vdd.n262 Vdd.n228 36.2255
R986 Vdd.n262 Vdd.n229 36.2255
R987 Vdd.n238 Vdd.n235 36.2255
R988 Vdd.n238 Vdd.n237 36.2255
R989 Vdd.n241 Vdd.n232 36.2255
R990 Vdd.n241 Vdd.n233 36.2255
R991 Vdd.n783 Vdd.n673 32.646
R992 Vdd.n1076 Vdd.n1075 29.3622
R993 Vdd.n1053 Vdd.n1052 29.3622
R994 Vdd.n47 Vdd.t968 27.3166
R995 Vdd.n46 Vdd.t960 27.3166
R996 Vdd.n133 Vdd.t973 27.3166
R997 Vdd.n132 Vdd.t971 27.3166
R998 Vdd.n514 Vdd.t959 27.3166
R999 Vdd.n513 Vdd.t995 27.3166
R1000 Vdd.n786 Vdd.t970 27.3166
R1001 Vdd.n784 Vdd.t986 27.3166
R1002 Vdd.n824 Vdd.t958 27.3166
R1003 Vdd.n822 Vdd.t977 27.3166
R1004 Vdd.n862 Vdd.t981 27.3166
R1005 Vdd.n860 Vdd.t966 27.3166
R1006 Vdd.n901 Vdd.t999 27.3166
R1007 Vdd.n899 Vdd.t978 27.3166
R1008 Vdd.n939 Vdd.t980 27.3166
R1009 Vdd.n937 Vdd.t976 27.3166
R1010 Vdd.n711 Vdd.t982 27.3166
R1011 Vdd.n709 Vdd.t974 27.3166
R1012 Vdd.n565 Vdd.t962 27.3166
R1013 Vdd.n564 Vdd.t996 27.3166
R1014 Vdd.n634 Vdd.t957 27.3166
R1015 Vdd.n633 Vdd.t985 27.3166
R1016 Vdd.n1 Vdd.t979 27.3166
R1017 Vdd.n0 Vdd.t975 27.3166
R1018 Vdd.n207 Vdd.t992 27.1302
R1019 Vdd.n206 Vdd.t984 27.1302
R1020 Vdd.n94 Vdd.t967 27.1302
R1021 Vdd.n93 Vdd.t961 27.1302
R1022 Vdd.n167 Vdd.t972 27.1302
R1023 Vdd.n166 Vdd.t965 27.1302
R1024 Vdd.n977 Vdd.t997 27.1302
R1025 Vdd.n976 Vdd.t989 27.1302
R1026 Vdd.n729 Vdd.t969 27.1302
R1027 Vdd.n728 Vdd.t956 27.1302
R1028 Vdd.n432 Vdd.t955 27.1302
R1029 Vdd.n431 Vdd.t993 27.1302
R1030 Vdd.n346 Vdd.t998 27.1302
R1031 Vdd.n345 Vdd.t990 27.1302
R1032 Vdd.n205 Vdd.t983 26.9438
R1033 Vdd.n92 Vdd.t988 26.9438
R1034 Vdd.n165 Vdd.t963 26.9438
R1035 Vdd.n975 Vdd.t987 26.9438
R1036 Vdd.n726 Vdd.t991 26.9438
R1037 Vdd.n430 Vdd.t964 26.9438
R1038 Vdd.n344 Vdd.t994 26.9438
R1039 Vdd.t747 Vdd.n1040 23.438
R1040 Vdd.n59 Vdd.t542 23.438
R1041 Vdd.n1068 Vdd.n1049 20.1255
R1042 Vdd.n1068 Vdd.n1050 20.1255
R1043 Vdd.n1070 Vdd.n1047 20.1255
R1044 Vdd.n1070 Vdd.n1048 20.1255
R1045 Vdd.n1077 Vdd.n1076 19.9167
R1046 Vdd.n1052 Vdd.n1051 19.9167
R1047 Vdd.n1027 Vdd.n1024 18.7255
R1048 Vdd.n1027 Vdd.n1025 18.7255
R1049 Vdd.n737 SARlogic_0.dffrs_13.resetb 18.2673
R1050 Vdd.n102 adc_PISO_0.dffrs_5.resetb 18.2415
R1051 Vdd.n175 adc_PISO_0.dffrs_4.resetb 18.2415
R1052 Vdd.n1087 adc_PISO_0.dffrs_3.resetb 18.2061
R1053 Vdd.n986 adc_PISO_0.dffrs_2.resetb 18.2061
R1054 Vdd.n673 adc_PISO_0.dffrs_0.resetb 18.2061
R1055 Vdd.n349 adc_PISO_0.dffrs_1.resetb 18.2061
R1056 Vdd.n68 Vdd.n49 18.0418
R1057 Vdd.n141 Vdd.n135 18.0418
R1058 Vdd.n522 Vdd.n516 18.0418
R1059 Vdd.n573 Vdd.n567 18.0418
R1060 Vdd.n642 Vdd.n636 18.0418
R1061 Vdd.n1114 Vdd.n1113 18.0418
R1062 Vdd.n789 Vdd.n788 18.0005
R1063 Vdd.n827 Vdd.n826 18.0005
R1064 Vdd.n865 Vdd.n864 18.0005
R1065 Vdd.n904 Vdd.n903 18.0005
R1066 Vdd.n942 Vdd.n941 18.0005
R1067 Vdd.n714 Vdd.n713 18.0005
R1068 Vdd.n208 Vdd.n206 17.6364
R1069 Vdd.n95 Vdd.n93 17.6364
R1070 Vdd.n168 Vdd.n166 17.6364
R1071 Vdd.n978 Vdd.n976 17.6364
R1072 Vdd.n433 Vdd.n431 17.6364
R1073 Vdd.n347 Vdd.n345 17.6364
R1074 Vdd.n1079 Vdd.n1078 14.6602
R1075 Vdd.n48 Vdd.n46 14.3609
R1076 Vdd.n134 Vdd.n132 14.3609
R1077 Vdd.n515 Vdd.n513 14.3609
R1078 Vdd.n566 Vdd.n564 14.3609
R1079 Vdd.n635 Vdd.n633 14.3609
R1080 Vdd.n2 Vdd.n0 14.3609
R1081 Vdd.n226 Vdd.n220 13.5842
R1082 Vdd.n522 Vdd.n521 13.5431
R1083 Vdd.n1113 Vdd.n7 13.5174
R1084 Vdd.n141 Vdd.n140 13.5174
R1085 Vdd.n642 Vdd.n641 13.5174
R1086 Vdd.n573 Vdd.n572 13.5174
R1087 Vdd.n714 Vdd.n708 13.5152
R1088 Vdd.n1112 Vdd.n1111 13.5005
R1089 Vdd.n1112 Vdd.n12 13.5005
R1090 Vdd.n1100 Vdd.n1099 13.5005
R1091 Vdd.n1106 Vdd.n1105 13.5005
R1092 Vdd.n1093 Vdd.n1092 13.5005
R1093 Vdd.n67 Vdd.n66 13.5005
R1094 Vdd.n79 Vdd.n78 13.5005
R1095 Vdd.n79 Vdd.n73 13.5005
R1096 Vdd.n91 Vdd.n90 13.5005
R1097 Vdd.n85 Vdd.n84 13.5005
R1098 Vdd.n102 Vdd.n101 13.5005
R1099 Vdd.n152 Vdd.n151 13.5005
R1100 Vdd.n152 Vdd.n146 13.5005
R1101 Vdd.n164 Vdd.n163 13.5005
R1102 Vdd.n158 Vdd.n157 13.5005
R1103 Vdd.n175 Vdd.n174 13.5005
R1104 Vdd.n226 Vdd.n225 13.5005
R1105 Vdd.n215 Vdd.n214 13.5005
R1106 Vdd.n1018 Vdd.n1017 13.5005
R1107 Vdd.n1018 Vdd.n1000 13.5005
R1108 Vdd.n1006 Vdd.n1005 13.5005
R1109 Vdd.n1012 Vdd.n1011 13.5005
R1110 Vdd.n994 Vdd.n993 13.5005
R1111 Vdd.n528 Vdd.n527 13.5005
R1112 Vdd.n534 Vdd.n533 13.5005
R1113 Vdd.n985 Vdd.n984 13.5005
R1114 Vdd.n771 Vdd.n770 13.5005
R1115 Vdd.n810 Vdd.n809 13.5005
R1116 Vdd.n848 Vdd.n847 13.5005
R1117 Vdd.n886 Vdd.n885 13.5005
R1118 Vdd.n925 Vdd.n924 13.5005
R1119 Vdd.n963 Vdd.n962 13.5005
R1120 Vdd.n771 Vdd.n688 13.5005
R1121 Vdd.n782 Vdd.n781 13.5005
R1122 Vdd.n810 Vdd.n414 13.5005
R1123 Vdd.n821 Vdd.n820 13.5005
R1124 Vdd.n848 Vdd.n384 13.5005
R1125 Vdd.n859 Vdd.n858 13.5005
R1126 Vdd.n886 Vdd.n354 13.5005
R1127 Vdd.n898 Vdd.n897 13.5005
R1128 Vdd.n925 Vdd.n318 13.5005
R1129 Vdd.n936 Vdd.n935 13.5005
R1130 Vdd.n963 Vdd.n288 13.5005
R1131 Vdd.n974 Vdd.n973 13.5005
R1132 Vdd.n771 Vdd.n765 13.5005
R1133 Vdd.n782 Vdd.n678 13.5005
R1134 Vdd.n810 Vdd.n804 13.5005
R1135 Vdd.n821 Vdd.n404 13.5005
R1136 Vdd.n848 Vdd.n842 13.5005
R1137 Vdd.n859 Vdd.n374 13.5005
R1138 Vdd.n886 Vdd.n880 13.5005
R1139 Vdd.n898 Vdd.n338 13.5005
R1140 Vdd.n925 Vdd.n919 13.5005
R1141 Vdd.n936 Vdd.n308 13.5005
R1142 Vdd.n963 Vdd.n957 13.5005
R1143 Vdd.n974 Vdd.n278 13.5005
R1144 Vdd.n771 Vdd.n693 13.5005
R1145 Vdd.n810 Vdd.n419 13.5005
R1146 Vdd.n848 Vdd.n389 13.5005
R1147 Vdd.n886 Vdd.n359 13.5005
R1148 Vdd.n925 Vdd.n323 13.5005
R1149 Vdd.n963 Vdd.n293 13.5005
R1150 Vdd.n771 Vdd.n760 13.5005
R1151 Vdd.n771 Vdd.n698 13.5005
R1152 Vdd.n810 Vdd.n799 13.5005
R1153 Vdd.n782 Vdd.n776 13.5005
R1154 Vdd.n810 Vdd.n424 13.5005
R1155 Vdd.n848 Vdd.n837 13.5005
R1156 Vdd.n821 Vdd.n815 13.5005
R1157 Vdd.n848 Vdd.n394 13.5005
R1158 Vdd.n886 Vdd.n875 13.5005
R1159 Vdd.n859 Vdd.n853 13.5005
R1160 Vdd.n886 Vdd.n364 13.5005
R1161 Vdd.n925 Vdd.n914 13.5005
R1162 Vdd.n898 Vdd.n892 13.5005
R1163 Vdd.n925 Vdd.n328 13.5005
R1164 Vdd.n963 Vdd.n952 13.5005
R1165 Vdd.n936 Vdd.n930 13.5005
R1166 Vdd.n963 Vdd.n298 13.5005
R1167 Vdd.n974 Vdd.n968 13.5005
R1168 Vdd.n771 Vdd.n755 13.5005
R1169 Vdd.n782 Vdd.n683 13.5005
R1170 Vdd.n810 Vdd.n794 13.5005
R1171 Vdd.n821 Vdd.n409 13.5005
R1172 Vdd.n848 Vdd.n832 13.5005
R1173 Vdd.n859 Vdd.n379 13.5005
R1174 Vdd.n886 Vdd.n870 13.5005
R1175 Vdd.n898 Vdd.n343 13.5005
R1176 Vdd.n925 Vdd.n909 13.5005
R1177 Vdd.n936 Vdd.n313 13.5005
R1178 Vdd.n963 Vdd.n947 13.5005
R1179 Vdd.n974 Vdd.n283 13.5005
R1180 Vdd.n771 Vdd.n703 13.5005
R1181 Vdd.n810 Vdd.n429 13.5005
R1182 Vdd.n848 Vdd.n399 13.5005
R1183 Vdd.n886 Vdd.n369 13.5005
R1184 Vdd.n925 Vdd.n333 13.5005
R1185 Vdd.n963 Vdd.n303 13.5005
R1186 Vdd.n725 Vdd.n724 13.5005
R1187 Vdd.n725 Vdd.n719 13.5005
R1188 Vdd.n743 Vdd.n742 13.5005
R1189 Vdd.n749 Vdd.n748 13.5005
R1190 Vdd.n737 Vdd.n736 13.5005
R1191 Vdd.n653 Vdd.n652 13.5005
R1192 Vdd.n653 Vdd.n647 13.5005
R1193 Vdd.n665 Vdd.n664 13.5005
R1194 Vdd.n659 Vdd.n658 13.5005
R1195 Vdd.n672 Vdd.n671 13.5005
R1196 Vdd.n584 Vdd.n583 13.5005
R1197 Vdd.n584 Vdd.n578 13.5005
R1198 Vdd.n596 Vdd.n595 13.5005
R1199 Vdd.n590 Vdd.n589 13.5005
R1200 Vdd.n603 Vdd.n602 13.5005
R1201 Vdd.n1084 Vdd.n1021 13.4987
R1202 Vdd.n209 Vdd.n205 13.4839
R1203 Vdd.n96 Vdd.n92 13.4839
R1204 Vdd.n169 Vdd.n165 13.4839
R1205 Vdd.n979 Vdd.n975 13.4839
R1206 Vdd.n434 Vdd.n430 13.4839
R1207 Vdd.n348 Vdd.n344 13.4839
R1208 Vdd.n1040 Vdd.n1034 12.6005
R1209 Vdd.n1044 Vdd.n1043 12.6005
R1210 Vdd.n1042 Vdd.n1041 12.6005
R1211 Vdd.n59 Vdd.n58 12.6005
R1212 Vdd.n57 Vdd.n56 12.6005
R1213 Vdd.n55 Vdd.n54 12.6005
R1214 Vdd.n730 SARlogic_0.dffrs_13.nand3_1.B 12.1571
R1215 Vdd.n1066 Vdd.n1065 12.136
R1216 Vdd.n1064 Vdd.n1063 12.136
R1217 Vdd.n1062 Vdd.n1061 12.136
R1218 Vdd.n1060 Vdd.n1059 12.136
R1219 Vdd.n1058 Vdd.n1057 12.136
R1220 Vdd.n1070 Vdd.n1046 11.111
R1221 Vdd.n1068 Vdd.n1067 11.111
R1222 Vdd.n208 Vdd.n207 10.5752
R1223 Vdd.n95 Vdd.n94 10.5752
R1224 Vdd.n168 Vdd.n167 10.5752
R1225 Vdd.n978 Vdd.n977 10.5752
R1226 Vdd.n433 Vdd.n432 10.5752
R1227 Vdd.n347 Vdd.n346 10.5752
R1228 Vdd.n1051 Vdd.n1021 9.86945
R1229 Vdd.n1056 Vdd.n1055 9.536
R1230 Vdd.n1074 Vdd.n1073 9.536
R1231 Vdd.n1078 Vdd.n1077 9.536
R1232 Vdd.n67 Vdd.n61 9.53505
R1233 Vdd.n787 Vdd.n785 9.22229
R1234 Vdd.n825 Vdd.n823 9.22229
R1235 Vdd.n863 Vdd.n861 9.22229
R1236 Vdd.n902 Vdd.n900 9.22229
R1237 Vdd.n940 Vdd.n938 9.22229
R1238 Vdd.n712 Vdd.n710 9.22229
R1239 Vdd.n731 Vdd.n727 7.75389
R1240 Vdd.n1055 Vdd.t67 7.4755
R1241 Vdd.n1073 Vdd.t57 7.4755
R1242 Vdd.n1077 Vdd.t59 7.4755
R1243 Vdd.n1051 Vdd.t53 7.4755
R1244 Vdd.n988 Vdd.n987 6.55364
R1245 Vdd.n7 Vdd.n4 6.4802
R1246 Vdd.n1111 Vdd.n1108 6.4802
R1247 Vdd.n12 Vdd.n9 6.4802
R1248 Vdd.n1099 Vdd.n1096 6.4802
R1249 Vdd.n1105 Vdd.n1102 6.4802
R1250 Vdd.n1092 Vdd.n1089 6.4802
R1251 Vdd.n66 Vdd.n63 6.4802
R1252 Vdd.n78 Vdd.n75 6.4802
R1253 Vdd.n73 Vdd.n70 6.4802
R1254 Vdd.n90 Vdd.n87 6.4802
R1255 Vdd.n84 Vdd.n81 6.4802
R1256 Vdd.n101 Vdd.n98 6.4802
R1257 Vdd.n140 Vdd.n137 6.4802
R1258 Vdd.n151 Vdd.n148 6.4802
R1259 Vdd.n146 Vdd.n143 6.4802
R1260 Vdd.n163 Vdd.n160 6.4802
R1261 Vdd.n157 Vdd.n154 6.4802
R1262 Vdd.n174 Vdd.n171 6.4802
R1263 Vdd.n220 Vdd.n217 6.4802
R1264 Vdd.n225 Vdd.n222 6.4802
R1265 Vdd.n214 Vdd.n211 6.4802
R1266 Vdd.n1017 Vdd.n1014 6.4802
R1267 Vdd.n1000 Vdd.n997 6.4802
R1268 Vdd.n1005 Vdd.n1002 6.4802
R1269 Vdd.n1011 Vdd.n1008 6.4802
R1270 Vdd.n993 Vdd.n990 6.4802
R1271 Vdd.n521 Vdd.n518 6.4802
R1272 Vdd.n527 Vdd.n524 6.4802
R1273 Vdd.n533 Vdd.n530 6.4802
R1274 Vdd.n984 Vdd.n981 6.4802
R1275 Vdd.n770 Vdd.n767 6.4802
R1276 Vdd.n809 Vdd.n806 6.4802
R1277 Vdd.n847 Vdd.n844 6.4802
R1278 Vdd.n885 Vdd.n882 6.4802
R1279 Vdd.n924 Vdd.n921 6.4802
R1280 Vdd.n962 Vdd.n959 6.4802
R1281 Vdd.n688 Vdd.n685 6.4802
R1282 Vdd.n781 Vdd.n778 6.4802
R1283 Vdd.n414 Vdd.n411 6.4802
R1284 Vdd.n820 Vdd.n817 6.4802
R1285 Vdd.n384 Vdd.n381 6.4802
R1286 Vdd.n858 Vdd.n855 6.4802
R1287 Vdd.n354 Vdd.n351 6.4802
R1288 Vdd.n897 Vdd.n894 6.4802
R1289 Vdd.n318 Vdd.n315 6.4802
R1290 Vdd.n935 Vdd.n932 6.4802
R1291 Vdd.n288 Vdd.n285 6.4802
R1292 Vdd.n973 Vdd.n970 6.4802
R1293 Vdd.n765 Vdd.n762 6.4802
R1294 Vdd.n678 Vdd.n675 6.4802
R1295 Vdd.n804 Vdd.n801 6.4802
R1296 Vdd.n404 Vdd.n401 6.4802
R1297 Vdd.n842 Vdd.n839 6.4802
R1298 Vdd.n374 Vdd.n371 6.4802
R1299 Vdd.n880 Vdd.n877 6.4802
R1300 Vdd.n338 Vdd.n335 6.4802
R1301 Vdd.n919 Vdd.n916 6.4802
R1302 Vdd.n308 Vdd.n305 6.4802
R1303 Vdd.n957 Vdd.n954 6.4802
R1304 Vdd.n278 Vdd.n275 6.4802
R1305 Vdd.n693 Vdd.n690 6.4802
R1306 Vdd.n419 Vdd.n416 6.4802
R1307 Vdd.n389 Vdd.n386 6.4802
R1308 Vdd.n359 Vdd.n356 6.4802
R1309 Vdd.n323 Vdd.n320 6.4802
R1310 Vdd.n293 Vdd.n290 6.4802
R1311 Vdd.n760 Vdd.n757 6.4802
R1312 Vdd.n698 Vdd.n695 6.4802
R1313 Vdd.n799 Vdd.n796 6.4802
R1314 Vdd.n776 Vdd.n773 6.4802
R1315 Vdd.n424 Vdd.n421 6.4802
R1316 Vdd.n837 Vdd.n834 6.4802
R1317 Vdd.n815 Vdd.n812 6.4802
R1318 Vdd.n394 Vdd.n391 6.4802
R1319 Vdd.n875 Vdd.n872 6.4802
R1320 Vdd.n853 Vdd.n850 6.4802
R1321 Vdd.n364 Vdd.n361 6.4802
R1322 Vdd.n914 Vdd.n911 6.4802
R1323 Vdd.n892 Vdd.n889 6.4802
R1324 Vdd.n328 Vdd.n325 6.4802
R1325 Vdd.n952 Vdd.n949 6.4802
R1326 Vdd.n930 Vdd.n927 6.4802
R1327 Vdd.n298 Vdd.n295 6.4802
R1328 Vdd.n968 Vdd.n965 6.4802
R1329 Vdd.n755 Vdd.n752 6.4802
R1330 Vdd.n683 Vdd.n680 6.4802
R1331 Vdd.n794 Vdd.n791 6.4802
R1332 Vdd.n409 Vdd.n406 6.4802
R1333 Vdd.n832 Vdd.n829 6.4802
R1334 Vdd.n379 Vdd.n376 6.4802
R1335 Vdd.n870 Vdd.n867 6.4802
R1336 Vdd.n343 Vdd.n340 6.4802
R1337 Vdd.n909 Vdd.n906 6.4802
R1338 Vdd.n313 Vdd.n310 6.4802
R1339 Vdd.n947 Vdd.n944 6.4802
R1340 Vdd.n283 Vdd.n280 6.4802
R1341 Vdd.n703 Vdd.n700 6.4802
R1342 Vdd.n429 Vdd.n426 6.4802
R1343 Vdd.n399 Vdd.n396 6.4802
R1344 Vdd.n369 Vdd.n366 6.4802
R1345 Vdd.n333 Vdd.n330 6.4802
R1346 Vdd.n303 Vdd.n300 6.4802
R1347 Vdd.n708 Vdd.n705 6.4802
R1348 Vdd.n724 Vdd.n721 6.4802
R1349 Vdd.n719 Vdd.n716 6.4802
R1350 Vdd.n742 Vdd.n739 6.4802
R1351 Vdd.n748 Vdd.n745 6.4802
R1352 Vdd.n736 Vdd.n733 6.4802
R1353 Vdd.n641 Vdd.n638 6.4802
R1354 Vdd.n652 Vdd.n649 6.4802
R1355 Vdd.n647 Vdd.n644 6.4802
R1356 Vdd.n664 Vdd.n661 6.4802
R1357 Vdd.n658 Vdd.n655 6.4802
R1358 Vdd.n671 Vdd.n668 6.4802
R1359 Vdd.n572 Vdd.n569 6.4802
R1360 Vdd.n583 Vdd.n580 6.4802
R1361 Vdd.n578 Vdd.n575 6.4802
R1362 Vdd.n595 Vdd.n592 6.4802
R1363 Vdd.n589 Vdd.n586 6.4802
R1364 Vdd.n602 Vdd.n599 6.4802
R1365 Vdd.n7 Vdd.n3 6.25878
R1366 Vdd.n1111 Vdd.n1107 6.25878
R1367 Vdd.n12 Vdd.n8 6.25878
R1368 Vdd.n1099 Vdd.n1095 6.25878
R1369 Vdd.n1105 Vdd.n1101 6.25878
R1370 Vdd.n1092 Vdd.n1088 6.25878
R1371 Vdd.n66 Vdd.n62 6.25878
R1372 Vdd.n78 Vdd.n74 6.25878
R1373 Vdd.n73 Vdd.n69 6.25878
R1374 Vdd.n90 Vdd.n86 6.25878
R1375 Vdd.n84 Vdd.n80 6.25878
R1376 Vdd.n101 Vdd.n97 6.25878
R1377 Vdd.n140 Vdd.n136 6.25878
R1378 Vdd.n151 Vdd.n147 6.25878
R1379 Vdd.n146 Vdd.n142 6.25878
R1380 Vdd.n163 Vdd.n159 6.25878
R1381 Vdd.n157 Vdd.n153 6.25878
R1382 Vdd.n174 Vdd.n170 6.25878
R1383 Vdd.n220 Vdd.n216 6.25878
R1384 Vdd.n225 Vdd.n221 6.25878
R1385 Vdd.n214 Vdd.n210 6.25878
R1386 Vdd.n1017 Vdd.n1013 6.25878
R1387 Vdd.n1000 Vdd.n996 6.25878
R1388 Vdd.n1005 Vdd.n1001 6.25878
R1389 Vdd.n1011 Vdd.n1007 6.25878
R1390 Vdd.n993 Vdd.n989 6.25878
R1391 Vdd.n521 Vdd.n517 6.25878
R1392 Vdd.n527 Vdd.n523 6.25878
R1393 Vdd.n533 Vdd.n529 6.25878
R1394 Vdd.n984 Vdd.n980 6.25878
R1395 Vdd.n770 Vdd.n766 6.25878
R1396 Vdd.n809 Vdd.n805 6.25878
R1397 Vdd.n847 Vdd.n843 6.25878
R1398 Vdd.n885 Vdd.n881 6.25878
R1399 Vdd.n924 Vdd.n920 6.25878
R1400 Vdd.n962 Vdd.n958 6.25878
R1401 Vdd.n688 Vdd.n684 6.25878
R1402 Vdd.n781 Vdd.n777 6.25878
R1403 Vdd.n414 Vdd.n410 6.25878
R1404 Vdd.n820 Vdd.n816 6.25878
R1405 Vdd.n384 Vdd.n380 6.25878
R1406 Vdd.n858 Vdd.n854 6.25878
R1407 Vdd.n354 Vdd.n350 6.25878
R1408 Vdd.n897 Vdd.n893 6.25878
R1409 Vdd.n318 Vdd.n314 6.25878
R1410 Vdd.n935 Vdd.n931 6.25878
R1411 Vdd.n288 Vdd.n284 6.25878
R1412 Vdd.n973 Vdd.n969 6.25878
R1413 Vdd.n765 Vdd.n761 6.25878
R1414 Vdd.n678 Vdd.n674 6.25878
R1415 Vdd.n804 Vdd.n800 6.25878
R1416 Vdd.n404 Vdd.n400 6.25878
R1417 Vdd.n842 Vdd.n838 6.25878
R1418 Vdd.n374 Vdd.n370 6.25878
R1419 Vdd.n880 Vdd.n876 6.25878
R1420 Vdd.n338 Vdd.n334 6.25878
R1421 Vdd.n919 Vdd.n915 6.25878
R1422 Vdd.n308 Vdd.n304 6.25878
R1423 Vdd.n957 Vdd.n953 6.25878
R1424 Vdd.n278 Vdd.n274 6.25878
R1425 Vdd.n693 Vdd.n689 6.25878
R1426 Vdd.n419 Vdd.n415 6.25878
R1427 Vdd.n389 Vdd.n385 6.25878
R1428 Vdd.n359 Vdd.n355 6.25878
R1429 Vdd.n323 Vdd.n319 6.25878
R1430 Vdd.n293 Vdd.n289 6.25878
R1431 Vdd.n760 Vdd.n756 6.25878
R1432 Vdd.n698 Vdd.n694 6.25878
R1433 Vdd.n799 Vdd.n795 6.25878
R1434 Vdd.n776 Vdd.n772 6.25878
R1435 Vdd.n424 Vdd.n420 6.25878
R1436 Vdd.n837 Vdd.n833 6.25878
R1437 Vdd.n815 Vdd.n811 6.25878
R1438 Vdd.n394 Vdd.n390 6.25878
R1439 Vdd.n875 Vdd.n871 6.25878
R1440 Vdd.n853 Vdd.n849 6.25878
R1441 Vdd.n364 Vdd.n360 6.25878
R1442 Vdd.n914 Vdd.n910 6.25878
R1443 Vdd.n892 Vdd.n888 6.25878
R1444 Vdd.n328 Vdd.n324 6.25878
R1445 Vdd.n952 Vdd.n948 6.25878
R1446 Vdd.n930 Vdd.n926 6.25878
R1447 Vdd.n298 Vdd.n294 6.25878
R1448 Vdd.n968 Vdd.n964 6.25878
R1449 Vdd.n755 Vdd.n751 6.25878
R1450 Vdd.n683 Vdd.n679 6.25878
R1451 Vdd.n794 Vdd.n790 6.25878
R1452 Vdd.n409 Vdd.n405 6.25878
R1453 Vdd.n832 Vdd.n828 6.25878
R1454 Vdd.n379 Vdd.n375 6.25878
R1455 Vdd.n870 Vdd.n866 6.25878
R1456 Vdd.n343 Vdd.n339 6.25878
R1457 Vdd.n909 Vdd.n905 6.25878
R1458 Vdd.n313 Vdd.n309 6.25878
R1459 Vdd.n947 Vdd.n943 6.25878
R1460 Vdd.n283 Vdd.n279 6.25878
R1461 Vdd.n703 Vdd.n699 6.25878
R1462 Vdd.n429 Vdd.n425 6.25878
R1463 Vdd.n399 Vdd.n395 6.25878
R1464 Vdd.n369 Vdd.n365 6.25878
R1465 Vdd.n333 Vdd.n329 6.25878
R1466 Vdd.n303 Vdd.n299 6.25878
R1467 Vdd.n708 Vdd.n704 6.25878
R1468 Vdd.n724 Vdd.n720 6.25878
R1469 Vdd.n719 Vdd.n715 6.25878
R1470 Vdd.n742 Vdd.n738 6.25878
R1471 Vdd.n748 Vdd.n744 6.25878
R1472 Vdd.n736 Vdd.n732 6.25878
R1473 Vdd.n641 Vdd.n637 6.25878
R1474 Vdd.n652 Vdd.n648 6.25878
R1475 Vdd.n647 Vdd.n643 6.25878
R1476 Vdd.n664 Vdd.n660 6.25878
R1477 Vdd.n658 Vdd.n654 6.25878
R1478 Vdd.n671 Vdd.n667 6.25878
R1479 Vdd.n572 Vdd.n568 6.25878
R1480 Vdd.n583 Vdd.n579 6.25878
R1481 Vdd.n578 Vdd.n574 6.25878
R1482 Vdd.n595 Vdd.n591 6.25878
R1483 Vdd.n589 Vdd.n585 6.25878
R1484 Vdd.n602 Vdd.n598 6.25878
R1485 Vdd.n209 Vdd.n208 5.93546
R1486 Vdd.n96 Vdd.n95 5.93546
R1487 Vdd.n169 Vdd.n168 5.93546
R1488 Vdd.n979 Vdd.n978 5.93546
R1489 Vdd.n731 Vdd.n730 5.93546
R1490 Vdd.n434 Vdd.n433 5.93546
R1491 Vdd.n348 Vdd.n347 5.93546
R1492 Vdd.n727 Vdd.n726 5.7305
R1493 SARlogic_0.dffrs_13.nand3_8.B Vdd.n729 5.47979
R1494 SARlogic_0.dffrs_13.nand3_1.B Vdd.n728 5.47979
R1495 Vdd.n7 Vdd.n6 5.44497
R1496 Vdd.n1111 Vdd.n1110 5.44497
R1497 Vdd.n12 Vdd.n11 5.44497
R1498 Vdd.n1099 Vdd.n1098 5.44497
R1499 Vdd.n1105 Vdd.n1104 5.44497
R1500 Vdd.n1092 Vdd.n1091 5.44497
R1501 Vdd.n66 Vdd.n65 5.44497
R1502 Vdd.n78 Vdd.n77 5.44497
R1503 Vdd.n73 Vdd.n72 5.44497
R1504 Vdd.n90 Vdd.n89 5.44497
R1505 Vdd.n84 Vdd.n83 5.44497
R1506 Vdd.n101 Vdd.n100 5.44497
R1507 Vdd.n140 Vdd.n139 5.44497
R1508 Vdd.n151 Vdd.n150 5.44497
R1509 Vdd.n146 Vdd.n145 5.44497
R1510 Vdd.n163 Vdd.n162 5.44497
R1511 Vdd.n157 Vdd.n156 5.44497
R1512 Vdd.n174 Vdd.n173 5.44497
R1513 Vdd.n220 Vdd.n219 5.44497
R1514 Vdd.n225 Vdd.n224 5.44497
R1515 Vdd.n214 Vdd.n213 5.44497
R1516 Vdd.n1017 Vdd.n1016 5.44497
R1517 Vdd.n1000 Vdd.n999 5.44497
R1518 Vdd.n1005 Vdd.n1004 5.44497
R1519 Vdd.n1011 Vdd.n1010 5.44497
R1520 Vdd.n993 Vdd.n992 5.44497
R1521 Vdd.n521 Vdd.n520 5.44497
R1522 Vdd.n527 Vdd.n526 5.44497
R1523 Vdd.n533 Vdd.n532 5.44497
R1524 Vdd.n984 Vdd.n983 5.44497
R1525 Vdd.n770 Vdd.n769 5.44497
R1526 Vdd.n809 Vdd.n808 5.44497
R1527 Vdd.n847 Vdd.n846 5.44497
R1528 Vdd.n885 Vdd.n884 5.44497
R1529 Vdd.n924 Vdd.n923 5.44497
R1530 Vdd.n962 Vdd.n961 5.44497
R1531 Vdd.n688 Vdd.n687 5.44497
R1532 Vdd.n781 Vdd.n780 5.44497
R1533 Vdd.n414 Vdd.n413 5.44497
R1534 Vdd.n820 Vdd.n819 5.44497
R1535 Vdd.n384 Vdd.n383 5.44497
R1536 Vdd.n858 Vdd.n857 5.44497
R1537 Vdd.n354 Vdd.n353 5.44497
R1538 Vdd.n897 Vdd.n896 5.44497
R1539 Vdd.n318 Vdd.n317 5.44497
R1540 Vdd.n935 Vdd.n934 5.44497
R1541 Vdd.n288 Vdd.n287 5.44497
R1542 Vdd.n973 Vdd.n972 5.44497
R1543 Vdd.n765 Vdd.n764 5.44497
R1544 Vdd.n678 Vdd.n677 5.44497
R1545 Vdd.n804 Vdd.n803 5.44497
R1546 Vdd.n404 Vdd.n403 5.44497
R1547 Vdd.n842 Vdd.n841 5.44497
R1548 Vdd.n374 Vdd.n373 5.44497
R1549 Vdd.n880 Vdd.n879 5.44497
R1550 Vdd.n338 Vdd.n337 5.44497
R1551 Vdd.n919 Vdd.n918 5.44497
R1552 Vdd.n308 Vdd.n307 5.44497
R1553 Vdd.n957 Vdd.n956 5.44497
R1554 Vdd.n278 Vdd.n277 5.44497
R1555 Vdd.n693 Vdd.n692 5.44497
R1556 Vdd.n419 Vdd.n418 5.44497
R1557 Vdd.n389 Vdd.n388 5.44497
R1558 Vdd.n359 Vdd.n358 5.44497
R1559 Vdd.n323 Vdd.n322 5.44497
R1560 Vdd.n293 Vdd.n292 5.44497
R1561 Vdd.n760 Vdd.n759 5.44497
R1562 Vdd.n698 Vdd.n697 5.44497
R1563 Vdd.n799 Vdd.n798 5.44497
R1564 Vdd.n776 Vdd.n775 5.44497
R1565 Vdd.n424 Vdd.n423 5.44497
R1566 Vdd.n837 Vdd.n836 5.44497
R1567 Vdd.n815 Vdd.n814 5.44497
R1568 Vdd.n394 Vdd.n393 5.44497
R1569 Vdd.n875 Vdd.n874 5.44497
R1570 Vdd.n853 Vdd.n852 5.44497
R1571 Vdd.n364 Vdd.n363 5.44497
R1572 Vdd.n914 Vdd.n913 5.44497
R1573 Vdd.n892 Vdd.n891 5.44497
R1574 Vdd.n328 Vdd.n327 5.44497
R1575 Vdd.n952 Vdd.n951 5.44497
R1576 Vdd.n930 Vdd.n929 5.44497
R1577 Vdd.n298 Vdd.n297 5.44497
R1578 Vdd.n968 Vdd.n967 5.44497
R1579 Vdd.n755 Vdd.n754 5.44497
R1580 Vdd.n683 Vdd.n682 5.44497
R1581 Vdd.n794 Vdd.n793 5.44497
R1582 Vdd.n409 Vdd.n408 5.44497
R1583 Vdd.n832 Vdd.n831 5.44497
R1584 Vdd.n379 Vdd.n378 5.44497
R1585 Vdd.n870 Vdd.n869 5.44497
R1586 Vdd.n343 Vdd.n342 5.44497
R1587 Vdd.n909 Vdd.n908 5.44497
R1588 Vdd.n313 Vdd.n312 5.44497
R1589 Vdd.n947 Vdd.n946 5.44497
R1590 Vdd.n283 Vdd.n282 5.44497
R1591 Vdd.n703 Vdd.n702 5.44497
R1592 Vdd.n429 Vdd.n428 5.44497
R1593 Vdd.n399 Vdd.n398 5.44497
R1594 Vdd.n369 Vdd.n368 5.44497
R1595 Vdd.n333 Vdd.n332 5.44497
R1596 Vdd.n303 Vdd.n302 5.44497
R1597 Vdd.n708 Vdd.n707 5.44497
R1598 Vdd.n724 Vdd.n723 5.44497
R1599 Vdd.n719 Vdd.n718 5.44497
R1600 Vdd.n742 Vdd.n741 5.44497
R1601 Vdd.n748 Vdd.n747 5.44497
R1602 Vdd.n736 Vdd.n735 5.44497
R1603 Vdd.n641 Vdd.n640 5.44497
R1604 Vdd.n652 Vdd.n651 5.44497
R1605 Vdd.n647 Vdd.n646 5.44497
R1606 Vdd.n664 Vdd.n663 5.44497
R1607 Vdd.n658 Vdd.n657 5.44497
R1608 Vdd.n671 Vdd.n670 5.44497
R1609 Vdd.n572 Vdd.n571 5.44497
R1610 Vdd.n583 Vdd.n582 5.44497
R1611 Vdd.n578 Vdd.n577 5.44497
R1612 Vdd.n595 Vdd.n594 5.44497
R1613 Vdd.n589 Vdd.n588 5.44497
R1614 Vdd.n602 Vdd.n601 5.44497
R1615 Vdd.n48 Vdd.n47 5.14711
R1616 Vdd.n134 Vdd.n133 5.14711
R1617 Vdd.n515 Vdd.n514 5.14711
R1618 Vdd.n787 Vdd.n786 5.14711
R1619 Vdd.n825 Vdd.n824 5.14711
R1620 Vdd.n863 Vdd.n862 5.14711
R1621 Vdd.n902 Vdd.n901 5.14711
R1622 Vdd.n940 Vdd.n939 5.14711
R1623 Vdd.n712 Vdd.n711 5.14711
R1624 Vdd.n566 Vdd.n565 5.14711
R1625 Vdd.n635 Vdd.n634 5.14711
R1626 Vdd.n2 Vdd.n1 5.14711
R1627 Vdd.n785 Vdd.n784 5.13907
R1628 Vdd.n823 Vdd.n822 5.13907
R1629 Vdd.n861 Vdd.n860 5.13907
R1630 Vdd.n900 Vdd.n899 5.13907
R1631 Vdd.n938 Vdd.n937 5.13907
R1632 Vdd.n710 Vdd.n709 5.13907
R1633 Vdd.n730 SARlogic_0.dffrs_13.nand3_8.B 5.09593
R1634 Vdd.n1085 Vdd.n1084 4.98176
R1635 Vdd.n1030 Vdd.t331 4.4205
R1636 Vdd.n1023 Vdd.t595 4.4205
R1637 Vdd.n988 Vdd.n273 4.3905
R1638 Vdd.n1041 Vdd.t752 3.38176
R1639 Vdd.n54 Vdd.t545 3.38176
R1640 Vdd.n191 Vdd.n190 2.49936
R1641 Vdd.n118 Vdd.n117 2.49936
R1642 Vdd.n256 Vdd.n255 2.49936
R1643 Vdd.n619 Vdd.n618 2.49936
R1644 Vdd.n550 Vdd.n549 2.49936
R1645 Vdd.n478 Vdd.n477 2.49936
R1646 Vdd.n1055 Vdd.n1054 2.1905
R1647 Vdd.n1073 Vdd.n1072 2.1905
R1648 Vdd.n1036 Vdd.n1035 2.16583
R1649 Vdd.n1038 Vdd.n1037 2.16583
R1650 Vdd.n53 Vdd.n52 2.16583
R1651 Vdd.n51 Vdd.n50 2.16583
R1652 Vdd.n1022 Vdd.t930 1.99236
R1653 Vdd.n190 Vdd.n179 1.93883
R1654 Vdd.n117 Vdd.n106 1.93883
R1655 Vdd.n255 Vdd.n244 1.93883
R1656 Vdd.n618 Vdd.n607 1.93883
R1657 Vdd.n549 Vdd.n538 1.93883
R1658 Vdd.n477 Vdd.n466 1.93883
R1659 Vdd.n1032 Vdd.t575 1.91107
R1660 Vdd.n994 Vdd.n988 1.89424
R1661 Vdd.n6 Vdd.t677 1.85637
R1662 Vdd.n1110 Vdd.t221 1.85637
R1663 Vdd.n11 Vdd.t698 1.85637
R1664 Vdd.n1098 Vdd.t237 1.85637
R1665 Vdd.n1104 Vdd.t591 1.85637
R1666 Vdd.n1091 Vdd.t217 1.85637
R1667 Vdd.n65 Vdd.t725 1.85637
R1668 Vdd.n77 Vdd.t193 1.85637
R1669 Vdd.n72 Vdd.t614 1.85637
R1670 Vdd.n89 Vdd.t179 1.85637
R1671 Vdd.n83 Vdd.t894 1.85637
R1672 Vdd.n100 Vdd.t115 1.85637
R1673 Vdd.n139 Vdd.t704 1.85637
R1674 Vdd.n150 Vdd.t820 1.85637
R1675 Vdd.n145 Vdd.t716 1.85637
R1676 Vdd.n162 Vdd.t529 1.85637
R1677 Vdd.n156 Vdd.t453 1.85637
R1678 Vdd.n173 Vdd.t810 1.85637
R1679 Vdd.n219 Vdd.t635 1.85637
R1680 Vdd.n224 Vdd.t85 1.85637
R1681 Vdd.n213 Vdd.t846 1.85637
R1682 Vdd.n1016 Vdd.t884 1.85637
R1683 Vdd.n999 Vdd.t848 1.85637
R1684 Vdd.n1004 Vdd.t345 1.85637
R1685 Vdd.n1010 Vdd.t559 1.85637
R1686 Vdd.n992 Vdd.t491 1.85637
R1687 Vdd.n520 Vdd.t620 1.85637
R1688 Vdd.n526 Vdd.t489 1.85637
R1689 Vdd.n532 Vdd.t858 1.85637
R1690 Vdd.n983 Vdd.t333 1.85637
R1691 Vdd.n769 Vdd.t814 1.85637
R1692 Vdd.n808 Vdd.t233 1.85637
R1693 Vdd.n846 Vdd.t371 1.85637
R1694 Vdd.n884 Vdd.t519 1.85637
R1695 Vdd.n923 Vdd.t169 1.85637
R1696 Vdd.n961 Vdd.t255 1.85637
R1697 Vdd.n687 Vdd.t469 1.85637
R1698 Vdd.n780 Vdd.t818 1.85637
R1699 Vdd.n413 Vdd.t455 1.85637
R1700 Vdd.n819 Vdd.t229 1.85637
R1701 Vdd.n383 Vdd.t129 1.85637
R1702 Vdd.n857 Vdd.t369 1.85637
R1703 Vdd.n353 Vdd.t285 1.85637
R1704 Vdd.n896 Vdd.t517 1.85637
R1705 Vdd.n317 Vdd.t123 1.85637
R1706 Vdd.n934 Vdd.t167 1.85637
R1707 Vdd.n287 Vdd.t243 1.85637
R1708 Vdd.n972 Vdd.t257 1.85637
R1709 Vdd.n764 Vdd.t381 1.85637
R1710 Vdd.n677 Vdd.t299 1.85637
R1711 Vdd.n803 Vdd.t579 1.85637
R1712 Vdd.n403 Vdd.t890 1.85637
R1713 Vdd.n841 Vdd.t91 1.85637
R1714 Vdd.n373 Vdd.t101 1.85637
R1715 Vdd.n879 Vdd.t904 1.85637
R1716 Vdd.n337 Vdd.t305 1.85637
R1717 Vdd.n918 Vdd.t291 1.85637
R1718 Vdd.n307 Vdd.t563 1.85637
R1719 Vdd.n956 Vdd.t77 1.85637
R1720 Vdd.n277 Vdd.t946 1.85637
R1721 Vdd.n692 Vdd.t351 1.85637
R1722 Vdd.n418 Vdd.t185 1.85637
R1723 Vdd.n388 Vdd.t187 1.85637
R1724 Vdd.n358 Vdd.t589 1.85637
R1725 Vdd.n322 Vdd.t319 1.85637
R1726 Vdd.n292 Vdd.t253 1.85637
R1727 Vdd.n759 Vdd.t710 1.85637
R1728 Vdd.n697 Vdd.t367 1.85637
R1729 Vdd.n798 Vdd.t617 1.85637
R1730 Vdd.n775 Vdd.t701 1.85637
R1731 Vdd.n423 Vdd.t872 1.85637
R1732 Vdd.n836 Vdd.t665 1.85637
R1733 Vdd.n814 Vdd.t659 1.85637
R1734 Vdd.n393 Vdd.t71 1.85637
R1735 Vdd.n874 Vdd.t713 1.85637
R1736 Vdd.n852 Vdd.t683 1.85637
R1737 Vdd.n363 Vdd.t223 1.85637
R1738 Vdd.n913 Vdd.t674 1.85637
R1739 Vdd.n891 Vdd.t731 1.85637
R1740 Vdd.n327 Vdd.t487 1.85637
R1741 Vdd.n951 Vdd.t719 1.85637
R1742 Vdd.n929 Vdd.t680 1.85637
R1743 Vdd.n297 Vdd.t830 1.85637
R1744 Vdd.n967 Vdd.t695 1.85637
R1745 Vdd.n754 Vdd.t33 1.85637
R1746 Vdd.n682 Vdd.t195 1.85637
R1747 Vdd.n793 Vdd.t147 1.85637
R1748 Vdd.n408 Vdd.t41 1.85637
R1749 Vdd.n831 Vdd.t495 1.85637
R1750 Vdd.n378 Vdd.t477 1.85637
R1751 Vdd.n869 Vdd.t383 1.85637
R1752 Vdd.n342 Vdd.t541 1.85637
R1753 Vdd.n908 Vdd.t109 1.85637
R1754 Vdd.n312 Vdd.t227 1.85637
R1755 Vdd.n946 Vdd.t742 1.85637
R1756 Vdd.n282 Vdd.t465 1.85637
R1757 Vdd.n702 Vdd.t105 1.85637
R1758 Vdd.n428 Vdd.t533 1.85637
R1759 Vdd.n398 Vdd.t918 1.85637
R1760 Vdd.n368 Vdd.t521 1.85637
R1761 Vdd.n332 Vdd.t457 1.85637
R1762 Vdd.n302 Vdd.t463 1.85637
R1763 Vdd.n707 Vdd.t780 1.85637
R1764 Vdd.n723 Vdd.t603 1.85637
R1765 Vdd.n718 Vdd.t778 1.85637
R1766 Vdd.n741 Vdd.t952 1.85637
R1767 Vdd.n747 Vdd.t824 1.85637
R1768 Vdd.n735 Vdd.t31 1.85637
R1769 Vdd.n640 Vdd.t623 1.85637
R1770 Vdd.n651 Vdd.t583 1.85637
R1771 Vdd.n646 Vdd.t662 1.85637
R1772 Vdd.n663 Vdd.t932 1.85637
R1773 Vdd.n657 Vdd.t75 1.85637
R1774 Vdd.n670 Vdd.t551 1.85637
R1775 Vdd.n571 Vdd.t608 1.85637
R1776 Vdd.n582 Vdd.t505 1.85637
R1777 Vdd.n577 Vdd.t629 1.85637
R1778 Vdd.n594 Vdd.t475 1.85637
R1779 Vdd.n588 Vdd.t844 1.85637
R1780 Vdd.n601 Vdd.t315 1.85637
R1781 Vdd.n1081 Vdd.n1033 1.83762
R1782 Vdd.n1083 Vdd.n1022 1.83762
R1783 Vdd.n1065 Vdd.t493 1.8205
R1784 Vdd.n1065 Vdd.t449 1.8205
R1785 Vdd.n1063 Vdd.t928 1.8205
R1786 Vdd.n1063 Vdd.t567 1.8205
R1787 Vdd.n1061 Vdd.t573 1.8205
R1788 Vdd.n1061 Vdd.t445 1.8205
R1789 Vdd.n1059 Vdd.t447 1.8205
R1790 Vdd.n1059 Vdd.t569 1.8205
R1791 Vdd.n1057 Vdd.t571 1.8205
R1792 Vdd.n1057 Vdd.t313 1.8205
R1793 Vdd.n450 Vdd.t375 1.80717
R1794 Vdd.n104 Vdd.n45 1.80479
R1795 Vdd.n177 Vdd.n29 1.80479
R1796 Vdd.n536 Vdd.n512 1.80479
R1797 Vdd.n605 Vdd.n496 1.80479
R1798 Vdd.n480 Vdd.n435 1.80479
R1799 Vdd.n234 Vdd.n13 1.80479
R1800 Vdd.n127 Vdd.n126 1.78583
R1801 Vdd.n200 Vdd.n199 1.78583
R1802 Vdd.n559 Vdd.n558 1.78583
R1803 Vdd.n628 Vdd.n627 1.78583
R1804 Vdd.n463 Vdd.n448 1.78583
R1805 Vdd.n260 Vdd.n259 1.78583
R1806 Vdd.n130 Vdd.t760 1.74654
R1807 Vdd.n203 Vdd.t922 1.74654
R1808 Vdd.n562 Vdd.t768 1.74654
R1809 Vdd.n631 Vdd.t920 1.74654
R1810 Vdd.n451 Vdd.t770 1.74654
R1811 Vdd.n268 Vdd.t758 1.74654
R1812 Vdd.n452 Vdd.n450 1.62809
R1813 Vdd.n1028 Vdd.n1027 1.5755
R1814 Vdd.n1030 Vdd.n1029 1.5755
R1815 Vdd.n1026 Vdd.n1023 1.5755
R1816 Vdd.n1069 Vdd.n1068 1.5755
R1817 Vdd.n1071 Vdd.n1070 1.5755
R1818 Vdd.n15 Vdd.t247 1.49467
R1819 Vdd.n187 Vdd.t197 1.49467
R1820 Vdd.n186 Vdd.t585 1.49467
R1821 Vdd.n31 Vdd.t451 1.49467
R1822 Vdd.n114 Vdd.t263 1.49467
R1823 Vdd.n113 Vdd.t948 1.49467
R1824 Vdd.n30 Vdd.t926 1.49467
R1825 Vdd.n14 Vdd.t766 1.49467
R1826 Vdd.n252 Vdd.t601 1.49467
R1827 Vdd.n251 Vdd.t309 1.49467
R1828 Vdd.n266 Vdd.t874 1.49467
R1829 Vdd.n265 Vdd.t772 1.49467
R1830 Vdd.n482 Vdd.t73 1.49467
R1831 Vdd.n615 Vdd.t756 1.49467
R1832 Vdd.n614 Vdd.t161 1.49467
R1833 Vdd.n498 Vdd.t852 1.49467
R1834 Vdd.n546 Vdd.t151 1.49467
R1835 Vdd.n545 Vdd.t97 1.49467
R1836 Vdd.n497 Vdd.t764 1.49467
R1837 Vdd.n481 Vdd.t762 1.49467
R1838 Vdd.n474 Vdd.t365 1.49467
R1839 Vdd.n473 Vdd.t301 1.49467
R1840 Vdd.n460 Vdd.t13 1.49467
R1841 Vdd.n459 Vdd.t924 1.49467
R1842 Vdd.n180 Vdd.t467 1.47383
R1843 Vdd.n107 Vdd.t503 1.47383
R1844 Vdd.n33 Vdd.t900 1.47383
R1845 Vdd.n34 Vdd.t902 1.47383
R1846 Vdd.n35 Vdd.t842 1.47383
R1847 Vdd.n32 Vdd.t347 1.47383
R1848 Vdd.n17 Vdd.t143 1.47383
R1849 Vdd.n18 Vdd.t141 1.47383
R1850 Vdd.n19 Vdd.t339 1.47383
R1851 Vdd.n16 Vdd.t812 1.47383
R1852 Vdd.n245 Vdd.t205 1.47383
R1853 Vdd.n608 Vdd.t593 1.47383
R1854 Vdd.n539 Vdd.t912 1.47383
R1855 Vdd.n500 Vdd.t886 1.47383
R1856 Vdd.n501 Vdd.t888 1.47383
R1857 Vdd.n502 Vdd.t209 1.47383
R1858 Vdd.n499 Vdd.t806 1.47383
R1859 Vdd.n484 Vdd.t135 1.47383
R1860 Vdd.n485 Vdd.t133 1.47383
R1861 Vdd.n486 Vdd.t235 1.47383
R1862 Vdd.n483 Vdd.t107 1.47383
R1863 Vdd.n467 Vdd.t515 1.47383
R1864 Vdd.n449 Vdd.t191 1.47383
R1865 Vdd.n447 Vdd.t139 1.47383
R1866 Vdd.n437 Vdd.t137 1.47383
R1867 Vdd.n436 Vdd.t776 1.47383
R1868 Vdd.n261 Vdd.t802 1.47383
R1869 Vdd.n230 Vdd.t119 1.47383
R1870 Vdd.n231 Vdd.t121 1.47383
R1871 Vdd.n242 Vdd.t577 1.47383
R1872 Vdd.n176 Vdd.n131 1.19311
R1873 Vdd.n1094 Vdd.n204 1.19311
R1874 Vdd.n597 Vdd.n563 1.19311
R1875 Vdd.n666 Vdd.n632 1.19311
R1876 Vdd.n270 Vdd.n269 1.19311
R1877 Vdd.n1035 Vdd.t750 1.13285
R1878 Vdd.n1035 Vdd.t754 1.13285
R1879 Vdd.n1037 Vdd.t597 1.13285
R1880 Vdd.n1037 Vdd.t748 1.13285
R1881 Vdd.n52 Vdd.t547 1.13285
R1882 Vdd.n52 Vdd.t549 1.13285
R1883 Vdd.n50 Vdd.t892 1.13285
R1884 Vdd.n50 Vdd.t543 1.13285
R1885 Vdd.n1082 Vdd.n1031 1.058
R1886 Vdd.n6 Vdd.n5 1.04105
R1887 Vdd.n1110 Vdd.n1109 1.04105
R1888 Vdd.n11 Vdd.n10 1.04105
R1889 Vdd.n1098 Vdd.n1097 1.04105
R1890 Vdd.n1104 Vdd.n1103 1.04105
R1891 Vdd.n1091 Vdd.n1090 1.04105
R1892 Vdd.n65 Vdd.n64 1.04105
R1893 Vdd.n77 Vdd.n76 1.04105
R1894 Vdd.n72 Vdd.n71 1.04105
R1895 Vdd.n89 Vdd.n88 1.04105
R1896 Vdd.n83 Vdd.n82 1.04105
R1897 Vdd.n100 Vdd.n99 1.04105
R1898 Vdd.n139 Vdd.n138 1.04105
R1899 Vdd.n150 Vdd.n149 1.04105
R1900 Vdd.n145 Vdd.n144 1.04105
R1901 Vdd.n162 Vdd.n161 1.04105
R1902 Vdd.n156 Vdd.n155 1.04105
R1903 Vdd.n173 Vdd.n172 1.04105
R1904 Vdd.n219 Vdd.n218 1.04105
R1905 Vdd.n224 Vdd.n223 1.04105
R1906 Vdd.n213 Vdd.n212 1.04105
R1907 Vdd.n1016 Vdd.n1015 1.04105
R1908 Vdd.n999 Vdd.n998 1.04105
R1909 Vdd.n1004 Vdd.n1003 1.04105
R1910 Vdd.n1010 Vdd.n1009 1.04105
R1911 Vdd.n992 Vdd.n991 1.04105
R1912 Vdd.n520 Vdd.n519 1.04105
R1913 Vdd.n526 Vdd.n525 1.04105
R1914 Vdd.n532 Vdd.n531 1.04105
R1915 Vdd.n983 Vdd.n982 1.04105
R1916 Vdd.n769 Vdd.n768 1.04105
R1917 Vdd.n808 Vdd.n807 1.04105
R1918 Vdd.n846 Vdd.n845 1.04105
R1919 Vdd.n884 Vdd.n883 1.04105
R1920 Vdd.n923 Vdd.n922 1.04105
R1921 Vdd.n961 Vdd.n960 1.04105
R1922 Vdd.n687 Vdd.n686 1.04105
R1923 Vdd.n780 Vdd.n779 1.04105
R1924 Vdd.n413 Vdd.n412 1.04105
R1925 Vdd.n819 Vdd.n818 1.04105
R1926 Vdd.n383 Vdd.n382 1.04105
R1927 Vdd.n857 Vdd.n856 1.04105
R1928 Vdd.n353 Vdd.n352 1.04105
R1929 Vdd.n896 Vdd.n895 1.04105
R1930 Vdd.n317 Vdd.n316 1.04105
R1931 Vdd.n934 Vdd.n933 1.04105
R1932 Vdd.n287 Vdd.n286 1.04105
R1933 Vdd.n972 Vdd.n971 1.04105
R1934 Vdd.n764 Vdd.n763 1.04105
R1935 Vdd.n677 Vdd.n676 1.04105
R1936 Vdd.n803 Vdd.n802 1.04105
R1937 Vdd.n403 Vdd.n402 1.04105
R1938 Vdd.n841 Vdd.n840 1.04105
R1939 Vdd.n373 Vdd.n372 1.04105
R1940 Vdd.n879 Vdd.n878 1.04105
R1941 Vdd.n337 Vdd.n336 1.04105
R1942 Vdd.n918 Vdd.n917 1.04105
R1943 Vdd.n307 Vdd.n306 1.04105
R1944 Vdd.n956 Vdd.n955 1.04105
R1945 Vdd.n277 Vdd.n276 1.04105
R1946 Vdd.n692 Vdd.n691 1.04105
R1947 Vdd.n418 Vdd.n417 1.04105
R1948 Vdd.n388 Vdd.n387 1.04105
R1949 Vdd.n358 Vdd.n357 1.04105
R1950 Vdd.n322 Vdd.n321 1.04105
R1951 Vdd.n292 Vdd.n291 1.04105
R1952 Vdd.n759 Vdd.n758 1.04105
R1953 Vdd.n697 Vdd.n696 1.04105
R1954 Vdd.n798 Vdd.n797 1.04105
R1955 Vdd.n775 Vdd.n774 1.04105
R1956 Vdd.n423 Vdd.n422 1.04105
R1957 Vdd.n836 Vdd.n835 1.04105
R1958 Vdd.n814 Vdd.n813 1.04105
R1959 Vdd.n393 Vdd.n392 1.04105
R1960 Vdd.n874 Vdd.n873 1.04105
R1961 Vdd.n852 Vdd.n851 1.04105
R1962 Vdd.n363 Vdd.n362 1.04105
R1963 Vdd.n913 Vdd.n912 1.04105
R1964 Vdd.n891 Vdd.n890 1.04105
R1965 Vdd.n327 Vdd.n326 1.04105
R1966 Vdd.n951 Vdd.n950 1.04105
R1967 Vdd.n929 Vdd.n928 1.04105
R1968 Vdd.n297 Vdd.n296 1.04105
R1969 Vdd.n967 Vdd.n966 1.04105
R1970 Vdd.n754 Vdd.n753 1.04105
R1971 Vdd.n682 Vdd.n681 1.04105
R1972 Vdd.n793 Vdd.n792 1.04105
R1973 Vdd.n408 Vdd.n407 1.04105
R1974 Vdd.n831 Vdd.n830 1.04105
R1975 Vdd.n378 Vdd.n377 1.04105
R1976 Vdd.n869 Vdd.n868 1.04105
R1977 Vdd.n342 Vdd.n341 1.04105
R1978 Vdd.n908 Vdd.n907 1.04105
R1979 Vdd.n312 Vdd.n311 1.04105
R1980 Vdd.n946 Vdd.n945 1.04105
R1981 Vdd.n282 Vdd.n281 1.04105
R1982 Vdd.n702 Vdd.n701 1.04105
R1983 Vdd.n428 Vdd.n427 1.04105
R1984 Vdd.n398 Vdd.n397 1.04105
R1985 Vdd.n368 Vdd.n367 1.04105
R1986 Vdd.n332 Vdd.n331 1.04105
R1987 Vdd.n302 Vdd.n301 1.04105
R1988 Vdd.n707 Vdd.n706 1.04105
R1989 Vdd.n723 Vdd.n722 1.04105
R1990 Vdd.n718 Vdd.n717 1.04105
R1991 Vdd.n741 Vdd.n740 1.04105
R1992 Vdd.n747 Vdd.n746 1.04105
R1993 Vdd.n735 Vdd.n734 1.04105
R1994 Vdd.n640 Vdd.n639 1.04105
R1995 Vdd.n651 Vdd.n650 1.04105
R1996 Vdd.n646 Vdd.n645 1.04105
R1997 Vdd.n663 Vdd.n662 1.04105
R1998 Vdd.n657 Vdd.n656 1.04105
R1999 Vdd.n670 Vdd.n669 1.04105
R2000 Vdd.n571 Vdd.n570 1.04105
R2001 Vdd.n582 Vdd.n581 1.04105
R2002 Vdd.n577 Vdd.n576 1.04105
R2003 Vdd.n594 Vdd.n593 1.04105
R2004 Vdd.n588 Vdd.n587 1.04105
R2005 Vdd.n601 Vdd.n600 1.04105
R2006 Vdd.n1031 Vdd.n1023 1.01373
R2007 Vdd.n1031 Vdd.n1030 0.979984
R2008 Vdd.n104 Vdd.n103 0.809622
R2009 Vdd.n177 Vdd.n176 0.809622
R2010 Vdd.n536 Vdd.n535 0.809622
R2011 Vdd.n605 Vdd.n604 0.809622
R2012 Vdd.n666 Vdd.n480 0.809622
R2013 Vdd.n1094 Vdd.n13 0.809622
R2014 Vdd.n183 Vdd.n180 0.788
R2015 Vdd.n184 Vdd.n183 0.788
R2016 Vdd.n186 Vdd.n185 0.788
R2017 Vdd.n110 Vdd.n107 0.788
R2018 Vdd.n111 Vdd.n110 0.788
R2019 Vdd.n113 Vdd.n112 0.788
R2020 Vdd.n41 Vdd.n34 0.788
R2021 Vdd.n42 Vdd.n41 0.788
R2022 Vdd.n43 Vdd.n35 0.788
R2023 Vdd.n44 Vdd.n43 0.788
R2024 Vdd.n39 Vdd.n33 0.788
R2025 Vdd.n124 Vdd.n32 0.788
R2026 Vdd.n125 Vdd.n124 0.788
R2027 Vdd.n123 Vdd.n30 0.788
R2028 Vdd.n25 Vdd.n18 0.788
R2029 Vdd.n26 Vdd.n25 0.788
R2030 Vdd.n27 Vdd.n19 0.788
R2031 Vdd.n28 Vdd.n27 0.788
R2032 Vdd.n23 Vdd.n17 0.788
R2033 Vdd.n197 Vdd.n16 0.788
R2034 Vdd.n198 Vdd.n197 0.788
R2035 Vdd.n196 Vdd.n14 0.788
R2036 Vdd.n248 Vdd.n245 0.788
R2037 Vdd.n249 Vdd.n248 0.788
R2038 Vdd.n251 Vdd.n250 0.788
R2039 Vdd.n611 Vdd.n608 0.788
R2040 Vdd.n612 Vdd.n611 0.788
R2041 Vdd.n614 Vdd.n613 0.788
R2042 Vdd.n542 Vdd.n539 0.788
R2043 Vdd.n543 Vdd.n542 0.788
R2044 Vdd.n545 Vdd.n544 0.788
R2045 Vdd.n508 Vdd.n501 0.788
R2046 Vdd.n509 Vdd.n508 0.788
R2047 Vdd.n510 Vdd.n502 0.788
R2048 Vdd.n511 Vdd.n510 0.788
R2049 Vdd.n506 Vdd.n500 0.788
R2050 Vdd.n556 Vdd.n499 0.788
R2051 Vdd.n557 Vdd.n556 0.788
R2052 Vdd.n555 Vdd.n497 0.788
R2053 Vdd.n492 Vdd.n485 0.788
R2054 Vdd.n493 Vdd.n492 0.788
R2055 Vdd.n494 Vdd.n486 0.788
R2056 Vdd.n495 Vdd.n494 0.788
R2057 Vdd.n490 Vdd.n484 0.788
R2058 Vdd.n625 Vdd.n483 0.788
R2059 Vdd.n626 Vdd.n625 0.788
R2060 Vdd.n624 Vdd.n481 0.788
R2061 Vdd.n470 Vdd.n467 0.788
R2062 Vdd.n471 Vdd.n470 0.788
R2063 Vdd.n473 Vdd.n472 0.788
R2064 Vdd.n456 Vdd.n449 0.788
R2065 Vdd.n457 Vdd.n456 0.788
R2066 Vdd.n459 Vdd.n458 0.788
R2067 Vdd.n444 Vdd.n437 0.788
R2068 Vdd.n445 Vdd.n444 0.788
R2069 Vdd.n442 Vdd.n436 0.788
R2070 Vdd.n443 Vdd.n442 0.788
R2071 Vdd.n447 Vdd.n446 0.788
R2072 Vdd.n262 Vdd.n261 0.788
R2073 Vdd.n263 Vdd.n262 0.788
R2074 Vdd.n265 Vdd.n264 0.788
R2075 Vdd.n238 Vdd.n231 0.788
R2076 Vdd.n239 Vdd.n238 0.788
R2077 Vdd.n242 Vdd.n241 0.788
R2078 Vdd.n241 Vdd.n240 0.788
R2079 Vdd.n236 Vdd.n230 0.788
R2080 Vdd.n49 Vdd.n48 0.754571
R2081 Vdd.n135 Vdd.n134 0.754571
R2082 Vdd.n516 Vdd.n515 0.754571
R2083 Vdd.n567 Vdd.n566 0.754571
R2084 Vdd.n636 Vdd.n635 0.754571
R2085 Vdd.n1114 Vdd.n2 0.754571
R2086 Vdd.n1080 Vdd.n1045 0.750875
R2087 Vdd.n3 Vdd.t239 0.7285
R2088 Vdd.n3 Vdd.t836 0.7285
R2089 Vdd.n1107 Vdd.t880 0.7285
R2090 Vdd.n1107 Vdd.t668 0.7285
R2091 Vdd.n8 Vdd.t337 0.7285
R2092 Vdd.n8 Vdd.t241 0.7285
R2093 Vdd.n1095 Vdd.t838 0.7285
R2094 Vdd.n1095 Vdd.t878 0.7285
R2095 Vdd.n1101 Vdd.t671 0.7285
R2096 Vdd.n1101 Vdd.t219 0.7285
R2097 Vdd.n1088 Vdd.t828 0.7285
R2098 Vdd.n1088 Vdd.t707 0.7285
R2099 Vdd.n62 Vdd.t175 0.7285
R2100 Vdd.n62 Vdd.t898 0.7285
R2101 Vdd.n74 Vdd.t862 0.7285
R2102 Vdd.n74 Vdd.t611 0.7285
R2103 Vdd.n69 Vdd.t513 0.7285
R2104 Vdd.n69 Vdd.t177 0.7285
R2105 Vdd.n86 Vdd.t896 0.7285
R2106 Vdd.n86 Vdd.t866 0.7285
R2107 Vdd.n80 Vdd.t653 0.7285
R2108 Vdd.n80 Vdd.t832 0.7285
R2109 Vdd.n97 Vdd.t834 0.7285
R2110 Vdd.n97 Vdd.t647 0.7285
R2111 Vdd.n136 Vdd.t525 0.7285
R2112 Vdd.n136 Vdd.t509 0.7285
R2113 Vdd.n147 Vdd.t876 0.7285
R2114 Vdd.n147 Vdd.t734 0.7285
R2115 Vdd.n142 Vdd.t605 0.7285
R2116 Vdd.n142 Vdd.t527 0.7285
R2117 Vdd.n159 Vdd.t511 0.7285
R2118 Vdd.n159 Vdd.t870 0.7285
R2119 Vdd.n153 Vdd.t740 0.7285
R2120 Vdd.n153 Vdd.t808 0.7285
R2121 Vdd.n170 Vdd.t501 0.7285
R2122 Vdd.n170 Vdd.t632 0.7285
R2123 Vdd.n216 Vdd.t481 0.7285
R2124 Vdd.n216 Vdd.t860 0.7285
R2125 Vdd.n221 Vdd.t656 0.7285
R2126 Vdd.n221 Vdd.t335 0.7285
R2127 Vdd.n210 Vdd.t343 0.7285
R2128 Vdd.n210 Vdd.t23 0.7285
R2129 Vdd.n1013 Vdd.t19 0.7285
R2130 Vdd.n1013 Vdd.t427 0.7285
R2131 Vdd.n996 Vdd.t153 0.7285
R2132 Vdd.n996 Vdd.t297 0.7285
R2133 Vdd.n1001 Vdd.t21 0.7285
R2134 Vdd.n1001 Vdd.t15 0.7285
R2135 Vdd.n1007 Vdd.t395 0.7285
R2136 Vdd.n1007 Vdd.t940 0.7285
R2137 Vdd.n989 Vdd.t11 0.7285
R2138 Vdd.n989 Vdd.t431 0.7285
R2139 Vdd.n517 Vdd.t856 0.7285
R2140 Vdd.n517 Vdd.t910 0.7285
R2141 Vdd.n523 Vdd.t273 0.7285
R2142 Vdd.n523 Vdd.t650 0.7285
R2143 Vdd.n529 Vdd.t329 0.7285
R2144 Vdd.n529 Vdd.t882 0.7285
R2145 Vdd.n980 Vdd.t267 0.7285
R2146 Vdd.n980 Vdd.t692 0.7285
R2147 Vdd.n766 Vdd.t379 0.7285
R2148 Vdd.n766 Vdd.t27 0.7285
R2149 Vdd.n805 Vdd.t303 0.7285
R2150 Vdd.n805 Vdd.t277 0.7285
R2151 Vdd.n843 Vdd.t87 0.7285
R2152 Vdd.n843 Vdd.t327 0.7285
R2153 Vdd.n881 Vdd.t906 0.7285
R2154 Vdd.n881 Vdd.t155 0.7285
R2155 Vdd.n920 Vdd.t287 0.7285
R2156 Vdd.n920 Vdd.t353 0.7285
R2157 Vdd.n958 Vdd.t81 0.7285
R2158 Vdd.n958 Vdd.t171 0.7285
R2159 Vdd.n684 Vdd.t163 0.7285
R2160 Vdd.n684 Vdd.t507 0.7285
R2161 Vdd.n777 Vdd.t341 0.7285
R2162 Vdd.n777 Vdd.t377 0.7285
R2163 Vdd.n410 Vdd.t99 0.7285
R2164 Vdd.n410 Vdd.t439 0.7285
R2165 Vdd.n816 Vdd.t265 0.7285
R2166 Vdd.n816 Vdd.t581 0.7285
R2167 Vdd.n380 Vdd.t307 0.7285
R2168 Vdd.n380 Vdd.t429 0.7285
R2169 Vdd.n854 Vdd.t131 0.7285
R2170 Vdd.n854 Vdd.t89 0.7285
R2171 Vdd.n350 Vdd.t565 0.7285
R2172 Vdd.n350 Vdd.t407 0.7285
R2173 Vdd.n893 Vdd.t822 0.7285
R2174 Vdd.n893 Vdd.t908 0.7285
R2175 Vdd.n314 Vdd.t944 0.7285
R2176 Vdd.n314 Vdd.t800 0.7285
R2177 Vdd.n931 Vdd.t127 0.7285
R2178 Vdd.n931 Vdd.t289 0.7285
R2179 Vdd.n284 Vdd.t557 0.7285
R2180 Vdd.n284 Vdd.t788 0.7285
R2181 Vdd.n969 Vdd.t245 0.7285
R2182 Vdd.n969 Vdd.t79 0.7285
R2183 Vdd.n761 Vdd.t25 0.7285
R2184 Vdd.n761 Vdd.t165 0.7285
R2185 Vdd.n674 Vdd.t435 0.7285
R2186 Vdd.n674 Vdd.t349 0.7285
R2187 Vdd.n800 Vdd.t279 0.7285
R2188 Vdd.n800 Vdd.t103 0.7285
R2189 Vdd.n400 Vdd.t415 0.7285
R2190 Vdd.n400 Vdd.t183 0.7285
R2191 Vdd.n838 Vdd.t325 0.7285
R2192 Vdd.n838 Vdd.t311 0.7285
R2193 Vdd.n370 Vdd.t397 0.7285
R2194 Vdd.n370 Vdd.t189 0.7285
R2195 Vdd.n876 Vdd.t157 0.7285
R2196 Vdd.n876 Vdd.t561 0.7285
R2197 Vdd.n334 Vdd.t401 0.7285
R2198 Vdd.n334 Vdd.t587 0.7285
R2199 Vdd.n915 Vdd.t355 0.7285
R2200 Vdd.n915 Vdd.t950 0.7285
R2201 Vdd.n304 Vdd.t391 0.7285
R2202 Vdd.n304 Vdd.t321 0.7285
R2203 Vdd.n953 Vdd.t173 0.7285
R2204 Vdd.n953 Vdd.t555 0.7285
R2205 Vdd.n274 Vdd.t784 0.7285
R2206 Vdd.n274 Vdd.t251 0.7285
R2207 Vdd.n689 Vdd.t363 0.7285
R2208 Vdd.n689 Vdd.t423 0.7285
R2209 Vdd.n415 Vdd.t357 0.7285
R2210 Vdd.n415 Vdd.t393 0.7285
R2211 Vdd.n385 Vdd.t261 0.7285
R2212 Vdd.n385 Vdd.t443 0.7285
R2213 Vdd.n355 Vdd.t361 0.7285
R2214 Vdd.n355 Vdd.t413 0.7285
R2215 Vdd.n319 Vdd.t259 0.7285
R2216 Vdd.n319 Vdd.t419 0.7285
R2217 Vdd.n289 Vdd.t359 0.7285
R2218 Vdd.n289 Vdd.t796 0.7285
R2219 Vdd.n756 Vdd.t35 0.7285
R2220 Vdd.n756 Vdd.t117 0.7285
R2221 Vdd.n694 Vdd.t47 0.7285
R2222 Vdd.n694 Vdd.t441 0.7285
R2223 Vdd.n795 Vdd.t149 0.7285
R2224 Vdd.n795 Vdd.t211 0.7285
R2225 Vdd.n772 Vdd.t231 0.7285
R2226 Vdd.n772 Vdd.t37 0.7285
R2227 Vdd.n420 Vdd.t3 0.7285
R2228 Vdd.n420 Vdd.t411 0.7285
R2229 Vdd.n833 Vdd.t499 0.7285
R2230 Vdd.n833 Vdd.t271 0.7285
R2231 Vdd.n811 Vdd.t373 0.7285
R2232 Vdd.n811 Vdd.t145 0.7285
R2233 Vdd.n390 Vdd.t61 0.7285
R2234 Vdd.n390 Vdd.t403 0.7285
R2235 Vdd.n871 Vdd.t385 0.7285
R2236 Vdd.n871 Vdd.t537 0.7285
R2237 Vdd.n849 Vdd.t840 0.7285
R2238 Vdd.n849 Vdd.t497 0.7285
R2239 Vdd.n360 Vdd.t43 0.7285
R2240 Vdd.n360 Vdd.t798 0.7285
R2241 Vdd.n910 Vdd.t111 0.7285
R2242 Vdd.n910 Vdd.t483 0.7285
R2243 Vdd.n888 Vdd.t181 0.7285
R2244 Vdd.n888 Vdd.t387 0.7285
R2245 Vdd.n324 Vdd.t55 0.7285
R2246 Vdd.n324 Vdd.t433 0.7285
R2247 Vdd.n948 Vdd.t746 0.7285
R2248 Vdd.n948 Vdd.t804 0.7285
R2249 Vdd.n926 Vdd.t942 0.7285
R2250 Vdd.n926 Vdd.t113 0.7285
R2251 Vdd.n294 Vdd.t7 0.7285
R2252 Vdd.n294 Vdd.t425 0.7285
R2253 Vdd.n964 Vdd.t850 0.7285
R2254 Vdd.n964 Vdd.t744 0.7285
R2255 Vdd.n751 Vdd.t125 0.7285
R2256 Vdd.n751 Vdd.t51 0.7285
R2257 Vdd.n679 Vdd.t405 0.7285
R2258 Vdd.n679 Vdd.t83 0.7285
R2259 Vdd.n790 Vdd.t213 0.7285
R2260 Vdd.n790 Vdd.t65 0.7285
R2261 Vdd.n405 Vdd.t417 0.7285
R2262 Vdd.n405 Vdd.t531 0.7285
R2263 Vdd.n828 Vdd.t269 0.7285
R2264 Vdd.n828 Vdd.t63 0.7285
R2265 Vdd.n375 Vdd.t786 0.7285
R2266 Vdd.n375 Vdd.t916 0.7285
R2267 Vdd.n866 Vdd.t535 0.7285
R2268 Vdd.n866 Vdd.t9 0.7285
R2269 Vdd.n339 Vdd.t790 0.7285
R2270 Vdd.n339 Vdd.t523 0.7285
R2271 Vdd.n905 Vdd.t485 0.7285
R2272 Vdd.n905 Vdd.t49 0.7285
R2273 Vdd.n309 Vdd.t782 0.7285
R2274 Vdd.n309 Vdd.t459 0.7285
R2275 Vdd.n943 Vdd.t207 0.7285
R2276 Vdd.n943 Vdd.t45 0.7285
R2277 Vdd.n279 Vdd.t421 0.7285
R2278 Vdd.n279 Vdd.t461 0.7285
R2279 Vdd.n699 Vdd.t826 0.7285
R2280 Vdd.n699 Vdd.t437 0.7285
R2281 Vdd.n425 Vdd.t774 0.7285
R2282 Vdd.n425 Vdd.t409 0.7285
R2283 Vdd.n395 Vdd.t39 0.7285
R2284 Vdd.n395 Vdd.t794 0.7285
R2285 Vdd.n365 Vdd.t479 0.7285
R2286 Vdd.n365 Vdd.t399 0.7285
R2287 Vdd.n329 Vdd.t539 0.7285
R2288 Vdd.n329 Vdd.t389 0.7285
R2289 Vdd.n299 Vdd.t225 0.7285
R2290 Vdd.n299 Vdd.t792 0.7285
R2291 Vdd.n704 Vdd.t954 0.7285
R2292 Vdd.n704 Vdd.t95 0.7285
R2293 Vdd.n720 Vdd.t69 0.7285
R2294 Vdd.n720 Vdd.t626 0.7285
R2295 Vdd.n715 Vdd.t816 0.7285
R2296 Vdd.n715 Vdd.t854 0.7285
R2297 Vdd.n738 Vdd.t93 0.7285
R2298 Vdd.n738 Vdd.t5 0.7285
R2299 Vdd.n744 Vdd.t728 0.7285
R2300 Vdd.n744 Vdd.t203 0.7285
R2301 Vdd.n732 Vdd.t17 0.7285
R2302 Vdd.n732 Vdd.t722 0.7285
R2303 Vdd.n637 Vdd.t936 0.7285
R2304 Vdd.n637 Vdd.t295 0.7285
R2305 Vdd.n648 Vdd.t275 0.7285
R2306 Vdd.n648 Vdd.t641 0.7285
R2307 Vdd.n643 Vdd.t1 0.7285
R2308 Vdd.n643 Vdd.t934 0.7285
R2309 Vdd.n660 Vdd.t293 0.7285
R2310 Vdd.n660 Vdd.t868 0.7285
R2311 Vdd.n654 Vdd.t737 0.7285
R2312 Vdd.n654 Vdd.t553 0.7285
R2313 Vdd.n667 Vdd.t199 0.7285
R2314 Vdd.n667 Vdd.t686 0.7285
R2315 Vdd.n568 Vdd.t471 0.7285
R2316 Vdd.n568 Vdd.t201 0.7285
R2317 Vdd.n579 Vdd.t938 0.7285
R2318 Vdd.n579 Vdd.t644 0.7285
R2319 Vdd.n574 Vdd.t159 0.7285
R2320 Vdd.n574 Vdd.t473 0.7285
R2321 Vdd.n591 Vdd.t914 0.7285
R2322 Vdd.n591 Vdd.t864 0.7285
R2323 Vdd.n585 Vdd.t638 0.7285
R2324 Vdd.n585 Vdd.t317 0.7285
R2325 Vdd.n598 Vdd.t215 0.7285
R2326 Vdd.n598 Vdd.t689 0.7285
R2327 Vdd.n788 SARlogic_0.dffrs_1.nand3_0.C 0.717607
R2328 Vdd.n826 SARlogic_0.dffrs_2.nand3_0.C 0.717607
R2329 Vdd.n864 SARlogic_0.dffrs_3.nand3_0.C 0.717607
R2330 Vdd.n903 SARlogic_0.dffrs_4.nand3_0.C 0.717607
R2331 Vdd.n941 SARlogic_0.dffrs_5.nand3_0.C 0.717607
R2332 Vdd.n713 SARlogic_0.dffrs_0.nand3_0.C 0.717607
R2333 Vdd.n1060 Vdd.n1058 0.667
R2334 Vdd.n1066 Vdd.n1064 0.662
R2335 Vdd.n1062 Vdd.n1060 0.643429
R2336 Vdd.n1064 Vdd.n1062 0.638429
R2337 Vdd.n1075 Vdd.n1074 0.58325
R2338 Vdd.n1056 Vdd.n1053 0.58325
R2339 Vdd.n189 Vdd.n180 0.561043
R2340 Vdd.n116 Vdd.n107 0.561043
R2341 Vdd.n120 Vdd.n33 0.561043
R2342 Vdd.n119 Vdd.n34 0.561043
R2343 Vdd.n105 Vdd.n35 0.561043
R2344 Vdd.n128 Vdd.n32 0.561043
R2345 Vdd.n193 Vdd.n17 0.561043
R2346 Vdd.n192 Vdd.n18 0.561043
R2347 Vdd.n178 Vdd.n19 0.561043
R2348 Vdd.n201 Vdd.n16 0.561043
R2349 Vdd.n254 Vdd.n245 0.561043
R2350 Vdd.n617 Vdd.n608 0.561043
R2351 Vdd.n548 Vdd.n539 0.561043
R2352 Vdd.n552 Vdd.n500 0.561043
R2353 Vdd.n551 Vdd.n501 0.561043
R2354 Vdd.n537 Vdd.n502 0.561043
R2355 Vdd.n560 Vdd.n499 0.561043
R2356 Vdd.n621 Vdd.n484 0.561043
R2357 Vdd.n620 Vdd.n485 0.561043
R2358 Vdd.n606 Vdd.n486 0.561043
R2359 Vdd.n629 Vdd.n483 0.561043
R2360 Vdd.n476 Vdd.n467 0.561043
R2361 Vdd.n462 Vdd.n449 0.561043
R2362 Vdd.n464 Vdd.n447 0.561043
R2363 Vdd.n465 Vdd.n437 0.561043
R2364 Vdd.n479 Vdd.n436 0.561043
R2365 Vdd.n261 Vdd.n227 0.561043
R2366 Vdd.n258 Vdd.n230 0.561043
R2367 Vdd.n257 Vdd.n231 0.561043
R2368 Vdd.n243 Vdd.n242 0.561043
R2369 Vdd.n131 Vdd.n129 0.490037
R2370 Vdd.n204 Vdd.n202 0.490037
R2371 Vdd.n563 Vdd.n561 0.490037
R2372 Vdd.n632 Vdd.n630 0.490037
R2373 Vdd.n269 Vdd.n267 0.490037
R2374 Vdd.n1058 Vdd.n1046 0.47525
R2375 Vdd.n1067 Vdd.n1066 0.47525
R2376 Vdd.n131 Vdd.n130 0.436534
R2377 Vdd.n204 Vdd.n203 0.436534
R2378 Vdd.n563 Vdd.n562 0.436534
R2379 Vdd.n632 Vdd.n631 0.436534
R2380 Vdd.n269 Vdd.n268 0.436534
R2381 Vdd.n461 Vdd.n453 0.415037
R2382 Vdd.n771 Vdd.n750 0.403945
R2383 Vdd.n452 Vdd.n451 0.3862
R2384 Vdd.n1080 Vdd.n1079 0.381816
R2385 Vdd.n1078 Vdd.n1075 0.34025
R2386 Vdd.n1074 Vdd.n1046 0.34025
R2387 Vdd.n1067 Vdd.n1056 0.34025
R2388 Vdd.n1084 Vdd.n1083 0.313132
R2389 Vdd.n1083 Vdd.n1082 0.289447
R2390 Vdd.n1082 Vdd.n1081 0.279974
R2391 Vdd.n1086 Vdd.n1085 0.265225
R2392 Vdd.n1081 Vdd.n1080 0.256289
R2393 Vdd.n189 Vdd.n188 0.255737
R2394 Vdd.n116 Vdd.n115 0.255737
R2395 Vdd.n129 Vdd.n128 0.255737
R2396 Vdd.n202 Vdd.n201 0.255737
R2397 Vdd.n254 Vdd.n253 0.255737
R2398 Vdd.n617 Vdd.n616 0.255737
R2399 Vdd.n548 Vdd.n547 0.255737
R2400 Vdd.n561 Vdd.n560 0.255737
R2401 Vdd.n630 Vdd.n629 0.255737
R2402 Vdd.n476 Vdd.n475 0.255737
R2403 Vdd.n462 Vdd.n461 0.255737
R2404 Vdd.n267 Vdd.n227 0.255737
R2405 Vdd.n271 Vdd.n215 0.236406
R2406 Vdd.n128 Vdd.n127 0.2165
R2407 Vdd.n201 Vdd.n200 0.2165
R2408 Vdd.n560 Vdd.n559 0.2165
R2409 Vdd.n629 Vdd.n628 0.2165
R2410 Vdd.n463 Vdd.n462 0.2165
R2411 Vdd.n259 Vdd.n227 0.2165
R2412 Vdd.n1032 comparator_no_offsetcal_0.x3.avdd 0.207699
R2413 Vdd.n1079 comparator_no_offsetcal_0.VDD 0.193526
R2414 Vdd.n987 Vdd.n986 0.165959
R2415 Vdd.n1085 Vdd 0.162037
R2416 Vdd.n58 Vdd.n57 0.154786
R2417 Vdd.n127 Vdd.n120 0.148424
R2418 Vdd.n200 Vdd.n193 0.148424
R2419 Vdd.n559 Vdd.n552 0.148424
R2420 Vdd.n628 Vdd.n621 0.148424
R2421 Vdd.n464 Vdd.n463 0.148424
R2422 Vdd.n259 Vdd.n258 0.148424
R2423 adc_PISO_0.dffrs_3.resetb Vdd.n209 0.136036
R2424 adc_PISO_0.dffrs_5.resetb Vdd.n96 0.136036
R2425 adc_PISO_0.dffrs_4.resetb Vdd.n169 0.136036
R2426 adc_PISO_0.dffrs_2.resetb Vdd.n979 0.136036
R2427 SARlogic_0.dffrs_13.resetb Vdd.n731 0.136036
R2428 adc_PISO_0.dffrs_0.resetb Vdd.n434 0.136036
R2429 adc_PISO_0.dffrs_1.resetb Vdd.n348 0.136036
R2430 Vdd.n1041 Vdd.n1036 0.1355
R2431 Vdd.n54 Vdd.n53 0.1355
R2432 Vdd.n453 Vdd.n452 0.124324
R2433 Vdd.n1039 Vdd.n1038 0.109786
R2434 Vdd.n1045 Vdd.n1034 0.103357
R2435 Vdd.n534 Vdd.n528 0.101647
R2436 Vdd.n1086 Vdd.n1020 0.0967961
R2437 Vdd.n1033 Vdd.n1032 0.0965492
R2438 Vdd.n986 Vdd.n985 0.0898578
R2439 Vdd.n988 Vdd.n272 0.0817571
R2440 Vdd.n60 Vdd.n51 0.0802199
R2441 Vdd.n535 Vdd.n534 0.0720596
R2442 Vdd.n1087 Vdd.n1086 0.0680047
R2443 Vdd.n887 Vdd.n349 0.0660636
R2444 Vdd.n190 Vdd.n189 0.0635
R2445 Vdd.n117 Vdd.n116 0.0635
R2446 Vdd.n255 Vdd.n254 0.0635
R2447 Vdd.n618 Vdd.n617 0.0635
R2448 Vdd.n549 Vdd.n548 0.0635
R2449 Vdd.n477 Vdd.n476 0.0635
R2450 Vdd.n270 Vdd.n226 0.0597785
R2451 Vdd.n528 Vdd.n522 0.0590321
R2452 Vdd.n1045 Vdd.n1044 0.0519286
R2453 Vdd.n1038 Vdd.n1034 0.0455
R2454 Vdd.n58 Vdd.n51 0.0455
R2455 Vdd.n785 SARlogic_0.dffrs_1.nand3_2.C 0.0455
R2456 Vdd.n823 SARlogic_0.dffrs_2.nand3_2.C 0.0455
R2457 Vdd.n861 SARlogic_0.dffrs_3.nand3_2.C 0.0455
R2458 Vdd.n900 SARlogic_0.dffrs_4.nand3_2.C 0.0455
R2459 Vdd.n938 SARlogic_0.dffrs_5.nand3_2.C 0.0455
R2460 Vdd.n710 SARlogic_0.dffrs_0.nand3_2.C 0.0455
R2461 Vdd.n727 SARlogic_0.dffrs_13.nand3_7.A 0.0455
R2462 Vdd.n120 Vdd.n119 0.0452384
R2463 Vdd.n193 Vdd.n192 0.0452384
R2464 Vdd.n552 Vdd.n551 0.0452384
R2465 Vdd.n621 Vdd.n620 0.0452384
R2466 Vdd.n465 Vdd.n464 0.0452384
R2467 Vdd.n258 Vdd.n257 0.0452384
R2468 Vdd.n85 Vdd.n79 0.0405727
R2469 Vdd.n158 Vdd.n152 0.0405727
R2470 Vdd.n590 Vdd.n584 0.0405727
R2471 Vdd.n659 Vdd.n653 0.0405727
R2472 Vdd.n1112 Vdd.n1106 0.0405727
R2473 SARlogic_0.dffrs_1.nand3_0.C Vdd.n787 0.0374643
R2474 SARlogic_0.dffrs_2.nand3_0.C Vdd.n825 0.0374643
R2475 SARlogic_0.dffrs_3.nand3_0.C Vdd.n863 0.0374643
R2476 SARlogic_0.dffrs_4.nand3_0.C Vdd.n902 0.0374643
R2477 SARlogic_0.dffrs_5.nand3_0.C Vdd.n940 0.0374643
R2478 SARlogic_0.dffrs_0.nand3_0.C Vdd.n712 0.0374643
R2479 Vdd.n1018 Vdd.n1012 0.0373206
R2480 Vdd.n603 Vdd.n349 0.0359182
R2481 Vdd.n673 Vdd.n672 0.0359182
R2482 Vdd.n1093 Vdd.n1087 0.0359182
R2483 Vdd.n743 Vdd.n737 0.0339767
R2484 Vdd.n49 adc_PISO_0.dffrs_5.setb 0.032
R2485 Vdd.n135 adc_PISO_0.dffrs_4.setb 0.032
R2486 Vdd.n516 adc_PISO_0.dffrs_2.setb 0.032
R2487 Vdd.n788 SARlogic_0.dffrs_1.setb 0.032
R2488 Vdd.n826 SARlogic_0.dffrs_2.setb 0.032
R2489 Vdd.n864 SARlogic_0.dffrs_3.setb 0.032
R2490 Vdd.n903 SARlogic_0.dffrs_4.setb 0.032
R2491 Vdd.n941 SARlogic_0.dffrs_5.setb 0.032
R2492 Vdd.n713 SARlogic_0.dffrs_0.setb 0.032
R2493 Vdd.n567 adc_PISO_0.dffrs_1.setb 0.032
R2494 Vdd.n636 adc_PISO_0.dffrs_0.setb 0.032
R2495 adc_PISO_0.dffrs_3.setb Vdd.n1114 0.032
R2496 Vdd.n750 Vdd.n725 0.0316083
R2497 Vdd.n188 Vdd.n186 0.0313054
R2498 Vdd.n188 Vdd.n187 0.0313054
R2499 Vdd.n115 Vdd.n113 0.0313054
R2500 Vdd.n115 Vdd.n114 0.0313054
R2501 Vdd.n129 Vdd.n30 0.0313054
R2502 Vdd.n129 Vdd.n31 0.0313054
R2503 Vdd.n202 Vdd.n14 0.0313054
R2504 Vdd.n202 Vdd.n15 0.0313054
R2505 Vdd.n253 Vdd.n251 0.0313054
R2506 Vdd.n253 Vdd.n252 0.0313054
R2507 Vdd.n616 Vdd.n614 0.0313054
R2508 Vdd.n616 Vdd.n615 0.0313054
R2509 Vdd.n547 Vdd.n545 0.0313054
R2510 Vdd.n547 Vdd.n546 0.0313054
R2511 Vdd.n561 Vdd.n497 0.0313054
R2512 Vdd.n561 Vdd.n498 0.0313054
R2513 Vdd.n630 Vdd.n481 0.0313054
R2514 Vdd.n630 Vdd.n482 0.0313054
R2515 Vdd.n475 Vdd.n473 0.0313054
R2516 Vdd.n475 Vdd.n474 0.0313054
R2517 Vdd.n461 Vdd.n459 0.0313054
R2518 Vdd.n461 Vdd.n460 0.0313054
R2519 Vdd.n267 Vdd.n265 0.0313054
R2520 Vdd.n267 Vdd.n266 0.0313054
R2521 Vdd.n118 Vdd.n105 0.0295407
R2522 Vdd.n191 Vdd.n178 0.0295407
R2523 Vdd.n550 Vdd.n537 0.0295407
R2524 Vdd.n619 Vdd.n606 0.0295407
R2525 Vdd.n479 Vdd.n478 0.0295407
R2526 Vdd.n256 Vdd.n243 0.0295407
R2527 Vdd.n103 Vdd.n91 0.0288636
R2528 Vdd.n176 Vdd.n164 0.0288636
R2529 Vdd.n666 Vdd.n665 0.0288636
R2530 Vdd.n1100 Vdd.n1094 0.0288636
R2531 Vdd.n597 Vdd.n596 0.0288455
R2532 Vdd.n1006 Vdd.n995 0.0286958
R2533 Vdd.n985 Vdd.n273 0.0279312
R2534 Vdd.n1020 Vdd.n215 0.0273926
R2535 Vdd.n79 Vdd.n68 0.0237
R2536 Vdd.n152 Vdd.n141 0.0237
R2537 Vdd.n584 Vdd.n573 0.0237
R2538 Vdd.n653 Vdd.n642 0.0237
R2539 Vdd.n1113 Vdd.n1112 0.0237
R2540 Vdd.n1044 Vdd.n1036 0.0197857
R2541 Vdd.n57 Vdd.n53 0.0197857
R2542 Vdd.n725 Vdd.n714 0.0192652
R2543 Vdd.n68 Vdd.n67 0.0173909
R2544 Vdd.n119 Vdd.n118 0.0161977
R2545 Vdd.n192 Vdd.n191 0.0161977
R2546 Vdd.n551 Vdd.n550 0.0161977
R2547 Vdd.n620 Vdd.n619 0.0161977
R2548 Vdd.n478 Vdd.n465 0.0161977
R2549 Vdd.n257 Vdd.n256 0.0161977
R2550 Vdd.n105 Vdd.n104 0.0129273
R2551 Vdd.n178 Vdd.n177 0.0129273
R2552 Vdd.n537 Vdd.n536 0.0129273
R2553 Vdd.n606 Vdd.n605 0.0129273
R2554 Vdd.n480 Vdd.n479 0.0129273
R2555 Vdd.n243 Vdd.n13 0.0129273
R2556 Vdd.n453 adc_PISO_0.avdd 0.0128676
R2557 Vdd.n103 Vdd.n102 0.0122273
R2558 Vdd.n176 Vdd.n175 0.0122273
R2559 Vdd.n604 Vdd.n603 0.0122273
R2560 Vdd.n672 Vdd.n666 0.0122273
R2561 Vdd.n1094 Vdd.n1093 0.0122273
R2562 Vdd.n995 Vdd.n994 0.0113078
R2563 Vdd.n1053 Vdd.n1021 0.0068
R2564 Vdd.n1020 Vdd.n1019 0.00613636
R2565 Vdd.n942 Vdd.n936 0.00505026
R2566 Vdd.n904 Vdd.n898 0.00505026
R2567 Vdd.n865 Vdd.n859 0.00505026
R2568 Vdd.n827 Vdd.n821 0.00505026
R2569 Vdd.n1019 Vdd.n1018 0.00441736
R2570 Vdd.n963 Vdd.n942 0.00430496
R2571 Vdd.n925 Vdd.n904 0.00430496
R2572 Vdd.n886 Vdd.n865 0.00430496
R2573 Vdd.n848 Vdd.n827 0.00430496
R2574 Vdd.n810 Vdd.n789 0.00430496
R2575 Vdd.n1039 comparator_no_offsetcal_0.x4.VDD 0.00371429
R2576 SARlogic_0.dffrs_5.vdd Vdd.n963 0.00349428
R2577 SARlogic_0.dffrs_4.vdd Vdd.n925 0.00349428
R2578 SARlogic_0.dffrs_3.vdd Vdd.n886 0.00349428
R2579 SARlogic_0.dffrs_2.vdd Vdd.n848 0.00349428
R2580 SARlogic_0.dffrs_1.vdd Vdd.n810 0.00349428
R2581 SARlogic_0.dffrs_0.vdd Vdd.n771 0.00349428
R2582 Vdd.n783 Vdd.n782 0.00291569
R2583 Vdd.n750 Vdd.n749 0.00285324
R2584 Vdd.n535 Vdd.n273 0.00265596
R2585 Vdd.n789 Vdd.n783 0.00263457
R2586 Vdd.n974 SARlogic_0.dffrs_5.vdd 0.00236325
R2587 Vdd.n936 SARlogic_0.dffrs_4.vdd 0.00236325
R2588 Vdd.n859 SARlogic_0.dffrs_2.vdd 0.00236325
R2589 Vdd.n821 SARlogic_0.dffrs_1.vdd 0.00236325
R2590 Vdd.n782 SARlogic_0.dffrs_0.vdd 0.00236325
R2591 Vdd.n271 Vdd.n270 0.00228481
R2592 Vdd.n61 osu_sc_buf_4_flat_0.VDD 0.00168943
R2593 Vdd.n898 Vdd.n887 0.0014349
R2594 Vdd.n887 SARlogic_0.dffrs_3.vdd 0.00142836
R2595 Vdd.n61 Vdd.n60 0.00129295
R2596 Vdd.n987 Vdd.n974 0.0008465
R2597 Vdd.n91 Vdd.n85 0.000518182
R2598 Vdd.n164 Vdd.n158 0.000518182
R2599 Vdd.n596 Vdd.n590 0.000518182
R2600 Vdd.n604 Vdd.n597 0.000518182
R2601 Vdd.n665 Vdd.n659 0.000518182
R2602 Vdd.n1106 Vdd.n1100 0.000518182
R2603 Vdd.n1012 Vdd.n1006 0.000517689
R2604 Vdd.n749 Vdd.n743 0.000515182
R2605 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t6 41.0041
R2606 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t5 40.6313
R2607 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t4 27.3166
R2608 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t7 26.9438
R2609 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d 17.5382
R2610 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d.n2 14.0582
R2611 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.t1 10.0473
R2612 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.t0 6.51042
R2613 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.n4 6.04952
R2614 SARlogic_0.dffrs_4.nand3_8.A SARlogic_0.dffrs_4.d.n0 5.7755
R2615 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_4.d.n1 5.13907
R2616 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n6 4.72925
R2617 SARlogic_0.dffrs_4.d SARlogic_0.dffrs_4.nand3_8.A 0.784786
R2618 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.n5 0.732092
R2619 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t2 0.7285
R2620 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t3 0.7285
R2621 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n3 0.166901
R2622 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_3.nand3_7.C 0.0455
R2623 Vss.n1117 Vss.n1116 9.36555e+06
R2624 Vss.n1117 Vss.n1052 2.41475e+06
R2625 Vss.n1116 Vss.n1078 2.41475e+06
R2626 Vss.n1468 Vss.n1467 1.11127e+06
R2627 Vss.n1466 Vss.n1465 1.11127e+06
R2628 Vss.n1472 Vss.n1471 653018
R2629 Vss.n1474 Vss.n1473 532071
R2630 Vss.n1470 Vss.n1469 511643
R2631 Vss.n1119 Vss.n232 267429
R2632 Vss.n105 Vss.n56 149958
R2633 Vss.n1120 Vss.n1119 134395
R2634 Vss.n1473 Vss.n1472 106786
R2635 Vss.n1471 Vss.n1470 106786
R2636 Vss.n247 Vss.n68 106554
R2637 Vss.n1475 Vss.n1474 101679
R2638 Vss.n1074 Vss.n1057 100518
R2639 Vss.n1477 Vss.n1476 100054
R2640 Vss.n1057 Vss.n1056 67692.9
R2641 Vss.n1056 Vss.n1053 67367.9
R2642 Vss.n1053 Vss.n232 56828.6
R2643 Vss.n1162 Vss.n433 50714
R2644 Vss.n1738 Vss.n115 50260.2
R2645 Vss.n1121 Vss.n1120 49525.3
R2646 Vss.n1862 Vss.n51 47256
R2647 Vss.n1477 Vss.n232 46428.6
R2648 Vss.n1476 Vss.n1475 45035.7
R2649 Vss.n459 Vss.n234 42464
R2650 Vss.n1829 Vss.n1828 41697.6
R2651 Vss.n1077 Vss.n1057 36083.3
R2652 Vss.n469 Vss.n233 32884
R2653 Vss.n1909 Vss.n11 31458.4
R2654 Vss.n1908 Vss.n1907 27213.5
R2655 Vss.n1828 Vss.n1827 26779.4
R2656 Vss.n1117 Vss.n1057 24300
R2657 Vss.n999 Vss.n998 24208.9
R2658 Vss.n1118 Vss.n1117 24183.3
R2659 Vss.n897 Vss.n896 22665.9
R2660 Vss.n669 Vss.n668 22665.9
R2661 Vss.n1056 Vss.n1055 21560.4
R2662 Vss.n1119 Vss.n1118 20400
R2663 Vss.t96 Vss.n106 18167.5
R2664 Vss.n810 Vss.n440 17546.4
R2665 Vss.n470 Vss.n469 17319
R2666 Vss.n998 Vss.n528 16547
R2667 Vss.n698 Vss.n11 16547
R2668 Vss.n1466 Vss.n245 16020.5
R2669 Vss.n1466 Vss.n191 16020.5
R2670 Vss.n669 Vss.n611 15733.7
R2671 Vss.n898 Vss.n897 15733.7
R2672 Vss.n1026 Vss.n529 15356.8
R2673 Vss.n469 Vss.n459 14805.6
R2674 Vss.n809 Vss.n808 13656.9
R2675 Vss.n1055 Vss.n154 13264.1
R2676 Vss.n530 Vss.n528 12982.5
R2677 Vss.n847 Vss.n782 11672.3
R2678 Vss.n1006 Vss.n514 11670.6
R2679 Vss.n1897 Vss.n1896 11568.1
R2680 Vss.n1484 Vss.n1481 11510.4
R2681 Vss.n1118 Vss.n1053 11510.4
R2682 Vss.n1752 Vss.n1749 11510.4
R2683 Vss.n1747 Vss.n1746 11510.4
R2684 Vss.n1006 Vss.n545 11510.4
R2685 Vss.n782 Vss.n595 11510.4
R2686 Vss.n1896 Vss.n16 11510.4
R2687 Vss.n1161 Vss.n440 11510.4
R2688 Vss.n1104 Vss.n1103 11412
R2689 Vss.n1073 Vss.n120 11108.6
R2690 Vss.n1023 Vss.n533 10562.5
R2691 Vss.n1828 Vss.n51 10357.6
R2692 Vss.n1862 Vss.t448 10202.1
R2693 Vss.n809 Vss.n531 10162.3
R2694 Vss.n1056 Vss.t35 9917.42
R2695 Vss.t337 Vss.n45 9747.75
R2696 Vss.n1470 Vss.n239 9694.18
R2697 Vss.n245 Vss.n241 9694.18
R2698 Vss.n1470 Vss.n241 9687.98
R2699 Vss.n1463 Vss.n191 9687.98
R2700 Vss.n1878 Vss.n1877 9213.04
R2701 Vss.n849 Vss.n848 9213.04
R2702 Vss.n1080 Vss.n119 7482.1
R2703 Vss.n685 Vss.n669 7082.44
R2704 Vss.n897 Vss.n574 7082.44
R2705 Vss.n501 Vss.n467 6961.73
R2706 Vss.n807 Vss.n527 6961.73
R2707 Vss.n842 Vss.n841 6961.73
R2708 Vss.n641 Vss.n640 6961.73
R2709 Vss.n37 Vss.n15 6921.73
R2710 Vss.n850 Vss.n847 6921.73
R2711 Vss.n247 Vss.n67 6841.13
R2712 Vss.n809 Vss.n529 6839.98
R2713 Vss.n1476 Vss.n233 6737.81
R2714 Vss.n1476 Vss.n234 6737.81
R2715 Vss.n1051 Vss.n1050 6663.38
R2716 Vss.n843 Vss.n784 6650
R2717 Vss.n643 Vss.n12 6650
R2718 Vss.n808 Vss.n515 6650
R2719 Vss.n1744 Vss.n1738 6375
R2720 Vss.n1863 Vss.n1862 6317.73
R2721 Vss.n531 Vss.n434 6190.48
R2722 Vss.n954 Vss.n514 6190.48
R2723 Vss.n1500 Vss.n155 6157.34
R2724 Vss.n1026 Vss.n1025 5894.95
R2725 Vss.n1048 Vss.n514 5875.76
R2726 Vss.n847 Vss.n592 5874.11
R2727 Vss.n1778 Vss.n1777 5751.62
R2728 Vss.n535 Vss.n360 5557.62
R2729 Vss.n962 Vss.n280 5557.62
R2730 Vss.n1397 Vss.n1396 5557.62
R2731 Vss.n1101 Vss.n1100 5557.62
R2732 Vss.n1707 Vss.n99 5557.62
R2733 Vss.n1571 Vss.n166 5557.62
R2734 Vss.n1570 Vss.n168 5557.62
R2735 Vss.n344 Vss.n310 5557.62
R2736 Vss.n1338 Vss.n1337 5557.62
R2737 Vss.n1719 Vss.n1718 5557.62
R2738 Vss.n1616 Vss.n1615 5557.62
R2739 Vss.n1214 Vss.n361 5557.62
R2740 Vss.n1184 Vss.n424 5557.62
R2741 Vss.n728 Vss.n727 5557.62
R2742 Vss.n841 Vss.n576 5551.58
R2743 Vss.n401 Vss.n361 5551.58
R2744 Vss.n1718 Vss.n1617 5551.58
R2745 Vss.n1399 Vss.n1397 5551.58
R2746 Vss.n1337 Vss.n1336 5551.58
R2747 Vss.n1396 Vss.n280 5551.58
R2748 Vss.n1707 Vss.n1706 5551.58
R2749 Vss.n503 Vss.n501 5551.58
R2750 Vss.n1033 Vss.n527 5551.58
R2751 Vss.n168 Vss.n83 5551.58
R2752 Vss.n1571 Vss.n1570 5551.58
R2753 Vss.n1338 Vss.n310 5551.58
R2754 Vss.n1719 Vss.n1616 5551.58
R2755 Vss.n1214 Vss.n360 5551.58
R2756 Vss.n1185 Vss.n1184 5551.58
R2757 Vss.n640 Vss.n614 5551.58
R2758 Vss.n729 Vss.n728 5551.58
R2759 Vss.n1910 Vss.n10 5159.25
R2760 Vss.n1087 Vss.n1052 5042.06
R2761 Vss.n1777 Vss.n1776 4925
R2762 Vss.n1831 Vss.n1830 4797.83
R2763 Vss.n1777 Vss.n106 4745.41
R2764 Vss.n1023 Vss.n1022 4485.19
R2765 Vss.n931 Vss.n362 4456.62
R2766 Vss.n1593 Vss.n1592 4448.54
R2767 Vss.n997 Vss.n533 4316.58
R2768 Vss.n726 Vss.n706 4273.71
R2769 Vss.n1025 Vss.n531 4229.5
R2770 Vss.n1078 Vss.n1077 4015.17
R2771 Vss.n1830 Vss.n45 3983.8
R2772 Vss.n533 Vss.n530 3889.63
R2773 Vss.n1025 Vss.n1024 3784.25
R2774 Vss.n684 Vss.n683 3765.76
R2775 Vss.n878 Vss.n877 3765.76
R2776 Vss.n727 Vss.n726 3568.02
R2777 Vss.n1854 Vss.t433 3463.67
R2778 Vss.n1049 Vss.n468 3419.7
R2779 Vss.n845 Vss.n844 3419.7
R2780 Vss.n1907 Vss.n13 3419.7
R2781 Vss.n1788 Vss.n98 3217.05
R2782 Vss.n1679 Vss.n1678 3214.99
R2783 Vss.n1745 Vss.n1744 3178.74
R2784 Vss.n1345 Vss.n308 3157.03
R2785 Vss.n1282 Vss.n325 3157.03
R2786 Vss.n949 Vss.n327 3157.03
R2787 Vss.n1531 Vss.n194 3157.03
R2788 Vss.n1510 Vss.n196 3157.03
R2789 Vss.n1248 Vss.n1247 3157.03
R2790 Vss.n976 Vss.n975 3157.03
R2791 Vss.n1438 Vss.n254 3157.03
R2792 Vss.n1802 Vss.n86 3157.03
R2793 Vss.n932 Vss.n534 3157.03
R2794 Vss.n1301 Vss.n267 3155.01
R2795 Vss.n379 Vss.n271 3155.01
R2796 Vss.n1282 Vss.n1281 3155.01
R2797 Vss.n248 Vss.n75 3155.01
R2798 Vss.n1531 Vss.n1530 3155.01
R2799 Vss.n1246 Vss.n254 3155.01
R2800 Vss.n1345 Vss.n309 3155.01
R2801 Vss.n1437 Vss.n1436 3155.01
R2802 Vss.n1804 Vss.n1803 3155.01
R2803 Vss.n157 Vss.n86 3148.94
R2804 Vss.n1596 Vss.n1595 3122.83
R2805 Vss.n1745 Vss.n120 3078.66
R2806 Vss.n1906 Vss.n14 3035.71
R2807 Vss.n1050 Vss.n467 2959.12
R2808 Vss.n808 Vss.n807 2959.12
R2809 Vss.n843 Vss.n842 2959.12
R2810 Vss.n641 Vss.n12 2959.12
R2811 Vss.t61 Vss.n1477 2954.55
R2812 Vss.n757 Vss.n756 2945.66
R2813 Vss.n1828 Vss.n45 2850.36
R2814 Vss.n1829 Vss.n67 2846.85
R2815 Vss.n1464 Vss.n247 2814.38
R2816 Vss.n1021 Vss.n536 2720.84
R2817 Vss.t337 Vss.n1867 2698.96
R2818 Vss.n1867 Vss.t433 2698.96
R2819 Vss.n1050 Vss.n1049 2677.48
R2820 Vss.n513 Vss.n468 2677.48
R2821 Vss.n844 Vss.n843 2677.48
R2822 Vss.n846 Vss.n845 2677.48
R2823 Vss.n1907 Vss.n12 2677.48
R2824 Vss.n612 Vss.n13 2677.48
R2825 Vss.n1771 Vss.n1770 2575.98
R2826 Vss.n1499 Vss.n1498 2567.94
R2827 Vss.n1101 Vss.n1052 2564.33
R2828 Vss.n1080 Vss.n1078 2536.1
R2829 Vss.n1744 Vss.t130 2437.5
R2830 Vss.n1077 Vss.n1076 2394.11
R2831 Vss.n1595 Vss.n154 2306.19
R2832 Vss.n1123 Vss.n1122 2267.8
R2833 Vss.n1047 Vss.n516 2257.8
R2834 Vss.n656 Vss.n655 2257.8
R2835 Vss.n811 Vss.n573 2257.8
R2836 Vss.n1595 Vss.n155 2253.62
R2837 Vss.n1074 Vss.n1073 2121.97
R2838 Vss.n1061 Vss.n1060 2096.57
R2839 Vss.n1746 Vss.n106 2047.72
R2840 Vss.n513 Vss.n512 2028.48
R2841 Vss.n613 Vss.n612 2027.23
R2842 Vss.n846 Vss.n575 2027.23
R2843 Vss.n1816 Vss.n1815 1972.34
R2844 Vss.n1818 Vss.n1816 1972.34
R2845 Vss.n1687 Vss.n84 1972.34
R2846 Vss.n1692 Vss.n1691 1953.93
R2847 Vss.n1693 Vss.n1692 1953.93
R2848 Vss.t89 Vss.n1747 1950
R2849 Vss.n1048 Vss.n1047 1943.45
R2850 Vss.n655 Vss.n592 1943.45
R2851 Vss.n811 Vss.n810 1943.45
R2852 Vss.n514 Vss.n513 1891.48
R2853 Vss.n612 Vss.n15 1890.32
R2854 Vss.n847 Vss.n846 1890.32
R2855 Vss.n962 Vss.n961 1883.67
R2856 Vss.n1509 Vss.n166 1883.67
R2857 Vss.n1471 Vss.n237 1883.67
R2858 Vss.n977 Vss.n344 1883.67
R2859 Vss.n1022 Vss.n535 1883.67
R2860 Vss.n1787 Vss.n99 1861.56
R2861 Vss.n1906 Vss.n1897 1849.33
R2862 Vss.n1075 Vss.n1074 1841.93
R2863 Vss.n1021 Vss.n1020 1775.77
R2864 Vss.n810 Vss.n809 1732.36
R2865 Vss.n84 Vss.n51 1726.87
R2866 Vss.t89 Vss.t96 1657.5
R2867 Vss.n1474 Vss.n234 1645.06
R2868 Vss.n1055 Vss.n155 1579.08
R2869 Vss.n1055 Vss.n1054 1476.63
R2870 Vss.n1509 Vss.n155 1450.15
R2871 Vss.n1122 Vss.n1121 1347.31
R2872 Vss.n920 Vss.n534 1336.79
R2873 Vss.n949 Vss.n948 1336.79
R2874 Vss.n976 Vss.n971 1336.79
R2875 Vss.n1249 Vss.n1248 1336.79
R2876 Vss.n1511 Vss.n1510 1336.79
R2877 Vss.n403 Vss.n271 1336.25
R2878 Vss.n1400 Vss.n267 1336.25
R2879 Vss.n1805 Vss.n1804 1336.25
R2880 Vss.n1426 Vss.n75 1336.25
R2881 Vss.n1789 Vss.n1788 1314.68
R2882 Vss.n1679 Vss.n1676 1314.15
R2883 Vss.n1854 Vss.n1853 1303.34
R2884 Vss.n1853 Vss.n1852 1223
R2885 Vss.n1073 Vss.n154 1218.08
R2886 Vss.n726 Vss.n725 1212.42
R2887 Vss.n1104 Vss.n119 1210.86
R2888 Vss.n978 Vss.n977 1201.62
R2889 Vss.n1021 Vss.n537 1200.6
R2890 Vss.n961 Vss.n949 1095.12
R2891 Vss.n1788 Vss.n1787 1095.12
R2892 Vss.n1510 Vss.n1509 1095.12
R2893 Vss.n977 Vss.n976 1095.12
R2894 Vss.n1022 Vss.n534 1095.12
R2895 Vss.n1416 Vss.n267 1094.63
R2896 Vss.n1410 Vss.n271 1094.63
R2897 Vss.n1692 Vss.n1679 1094.63
R2898 Vss.n1816 Vss.n75 1094.63
R2899 Vss.n1804 Vss.n84 1094.63
R2900 Vss.n1746 Vss.n1745 1066.44
R2901 Vss.n1509 Vss.n1508 1055.77
R2902 Vss.n1025 Vss.n530 996.898
R2903 Vss.n1595 Vss.n1593 933.769
R2904 Vss.n1694 Vss.n56 928.572
R2905 Vss.n1201 Vss.n362 927.706
R2906 Vss.n1121 Vss.n1051 920.491
R2907 Vss.n727 Vss.n10 897.806
R2908 Vss.n1465 Vss.n1464 885.807
R2909 Vss.n999 Vss.n989 873.918
R2910 Vss.n742 Vss.n14 873.918
R2911 Vss.n1771 Vss.t553 857.144
R2912 Vss.n1775 Vss.t553 857.144
R2913 Vss.t86 Vss.n602 849.126
R2914 Vss.n866 Vss.t73 849.126
R2915 Vss.t130 Vss.n1739 847.827
R2916 Vss.n1749 Vss.t89 847.827
R2917 Vss.n1770 Vss.t96 847.827
R2918 Vss.t61 Vss.n231 847.827
R2919 Vss.n1498 Vss.t35 847.827
R2920 Vss.t558 Vss.n1499 847.827
R2921 Vss.n1500 Vss.t558 847.827
R2922 Vss.t666 Vss.n37 847.827
R2923 Vss.n1878 Vss.t666 847.827
R2924 Vss.n683 Vss.t257 847.827
R2925 Vss.n680 Vss.t257 847.827
R2926 Vss.n679 Vss.t181 847.827
R2927 Vss.n676 Vss.t181 847.827
R2928 Vss.n675 Vss.t86 847.827
R2929 Vss.n850 Vss.t560 847.827
R2930 Vss.t560 Vss.n849 847.827
R2931 Vss.n877 Vss.t437 847.827
R2932 Vss.n874 Vss.t437 847.827
R2933 Vss.n873 Vss.t11 847.827
R2934 Vss.t11 Vss.n872 847.827
R2935 Vss.t73 Vss.n583 847.827
R2936 Vss.n1100 Vss.n1099 832.75
R2937 Vss.n1100 Vss.n1079 832.75
R2938 Vss.n364 Vss.n361 832.22
R2939 Vss.n1337 Vss.n311 832.22
R2940 Vss.n1397 Vss.n278 832.22
R2941 Vss.n1272 Vss.n280 832.22
R2942 Vss.n1708 Vss.n1707 832.22
R2943 Vss.n501 Vss.n471 832.22
R2944 Vss.n1453 Vss.n168 832.22
R2945 Vss.n1571 Vss.n167 832.22
R2946 Vss.n973 Vss.n310 832.22
R2947 Vss.n1718 Vss.n1618 832.22
R2948 Vss.n1616 Vss.n143 832.22
R2949 Vss.n934 Vss.n360 832.22
R2950 Vss.n796 Vss.n527 832.22
R2951 Vss.n1184 Vss.n425 832.22
R2952 Vss.n841 Vss.n786 832.22
R2953 Vss.n640 Vss.n638 832.22
R2954 Vss.n728 Vss.n696 832.22
R2955 Vss.n378 Vss.n361 832.101
R2956 Vss.n1337 Vss.n312 832.101
R2957 Vss.n1397 Vss.n279 832.101
R2958 Vss.n1260 Vss.n280 832.101
R2959 Vss.n1707 Vss.n1626 832.101
R2960 Vss.n501 Vss.n500 832.101
R2961 Vss.n178 Vss.n168 832.101
R2962 Vss.n1573 Vss.n1571 832.101
R2963 Vss.n346 Vss.n310 832.101
R2964 Vss.n1718 Vss.n1717 832.101
R2965 Vss.n1616 Vss.n144 832.101
R2966 Vss.n360 Vss.n359 832.101
R2967 Vss.n527 Vss.n526 832.101
R2968 Vss.n1184 Vss.n1183 832.101
R2969 Vss.n841 Vss.n840 832.101
R2970 Vss.n640 Vss.n639 832.101
R2971 Vss.n728 Vss.n697 832.101
R2972 Vss.n1022 Vss.n1021 829.364
R2973 Vss.n1463 Vss.n1462 814.398
R2974 Vss.n241 Vss.n240 814.398
R2975 Vss.n1054 Vss.t139 812.5
R2976 Vss.n1596 Vss.t422 812.5
R2977 Vss.n1877 Vss.t264 812.5
R2978 Vss.n848 Vss.t70 812.5
R2979 Vss.n1134 Vss.n1133 798.088
R2980 Vss.n689 Vss.n11 767.827
R2981 Vss.n1747 Vss.n118 755.625
R2982 Vss.n977 Vss.n557 750.922
R2983 Vss.n1123 Vss.n233 748.735
R2984 Vss.n1061 Vss.t33 732.843
R2985 Vss.n1060 Vss.t227 732.843
R2986 Vss.n1072 Vss.t671 732.843
R2987 Vss.t89 Vss.t96 720.653
R2988 Vss.n680 Vss.n679 720.653
R2989 Vss.n676 Vss.n675 720.653
R2990 Vss.n874 Vss.n873 720.653
R2991 Vss.n872 Vss.n583 720.653
R2992 Vss.n1829 Vss.n1826 702.332
R2993 Vss.n1248 Vss.n237 698.639
R2994 Vss.n503 Vss.n502 693.082
R2995 Vss.n619 Vss.n614 692.747
R2996 Vss.n884 Vss.n576 692.747
R2997 Vss.n1827 Vss.t348 676.471
R2998 Vss.n1867 Vss.t348 676.471
R2999 Vss.n1867 Vss.t286 676.471
R3000 Vss.n1863 Vss.t286 676.471
R3001 Vss.n1020 Vss.t159 670.104
R3002 Vss.t159 Vss.n1019 670.104
R3003 Vss.n1016 Vss.t451 670.104
R3004 Vss.n549 Vss.t451 670.104
R3005 Vss.n550 Vss.t632 670.104
R3006 Vss.n989 Vss.t632 670.104
R3007 Vss.n756 Vss.t609 670.104
R3008 Vss.n750 Vss.t609 670.104
R3009 Vss.n749 Vss.t215 670.104
R3010 Vss.n746 Vss.t215 670.104
R3011 Vss.n745 Vss.t645 670.104
R3012 Vss.t645 Vss.n742 670.104
R3013 Vss.n1063 Vss.n1057 667.231
R3014 Vss.n999 Vss.n516 665.564
R3015 Vss.n656 Vss.n611 665.564
R3016 Vss.n898 Vss.n573 665.564
R3017 Vss.n1468 Vss.n241 662.646
R3018 Vss.n504 Vss.n503 662.074
R3019 Vss.n1907 Vss.n1906 661.894
R3020 Vss.n667 Vss.n614 661.665
R3021 Vss.n895 Vss.n576 661.665
R3022 Vss.t139 Vss.t529 650
R3023 Vss.t529 Vss.t422 650
R3024 Vss.t503 Vss.t582 650
R3025 Vss.t471 Vss.t150 650
R3026 Vss.t251 Vss.n537 642.183
R3027 Vss.n689 Vss.t603 642.183
R3028 Vss.n740 Vss.t599 642.183
R3029 Vss.t665 Vss.n1478 624
R3030 Vss.n1479 Vss.t556 624
R3031 Vss.n1478 Vss.t61 624
R3032 Vss.n1479 Vss.t37 624
R3033 Vss.n1776 Vss.n1775 607.144
R3034 Vss.n1743 Vss.t562 590.91
R3035 Vss.t130 Vss.n1743 590.91
R3036 Vss.t579 Vss.n1000 590.909
R3037 Vss.n1004 Vss.t579 590.909
R3038 Vss.t549 Vss.n1004 590.909
R3039 Vss.n1006 Vss.t557 590.909
R3040 Vss.t613 Vss.n1006 590.909
R3041 Vss.n1007 Vss.t620 590.909
R3042 Vss.n610 Vss.t584 590.909
R3043 Vss.t584 Vss.n609 590.909
R3044 Vss.n609 Vss.t550 590.909
R3045 Vss.n782 Vss.t563 590.909
R3046 Vss.n782 Vss.t179 590.909
R3047 Vss.t444 Vss.n591 590.909
R3048 Vss.n26 Vss.t270 590.909
R3049 Vss.t270 Vss.n25 590.909
R3050 Vss.n25 Vss.t661 590.909
R3051 Vss.n1896 Vss.t548 590.909
R3052 Vss.n1896 Vss.t340 590.909
R3053 Vss.t344 Vss.n1895 590.909
R3054 Vss.t20 Vss.n899 590.909
R3055 Vss.n900 Vss.t20 590.909
R3056 Vss.n900 Vss.t555 590.909
R3057 Vss.t664 Vss.n440 590.909
R3058 Vss.t47 Vss.n440 590.909
R3059 Vss.n904 Vss.t627 590.909
R3060 Vss.t421 Vss.t515 586.274
R3061 Vss.t33 Vss.t421 586.274
R3062 Vss.t227 Vss.t186 586.274
R3063 Vss.t186 Vss.t671 586.274
R3064 Vss.n1309 Vss.t123 582.165
R3065 Vss.t512 Vss.n311 582.165
R3066 Vss.n374 Vss.t189 582.165
R3067 Vss.t491 Vss.n278 582.165
R3068 Vss.n1273 Vss.t78 582.165
R3069 Vss.t119 Vss.n1272 582.165
R3070 Vss.n1087 Vss.t0 582.165
R3071 Vss.n1099 Vss.t479 582.165
R3072 Vss.t439 Vss.n1115 582.165
R3073 Vss.n1709 Vss.t598 582.165
R3074 Vss.t573 Vss.n1708 582.165
R3075 Vss.n478 Vss.t113 582.165
R3076 Vss.t465 Vss.n471 582.165
R3077 Vss.n1454 Vss.t292 582.165
R3078 Vss.t477 Vss.n1453 582.165
R3079 Vss.n1522 Vss.t198 582.165
R3080 Vss.t161 Vss.n167 582.165
R3081 Vss.n345 Vss.t81 582.165
R3082 Vss.t288 Vss.n242 582.165
R3083 Vss.n974 Vss.t594 582.165
R3084 Vss.t399 Vss.n973 582.165
R3085 Vss.n1439 Vss.t608 582.165
R3086 Vss.t493 Vss.n246 582.165
R3087 Vss.n1801 Vss.t622 582.165
R3088 Vss.n1618 Vss.t499 582.165
R3089 Vss.n1591 Vss.t265 582.165
R3090 Vss.t586 Vss.n143 582.165
R3091 Vss.t176 Vss.n933 582.165
R3092 Vss.n934 Vss.t680 582.165
R3093 Vss.n416 Vss.t619 582.165
R3094 Vss.n364 Vss.t495 582.165
R3095 Vss.n797 Vss.t366 582.165
R3096 Vss.t467 Vss.n796 582.165
R3097 Vss.n1163 Vss.t110 582.165
R3098 Vss.t617 Vss.n425 582.165
R3099 Vss.t259 Vss.n783 582.165
R3100 Vss.n786 Vss.t497 582.165
R3101 Vss.n626 Vss.t460 582.165
R3102 Vss.n638 Vss.t504 582.165
R3103 Vss.n725 Vss.t388 582.165
R3104 Vss.t520 Vss.n696 582.165
R3105 Vss.t267 Vss.n532 581.712
R3106 Vss.n920 Vss.t615 581.712
R3107 Vss.n558 Vss.t42 581.712
R3108 Vss.n948 Vss.t190 581.712
R3109 Vss.t275 Vss.n282 581.712
R3110 Vss.n1347 Vss.t224 581.712
R3111 Vss.t66 Vss.n283 581.712
R3112 Vss.n306 Vss.t461 581.712
R3113 Vss.n357 Vss.t117 581.712
R3114 Vss.t39 Vss.n323 581.712
R3115 Vss.n404 Vss.t146 581.712
R3116 Vss.t532 Vss.n403 581.712
R3117 Vss.n358 Vss.t534 581.712
R3118 Vss.n1284 Vss.t487 581.712
R3119 Vss.t24 Vss.n378 581.712
R3120 Vss.n380 Vss.t299 581.712
R3121 Vss.n1335 Vss.t411 581.712
R3122 Vss.n1331 Vss.t297 581.712
R3123 Vss.n1401 Vss.t367 581.712
R3124 Vss.t63 Vss.n1400 581.712
R3125 Vss.n312 Vss.t26 581.712
R3126 Vss.t154 Vss.n255 581.712
R3127 Vss.t30 Vss.n279 581.712
R3128 Vss.n1302 Vss.t369 581.712
R3129 Vss.t682 Vss.n1260 581.712
R3130 Vss.n1261 Vss.t75 581.712
R3131 Vss.n963 Vss.t222 581.712
R3132 Vss.n971 Vss.t121 581.712
R3133 Vss.n1250 Vss.t650 581.712
R3134 Vss.t592 Vss.n1249 581.712
R3135 Vss.n1102 Vss.t670 581.712
R3136 Vss.n1105 Vss.t526 581.712
R3137 Vss.n137 Vss.t9 581.712
R3138 Vss.t295 Vss.n121 581.712
R3139 Vss.n1790 Vss.t377 581.712
R3140 Vss.t483 Vss.n1789 581.712
R3141 Vss.n1672 Vss.t68 581.712
R3142 Vss.n1676 Vss.t14 581.712
R3143 Vss.n1705 Vss.t72 581.712
R3144 Vss.n1628 Vss.t601 581.712
R3145 Vss.t625 Vss.n1642 581.712
R3146 Vss.n1643 Vss.t332 581.712
R3147 Vss.t5 Vss.n1626 581.712
R3148 Vss.n1655 Vss.t457 581.712
R3149 Vss.n500 Vss.t188 581.712
R3150 Vss.t380 Vss.n465 581.712
R3151 Vss.n488 Vss.t359 581.712
R3152 Vss.t517 Vss.n466 581.712
R3153 Vss.n502 Vss.t140 581.712
R3154 Vss.n1124 Vss.t361 581.712
R3155 Vss.t206 Vss.n1034 581.712
R3156 Vss.n1035 Vss.t392 581.712
R3157 Vss.n205 Vss.t233 581.712
R3158 Vss.t623 Vss.n156 581.712
R3159 Vss.n238 Vss.t49 581.712
R3160 Vss.n1511 Vss.t290 581.712
R3161 Vss.t207 Vss.n170 581.712
R3162 Vss.n1549 Vss.t234 581.712
R3163 Vss.t104 Vss.n171 581.712
R3164 Vss.n1546 Vss.t506 581.712
R3165 Vss.n1367 Vss.t249 581.712
R3166 Vss.t51 Vss.n192 581.712
R3167 Vss.n1534 Vss.t373 581.712
R3168 Vss.t524 Vss.n1533 581.712
R3169 Vss.n1806 Vss.t22 581.712
R3170 Vss.t102 Vss.n1805 581.712
R3171 Vss.n1462 Vss.t32 581.712
R3172 Vss.n249 Vss.t395 581.712
R3173 Vss.n1427 Vss.t201 581.712
R3174 Vss.t374 Vss.n1426 581.712
R3175 Vss.n178 Vss.t23 581.712
R3176 Vss.t397 Vss.n85 581.712
R3177 Vss.n1573 Vss.t56 581.712
R3178 Vss.t346 Vss.n1572 581.712
R3179 Vss.n240 Vss.t236 581.712
R3180 Vss.n1529 Vss.t79 581.712
R3181 Vss.n346 Vss.t431 581.712
R3182 Vss.n1245 Vss.t220 581.712
R3183 Vss.n1353 Vss.t112 581.712
R3184 Vss.t648 Vss.n291 581.712
R3185 Vss.n292 Vss.t302 581.712
R3186 Vss.n1383 Vss.t485 581.712
R3187 Vss.n1717 Vss.t29 581.712
R3188 Vss.n1677 Vss.t284 581.712
R3189 Vss.n144 Vss.t634 581.712
R3190 Vss.t357 Vss.n123 581.712
R3191 Vss.n1732 Vss.t294 581.712
R3192 Vss.t588 Vss.n124 581.712
R3193 Vss.n359 Vss.t426 581.712
R3194 Vss.n1280 Vss.t173 581.712
R3195 Vss.n1189 Vss.t7 581.712
R3196 Vss.t268 Vss.n1188 581.712
R3197 Vss.n806 Vss.t391 581.712
R3198 Vss.n787 Vss.t522 581.712
R3199 Vss.n526 Vss.t626 581.712
R3200 Vss.n1046 Vss.t371 581.712
R3201 Vss.n1183 Vss.t99 581.712
R3202 Vss.n930 Vss.t630 581.712
R3203 Vss.t171 Vss.n785 581.712
R3204 Vss.n830 Vss.t489 581.712
R3205 Vss.n840 Vss.t204 581.712
R3206 Vss.n812 Vss.t152 581.712
R3207 Vss.t406 Vss.n642 581.712
R3208 Vss.n644 Vss.t501 581.712
R3209 Vss.n639 Vss.t202 581.712
R3210 Vss.n654 Vss.t590 581.712
R3211 Vss.n9 Vss.t163 581.712
R3212 Vss.n1911 Vss.t509 581.712
R3213 Vss.n730 Vss.t644 581.712
R3214 Vss.t165 Vss.n7 581.712
R3215 Vss.n697 Vss.t675 581.712
R3216 Vss.t606 Vss.n8 581.712
R3217 Vss.t384 Vss.n619 581.712
R3218 Vss.n657 Vss.t404 581.712
R3219 Vss.t604 Vss.n884 581.712
R3220 Vss.n885 Vss.t169 581.712
R3221 Vss.n1019 Vss.n1016 569.588
R3222 Vss.n550 Vss.n549 569.588
R3223 Vss.n750 Vss.n749 569.588
R3224 Vss.n746 Vss.n745 569.588
R3225 Vss.t582 Vss.n685 561.686
R3226 Vss.t150 Vss.n574 561.686
R3227 Vss.n558 Vss.n535 548.236
R3228 Vss.n963 Vss.n962 548.236
R3229 Vss.n1250 Vss.n344 548.236
R3230 Vss.n1642 Vss.n99 548.236
R3231 Vss.n205 Vss.n166 548.236
R3232 Vss.n1336 Vss.n1335 548.058
R3233 Vss.n1401 Vss.n1399 548.058
R3234 Vss.n1672 Vss.n1617 548.058
R3235 Vss.n1706 Vss.n1705 548.058
R3236 Vss.n1034 Vss.n1033 548.058
R3237 Vss.n1806 Vss.n83 548.058
R3238 Vss.n730 Vss.n729 548.058
R3239 Vss.t556 Vss.t665 530.4
R3240 Vss.t37 Vss.t35 530.4
R3241 Vss.n1745 Vss.n119 522.33
R3242 Vss.t199 Vss.t464 513.746
R3243 Vss.t464 Vss.t251 513.746
R3244 Vss.t603 Vss.t511 513.746
R3245 Vss.t511 Vss.t599 513.746
R3246 Vss.t562 Vss.t668 502.274
R3247 Vss.t557 Vss.t549 502.274
R3248 Vss.t620 Vss.t613 502.274
R3249 Vss.t550 Vss.t563 502.274
R3250 Vss.t179 Vss.t444 502.274
R3251 Vss.t661 Vss.t548 502.274
R3252 Vss.t340 Vss.t344 502.274
R3253 Vss.t555 Vss.t664 502.274
R3254 Vss.t627 Vss.t47 502.274
R3255 Vss.n1336 Vss.n1329 484.702
R3256 Vss.n1399 Vss.n1398 484.702
R3257 Vss.n1706 Vss.n1627 484.702
R3258 Vss.n1033 Vss.n1032 484.702
R3259 Vss.n83 Vss.n82 484.702
R3260 Vss.n1665 Vss.n1617 484.702
R3261 Vss.n729 Vss.n695 484.702
R3262 Vss.t123 Vss.t301 465.733
R3263 Vss.t301 Vss.t512 465.733
R3264 Vss.t189 Vss.t65 465.733
R3265 Vss.t65 Vss.t491 465.733
R3266 Vss.t78 Vss.t223 465.733
R3267 Vss.t223 Vss.t119 465.733
R3268 Vss.t0 Vss.t673 465.733
R3269 Vss.t673 Vss.t479 465.733
R3270 Vss.t674 Vss.t470 465.733
R3271 Vss.t470 Vss.t439 465.733
R3272 Vss.t598 Vss.t686 465.733
R3273 Vss.t686 Vss.t573 465.733
R3274 Vss.t113 Vss.t360 465.733
R3275 Vss.t360 Vss.t465 465.733
R3276 Vss.t292 Vss.t105 465.733
R3277 Vss.t105 Vss.t477 465.733
R3278 Vss.t198 Vss.t232 465.733
R3279 Vss.t232 Vss.t161 465.733
R3280 Vss.t81 Vss.t50 465.733
R3281 Vss.t50 Vss.t288 465.733
R3282 Vss.t594 Vss.t647 465.733
R3283 Vss.t647 Vss.t399 465.733
R3284 Vss.t608 Vss.t376 465.733
R3285 Vss.t376 Vss.t493 465.733
R3286 Vss.t16 Vss.t622 465.733
R3287 Vss.t499 Vss.t16 465.733
R3288 Vss.t265 Vss.t293 465.733
R3289 Vss.t293 Vss.t586 465.733
R3290 Vss.t41 Vss.t176 465.733
R3291 Vss.t680 Vss.t41 465.733
R3292 Vss.t535 Vss.t619 465.733
R3293 Vss.t495 Vss.t535 465.733
R3294 Vss.t366 Vss.t394 465.733
R3295 Vss.t394 Vss.t467 465.733
R3296 Vss.t110 Vss.t266 465.733
R3297 Vss.t266 Vss.t617 465.733
R3298 Vss.t172 Vss.t259 465.733
R3299 Vss.t497 Vss.t172 465.733
R3300 Vss.t460 Vss.t407 465.733
R3301 Vss.t407 Vss.t504 465.733
R3302 Vss.t388 Vss.t164 465.733
R3303 Vss.t164 Vss.t520 465.733
R3304 Vss.t8 Vss.t267 465.37
R3305 Vss.t615 Vss.t8 465.37
R3306 Vss.t42 Vss.t118 465.37
R3307 Vss.t118 Vss.t190 465.37
R3308 Vss.t683 Vss.t275 465.37
R3309 Vss.t224 Vss.t683 465.37
R3310 Vss.t368 Vss.t66 465.37
R3311 Vss.t461 Vss.t368 465.37
R3312 Vss.t117 Vss.t53 465.37
R3313 Vss.t53 Vss.t39 465.37
R3314 Vss.t146 Vss.t27 465.37
R3315 Vss.t27 Vss.t532 465.37
R3316 Vss.t534 Vss.t145 465.37
R3317 Vss.t145 Vss.t487 465.37
R3318 Vss.t335 Vss.t24 465.37
R3319 Vss.t299 Vss.t335 465.37
R3320 Vss.t6 Vss.t411 465.37
R3321 Vss.t297 Vss.t6 465.37
R3322 Vss.t367 Vss.t4 465.37
R3323 Vss.t4 Vss.t63 465.37
R3324 Vss.t26 Vss.t327 465.37
R3325 Vss.t327 Vss.t154 465.37
R3326 Vss.t309 Vss.t30 465.37
R3327 Vss.t369 Vss.t309 465.37
R3328 Vss.t328 Vss.t682 465.37
R3329 Vss.t75 Vss.t328 465.37
R3330 Vss.t222 Vss.t276 465.37
R3331 Vss.t276 Vss.t121 465.37
R3332 Vss.t650 Vss.t111 465.37
R3333 Vss.t111 Vss.t592 465.37
R3334 Vss.t670 Vss.t226 465.37
R3335 Vss.t226 Vss.t526 465.37
R3336 Vss.t9 Vss.t638 465.37
R3337 Vss.t638 Vss.t295 465.37
R3338 Vss.t377 Vss.t69 465.37
R3339 Vss.t69 Vss.t483 465.37
R3340 Vss.t68 Vss.t1 465.37
R3341 Vss.t1 Vss.t14 465.37
R3342 Vss.t31 Vss.t72 465.37
R3343 Vss.t601 Vss.t31 465.37
R3344 Vss.t71 Vss.t625 465.37
R3345 Vss.t332 Vss.t71 465.37
R3346 Vss.t528 Vss.t5 465.37
R3347 Vss.t457 Vss.t528 465.37
R3348 Vss.t188 Vss.t473 465.37
R3349 Vss.t473 Vss.t380 465.37
R3350 Vss.t359 Vss.t657 465.37
R3351 Vss.t657 Vss.t517 465.37
R3352 Vss.t140 Vss.t676 465.37
R3353 Vss.t676 Vss.t361 465.37
R3354 Vss.t205 Vss.t206 465.37
R3355 Vss.t392 Vss.t205 465.37
R3356 Vss.t233 Vss.t208 465.37
R3357 Vss.t208 Vss.t623 465.37
R3358 Vss.t49 Vss.t250 465.37
R3359 Vss.t250 Vss.t290 465.37
R3360 Vss.t55 Vss.t207 465.37
R3361 Vss.t234 Vss.t55 465.37
R3362 Vss.t147 Vss.t104 465.37
R3363 Vss.t506 Vss.t147 465.37
R3364 Vss.t249 Vss.t238 465.37
R3365 Vss.t238 Vss.t51 465.37
R3366 Vss.t373 Vss.t200 465.37
R3367 Vss.t200 Vss.t524 465.37
R3368 Vss.t22 Vss.t25 465.37
R3369 Vss.t25 Vss.t102 465.37
R3370 Vss.t568 Vss.t32 465.37
R3371 Vss.t395 Vss.t568 465.37
R3372 Vss.t201 Vss.t28 465.37
R3373 Vss.t28 Vss.t374 465.37
R3374 Vss.t23 Vss.t572 465.37
R3375 Vss.t572 Vss.t397 465.37
R3376 Vss.t56 Vss.t313 465.37
R3377 Vss.t313 Vss.t346 465.37
R3378 Vss.t236 Vss.t308 465.37
R3379 Vss.t308 Vss.t79 465.37
R3380 Vss.t431 Vss.t569 465.37
R3381 Vss.t569 Vss.t220 465.37
R3382 Vss.t112 Vss.t432 465.37
R3383 Vss.t432 Vss.t648 465.37
R3384 Vss.t302 Vss.t412 465.37
R3385 Vss.t412 Vss.t485 465.37
R3386 Vss.t314 Vss.t29 465.37
R3387 Vss.t284 Vss.t314 465.37
R3388 Vss.t634 Vss.t331 465.37
R3389 Vss.t331 Vss.t357 465.37
R3390 Vss.t294 Vss.t10 465.37
R3391 Vss.t10 Vss.t588 465.37
R3392 Vss.t426 Vss.t318 465.37
R3393 Vss.t318 Vss.t173 465.37
R3394 Vss.t7 Vss.t92 465.37
R3395 Vss.t92 Vss.t268 465.37
R3396 Vss.t651 Vss.t391 465.37
R3397 Vss.t522 Vss.t651 465.37
R3398 Vss.t626 Vss.t474 465.37
R3399 Vss.t474 Vss.t371 465.37
R3400 Vss.t303 Vss.t99 465.37
R3401 Vss.t630 Vss.t303 465.37
R3402 Vss.t605 Vss.t171 465.37
R3403 Vss.t489 Vss.t605 465.37
R3404 Vss.t481 Vss.t204 465.37
R3405 Vss.t152 Vss.t481 465.37
R3406 Vss.t385 Vss.t406 465.37
R3407 Vss.t501 Vss.t385 465.37
R3408 Vss.t202 Vss.t514 465.37
R3409 Vss.t514 Vss.t590 465.37
R3410 Vss.t163 Vss.t639 465.37
R3411 Vss.t639 Vss.t509 465.37
R3412 Vss.t644 Vss.t677 465.37
R3413 Vss.t677 Vss.t165 465.37
R3414 Vss.t675 Vss.t519 465.37
R3415 Vss.t519 Vss.t606 465.37
R3416 Vss.t187 Vss.t384 465.37
R3417 Vss.t404 Vss.t187 465.37
R3418 Vss.t203 Vss.t604 465.37
R3419 Vss.t169 Vss.t203 465.37
R3420 Vss.n504 Vss.t611 462.849
R3421 Vss.t342 Vss.n667 462.562
R3422 Vss.t177 Vss.n895 462.562
R3423 Vss.n1410 Vss.n270 443.358
R3424 Vss.n1411 Vss.n1410 443.358
R3425 Vss.n1416 Vss.n1415 443.358
R3426 Vss.n1418 Vss.n1416 443.358
R3427 Vss.n1282 Vss.n326 435.214
R3428 Vss.n1531 Vss.n195 435.214
R3429 Vss.n1345 Vss.n1344 435.214
R3430 Vss.n297 Vss.n254 435.214
R3431 Vss.n142 Vss.n86 435.012
R3432 Vss.n1832 Vss.n58 414.478
R3433 Vss.n1283 Vss.n1282 404.991
R3434 Vss.n1532 Vss.n1531 404.991
R3435 Vss.n1346 Vss.n1345 404.991
R3436 Vss.n1384 Vss.n254 404.991
R3437 Vss.n1548 Vss.n86 404.803
R3438 Vss.n998 Vss.n997 402.062
R3439 Vss.t540 Vss.t538 384.214
R3440 Vss.n765 Vss.n764 383.418
R3441 Vss.n766 Vss.n765 383.418
R3442 Vss.n858 Vss.n857 383.418
R3443 Vss.n862 Vss.n858 383.418
R3444 Vss.n1908 Vss.n0 377.236
R3445 Vss.t629 Vss.t469 370.279
R3446 Vss.t611 Vss.t629 370.279
R3447 Vss.t516 Vss.t581 370.05
R3448 Vss.t581 Vss.t342 370.05
R3449 Vss.t482 Vss.t149 370.05
R3450 Vss.t149 Vss.t177 370.05
R3451 Vss.n765 Vss.t503 367.392
R3452 Vss.n858 Vss.t471 367.392
R3453 Vss.n1116 Vss.n1079 367.017
R3454 Vss.n512 Vss.n470 366.255
R3455 Vss.n1394 Vss.t193 366.243
R3456 Vss.n307 Vss.t245 366.243
R3457 Vss.n1216 Vss.t279 366.243
R3458 Vss.t183 Vss.n324 366.243
R3459 Vss.n1568 Vss.t278 366.243
R3460 Vss.n1547 Vss.t124 366.243
R3461 Vss.n244 Vss.t277 366.243
R3462 Vss.t128 Vss.n193 366.243
R3463 Vss.n1386 Vss.t77 366.243
R3464 Vss.t441 Vss.n1385 366.243
R3465 Vss.n668 Vss.n613 366.027
R3466 Vss.n896 Vss.n575 366.027
R3467 Vss.n1559 Vss.t192 365.705
R3468 Vss.t273 Vss.n122 365.705
R3469 Vss.t668 Vss.n118 361.933
R3470 Vss.t448 Vss.n52 350.313
R3471 Vss.t319 Vss.n268 338.849
R3472 Vss.n1329 Vss.t655 338.849
R3473 Vss.n1409 Vss.t311 338.849
R3474 Vss.n1398 Vss.t157 338.849
R3475 Vss.n1684 Vss.t472 338.849
R3476 Vss.t595 Vss.n1627 338.849
R3477 Vss.n1027 Vss.t476 338.849
R3478 Vss.n1814 Vss.t320 338.849
R3479 Vss.n82 Vss.t18 338.849
R3480 Vss.t321 Vss.n1664 338.849
R3481 Vss.n1665 Vss.t132 338.849
R3482 Vss.n706 Vss.t475 338.849
R3483 Vss.t640 Vss.n695 338.849
R3484 Vss.n758 Vss.n757 330.211
R3485 Vss.n1749 Vss.n118 328.534
R3486 Vss.n1048 Vss.n515 314.351
R3487 Vss.n643 Vss.n592 314.351
R3488 Vss.n810 Vss.n784 314.351
R3489 Vss.n1076 Vss.n1075 307.647
R3490 Vss.t334 Vss.t193 292.995
R3491 Vss.t245 Vss.t334 292.995
R3492 Vss.t279 Vss.t329 292.995
R3493 Vss.t329 Vss.t183 292.995
R3494 Vss.t567 Vss.t278 292.995
R3495 Vss.t124 Vss.t567 292.995
R3496 Vss.t277 Vss.t315 292.995
R3497 Vss.t315 Vss.t128 292.995
R3498 Vss.t77 Vss.t575 292.995
R3499 Vss.t575 Vss.t441 292.995
R3500 Vss.t192 Vss.t305 292.565
R3501 Vss.t305 Vss.t273 292.565
R3502 Vss.n765 Vss.t264 282.61
R3503 Vss.n858 Vss.t70 282.61
R3504 Vss.t536 Vss.n1856 282.512
R3505 Vss.n1826 Vss.t17 282.289
R3506 Vss.n1815 Vss.t658 282.289
R3507 Vss.n1818 Vss.t564 282.289
R3508 Vss.t409 Vss.n1817 282.289
R3509 Vss.n1687 Vss.t597 282.289
R3510 Vss.n1691 Vss.t43 282.289
R3511 Vss.t101 Vss.n1693 282.289
R3512 Vss.n1695 Vss.t141 282.289
R3513 Vss.t401 Vss.t319 271.079
R3514 Vss.t655 Vss.t401 271.079
R3515 Vss.t350 Vss.t311 271.079
R3516 Vss.t157 Vss.t350 271.079
R3517 Vss.t472 Vss.t13 271.079
R3518 Vss.t13 Vss.t595 271.079
R3519 Vss.t476 Vss.t253 271.079
R3520 Vss.t253 Vss.t45 271.079
R3521 Vss.t408 Vss.t320 271.079
R3522 Vss.t18 Vss.t408 271.079
R3523 Vss.t60 Vss.t321 271.079
R3524 Vss.t132 Vss.t60 271.079
R3525 Vss.t67 Vss.t640 271.079
R3526 Vss.n1786 Vss.n100 266.082
R3527 Vss.n1857 Vss.t536 259.911
R3528 Vss.n100 Vss.n56 250.827
R3529 Vss.n685 Vss.n684 250.815
R3530 Vss.n878 Vss.n574 250.815
R3531 Vss.n1201 Vss.n1200 247.475
R3532 Vss.t448 Vss.n1861 246.108
R3533 Vss.n1817 Vss.n51 245.469
R3534 Vss.n998 Vss.t199 240.12
R3535 Vss.n1469 Vss.n1468 232.143
R3536 Vss.n1467 Vss.n1466 232.143
R3537 Vss.n1473 Vss.n235 229.095
R3538 Vss.n1485 Vss.t446 228.071
R3539 Vss.n1485 Vss.t114 228.071
R3540 Vss.t637 Vss.n1484 228.071
R3541 Vss.n1484 Vss.t544 228.071
R3542 Vss.n1508 Vss.t546 228.071
R3543 Vss.t652 Vss.n536 228.004
R3544 Vss.n960 Vss.t54 228.004
R3545 Vss.t57 Vss.n545 228.004
R3546 Vss.t108 Vss.n545 228.004
R3547 Vss.n955 Vss.t106 228.004
R3548 Vss.t542 Vss.n1854 226.008
R3549 Vss.t324 Vss.t17 225.832
R3550 Vss.t658 Vss.t324 225.832
R3551 Vss.t564 Vss.t570 225.832
R3552 Vss.t570 Vss.t409 225.832
R3553 Vss.t597 Vss.t310 225.832
R3554 Vss.t310 Vss.t43 225.832
R3555 Vss.t141 Vss.t508 225.832
R3556 Vss.n1738 Vss.n1737 225.304
R3557 Vss.n698 Vss.t67 220.988
R3558 Vss.n1103 Vss.n1101 219.055
R3559 Vss.n1116 Vss.t674 215.149
R3560 Vss.n1032 Vss.n528 213.623
R3561 Vss.n1739 Vss.n1738 211.958
R3562 Vss.n1475 Vss.n231 211.958
R3563 Vss.n1843 Vss.n64 205.139
R3564 Vss.n1845 Vss.n64 205.139
R3565 Vss.n1845 Vss.n1844 205.139
R3566 Vss.n1844 Vss.n1843 205.139
R3567 Vss.n1436 Vss.n1435 200.773
R3568 Vss.t114 Vss.t637 193.861
R3569 Vss.t544 Vss.t546 193.861
R3570 Vss.t54 Vss.t57 193.804
R3571 Vss.t106 Vss.t108 193.804
R3572 Vss.n1842 Vss.n1831 193.476
R3573 Vss.n1852 Vss.n57 193.476
R3574 Vss.n239 Vss.n236 191.959
R3575 Vss.n1076 Vss.n1072 191.177
R3576 Vss.n1436 Vss.n256 186.831
R3577 Vss.n1910 Vss.n1909 181.153
R3578 Vss.n953 Vss.t551 179.683
R3579 Vss.n978 Vss.t551 179.683
R3580 Vss.t167 Vss.n1134 179.683
R3581 Vss.n1143 Vss.t167 179.683
R3582 Vss.n1139 Vss.t218 179.683
R3583 Vss.n1138 Vss.t82 179.683
R3584 Vss.t82 Vss.n235 179.683
R3585 Vss.n1416 Vss.n268 178.264
R3586 Vss.n1410 Vss.n1409 178.264
R3587 Vss.n1816 Vss.n1814 178.264
R3588 Vss.n1664 Vss.n84 178.264
R3589 Vss.n557 Vss.t148 172.196
R3590 Vss.t84 Vss.n1736 170.268
R3591 Vss.n1737 Vss.t84 170.268
R3592 Vss.n1075 Vss.n120 168.581
R3593 Vss.n955 Vss.n954 167.056
R3594 Vss.n1835 Vss.n1834 166.989
R3595 Vss.n1850 Vss.n59 166.989
R3596 Vss.n961 Vss.n960 166.254
R3597 Vss.n1396 Vss.n281 165.725
R3598 Vss.n1570 Vss.n169 165.725
R3599 Vss.n1339 Vss.n1338 165.725
R3600 Vss.n1214 Vss.n1213 165.725
R3601 Vss.n1720 Vss.n1719 165.648
R3602 Vss.n844 Vss.n592 161.839
R3603 Vss.n1049 Vss.n1048 160.189
R3604 Vss.n1692 Vss.n1684 156.166
R3605 Vss.n954 Vss.n953 154.976
R3606 Vss.n1143 Vss.n1142 152.731
R3607 Vss.n1139 Vss.n1138 152.731
R3608 Vss.n1309 Vss.n308 151.869
R3609 Vss.n374 Vss.n325 151.869
R3610 Vss.n1273 Vss.n327 151.869
R3611 Vss.n1115 Vss.n1080 151.869
R3612 Vss.n1709 Vss.n98 151.869
R3613 Vss.n478 Vss.n468 151.869
R3614 Vss.n1454 Vss.n194 151.869
R3615 Vss.n1522 Vss.n196 151.869
R3616 Vss.n1247 Vss.n345 151.869
R3617 Vss.n1469 Vss.n242 151.869
R3618 Vss.n975 Vss.n974 151.869
R3619 Vss.n1439 Vss.n1438 151.869
R3620 Vss.n1465 Vss.n246 151.869
R3621 Vss.n1802 Vss.n1801 151.869
R3622 Vss.n1592 Vss.n1591 151.869
R3623 Vss.n933 Vss.n932 151.869
R3624 Vss.n1201 Vss.n416 151.869
R3625 Vss.n797 Vss.n529 151.869
R3626 Vss.n1163 Vss.n1162 151.869
R3627 Vss.n845 Vss.n783 151.869
R3628 Vss.n626 Vss.n13 151.869
R3629 Vss.n1023 Vss.n532 151.751
R3630 Vss.n1395 Vss.n282 151.751
R3631 Vss.n1347 Vss.n1346 151.751
R3632 Vss.n1395 Vss.n283 151.751
R3633 Vss.n1346 Vss.n306 151.751
R3634 Vss.n1215 Vss.n357 151.751
R3635 Vss.n1283 Vss.n323 151.751
R3636 Vss.n404 Vss.n402 151.751
R3637 Vss.n1215 Vss.n358 151.751
R3638 Vss.n1284 Vss.n1283 151.751
R3639 Vss.n380 Vss.n379 151.751
R3640 Vss.n1331 Vss.n256 151.751
R3641 Vss.n1437 Vss.n255 151.751
R3642 Vss.n1302 Vss.n1301 151.751
R3643 Vss.n1261 Vss.n309 151.751
R3644 Vss.n1103 Vss.n1102 151.751
R3645 Vss.n1105 Vss.n1104 151.751
R3646 Vss.n137 Vss.n97 151.751
R3647 Vss.n1738 Vss.n121 151.751
R3648 Vss.n1790 Vss.n97 151.751
R3649 Vss.n1628 Vss.n56 151.751
R3650 Vss.n1643 Vss.n56 151.751
R3651 Vss.n1655 Vss.n56 151.751
R3652 Vss.n1122 Vss.n465 151.751
R3653 Vss.n488 Vss.n467 151.751
R3654 Vss.n1051 Vss.n466 151.751
R3655 Vss.n1124 Vss.n1123 151.751
R3656 Vss.n1035 Vss.n516 151.751
R3657 Vss.n1593 Vss.n156 151.751
R3658 Vss.n1470 Vss.n238 151.751
R3659 Vss.n1569 Vss.n170 151.751
R3660 Vss.n1549 Vss.n1548 151.751
R3661 Vss.n1569 Vss.n171 151.751
R3662 Vss.n1548 Vss.n1546 151.751
R3663 Vss.n1367 Vss.n245 151.751
R3664 Vss.n1532 Vss.n192 151.751
R3665 Vss.n1534 Vss.n191 151.751
R3666 Vss.n1533 Vss.n1532 151.751
R3667 Vss.n249 Vss.n248 151.751
R3668 Vss.n1427 Vss.n67 151.751
R3669 Vss.n1803 Vss.n85 151.751
R3670 Vss.n1572 Vss.n157 151.751
R3671 Vss.n1530 Vss.n1529 151.751
R3672 Vss.n1246 Vss.n1245 151.751
R3673 Vss.n1353 Vss.n290 151.751
R3674 Vss.n1384 Vss.n291 151.751
R3675 Vss.n292 Vss.n290 151.751
R3676 Vss.n1384 Vss.n1383 151.751
R3677 Vss.n1678 Vss.n1677 151.751
R3678 Vss.n1738 Vss.n123 151.751
R3679 Vss.n1733 Vss.n1732 151.751
R3680 Vss.n1738 Vss.n124 151.751
R3681 Vss.n1281 Vss.n1280 151.751
R3682 Vss.n1189 Vss.n1187 151.751
R3683 Vss.n1188 Vss.n362 151.751
R3684 Vss.n807 Vss.n806 151.751
R3685 Vss.n787 Vss.n515 151.751
R3686 Vss.n1047 Vss.n1046 151.751
R3687 Vss.n931 Vss.n930 151.751
R3688 Vss.n842 Vss.n785 151.751
R3689 Vss.n830 Vss.n784 151.751
R3690 Vss.n812 Vss.n811 151.751
R3691 Vss.n642 Vss.n641 151.751
R3692 Vss.n644 Vss.n643 151.751
R3693 Vss.n655 Vss.n654 151.751
R3694 Vss.n10 Vss.n9 151.751
R3695 Vss.n1911 Vss.n1910 151.751
R3696 Vss.n1910 Vss.n7 151.751
R3697 Vss.n1910 Vss.n8 151.751
R3698 Vss.n657 Vss.n656 151.751
R3699 Vss.n885 Vss.n573 151.751
R3700 Vss.n1000 Vss.n999 147.727
R3701 Vss.n1007 Vss.n514 147.727
R3702 Vss.n611 Vss.n610 147.727
R3703 Vss.n847 Vss.n591 147.727
R3704 Vss.n26 Vss.n14 147.727
R3705 Vss.n1895 Vss.n15 147.727
R3706 Vss.n899 Vss.n898 147.727
R3707 Vss.n904 Vss.n531 147.727
R3708 Vss.n1142 Vss.n237 143.746
R3709 Vss.t148 Vss.t463 137.756
R3710 Vss.t463 Vss.t242 137.756
R3711 Vss.n1396 Vss.n1395 135.501
R3712 Vss.n1570 Vss.n1569 135.501
R3713 Vss.n1338 Vss.n290 135.501
R3714 Vss.n1215 Vss.n1214 135.501
R3715 Vss.n1719 Vss.n97 135.439
R3716 Vss.n1743 Vss.n1742 129.76
R3717 Vss.t45 Vss.n528 125.228
R3718 Vss.n1857 Vss.t540 124.305
R3719 Vss.n1694 Vss.t101 120.279
R3720 Vss.t662 Vss.n446 119.157
R3721 Vss.n447 Vss.t662 119.157
R3722 Vss.n1840 Vss.n1839 118.222
R3723 Vss.n326 Vss.t323 115.856
R3724 Vss.t427 Vss.n281 115.856
R3725 Vss.n195 Vss.t304 115.856
R3726 Vss.t635 Vss.n169 115.856
R3727 Vss.n1344 Vss.t330 115.856
R3728 Vss.n1339 Vss.t239 115.856
R3729 Vss.n297 Vss.t326 115.856
R3730 Vss.t58 Vss.n243 115.856
R3731 Vss.n1202 Vss.t307 115.856
R3732 Vss.n1213 Vss.t255 115.856
R3733 Vss.t576 Vss.n142 115.802
R3734 Vss.n1720 Vss.t230 115.802
R3735 Vss.n1594 Vss.t565 114.944
R3736 Vss.n1610 Vss.t565 114.944
R3737 Vss.t247 Vss.n1614 114.944
R3738 Vss.t242 Vss.n459 113.799
R3739 Vss.n447 Vss.n424 113.695
R3740 Vss.n1478 Vss.n230 113.215
R3741 Vss.n1024 Vss.n1023 108.731
R3742 Vss.t382 Vss.t175 108.138
R3743 Vss.t211 Vss.t459 108.138
R3744 Vss.t260 Vss.t436 108.138
R3745 Vss.t214 Vss.t435 108.138
R3746 Vss.t336 Vss.t209 108.138
R3747 Vss.t669 Vss.t261 108.138
R3748 Vss.t339 Vss.t213 108.138
R3749 Vss.t685 Vss.t217 108.138
R3750 Vss.t508 Vss.n1694 105.552
R3751 Vss.n1909 Vss.n1908 103.79
R3752 Vss.n446 Vss.n434 102.773
R3753 Vss.n1856 Vss.t542 101.704
R3754 Vss.t2 Vss.t210 99.0183
R3755 Vss.t263 Vss.t2 99.0183
R3756 Vss.n1614 Vss.n1610 97.7016
R3757 Vss.n1906 Vss.t417 97.5981
R3758 Vss.t469 Vss.n470 96.5949
R3759 Vss.n668 Vss.t516 96.5352
R3760 Vss.n896 Vss.t482 96.5352
R3761 Vss.n1395 Vss.n1394 95.5419
R3762 Vss.n1346 Vss.n307 95.5419
R3763 Vss.n1216 Vss.n1215 95.5419
R3764 Vss.n1283 Vss.n324 95.5419
R3765 Vss.n1569 Vss.n1568 95.5419
R3766 Vss.n1548 Vss.n1547 95.5419
R3767 Vss.n1466 Vss.n244 95.5419
R3768 Vss.n1532 Vss.n193 95.5419
R3769 Vss.n1386 Vss.n290 95.5419
R3770 Vss.n1385 Vss.n1384 95.5419
R3771 Vss.n1559 Vss.n97 95.4017
R3772 Vss.n1738 Vss.n122 95.4017
R3773 Vss.t323 Vss.t244 92.6849
R3774 Vss.t244 Vss.t427 92.6849
R3775 Vss.t304 Vss.t126 92.6849
R3776 Vss.t126 Vss.t635 92.6849
R3777 Vss.t443 Vss.t330 92.6849
R3778 Vss.t239 Vss.t443 92.6849
R3779 Vss.t326 Vss.t127 92.6849
R3780 Vss.t127 Vss.t58 92.6849
R3781 Vss.t307 Vss.t185 92.6849
R3782 Vss.t185 Vss.t255 92.6849
R3783 Vss.t272 Vss.t576 92.6419
R3784 Vss.t230 Vss.t272 92.6419
R3785 Vss.t175 Vss.t211 89.8983
R3786 Vss.t459 Vss.t260 89.8983
R3787 Vss.t436 Vss.t214 89.8983
R3788 Vss.t435 Vss.t262 89.8983
R3789 Vss.t212 Vss.t336 89.8983
R3790 Vss.t209 Vss.t669 89.8983
R3791 Vss.t261 Vss.t339 89.8983
R3792 Vss.t213 Vss.t685 89.8983
R3793 Vss.n1027 Vss.n1026 88.3958
R3794 Vss.n856 Vss.n586 87.3061
R3795 Vss.n856 Vss.n587 87.3061
R3796 Vss.n763 Vss.n686 87.3061
R3797 Vss.n763 Vss.n762 87.3061
R3798 Vss.n905 Vss.n570 87.3061
R3799 Vss.n905 Vss.n903 87.3061
R3800 Vss.n956 Vss.n952 87.3061
R3801 Vss.n957 Vss.n956 87.3061
R3802 Vss.n1507 Vss.n213 87.3061
R3803 Vss.n1507 Vss.n214 87.3061
R3804 Vss.n1497 Vss.n217 87.3061
R3805 Vss.n1497 Vss.n218 87.3061
R3806 Vss.n1769 Vss.n107 87.3061
R3807 Vss.n1769 Vss.n108 87.3061
R3808 Vss.n1785 Vss.n101 87.3061
R3809 Vss.n1785 Vss.n102 87.3061
R3810 Vss.n1008 Vss.n543 87.3061
R3811 Vss.n1008 Vss.n544 87.3061
R3812 Vss.n441 Vss.n433 87.3061
R3813 Vss.n442 Vss.n433 87.3061
R3814 Vss.n777 Vss.n596 87.3061
R3815 Vss.n777 Vss.n597 87.3061
R3816 Vss.n1894 Vss.n18 87.3061
R3817 Vss.n1894 Vss.n19 87.3061
R3818 Vss.n1595 Vss.n1594 86.8248
R3819 Vss.n1842 Vss.t382 80.7782
R3820 Vss.n1841 Vss.t134 80.7782
R3821 Vss.n1838 Vss.t356 80.7782
R3822 Vss.t217 Vss.n57 80.7782
R3823 Vss.n1835 Vss.n59 80.5005
R3824 Vss.n401 Vss.n400 76.452
R3825 Vss.n1695 Vss.n56 73.641
R3826 Vss.n1162 Vss.n434 72.984
R3827 Vss.t419 Vss.t415 72.1379
R3828 Vss.t450 Vss.t134 69.0524
R3829 Vss.t356 Vss.t386 69.0524
R3830 Vss.n604 Vss.n603 67.4727
R3831 Vss.n605 Vss.n603 67.4727
R3832 Vss.n688 Vss.n31 67.4727
R3833 Vss.n761 Vss.n31 67.4727
R3834 Vss.n572 Vss.n567 67.4727
R3835 Vss.n902 Vss.n567 67.4727
R3836 Vss.n950 Vss.n552 67.4727
R3837 Vss.n958 Vss.n552 67.4727
R3838 Vss.n226 Vss.n225 67.4727
R3839 Vss.n227 Vss.n225 67.4727
R3840 Vss.n228 Vss.n221 67.4727
R3841 Vss.n229 Vss.n221 67.4727
R3842 Vss.n1740 Vss.n111 67.4727
R3843 Vss.n1741 Vss.n111 67.4727
R3844 Vss.n116 Vss.n115 67.4727
R3845 Vss.n117 Vss.n115 67.4727
R3846 Vss.n1001 Vss.n540 67.4727
R3847 Vss.n1002 Vss.n540 67.4727
R3848 Vss.n863 Vss.n584 67.4727
R3849 Vss.n863 Vss.n585 67.4727
R3850 Vss.n606 Vss.n599 67.4727
R3851 Vss.n607 Vss.n599 67.4727
R3852 Vss.n27 Vss.n22 67.4727
R3853 Vss.n27 Vss.n23 67.4727
R3854 Vss.n1733 Vss.n125 67.0503
R3855 Vss.n1897 Vss.n15 66.9416
R3856 Vss.t515 Vss.n1057 66.9123
R3857 Vss.n604 Vss.n586 66.5005
R3858 Vss.n605 Vss.n587 66.5005
R3859 Vss.n688 Vss.n686 66.5005
R3860 Vss.n762 Vss.n761 66.5005
R3861 Vss.n572 Vss.n570 66.5005
R3862 Vss.n903 Vss.n902 66.5005
R3863 Vss.n952 Vss.n950 66.5005
R3864 Vss.n958 Vss.n957 66.5005
R3865 Vss.n226 Vss.n213 66.5005
R3866 Vss.n227 Vss.n214 66.5005
R3867 Vss.n228 Vss.n217 66.5005
R3868 Vss.n229 Vss.n218 66.5005
R3869 Vss.n1740 Vss.n107 66.5005
R3870 Vss.n1741 Vss.n108 66.5005
R3871 Vss.n116 Vss.n101 66.5005
R3872 Vss.n117 Vss.n102 66.5005
R3873 Vss.n1001 Vss.n543 66.5005
R3874 Vss.n1002 Vss.n544 66.5005
R3875 Vss.n584 Vss.n441 66.5005
R3876 Vss.n585 Vss.n442 66.5005
R3877 Vss.n606 Vss.n596 66.5005
R3878 Vss.n607 Vss.n597 66.5005
R3879 Vss.n22 Vss.n18 66.5005
R3880 Vss.n23 Vss.n19 66.5005
R3881 Vss.n1900 Vss.t642 65.7728
R3882 Vss.n47 Vss.n46 65.5283
R3883 Vss.n1864 Vss.n46 65.5283
R3884 Vss.n1865 Vss.n1864 65.5283
R3885 Vss.n1865 Vss.n47 65.5283
R3886 Vss.n396 Vss.t156 63.4555
R3887 Vss.t530 Vss.n270 63.4555
R3888 Vss.n1411 Vss.t654 63.4555
R3889 Vss.n1415 Vss.t351 63.4555
R3890 Vss.n1418 Vss.t363 63.4555
R3891 Vss.t402 Vss.n1417 63.4555
R3892 Vss.n1481 Vss.n1479 62.511
R3893 Vss.n402 Vss.n401 62.5094
R3894 Vss.n1615 Vss.n125 61.7821
R3895 Vss.n961 Vss.t652 61.7514
R3896 Vss.n405 Vss.n389 61.0571
R3897 Vss.n1285 Vss.n322 61.0571
R3898 Vss.n381 Vss.n370 61.0571
R3899 Vss.n1106 Vss.n1086 61.0571
R3900 Vss.n1704 Vss.n1629 61.0571
R3901 Vss.n1644 Vss.n1641 61.0571
R3902 Vss.n490 Vss.n489 61.0571
R3903 Vss.n1031 Vss.n1028 61.0571
R3904 Vss.n1528 Vss.n197 61.0571
R3905 Vss.n1731 Vss.n126 61.0571
R3906 Vss.n805 Vss.n788 61.0571
R3907 Vss.n1165 Vss.n1164 61.0571
R3908 Vss.n831 Vss.n829 61.0571
R3909 Vss.n645 Vss.n625 61.0571
R3910 Vss.n739 Vss.n690 61.0561
R3911 Vss.n886 Vss.n580 61.0561
R3912 Vss.n894 Vss.n577 61.0561
R3913 Vss.n879 Vss.n582 61.0561
R3914 Vss.n1876 Vss.n38 61.0561
R3915 Vss.n839 Vss.n813 61.0561
R3916 Vss.n822 Vss.n821 61.0561
R3917 Vss.n1182 Vss.n426 61.0561
R3918 Vss.n1045 Vss.n517 61.0561
R3919 Vss.n798 Vss.n795 61.0561
R3920 Vss.n996 Vss.n990 61.0561
R3921 Vss.n921 Vss.n919 61.0561
R3922 Vss.n1199 Vss.n417 61.0561
R3923 Vss.n415 Vss.n365 61.0561
R3924 Vss.n399 Vss.n397 61.0561
R3925 Vss.n1212 Vss.n1203 61.0561
R3926 Vss.n1279 Vss.n328 61.0561
R3927 Vss.n935 Vss.n929 61.0561
R3928 Vss.n1582 Vss.n1581 61.0561
R3929 Vss.n1590 Vss.n158 61.0561
R3930 Vss.n1721 Vss.n141 61.0561
R3931 Vss.n1716 Vss.n1619 61.0561
R3932 Vss.n1800 Vss.n87 61.0561
R3933 Vss.n1666 Vss.n1663 61.0561
R3934 Vss.n1696 Vss.n1639 61.0561
R3935 Vss.n1690 Vss.n1688 61.0561
R3936 Vss.n1819 Vss.n74 61.0561
R3937 Vss.n1825 Vss.n69 61.0561
R3938 Vss.n1434 Vss.n258 61.0561
R3939 Vss.n1441 Vss.n1440 61.0561
R3940 Vss.n299 Vss.n298 61.0561
R3941 Vss.n1387 Vss.n289 61.0561
R3942 Vss.n1382 Vss.n293 61.0561
R3943 Vss.n1355 Vss.n1354 61.0561
R3944 Vss.n1343 Vss.n1340 61.0561
R3945 Vss.n1244 Vss.n347 61.0561
R3946 Vss.n972 Vss.n336 61.0561
R3947 Vss.n970 Vss.n964 61.0561
R3948 Vss.n947 Vss.n559 61.0561
R3949 Vss.n1224 Vss.n1223 61.0561
R3950 Vss.n1393 Vss.n284 61.0561
R3951 Vss.n1294 Vss.n1293 61.0561
R3952 Vss.n1348 Vss.n305 61.0561
R3953 Vss.n1217 Vss.n356 61.0561
R3954 Vss.n1206 Vss.n1205 61.0561
R3955 Vss.n1304 Vss.n1303 61.0561
R3956 Vss.n375 Vss.n373 61.0561
R3957 Vss.n1408 Vss.n272 61.0561
R3958 Vss.n1419 Vss.n266 61.0561
R3959 Vss.n1414 Vss.n1412 61.0561
R3960 Vss.n395 Vss.n390 61.0561
R3961 Vss.n1328 Vss.n313 61.0561
R3962 Vss.n1334 Vss.n1332 61.0561
R3963 Vss.n1402 Vss.n277 61.0561
R3964 Vss.n1317 Vss.n1315 61.0561
R3965 Vss.n1311 Vss.n1310 61.0561
R3966 Vss.n1262 Vss.n334 61.0561
R3967 Vss.n1274 Vss.n1271 61.0561
R3968 Vss.n1132 Vss.n460 61.0561
R3969 Vss.n1251 Vss.n343 61.0561
R3970 Vss.n1239 Vss.n1238 61.0561
R3971 Vss.n1597 Vss.n153 61.0561
R3972 Vss.n1114 Vss.n1081 61.0561
R3973 Vss.n1098 Vss.n1088 61.0561
R3974 Vss.n1071 Vss.n1058 61.0561
R3975 Vss.n1063 Vss.n1062 61.0561
R3976 Vss.n1560 Vss.n1558 61.0561
R3977 Vss.n138 Vss.n136 61.0561
R3978 Vss.n1791 Vss.n96 61.0561
R3979 Vss.n1683 Vss.n1680 61.0561
R3980 Vss.n1675 Vss.n1673 61.0561
R3981 Vss.n1656 Vss.n1654 61.0561
R3982 Vss.n1710 Vss.n1625 61.0561
R3983 Vss.n511 Vss.n505 61.0561
R3984 Vss.n1125 Vss.n464 61.0561
R3985 Vss.n499 Vss.n472 61.0561
R3986 Vss.n480 Vss.n479 61.0561
R3987 Vss.n1036 Vss.n525 61.0561
R3988 Vss.n206 Vss.n204 61.0561
R3989 Vss.n1512 Vss.n212 61.0561
R3990 Vss.n1359 Vss.n1358 61.0561
R3991 Vss.n1567 Vss.n172 61.0561
R3992 Vss.n1545 Vss.n177 61.0561
R3993 Vss.n1550 Vss.n176 61.0561
R3994 Vss.n1375 Vss.n1374 61.0561
R3995 Vss.n1535 Vss.n190 61.0561
R3996 Vss.n1368 Vss.n1366 61.0561
R3997 Vss.n180 Vss.n179 61.0561
R3998 Vss.n1455 Vss.n1452 61.0561
R3999 Vss.n1813 Vss.n76 61.0561
R4000 Vss.n1807 Vss.n81 61.0561
R4001 Vss.n1428 Vss.n1425 61.0561
R4002 Vss.n1461 Vss.n250 61.0561
R4003 Vss.n1574 Vss.n165 61.0561
R4004 Vss.n1523 Vss.n1521 61.0561
R4005 Vss.n1190 Vss.n422 61.0561
R4006 Vss.n438 Vss.n435 61.0561
R4007 Vss.n658 Vss.n617 61.0561
R4008 Vss.n666 Vss.n615 61.0561
R4009 Vss.n653 Vss.n620 61.0561
R4010 Vss.n637 Vss.n627 61.0561
R4011 Vss.n1912 Vss.n6 61.0561
R4012 Vss.n705 Vss.n699 61.0561
R4013 Vss.n732 Vss.n731 61.0561
R4014 Vss.n716 Vss.n715 61.0561
R4015 Vss.n724 Vss.n707 61.0561
R4016 Vss.n1753 Vss.t389 60.019
R4017 Vss.n1753 Vss.t228 60.019
R4018 Vss.t229 Vss.n1752 60.019
R4019 Vss.n1752 Vss.t280 60.019
R4020 Vss.t282 Vss.n1786 60.019
R4021 Vss.n1133 Vss.n459 58.3972
R4022 Vss.n1472 Vss.n236 57.018
R4023 Vss.n1738 Vss.t389 54.0171
R4024 Vss.n1435 Vss.t571 53.4468
R4025 Vss.n257 Vss.t364 53.4468
R4026 Vss.t306 Vss.n363 53.4468
R4027 Vss.n400 Vss.t354 53.4468
R4028 Vss.n1615 Vss.t247 53.1614
R4029 Vss.n1905 Vss.t413 53.0427
R4030 Vss.t228 Vss.t229 51.0162
R4031 Vss.t156 Vss.t322 50.7645
R4032 Vss.t322 Vss.t530 50.7645
R4033 Vss.t654 Vss.t316 50.7645
R4034 Vss.t316 Vss.t351 50.7645
R4035 Vss.t363 Vss.t317 50.7645
R4036 Vss.t317 Vss.t402 50.7645
R4037 Vss.t475 Vss.n698 50.0912
R4038 Vss.n1901 Vss.t413 48.7993
R4039 Vss.n1736 Vss.n1733 45.4054
R4040 Vss.n1185 Vss.n423 45.3808
R4041 Vss.n1735 Vss.n114 44.1404
R4042 Vss.n678 Vss.n677 44.1404
R4043 Vss.n674 Vss.n602 44.1404
R4044 Vss.n744 Vss.n30 44.1394
R4045 Vss.n748 Vss.n747 44.1394
R4046 Vss.n755 Vss.n751 44.1394
R4047 Vss.n867 Vss.n866 44.1394
R4048 Vss.n871 Vss.n565 44.1394
R4049 Vss.n876 Vss.n875 44.1394
R4050 Vss.n851 Vss.n590 44.1394
R4051 Vss.n682 Vss.n681 44.1394
R4052 Vss.n1879 Vss.n36 44.1394
R4053 Vss.n448 Vss.n445 44.1394
R4054 Vss.n988 Vss.n551 44.1394
R4055 Vss.n1015 Vss.n538 44.1394
R4056 Vss.n1018 Vss.n451 44.1394
R4057 Vss.n1613 Vss.n1612 44.1394
R4058 Vss.n1609 Vss.n145 44.1394
R4059 Vss.n1137 Vss.n224 44.1394
R4060 Vss.n1141 Vss.n1140 44.1394
R4061 Vss.n1144 Vss.n458 44.1394
R4062 Vss.n979 Vss.n556 44.1394
R4063 Vss.n1501 Vss.n216 44.1394
R4064 Vss.n1774 Vss.n1772 44.1394
R4065 Vss.n1779 Vss.n105 44.1394
R4066 Vss.t660 Vss.t571 42.7575
R4067 Vss.t364 Vss.t660 42.7575
R4068 Vss.t353 Vss.t306 42.7575
R4069 Vss.t354 Vss.t353 42.7575
R4070 Vss.n1174 Vss.t691 41.0041
R4071 Vss.n1195 Vss.t687 41.0041
R4072 Vss.n1636 Vss.t690 41.0041
R4073 Vss.n1175 Vss.t689 40.8177
R4074 Vss.n1787 Vss.t280 38.0122
R4075 Vss.n1187 Vss.n1185 37.1047
R4076 Vss.n239 Vss.t446 36.1116
R4077 Vss.t642 Vss.n0 36.0692
R4078 Vss.t218 Vss.n237 35.9369
R4079 Vss.n1186 Vss.t94 35.0024
R4080 Vss.n1200 Vss.t678 35.0024
R4081 Vss.n1765 Vss.t688 34.1066
R4082 Vss.t538 Vss.n52 33.9022
R4083 Vss.n439 Vss.t325 31.7253
R4084 Vss.t424 Vss.n423 31.7253
R4085 Vss.n757 Vss.n740 30.7136
R4086 Vss.n65 Vss.n64 30.5283
R4087 Vss.n1844 Vss.n65 30.5283
R4088 Vss.n1467 Vss.n243 30.2237
R4089 Vss.n1202 Vss.n1201 30.2237
R4090 Vss.n1858 Vss.n1857 29.4859
R4091 Vss.t94 Vss.t312 28.002
R4092 Vss.t312 Vss.t678 28.002
R4093 Vss.n1856 Vss.n1855 27.3737
R4094 Vss.t262 Vss.n1841 27.3607
R4095 Vss.n1838 Vss.t212 27.3607
R4096 Vss.n1175 Vss.t91 27.1302
R4097 Vss.n1174 Vss.t98 26.9438
R4098 Vss.n1195 Vss.t93 26.9438
R4099 Vss.n1636 Vss.t100 26.9438
R4100 Vss.t325 Vss.t383 25.3804
R4101 Vss.t383 Vss.t424 25.3804
R4102 Vss.n1778 Vss.t115 24.9198
R4103 Vss.n1024 Vss.n424 24.8248
R4104 Vss.t378 Vss.n758 24.1401
R4105 Vss.n759 Vss.t378 24.1401
R4106 Vss.n759 Vss.t684 24.1401
R4107 Vss.t254 Vss.n16 24.1401
R4108 Vss.t194 Vss.n16 24.1401
R4109 Vss.n764 Vss.t196 24.1401
R4110 Vss.t577 Vss.n766 24.1401
R4111 Vss.n767 Vss.t577 24.1401
R4112 Vss.n767 Vss.t430 24.1401
R4113 Vss.t429 Vss.n595 24.1401
R4114 Vss.n595 Vss.t137 24.1401
R4115 Vss.n857 Vss.t135 24.1401
R4116 Vss.n862 Vss.t143 24.1401
R4117 Vss.t143 Vss.n861 24.1401
R4118 Vss.n861 Vss.t241 24.1401
R4119 Vss.n1161 Vss.t237 24.1401
R4120 Vss.t453 Vss.n1161 24.1401
R4121 Vss.n1901 Vss.t419 23.3391
R4122 Vss.t210 Vss.t450 20.8464
R4123 Vss.t386 Vss.t263 20.8464
R4124 Vss.n594 Vss.n586 20.8061
R4125 Vss.n594 Vss.n587 20.8061
R4126 Vss.n768 Vss.n604 20.8061
R4127 Vss.n768 Vss.n605 20.8061
R4128 Vss.n687 Vss.n686 20.8061
R4129 Vss.n762 Vss.n687 20.8061
R4130 Vss.n760 Vss.n688 20.8061
R4131 Vss.n761 Vss.n760 20.8061
R4132 Vss.n571 Vss.n570 20.8061
R4133 Vss.n903 Vss.n571 20.8061
R4134 Vss.n901 Vss.n572 20.8061
R4135 Vss.n902 Vss.n901 20.8061
R4136 Vss.n952 Vss.n951 20.8061
R4137 Vss.n957 Vss.n951 20.8061
R4138 Vss.n959 Vss.n950 20.8061
R4139 Vss.n959 Vss.n958 20.8061
R4140 Vss.n1483 Vss.n213 20.8061
R4141 Vss.n1483 Vss.n214 20.8061
R4142 Vss.n1486 Vss.n226 20.8061
R4143 Vss.n1486 Vss.n227 20.8061
R4144 Vss.n1480 Vss.n217 20.8061
R4145 Vss.n1480 Vss.n218 20.8061
R4146 Vss.n230 Vss.n228 20.8061
R4147 Vss.n230 Vss.n229 20.8061
R4148 Vss.n1748 Vss.n107 20.8061
R4149 Vss.n1748 Vss.n108 20.8061
R4150 Vss.n1742 Vss.n1740 20.8061
R4151 Vss.n1742 Vss.n1741 20.8061
R4152 Vss.n1866 Vss.n46 20.8061
R4153 Vss.n1866 Vss.n1865 20.8061
R4154 Vss.n1751 Vss.n101 20.8061
R4155 Vss.n1751 Vss.n102 20.8061
R4156 Vss.n1754 Vss.n116 20.8061
R4157 Vss.n1754 Vss.n117 20.8061
R4158 Vss.n1003 Vss.n1001 20.8061
R4159 Vss.n1003 Vss.n1002 20.8061
R4160 Vss.n1005 Vss.n543 20.8061
R4161 Vss.n1005 Vss.n544 20.8061
R4162 Vss.n860 Vss.n584 20.8061
R4163 Vss.n860 Vss.n585 20.8061
R4164 Vss.n1160 Vss.n441 20.8061
R4165 Vss.n1160 Vss.n442 20.8061
R4166 Vss.n781 Vss.n596 20.8061
R4167 Vss.n781 Vss.n597 20.8061
R4168 Vss.n608 Vss.n606 20.8061
R4169 Vss.n608 Vss.n607 20.8061
R4170 Vss.n18 Vss.n17 20.8061
R4171 Vss.n19 Vss.n17 20.8061
R4172 Vss.n24 Vss.n22 20.8061
R4173 Vss.n24 Vss.n23 20.8061
R4174 Vss.t684 Vss.t254 20.5192
R4175 Vss.t196 Vss.t194 20.5192
R4176 Vss.t430 Vss.t429 20.5192
R4177 Vss.t137 Vss.t135 20.5192
R4178 Vss.t241 Vss.t237 20.5192
R4179 Vss.t455 Vss.t453 20.5192
R4180 Vss.n1830 Vss.n1829 19.8869
R4181 Vss.n1764 Vss.t88 19.673
R4182 Vss.n1764 Vss.t95 19.4007
R4183 Vss.t417 Vss.n1905 19.0957
R4184 Vss.n1839 Vss.n59 18.8616
R4185 Vss.n1840 Vss.n1835 18.8616
R4186 Vss.t115 Vss.n56 18.5862
R4187 Vss.n63 comparator_no_offsetcal_0.x3.avss 17.8218
R4188 Vss.n1859 Vss.n52 17.4164
R4189 Vss.n1870 comparator_no_offsetcal_0.x5.avss 16.7565
R4190 Vss.n402 Vss.n396 16.554
R4191 Vss.n1417 Vss.n256 16.554
R4192 Vss.n1776 Vss.n100 16.1938
R4193 Vss.n257 Vss.n68 15.5696
R4194 Vss.n1162 Vss.t455 14.6854
R4195 Vss.n1767 Vss.n1766 14.6135
R4196 Vss.n1201 Vss.n363 13.943
R4197 Vss.n1637 SARlogic_0.dffrs_13.d 13.7563
R4198 Vss.n1177 SARlogic_0.dffrs_12.clk 13.599
R4199 Vss.n1196 SARlogic_0.dffrs_12.d 13.599
R4200 Vss.n1787 Vss.t282 13.0045
R4201 Vss.n1837 Vss.n1836 11.0305
R4202 Vss.n1900 Vss.n1899 10.4005
R4203 Vss.n1902 Vss.n1901 10.4005
R4204 Vss.n1905 Vss.n1904 10.4005
R4205 Vss.n1917 Vss.n0 10.4005
R4206 Vss.n1187 Vss.n1186 9.13142
R4207 Vss.n1871 Vss.n1870 9.05474
R4208 Vss.n1698 Vss.n1637 9.04466
R4209 Vss.n1197 Vss.n1196 9.04027
R4210 Vss.n394 Vss.n387 9.03475
R4211 Vss.n1193 Vss.n418 9.03475
R4212 Vss.n838 Vss.n837 9.0005
R4213 Vss.n581 Vss.n579 9.0005
R4214 Vss.n890 Vss.n889 9.0005
R4215 Vss.n519 Vss.n518 9.0005
R4216 Vss.n918 Vss.n917 9.0005
R4217 Vss.n1277 Vss.n1276 9.0005
R4218 Vss.n295 Vss.n294 9.0005
R4219 Vss.n407 Vss.n406 9.0005
R4220 Vss.n321 Vss.n319 9.0005
R4221 Vss.n385 Vss.n384 9.0005
R4222 Vss.n414 Vss.n413 9.0005
R4223 Vss.n412 Vss.n367 9.0005
R4224 Vss.n1321 Vss.n1320 9.0005
R4225 Vss.n1314 Vss.n1313 9.0005
R4226 Vss.n1266 Vss.n1265 9.0005
R4227 Vss.n966 Vss.n965 9.0005
R4228 Vss.n1269 Vss.n1268 9.0005
R4229 Vss.n348 Vss.n338 9.0005
R4230 Vss.n1257 Vss.n1256 9.0005
R4231 Vss.n1253 Vss.n1252 9.0005
R4232 Vss.n1066 Vss.n152 9.0005
R4233 Vss.n1068 Vss.n1067 9.0005
R4234 Vss.n1085 Vss.n1084 9.0005
R4235 Vss.n1109 Vss.n1108 9.0005
R4236 Vss.n1090 Vss.n1089 9.0005
R4237 Vss.n1096 Vss.n1095 9.0005
R4238 Vss.n1083 Vss.n1082 9.0005
R4239 Vss.n1112 Vss.n1111 9.0005
R4240 Vss.n1069 Vss.n151 9.0005
R4241 Vss.n1600 Vss.n1599 9.0005
R4242 Vss.n1653 Vss.n1652 9.0005
R4243 Vss.n1635 Vss.n1631 9.0005
R4244 Vss.n1648 Vss.n1647 9.0005
R4245 Vss.n1646 Vss.n1640 9.0005
R4246 Vss.n1659 Vss.n1658 9.0005
R4247 Vss.n1650 Vss.n1623 9.0005
R4248 Vss.n507 Vss.n461 9.0005
R4249 Vss.n487 Vss.n486 9.0005
R4250 Vss.n493 Vss.n492 9.0005
R4251 Vss.n477 Vss.n476 9.0005
R4252 Vss.n483 Vss.n482 9.0005
R4253 Vss.n498 Vss.n473 9.0005
R4254 Vss.n497 Vss.n495 9.0005
R4255 Vss.n1130 Vss.n1129 9.0005
R4256 Vss.n508 Vss.n463 9.0005
R4257 Vss.n1128 Vss.n1127 9.0005
R4258 Vss.n995 Vss.n994 9.0005
R4259 Vss.n993 Vss.n524 9.0005
R4260 Vss.n1039 Vss.n1038 9.0005
R4261 Vss.n992 Vss.n523 9.0005
R4262 Vss.n1541 Vss.n1540 9.0005
R4263 Vss.n184 Vss.n183 9.0005
R4264 Vss.n1450 Vss.n1449 9.0005
R4265 Vss.n199 Vss.n198 9.0005
R4266 Vss.n1236 Vss.n1235 9.0005
R4267 Vss.n1730 Vss.n1729 9.0005
R4268 Vss.n1728 Vss.n128 9.0005
R4269 Vss.n1588 Vss.n1586 9.0005
R4270 Vss.n1584 Vss.n1583 9.0005
R4271 Vss.n1579 Vss.n130 9.0005
R4272 Vss.n134 Vss.n131 9.0005
R4273 Vss.n1556 Vss.n1555 9.0005
R4274 Vss.n1714 Vss.n1712 9.0005
R4275 Vss.n1712 Vss.n1711 9.0005
R4276 Vss.n1620 Vss.n94 9.0005
R4277 Vss.n1700 Vss.n1638 9.0005
R4278 Vss.n1700 Vss.n1699 9.0005
R4279 Vss.n1702 Vss.n1633 9.0005
R4280 Vss.n1703 Vss.n1702 9.0005
R4281 Vss.n1685 Vss.n72 9.0005
R4282 Vss.n1686 Vss.n1685 9.0005
R4283 Vss.n1670 Vss.n79 9.0005
R4284 Vss.n1671 Vss.n1670 9.0005
R4285 Vss.n182 Vss.n88 9.0005
R4286 Vss.n1799 Vss.n88 9.0005
R4287 Vss.n1543 Vss.n1542 9.0005
R4288 Vss.n1798 Vss.n1796 9.0005
R4289 Vss.n1715 Vss.n91 9.0005
R4290 Vss.n1793 Vss.n1792 9.0005
R4291 Vss.n1565 Vss.n1563 9.0005
R4292 Vss.n1562 Vss.n1561 9.0005
R4293 Vss.n1553 Vss.n1552 9.0005
R4294 Vss.n140 Vss.n139 9.0005
R4295 Vss.n163 Vss.n162 9.0005
R4296 Vss.n1589 Vss.n159 9.0005
R4297 Vss.n202 Vss.n160 9.0005
R4298 Vss.n1519 Vss.n1518 9.0005
R4299 Vss.n1576 Vss.n1575 9.0005
R4300 Vss.n208 Vss.n207 9.0005
R4301 Vss.n1232 Vss.n211 9.0005
R4302 Vss.n1526 Vss.n1525 9.0005
R4303 Vss.n1525 Vss.n1524 9.0005
R4304 Vss.n1515 Vss.n1514 9.0005
R4305 Vss.n1372 Vss.n173 9.0005
R4306 Vss.n1566 Vss.n173 9.0005
R4307 Vss.n1364 Vss.n1363 9.0005
R4308 Vss.n1363 Vss.n175 9.0005
R4309 Vss.n1459 Vss.n1457 9.0005
R4310 Vss.n1457 Vss.n1456 9.0005
R4311 Vss.n188 Vss.n186 9.0005
R4312 Vss.n1823 Vss.n1821 9.0005
R4313 Vss.n1821 Vss.n1820 9.0005
R4314 Vss.n1809 Vss.n78 9.0005
R4315 Vss.n1809 Vss.n1808 9.0005
R4316 Vss.n264 Vss.n70 9.0005
R4317 Vss.n1824 Vss.n70 9.0005
R4318 Vss.n1430 Vss.n260 9.0005
R4319 Vss.n1430 Vss.n1429 9.0005
R4320 Vss.n1319 Vss.n1316 9.0005
R4321 Vss.n1316 Vss.n253 9.0005
R4322 Vss.n1380 Vss.n1379 9.0005
R4323 Vss.n1444 Vss.n1443 9.0005
R4324 Vss.n1460 Vss.n1446 9.0005
R4325 Vss.n1537 Vss.n1536 9.0005
R4326 Vss.n1377 Vss.n287 9.0005
R4327 Vss.n1377 Vss.n1376 9.0005
R4328 Vss.n1370 Vss.n1357 9.0005
R4329 Vss.n1370 Vss.n1369 9.0005
R4330 Vss.n1242 Vss.n1241 9.0005
R4331 Vss.n1241 Vss.n1240 9.0005
R4332 Vss.n349 Vss.n341 9.0005
R4333 Vss.n1264 Vss.n1259 9.0005
R4334 Vss.n1259 Vss.n1258 9.0005
R4335 Vss.n968 Vss.n967 9.0005
R4336 Vss.n1391 Vss.n1389 9.0005
R4337 Vss.n1389 Vss.n1388 9.0005
R4338 Vss.n1351 Vss.n1350 9.0005
R4339 Vss.n1352 Vss.n1351 9.0005
R4340 Vss.n1299 Vss.n314 9.0005
R4341 Vss.n1308 Vss.n314 9.0005
R4342 Vss.n1291 Vss.n316 9.0005
R4343 Vss.n1421 Vss.n263 9.0005
R4344 Vss.n1421 Vss.n1420 9.0005
R4345 Vss.n275 Vss.n262 9.0005
R4346 Vss.n1333 Vss.n262 9.0005
R4347 Vss.n393 Vss.n391 9.0005
R4348 Vss.n391 Vss.n269 9.0005
R4349 Vss.n1404 Vss.n274 9.0005
R4350 Vss.n1404 Vss.n1403 9.0005
R4351 Vss.n383 Vss.n377 9.0005
R4352 Vss.n377 Vss.n376 9.0005
R4353 Vss.n1288 Vss.n1287 9.0005
R4354 Vss.n371 Vss.n318 9.0005
R4355 Vss.n1306 Vss.n1305 9.0005
R4356 Vss.n1296 Vss.n1295 9.0005
R4357 Vss.n354 Vss.n285 9.0005
R4358 Vss.n1392 Vss.n285 9.0005
R4359 Vss.n1222 Vss.n352 9.0005
R4360 Vss.n1222 Vss.n304 9.0005
R4361 Vss.n1276 Vss.n1275 9.0005
R4362 Vss.n945 Vss.n944 9.0005
R4363 Vss.n943 Vss.n942 9.0005
R4364 Vss.n939 Vss.n329 9.0005
R4365 Vss.n938 Vss.n937 9.0005
R4366 Vss.n804 Vss.n803 9.0005
R4367 Vss.n790 Vss.n520 9.0005
R4368 Vss.n1043 Vss.n1042 9.0005
R4369 Vss.n800 Vss.n799 9.0005
R4370 Vss.n793 Vss.n792 9.0005
R4371 Vss.n432 Vss.n431 9.0005
R4372 Vss.n1168 Vss.n1167 9.0005
R4373 Vss.n1181 Vss.n427 9.0005
R4374 Vss.n1192 Vss.n1191 9.0005
R4375 Vss.n1172 Vss.n420 9.0005
R4376 Vss.n1180 Vss.n1178 9.0005
R4377 Vss.n924 Vss.n923 9.0005
R4378 Vss.n1219 Vss.n1218 9.0005
R4379 Vss.n1208 Vss.n1207 9.0005
R4380 Vss.n928 Vss.n927 9.0005
R4381 Vss.n882 Vss.n881 9.0005
R4382 Vss.n888 Vss.n883 9.0005
R4383 Vss.n828 Vss.n827 9.0005
R4384 Vss.n834 Vss.n833 9.0005
R4385 Vss.n836 Vss.n815 9.0005
R4386 Vss.n824 Vss.n823 9.0005
R4387 Vss.n819 Vss.n818 9.0005
R4388 Vss.n622 Vss.n621 9.0005
R4389 Vss.n662 Vss.n661 9.0005
R4390 Vss.n660 Vss.n618 9.0005
R4391 Vss.n624 Vss.n623 9.0005
R4392 Vss.n648 Vss.n647 9.0005
R4393 Vss.n651 Vss.n650 9.0005
R4394 Vss.n629 Vss.n628 9.0005
R4395 Vss.n635 Vss.n634 9.0005
R4396 Vss.n702 Vss.n694 9.0005
R4397 Vss.n5 Vss.n4 9.0005
R4398 Vss.n1915 Vss.n1914 9.0005
R4399 Vss.n723 Vss.n708 9.0005
R4400 Vss.n722 Vss.n720 9.0005
R4401 Vss.n718 Vss.n717 9.0005
R4402 Vss.n713 Vss.n712 9.0005
R4403 Vss.n735 Vss.n734 9.0005
R4404 Vss.n701 Vss.n691 9.0005
R4405 Vss.n737 Vss.n736 9.0005
R4406 Vss.n1855 Vss.t543 8.70131
R4407 Vss.n1904 Vss.t418 8.70131
R4408 Vss.n1162 Vss.n439 8.27654
R4409 Vss.n1592 Vss.n157 8.08508
R4410 Vss.n200 Vss.n147 8.05717
R4411 Vss.n1847 Vss.n1846 7.7564
R4412 Vss.n66 Vss.n43 7.59387
R4413 Vss.n1464 Vss.n1463 7.29099
R4414 Vss.n1917 Vss.n1916 7.12485
R4415 Vss.n892 Vss.n577 6.9012
R4416 Vss.n1210 Vss.n1203 6.9012
R4417 Vss.n1723 Vss.n141 6.9012
R4418 Vss.n1668 Vss.n1663 6.9012
R4419 Vss.n1434 Vss.n1433 6.9012
R4420 Vss.n301 Vss.n298 6.9012
R4421 Vss.n1343 Vss.n1342 6.9012
R4422 Vss.n1226 Vss.n1223 6.9012
R4423 Vss.n1408 Vss.n1407 6.9012
R4424 Vss.n397 Vss.n386 6.9012
R4425 Vss.n1326 Vss.n313 6.9012
R4426 Vss.n1064 Vss.n1063 6.9012
R4427 Vss.n1683 Vss.n1682 6.9012
R4428 Vss.n511 Vss.n510 6.9012
R4429 Vss.n1029 Vss.n1028 6.9012
R4430 Vss.n1361 Vss.n1358 6.9012
R4431 Vss.n1813 Vss.n1812 6.9012
R4432 Vss.n438 Vss.n437 6.9012
R4433 Vss.n664 Vss.n615 6.9012
R4434 Vss.n705 Vss.n704 6.9012
R4435 Vss.n1876 Vss.n1875 6.90005
R4436 Vss.n1834 Vss.n60 6.64904
R4437 Vss.n1860 Vss.n53 6.5795
R4438 Vss.n55 Vss.n54 6.5795
R4439 Vss.n2 Vss.n1 6.5795
R4440 Vss.n1903 Vss.n1898 6.5795
R4441 Vss.n839 Vss.n838 6.46296
R4442 Vss.n889 Vss.n580 6.46296
R4443 Vss.n1182 Vss.n1181 6.46296
R4444 Vss.n518 Vss.n517 6.46296
R4445 Vss.n329 Vss.n328 6.46296
R4446 Vss.n1583 Vss.n1582 6.46296
R4447 Vss.n1590 Vss.n1589 6.46296
R4448 Vss.n1716 Vss.n1715 6.46296
R4449 Vss.n1800 Vss.n1799 6.46296
R4450 Vss.n1440 Vss.n253 6.46296
R4451 Vss.n1354 Vss.n1352 6.46296
R4452 Vss.n305 Vss.n304 6.46296
R4453 Vss.n1207 Vss.n1206 6.46296
R4454 Vss.n1305 Vss.n1304 6.46296
R4455 Vss.n376 Vss.n375 6.46296
R4456 Vss.n406 Vss.n405 6.46296
R4457 Vss.n384 Vss.n370 6.46296
R4458 Vss.n415 Vss.n414 6.46296
R4459 Vss.n1334 Vss.n1333 6.46296
R4460 Vss.n1403 Vss.n1402 6.46296
R4461 Vss.n1320 Vss.n1315 6.46296
R4462 Vss.n1310 Vss.n1308 6.46296
R4463 Vss.n1265 Vss.n334 6.46296
R4464 Vss.n1275 Vss.n1274 6.46296
R4465 Vss.n348 Vss.n347 6.46296
R4466 Vss.n1258 Vss.n336 6.46296
R4467 Vss.n1082 Vss.n1081 6.46296
R4468 Vss.n1089 Vss.n1088 6.46296
R4469 Vss.n1068 Vss.n1058 6.46296
R4470 Vss.n139 Vss.n138 6.46296
R4471 Vss.n1673 Vss.n1671 6.46296
R4472 Vss.n1654 Vss.n1653 6.46296
R4473 Vss.n1704 Vss.n1703 6.46296
R4474 Vss.n1711 Vss.n1710 6.46296
R4475 Vss.n499 Vss.n498 6.46296
R4476 Vss.n479 Vss.n477 6.46296
R4477 Vss.n464 Vss.n463 6.46296
R4478 Vss.n525 Vss.n524 6.46296
R4479 Vss.n176 Vss.n175 6.46296
R4480 Vss.n1369 Vss.n1368 6.46296
R4481 Vss.n183 Vss.n179 6.46296
R4482 Vss.n1456 Vss.n1455 6.46296
R4483 Vss.n1808 Vss.n1807 6.46296
R4484 Vss.n1429 Vss.n1428 6.46296
R4485 Vss.n1461 Vss.n1460 6.46296
R4486 Vss.n1575 Vss.n1574 6.46296
R4487 Vss.n1524 Vss.n1523 6.46296
R4488 Vss.n198 Vss.n197 6.46296
R4489 Vss.n1240 Vss.n1239 6.46296
R4490 Vss.n929 Vss.n928 6.46296
R4491 Vss.n1191 Vss.n1190 6.46296
R4492 Vss.n799 Vss.n798 6.46296
R4493 Vss.n1164 Vss.n432 6.46296
R4494 Vss.n823 Vss.n822 6.46296
R4495 Vss.n621 Vss.n620 6.46296
R4496 Vss.n661 Vss.n617 6.46296
R4497 Vss.n628 Vss.n627 6.46296
R4498 Vss.n731 Vss.n694 6.46296
R4499 Vss.n717 Vss.n716 6.46296
R4500 Vss.n724 Vss.n723 6.46296
R4501 Vss.n691 Vss.n690 6.4618
R4502 Vss.n582 Vss.n581 6.4618
R4503 Vss.n919 Vss.n918 6.4618
R4504 Vss.n418 Vss.n417 6.4618
R4505 Vss.n1688 Vss.n1686 6.4618
R4506 Vss.n1820 Vss.n1819 6.4618
R4507 Vss.n1825 Vss.n1824 6.4618
R4508 Vss.n1388 Vss.n1387 6.4618
R4509 Vss.n294 Vss.n293 6.4618
R4510 Vss.n943 Vss.n559 6.4618
R4511 Vss.n1393 Vss.n1392 6.4618
R4512 Vss.n1295 Vss.n1294 6.4618
R4513 Vss.n1218 Vss.n1217 6.4618
R4514 Vss.n1420 Vss.n1419 6.4618
R4515 Vss.n1412 Vss.n269 6.4618
R4516 Vss.n322 Vss.n321 6.4618
R4517 Vss.n395 Vss.n394 6.4618
R4518 Vss.n966 Vss.n964 6.4618
R4519 Vss.n1252 Vss.n1251 6.4618
R4520 Vss.n153 Vss.n152 6.4618
R4521 Vss.n1086 Vss.n1085 6.4618
R4522 Vss.n1561 Vss.n1560 6.4618
R4523 Vss.n1792 Vss.n1791 6.4618
R4524 Vss.n1699 Vss.n1639 6.4618
R4525 Vss.n1647 Vss.n1641 6.4618
R4526 Vss.n461 Vss.n460 6.4618
R4527 Vss.n489 Vss.n487 6.4618
R4528 Vss.n996 Vss.n995 6.4618
R4529 Vss.n207 Vss.n206 6.4618
R4530 Vss.n212 Vss.n211 6.4618
R4531 Vss.n1567 Vss.n1566 6.4618
R4532 Vss.n1541 Vss.n177 6.4618
R4533 Vss.n1376 Vss.n1375 6.4618
R4534 Vss.n1536 Vss.n1535 6.4618
R4535 Vss.n1731 Vss.n1730 6.4618
R4536 Vss.n805 Vss.n804 6.4618
R4537 Vss.n829 Vss.n828 6.4618
R4538 Vss.n625 Vss.n624 6.4618
R4539 Vss.n6 Vss.n5 6.4618
R4540 Vss.t415 Vss.n1900 6.36556
R4541 Vss.n1846 Vss.n1845 6.33584
R4542 Vss.n1843 Vss.n66 6.32806
R4543 Vss.n1839 Vss.n1837 6.23383
R4544 SARlogic_0.dffrs_12.nand3_1.A Vss.n1174 5.7755
R4545 SARlogic_0.dffrs_12.nand3_8.A Vss.n1195 5.7755
R4546 SARlogic_0.dffrs_13.nand3_8.A Vss.n1636 5.7755
R4547 SARlogic_0.dffrs_12.nand3_6.B Vss.n1175 5.47979
R4548 Vss.n893 Vss.n892 5.47239
R4549 Vss.n1211 Vss.n1210 5.47239
R4550 Vss.n1723 Vss.n1722 5.47239
R4551 Vss.n1668 Vss.n1667 5.47239
R4552 Vss.n1433 Vss.n1432 5.47239
R4553 Vss.n301 Vss.n300 5.47239
R4554 Vss.n1342 Vss.n1341 5.47239
R4555 Vss.n1226 Vss.n1225 5.47239
R4556 Vss.n1407 Vss.n1406 5.47239
R4557 Vss.n398 Vss.n386 5.47239
R4558 Vss.n1327 Vss.n1326 5.47239
R4559 Vss.n1064 Vss.n1059 5.47239
R4560 Vss.n1682 Vss.n1681 5.47239
R4561 Vss.n510 Vss.n506 5.47239
R4562 Vss.n1030 Vss.n1029 5.47239
R4563 Vss.n1361 Vss.n1360 5.47239
R4564 Vss.n1812 Vss.n1811 5.47239
R4565 Vss.n437 Vss.n436 5.47239
R4566 Vss.n665 Vss.n664 5.47239
R4567 Vss.n1875 Vss.n39 5.47239
R4568 Vss.n704 Vss.n700 5.47239
R4569 Vss.n1766 Vss.n1765 5.18044
R4570 Vss.n738 Vss.n737 5.03414
R4571 Vss.n820 Vss.n819 5.03414
R4572 Vss.n815 Vss.n814 5.03414
R4573 Vss.n881 Vss.n880 5.03414
R4574 Vss.n888 Vss.n887 5.03414
R4575 Vss.n1180 Vss.n1179 5.03414
R4576 Vss.n794 Vss.n793 5.03414
R4577 Vss.n1044 Vss.n1043 5.03414
R4578 Vss.n923 Vss.n922 5.03414
R4579 Vss.n1198 Vss.n1197 5.03414
R4580 Vss.n937 Vss.n936 5.03414
R4581 Vss.n1278 Vss.n1277 5.03414
R4582 Vss.n1580 Vss.n1579 5.03414
R4583 Vss.n1588 Vss.n1587 5.03414
R4584 Vss.n1714 Vss.n1713 5.03414
R4585 Vss.n1798 Vss.n1797 5.03414
R4586 Vss.n1689 Vss.n1638 5.03414
R4587 Vss.n73 Vss.n72 5.03414
R4588 Vss.n1823 Vss.n1822 5.03414
R4589 Vss.n1443 Vss.n1442 5.03414
R4590 Vss.n288 Vss.n287 5.03414
R4591 Vss.n1381 Vss.n1380 5.03414
R4592 Vss.n1357 Vss.n1356 5.03414
R4593 Vss.n946 Vss.n945 5.03414
R4594 Vss.n1391 Vss.n1390 5.03414
R4595 Vss.n1292 Vss.n1291 5.03414
R4596 Vss.n1350 Vss.n1349 5.03414
R4597 Vss.n355 Vss.n354 5.03414
R4598 Vss.n1204 Vss.n352 5.03414
R4599 Vss.n1300 Vss.n1299 5.03414
R4600 Vss.n372 Vss.n371 5.03414
R4601 Vss.n265 Vss.n264 5.03414
R4602 Vss.n1413 Vss.n263 5.03414
R4603 Vss.n393 Vss.n392 5.03414
R4604 Vss.n388 Vss.n274 5.03414
R4605 Vss.n1287 Vss.n1286 5.03414
R4606 Vss.n383 Vss.n382 5.03414
R4607 Vss.n367 Vss.n366 5.03414
R4608 Vss.n1330 Vss.n260 5.03414
R4609 Vss.n276 Vss.n275 5.03414
R4610 Vss.n1313 Vss.n1312 5.03414
R4611 Vss.n1319 Vss.n1318 5.03414
R4612 Vss.n1270 Vss.n1269 5.03414
R4613 Vss.n1264 Vss.n1263 5.03414
R4614 Vss.n969 Vss.n968 5.03414
R4615 Vss.n342 Vss.n341 5.03414
R4616 Vss.n1243 Vss.n1242 5.03414
R4617 Vss.n1257 Vss.n337 5.03414
R4618 Vss.n1237 Vss.n1236 5.03414
R4619 Vss.n1599 Vss.n1598 5.03414
R4620 Vss.n1113 Vss.n1112 5.03414
R4621 Vss.n1097 Vss.n1096 5.03414
R4622 Vss.n1070 Vss.n1069 5.03414
R4623 Vss.n1108 Vss.n1107 5.03414
R4624 Vss.n1557 Vss.n1556 5.03414
R4625 Vss.n135 Vss.n134 5.03414
R4626 Vss.n95 Vss.n94 5.03414
R4627 Vss.n1674 Vss.n1633 5.03414
R4628 Vss.n1624 Vss.n1623 5.03414
R4629 Vss.n1658 Vss.n1657 5.03414
R4630 Vss.n1631 Vss.n1630 5.03414
R4631 Vss.n1698 Vss.n1697 5.03414
R4632 Vss.n1646 Vss.n1645 5.03414
R4633 Vss.n1127 Vss.n1126 5.03414
R4634 Vss.n1131 Vss.n1130 5.03414
R4635 Vss.n497 Vss.n496 5.03414
R4636 Vss.n482 Vss.n481 5.03414
R4637 Vss.n492 Vss.n491 5.03414
R4638 Vss.n992 Vss.n991 5.03414
R4639 Vss.n1038 Vss.n1037 5.03414
R4640 Vss.n203 Vss.n202 5.03414
R4641 Vss.n1514 Vss.n1513 5.03414
R4642 Vss.n1565 Vss.n1564 5.03414
R4643 Vss.n1544 Vss.n1543 5.03414
R4644 Vss.n1552 Vss.n1551 5.03414
R4645 Vss.n1373 Vss.n1372 5.03414
R4646 Vss.n189 Vss.n188 5.03414
R4647 Vss.n1365 Vss.n1364 5.03414
R4648 Vss.n1451 Vss.n1450 5.03414
R4649 Vss.n182 Vss.n181 5.03414
R4650 Vss.n80 Vss.n79 5.03414
R4651 Vss.n1424 Vss.n78 5.03414
R4652 Vss.n1459 Vss.n1458 5.03414
R4653 Vss.n164 Vss.n163 5.03414
R4654 Vss.n1520 Vss.n1519 5.03414
R4655 Vss.n1527 Vss.n1526 5.03414
R4656 Vss.n128 Vss.n127 5.03414
R4657 Vss.n421 Vss.n420 5.03414
R4658 Vss.n790 Vss.n789 5.03414
R4659 Vss.n1167 Vss.n1166 5.03414
R4660 Vss.n833 Vss.n832 5.03414
R4661 Vss.n636 Vss.n635 5.03414
R4662 Vss.n652 Vss.n651 5.03414
R4663 Vss.n660 Vss.n659 5.03414
R4664 Vss.n647 Vss.n646 5.03414
R4665 Vss.n1914 Vss.n1913 5.03414
R4666 Vss.n734 Vss.n733 5.03414
R4667 Vss.n714 Vss.n713 5.03414
R4668 Vss.n722 Vss.n721 5.03414
R4669 Vss.n1734 Vss.t85 4.84702
R4670 Vss.n1611 Vss.t248 4.84702
R4671 Vss.n868 Vss.t74 4.84702
R4672 Vss.n870 Vss.t12 4.84702
R4673 Vss.n548 Vss.t633 4.84702
R4674 Vss.n546 Vss.t452 4.84702
R4675 Vss.n1136 Vss.t83 4.84702
R4676 Vss.n1135 Vss.t219 4.84702
R4677 Vss.n743 Vss.t646 4.84702
R4678 Vss.n741 Vss.t216 4.84702
R4679 Vss.n673 Vss.t87 4.84702
R4680 Vss.n672 Vss.t182 4.84702
R4681 Vss.n1853 Vss.n56 4.79462
R4682 Vss.n738 Vss.t600 4.7885
R4683 Vss.n589 Vss.t561 4.7885
R4684 Vss.n671 Vss.t258 4.7885
R4685 Vss.n820 Vss.t498 4.7885
R4686 Vss.n814 Vss.t153 4.7885
R4687 Vss.n880 Vss.t151 4.7885
R4688 Vss.n887 Vss.t170 4.7885
R4689 Vss.n893 Vss.t178 4.7885
R4690 Vss.n1179 Vss.t631 4.7885
R4691 Vss.n794 Vss.t468 4.7885
R4692 Vss.n1044 Vss.t372 4.7885
R4693 Vss.n922 Vss.t616 4.7885
R4694 Vss.n1198 Vss.t679 4.7885
R4695 Vss.n1211 Vss.t256 4.7885
R4696 Vss.n936 Vss.t681 4.7885
R4697 Vss.n1278 Vss.t174 4.7885
R4698 Vss.n1580 Vss.t358 4.7885
R4699 Vss.n1587 Vss.t587 4.7885
R4700 Vss.n1722 Vss.t231 4.7885
R4701 Vss.n1713 Vss.t285 4.7885
R4702 Vss.n1797 Vss.t500 4.7885
R4703 Vss.n1667 Vss.t133 4.7885
R4704 Vss.n1689 Vss.t44 4.7885
R4705 Vss.n73 Vss.t410 4.7885
R4706 Vss.n1822 Vss.t659 4.7885
R4707 Vss.n1432 Vss.t365 4.7885
R4708 Vss.n1442 Vss.t494 4.7885
R4709 Vss.n300 Vss.t59 4.7885
R4710 Vss.n288 Vss.t442 4.7885
R4711 Vss.n1381 Vss.t486 4.7885
R4712 Vss.n1356 Vss.t649 4.7885
R4713 Vss.n1341 Vss.t240 4.7885
R4714 Vss.n946 Vss.t191 4.7885
R4715 Vss.n1225 Vss.t428 4.7885
R4716 Vss.n1390 Vss.t246 4.7885
R4717 Vss.n1292 Vss.t462 4.7885
R4718 Vss.n1349 Vss.t225 4.7885
R4719 Vss.n355 Vss.t184 4.7885
R4720 Vss.n1204 Vss.t40 4.7885
R4721 Vss.n1300 Vss.t370 4.7885
R4722 Vss.n372 Vss.t492 4.7885
R4723 Vss.n1406 Vss.t158 4.7885
R4724 Vss.n265 Vss.t403 4.7885
R4725 Vss.n1413 Vss.t352 4.7885
R4726 Vss.n392 Vss.t531 4.7885
R4727 Vss.n388 Vss.t533 4.7885
R4728 Vss.n398 Vss.t355 4.7885
R4729 Vss.n1286 Vss.t488 4.7885
R4730 Vss.n382 Vss.t300 4.7885
R4731 Vss.n366 Vss.t496 4.7885
R4732 Vss.n1327 Vss.t656 4.7885
R4733 Vss.n1330 Vss.t298 4.7885
R4734 Vss.n276 Vss.t64 4.7885
R4735 Vss.n1312 Vss.t513 4.7885
R4736 Vss.n1318 Vss.t155 4.7885
R4737 Vss.n1270 Vss.t120 4.7885
R4738 Vss.n1263 Vss.t76 4.7885
R4739 Vss.n969 Vss.t122 4.7885
R4740 Vss.n342 Vss.t593 4.7885
R4741 Vss.n1243 Vss.t221 4.7885
R4742 Vss.n337 Vss.t400 4.7885
R4743 Vss.n1237 Vss.t289 4.7885
R4744 Vss.n1598 Vss.t423 4.7885
R4745 Vss.n1113 Vss.t440 4.7885
R4746 Vss.n1097 Vss.t480 4.7885
R4747 Vss.n1059 Vss.t34 4.7885
R4748 Vss.n1070 Vss.t672 4.7885
R4749 Vss.n1107 Vss.t527 4.7885
R4750 Vss.n1608 Vss.t566 4.7885
R4751 Vss.n1557 Vss.t274 4.7885
R4752 Vss.n135 Vss.t296 4.7885
R4753 Vss.n110 Vss.t131 4.7885
R4754 Vss.n109 Vss.t90 4.7885
R4755 Vss.n1768 Vss.t97 4.7885
R4756 Vss.n48 Vss.t349 4.7885
R4757 Vss.n50 Vss.t287 4.7885
R4758 Vss.n95 Vss.t484 4.7885
R4759 Vss.n1681 Vss.t596 4.7885
R4760 Vss.n1674 Vss.t15 4.7885
R4761 Vss.n1624 Vss.t574 4.7885
R4762 Vss.n1657 Vss.t458 4.7885
R4763 Vss.n1630 Vss.t602 4.7885
R4764 Vss.n1697 Vss.t142 4.7885
R4765 Vss.n1780 Vss.t116 4.7885
R4766 Vss.n1755 Vss.t390 4.7885
R4767 Vss.n1750 Vss.t281 4.7885
R4768 Vss.n1784 Vss.t283 4.7885
R4769 Vss.n1773 Vss.t554 4.7885
R4770 Vss.n1645 Vss.t333 4.7885
R4771 Vss.n1502 Vss.t559 4.7885
R4772 Vss.n1487 Vss.t447 4.7885
R4773 Vss.n1482 Vss.t545 4.7885
R4774 Vss.n1506 Vss.t547 4.7885
R4775 Vss.n542 Vss.t614 4.7885
R4776 Vss.n541 Vss.t580 4.7885
R4777 Vss.n1126 Vss.t362 4.7885
R4778 Vss.n506 Vss.t612 4.7885
R4779 Vss.n1131 Vss.t243 4.7885
R4780 Vss.n496 Vss.t381 4.7885
R4781 Vss.n481 Vss.t466 4.7885
R4782 Vss.n491 Vss.t518 4.7885
R4783 Vss.n1009 Vss.t621 4.7885
R4784 Vss.n991 Vss.t252 4.7885
R4785 Vss.n1037 Vss.t393 4.7885
R4786 Vss.n1030 Vss.t46 4.7885
R4787 Vss.n568 Vss.t21 4.7885
R4788 Vss.n569 Vss.t48 4.7885
R4789 Vss.n906 Vss.t628 4.7885
R4790 Vss.n564 Vss.t438 4.7885
R4791 Vss.n859 Vss.t144 4.7885
R4792 Vss.n1159 Vss.t454 4.7885
R4793 Vss.n444 Vss.t456 4.7885
R4794 Vss.n449 Vss.t663 4.7885
R4795 Vss.n1017 Vss.t160 4.7885
R4796 Vss.n553 Vss.t653 4.7885
R4797 Vss.n554 Vss.t109 4.7885
R4798 Vss.n555 Vss.t107 4.7885
R4799 Vss.n980 Vss.t552 4.7885
R4800 Vss.n1145 Vss.t168 4.7885
R4801 Vss.n220 Vss.t62 4.7885
R4802 Vss.n219 Vss.t38 4.7885
R4803 Vss.n1496 Vss.t36 4.7885
R4804 Vss.n203 Vss.t624 4.7885
R4805 Vss.n1513 Vss.t291 4.7885
R4806 Vss.n1360 Vss.t636 4.7885
R4807 Vss.n1564 Vss.t125 4.7885
R4808 Vss.n1544 Vss.t507 4.7885
R4809 Vss.n1551 Vss.t235 4.7885
R4810 Vss.n1373 Vss.t129 4.7885
R4811 Vss.n189 Vss.t525 4.7885
R4812 Vss.n1365 Vss.t52 4.7885
R4813 Vss.n1451 Vss.t478 4.7885
R4814 Vss.n181 Vss.t398 4.7885
R4815 Vss.n1811 Vss.t19 4.7885
R4816 Vss.n80 Vss.t103 4.7885
R4817 Vss.n1424 Vss.t375 4.7885
R4818 Vss.n1458 Vss.t396 4.7885
R4819 Vss.n164 Vss.t347 4.7885
R4820 Vss.n1520 Vss.t162 4.7885
R4821 Vss.n1527 Vss.t80 4.7885
R4822 Vss.n127 Vss.t589 4.7885
R4823 Vss.n421 Vss.t269 4.7885
R4824 Vss.n436 Vss.t425 4.7885
R4825 Vss.n789 Vss.t523 4.7885
R4826 Vss.n1166 Vss.t618 4.7885
R4827 Vss.n832 Vss.t490 4.7885
R4828 Vss.n598 Vss.t585 4.7885
R4829 Vss.n780 Vss.t180 4.7885
R4830 Vss.n778 Vss.t445 4.7885
R4831 Vss.n1880 Vss.t667 4.7885
R4832 Vss.n32 Vss.t379 4.7885
R4833 Vss.n33 Vss.t195 4.7885
R4834 Vss.n34 Vss.t197 4.7885
R4835 Vss.n752 Vss.t610 4.7885
R4836 Vss.n21 Vss.t271 4.7885
R4837 Vss.n20 Vss.t341 4.7885
R4838 Vss.n1893 Vss.t345 4.7885
R4839 Vss.n636 Vss.t505 4.7885
R4840 Vss.n652 Vss.t591 4.7885
R4841 Vss.n659 Vss.t405 4.7885
R4842 Vss.n665 Vss.t343 4.7885
R4843 Vss.n39 Vss.t583 4.7885
R4844 Vss.n646 Vss.t502 4.7885
R4845 Vss.n1913 Vss.t510 4.7885
R4846 Vss.n733 Vss.t166 4.7885
R4847 Vss.n700 Vss.t641 4.7885
R4848 Vss.n714 Vss.t607 4.7885
R4849 Vss.n721 Vss.t521 4.7885
R4850 Vss.n769 Vss.t578 4.7885
R4851 Vss.n593 Vss.t138 4.7885
R4852 Vss.n855 Vss.t136 4.7885
R4853 Vss.n892 Vss.n891 4.28213
R4854 Vss.n408 Vss.n386 4.28213
R4855 Vss.n1065 Vss.n1064 4.28213
R4856 Vss.n510 Vss.n509 4.28213
R4857 Vss.n1029 Vss.n522 4.28213
R4858 Vss.n1682 Vss.n1632 4.28213
R4859 Vss.n1669 Vss.n1668 4.28213
R4860 Vss.n1724 Vss.n1723 4.28213
R4861 Vss.n1362 Vss.n1361 4.28213
R4862 Vss.n1812 Vss.n1810 4.28213
R4863 Vss.n1433 Vss.n1431 4.28213
R4864 Vss.n302 Vss.n301 4.28213
R4865 Vss.n1342 Vss.n303 4.28213
R4866 Vss.n1326 Vss.n1325 4.28213
R4867 Vss.n1407 Vss.n1405 4.28213
R4868 Vss.n1227 Vss.n1226 4.28213
R4869 Vss.n437 Vss.n419 4.28213
R4870 Vss.n1210 Vss.n1209 4.28213
R4871 Vss.n664 Vss.n663 4.28213
R4872 Vss.n1875 Vss.n1874 4.28213
R4873 Vss.n704 Vss.n703 4.28213
R4874 Vss.n1850 Vss.n1849 3.8722
R4875 Vss.n1832 Vss.n66 3.52248
R4876 Vss.n1846 Vss.n58 3.51469
R4877 Vss.n1761 Vss.n1760 3.51467
R4878 Vss.n1013 Vss.n1012 3.51467
R4879 Vss.n910 Vss.n909 3.51467
R4880 Vss.n1493 Vss.n1492 3.51467
R4881 Vss.n1890 Vss.n1889 3.51467
R4882 Vss.n775 Vss.n774 3.51467
R4883 Vss.n1868 Vss.t337 3.46717
R4884 Vss.n61 Vss.t433 3.46717
R4885 Vss.n1869 Vss.t338 2.9111
R4886 Vss.n62 Vss.t434 2.9111
R4887 Vss.n1120 Vss.n1052 2.83255
R4888 Vss.n1602 Vss.n150 2.45741
R4889 Vss.n1603 Vss.n1602 2.21573
R4890 Vss.n1176 SARlogic_0.dffrs_12.nand3_6.B 2.17818
R4891 Vss.n1678 Vss.n98 2.06007
R4892 Vss.n1761 Vss.n111 2.06002
R4893 Vss.n1012 Vss.n540 2.06002
R4894 Vss.n909 Vss.n567 2.06002
R4895 Vss.n1493 Vss.n221 2.06002
R4896 Vss.n775 Vss.n599 2.06002
R4897 Vss.n1890 Vss.n27 2.06002
R4898 Vss.n1836 Vss.t3 2.048
R4899 Vss.n1836 Vss.t387 2.048
R4900 Vss.n53 Vss.t449 2.03874
R4901 Vss.n53 Vss.t539 2.03874
R4902 Vss.n54 Vss.t541 2.03874
R4903 Vss.n54 Vss.t537 2.03874
R4904 Vss.n1 Vss.t643 2.03874
R4905 Vss.n1 Vss.t416 2.03874
R4906 Vss.n1898 Vss.t420 2.03874
R4907 Vss.n1898 Vss.t414 2.03874
R4908 Vss.n1301 Vss.n308 2.02164
R4909 Vss.n379 Vss.n325 2.02164
R4910 Vss.n1281 Vss.n327 2.02164
R4911 Vss.n248 Vss.n194 2.02164
R4912 Vss.n1530 Vss.n196 2.02164
R4913 Vss.n1247 Vss.n1246 2.02164
R4914 Vss.n975 Vss.n309 2.02164
R4915 Vss.n1438 Vss.n1437 2.02164
R4916 Vss.n1803 Vss.n1802 2.02164
R4917 Vss.n932 Vss.n931 2.02164
R4918 Vss.n755 Vss.n754 1.92616
R4919 Vss.n682 Vss.n35 1.90702
R4920 Vss.n146 Vss.n145 1.90702
R4921 Vss.n1613 Vss.n112 1.90702
R4922 Vss.n1757 Vss.n115 1.90702
R4923 Vss.n1772 Vss.n104 1.90702
R4924 Vss.n1781 Vss.n105 1.90702
R4925 Vss.n1758 Vss.n114 1.90702
R4926 Vss.n1503 Vss.n216 1.90702
R4927 Vss.n1489 Vss.n225 1.90702
R4928 Vss.n876 Vss.n563 1.90702
R4929 Vss.n911 Vss.n565 1.90702
R4930 Vss.n866 Vss.n865 1.90702
R4931 Vss.n864 Vss.n863 1.90702
R4932 Vss.n450 Vss.n445 1.90702
R4933 Vss.n1155 Vss.n451 1.90702
R4934 Vss.n1015 Vss.n1014 1.90702
R4935 Vss.n988 Vss.n987 1.90702
R4936 Vss.n986 Vss.n552 1.90702
R4937 Vss.n981 Vss.n556 1.90702
R4938 Vss.n458 Vss.n457 1.90702
R4939 Vss.n1141 Vss.n222 1.90702
R4940 Vss.n1490 Vss.n224 1.90702
R4941 Vss.n1881 Vss.n36 1.90702
R4942 Vss.n1886 Vss.n31 1.90702
R4943 Vss.n748 Vss.n28 1.90702
R4944 Vss.n1887 Vss.n30 1.90702
R4945 Vss.n678 Vss.n600 1.90702
R4946 Vss.n772 Vss.n602 1.90702
R4947 Vss.n771 Vss.n603 1.90702
R4948 Vss.n852 Vss.n851 1.90702
R4949 Vss.n1841 Vss.n1840 1.73383
R4950 Vss.n1839 Vss.n1838 1.73383
R4951 Vss.n1868 Vss.n44 1.70279
R4952 Vss.n61 Vss.n44 1.62925
R4953 Vss.n1829 Vss.n68 1.62713
R4954 Vss.n1766 adc_PISO_0.2inmux_0.Bit 1.54251
R4955 Vss.n1176 SARlogic_0.dffrs_12.nand3_1.A 1.34729
R4956 Vss.n919 Vss.n532 1.3005
R4957 Vss.n922 Vss.n921 1.3005
R4958 Vss.n921 Vss.n920 1.3005
R4959 Vss.n559 Vss.n558 1.3005
R4960 Vss.n947 Vss.n946 1.3005
R4961 Vss.n948 Vss.n947 1.3005
R4962 Vss.n305 Vss.n282 1.3005
R4963 Vss.n1349 Vss.n1348 1.3005
R4964 Vss.n1348 Vss.n1347 1.3005
R4965 Vss.n1294 Vss.n283 1.3005
R4966 Vss.n1293 Vss.n1292 1.3005
R4967 Vss.n1293 Vss.n306 1.3005
R4968 Vss.n1394 Vss.n1393 1.3005
R4969 Vss.n1390 Vss.n284 1.3005
R4970 Vss.n307 Vss.n284 1.3005
R4971 Vss.n1206 Vss.n357 1.3005
R4972 Vss.n1205 Vss.n1204 1.3005
R4973 Vss.n1205 Vss.n323 1.3005
R4974 Vss.n1217 Vss.n1216 1.3005
R4975 Vss.n356 Vss.n355 1.3005
R4976 Vss.n356 Vss.n324 1.3005
R4977 Vss.n389 Vss.n388 1.3005
R4978 Vss.n403 Vss.n389 1.3005
R4979 Vss.n405 Vss.n404 1.3005
R4980 Vss.n1286 Vss.n1285 1.3005
R4981 Vss.n1285 Vss.n1284 1.3005
R4982 Vss.n358 Vss.n322 1.3005
R4983 Vss.n382 Vss.n381 1.3005
R4984 Vss.n381 Vss.n380 1.3005
R4985 Vss.n378 Vss.n370 1.3005
R4986 Vss.n1335 Vss.n1334 1.3005
R4987 Vss.n1332 Vss.n1330 1.3005
R4988 Vss.n1332 Vss.n1331 1.3005
R4989 Vss.n1402 Vss.n1401 1.3005
R4990 Vss.n277 Vss.n276 1.3005
R4991 Vss.n1400 Vss.n277 1.3005
R4992 Vss.n1310 Vss.n1309 1.3005
R4993 Vss.n1312 Vss.n1311 1.3005
R4994 Vss.n1311 Vss.n311 1.3005
R4995 Vss.n1315 Vss.n312 1.3005
R4996 Vss.n1318 Vss.n1317 1.3005
R4997 Vss.n1317 Vss.n255 1.3005
R4998 Vss.n313 Vss.n268 1.3005
R4999 Vss.n1328 Vss.n1327 1.3005
R5000 Vss.n1329 Vss.n1328 1.3005
R5001 Vss.n396 Vss.n395 1.3005
R5002 Vss.n392 Vss.n390 1.3005
R5003 Vss.n390 Vss.n270 1.3005
R5004 Vss.n1412 Vss.n1411 1.3005
R5005 Vss.n1414 Vss.n1413 1.3005
R5006 Vss.n1415 Vss.n1414 1.3005
R5007 Vss.n1419 Vss.n1418 1.3005
R5008 Vss.n266 Vss.n265 1.3005
R5009 Vss.n1417 Vss.n266 1.3005
R5010 Vss.n1409 Vss.n1408 1.3005
R5011 Vss.n1406 Vss.n272 1.3005
R5012 Vss.n1398 Vss.n272 1.3005
R5013 Vss.n375 Vss.n374 1.3005
R5014 Vss.n373 Vss.n372 1.3005
R5015 Vss.n373 Vss.n278 1.3005
R5016 Vss.n1304 Vss.n279 1.3005
R5017 Vss.n1303 Vss.n1300 1.3005
R5018 Vss.n1303 Vss.n1302 1.3005
R5019 Vss.n1274 Vss.n1273 1.3005
R5020 Vss.n1271 Vss.n1270 1.3005
R5021 Vss.n1272 Vss.n1271 1.3005
R5022 Vss.n1260 Vss.n334 1.3005
R5023 Vss.n1263 Vss.n1262 1.3005
R5024 Vss.n1262 Vss.n1261 1.3005
R5025 Vss.n1223 Vss.n326 1.3005
R5026 Vss.n1225 Vss.n1224 1.3005
R5027 Vss.n1224 Vss.n281 1.3005
R5028 Vss.n964 Vss.n963 1.3005
R5029 Vss.n970 Vss.n969 1.3005
R5030 Vss.n971 Vss.n970 1.3005
R5031 Vss.n1251 Vss.n1250 1.3005
R5032 Vss.n343 Vss.n342 1.3005
R5033 Vss.n1249 Vss.n343 1.3005
R5034 Vss.n1062 Vss.n1059 1.3005
R5035 Vss.n1062 Vss.n1061 1.3005
R5036 Vss.n1060 Vss.n1058 1.3005
R5037 Vss.n1071 Vss.n1070 1.3005
R5038 Vss.n1072 Vss.n1071 1.3005
R5039 Vss.n1088 Vss.n1087 1.3005
R5040 Vss.n1098 Vss.n1097 1.3005
R5041 Vss.n1099 Vss.n1098 1.3005
R5042 Vss.n1081 Vss.n1079 1.3005
R5043 Vss.n1114 Vss.n1113 1.3005
R5044 Vss.n1115 Vss.n1114 1.3005
R5045 Vss.n1107 Vss.n1106 1.3005
R5046 Vss.n1106 Vss.n1105 1.3005
R5047 Vss.n1102 Vss.n1086 1.3005
R5048 Vss.n138 Vss.n137 1.3005
R5049 Vss.n136 Vss.n135 1.3005
R5050 Vss.n136 Vss.n121 1.3005
R5051 Vss.n1560 Vss.n1559 1.3005
R5052 Vss.n1558 Vss.n1557 1.3005
R5053 Vss.n1558 Vss.n122 1.3005
R5054 Vss.n48 Vss.n47 1.3005
R5055 Vss.n1827 Vss.n47 1.3005
R5056 Vss.n1867 Vss.n1866 1.3005
R5057 Vss.n1864 Vss.n50 1.3005
R5058 Vss.n1864 Vss.n1863 1.3005
R5059 Vss.n1791 Vss.n1790 1.3005
R5060 Vss.n96 Vss.n95 1.3005
R5061 Vss.n1789 Vss.n96 1.3005
R5062 Vss.n1673 Vss.n1672 1.3005
R5063 Vss.n1675 Vss.n1674 1.3005
R5064 Vss.n1676 Vss.n1675 1.3005
R5065 Vss.n1630 Vss.n1629 1.3005
R5066 Vss.n1629 Vss.n1628 1.3005
R5067 Vss.n1705 Vss.n1704 1.3005
R5068 Vss.n1780 Vss.n1779 1.3005
R5069 Vss.n1779 Vss.n1778 1.3005
R5070 Vss.n1645 Vss.n1644 1.3005
R5071 Vss.n1644 Vss.n1643 1.3005
R5072 Vss.n1642 Vss.n1641 1.3005
R5073 Vss.n1710 Vss.n1709 1.3005
R5074 Vss.n1625 Vss.n1624 1.3005
R5075 Vss.n1708 Vss.n1625 1.3005
R5076 Vss.n1654 Vss.n1626 1.3005
R5077 Vss.n1657 Vss.n1656 1.3005
R5078 Vss.n1656 Vss.n1655 1.3005
R5079 Vss.n1684 Vss.n1683 1.3005
R5080 Vss.n1681 Vss.n1680 1.3005
R5081 Vss.n1680 Vss.n1627 1.3005
R5082 Vss.n1755 Vss.n1754 1.3005
R5083 Vss.n1754 Vss.n1753 1.3005
R5084 Vss.n1751 Vss.n1750 1.3005
R5085 Vss.n1752 Vss.n1751 1.3005
R5086 Vss.n1785 Vss.n1784 1.3005
R5087 Vss.n1786 Vss.n1785 1.3005
R5088 Vss.n1772 Vss.n1771 1.3005
R5089 Vss.n1774 Vss.n1773 1.3005
R5090 Vss.n1775 Vss.n1774 1.3005
R5091 Vss.n1739 Vss.n111 1.3005
R5092 Vss.n1742 Vss.n110 1.3005
R5093 Vss.n1748 Vss.n109 1.3005
R5094 Vss.n1749 Vss.n1748 1.3005
R5095 Vss.n1769 Vss.n1768 1.3005
R5096 Vss.n1770 Vss.n1769 1.3005
R5097 Vss.n1735 Vss.n1734 1.3005
R5098 Vss.n1736 Vss.n1735 1.3005
R5099 Vss.n1737 Vss.n114 1.3005
R5100 Vss.n479 Vss.n478 1.3005
R5101 Vss.n481 Vss.n480 1.3005
R5102 Vss.n480 Vss.n471 1.3005
R5103 Vss.n500 Vss.n499 1.3005
R5104 Vss.n496 Vss.n472 1.3005
R5105 Vss.n472 Vss.n465 1.3005
R5106 Vss.n491 Vss.n490 1.3005
R5107 Vss.n490 Vss.n466 1.3005
R5108 Vss.n489 Vss.n488 1.3005
R5109 Vss.n502 Vss.n464 1.3005
R5110 Vss.n1126 Vss.n1125 1.3005
R5111 Vss.n1125 Vss.n1124 1.3005
R5112 Vss.n512 Vss.n511 1.3005
R5113 Vss.n506 Vss.n505 1.3005
R5114 Vss.n505 Vss.n504 1.3005
R5115 Vss.n1003 Vss.n541 1.3005
R5116 Vss.n1004 Vss.n1003 1.3005
R5117 Vss.n1000 Vss.n540 1.3005
R5118 Vss.n1005 Vss.n542 1.3005
R5119 Vss.n1006 Vss.n1005 1.3005
R5120 Vss.n1009 Vss.n1008 1.3005
R5121 Vss.n1008 Vss.n1007 1.3005
R5122 Vss.n1034 Vss.n525 1.3005
R5123 Vss.n1037 Vss.n1036 1.3005
R5124 Vss.n1036 Vss.n1035 1.3005
R5125 Vss.n1031 Vss.n1030 1.3005
R5126 Vss.n1032 Vss.n1031 1.3005
R5127 Vss.n1028 Vss.n1027 1.3005
R5128 Vss.n444 Vss.n433 1.3005
R5129 Vss.n231 Vss.n221 1.3005
R5130 Vss.n230 Vss.n220 1.3005
R5131 Vss.n1480 Vss.n219 1.3005
R5132 Vss.n1481 Vss.n1480 1.3005
R5133 Vss.n1497 Vss.n1496 1.3005
R5134 Vss.n1498 Vss.n1497 1.3005
R5135 Vss.n1499 Vss.n216 1.3005
R5136 Vss.n1502 Vss.n1501 1.3005
R5137 Vss.n1501 Vss.n1500 1.3005
R5138 Vss.n1054 Vss.n153 1.3005
R5139 Vss.n1598 Vss.n1597 1.3005
R5140 Vss.n1597 Vss.n1596 1.3005
R5141 Vss.n206 Vss.n205 1.3005
R5142 Vss.n204 Vss.n203 1.3005
R5143 Vss.n204 Vss.n156 1.3005
R5144 Vss.n238 Vss.n212 1.3005
R5145 Vss.n1513 Vss.n1512 1.3005
R5146 Vss.n1512 Vss.n1511 1.3005
R5147 Vss.n176 Vss.n170 1.3005
R5148 Vss.n1551 Vss.n1550 1.3005
R5149 Vss.n1550 Vss.n1549 1.3005
R5150 Vss.n177 Vss.n171 1.3005
R5151 Vss.n1545 Vss.n1544 1.3005
R5152 Vss.n1546 Vss.n1545 1.3005
R5153 Vss.n1568 Vss.n1567 1.3005
R5154 Vss.n1564 Vss.n172 1.3005
R5155 Vss.n1547 Vss.n172 1.3005
R5156 Vss.n1368 Vss.n1367 1.3005
R5157 Vss.n1366 Vss.n1365 1.3005
R5158 Vss.n1366 Vss.n192 1.3005
R5159 Vss.n1535 Vss.n1534 1.3005
R5160 Vss.n190 Vss.n189 1.3005
R5161 Vss.n1533 Vss.n190 1.3005
R5162 Vss.n1375 Vss.n244 1.3005
R5163 Vss.n1374 Vss.n1373 1.3005
R5164 Vss.n1374 Vss.n193 1.3005
R5165 Vss.n1807 Vss.n1806 1.3005
R5166 Vss.n81 Vss.n80 1.3005
R5167 Vss.n1805 Vss.n81 1.3005
R5168 Vss.n1462 Vss.n1461 1.3005
R5169 Vss.n1458 Vss.n250 1.3005
R5170 Vss.n250 Vss.n249 1.3005
R5171 Vss.n1428 Vss.n1427 1.3005
R5172 Vss.n1425 Vss.n1424 1.3005
R5173 Vss.n1426 Vss.n1425 1.3005
R5174 Vss.n1814 Vss.n1813 1.3005
R5175 Vss.n1811 Vss.n76 1.3005
R5176 Vss.n82 Vss.n76 1.3005
R5177 Vss.n1455 Vss.n1454 1.3005
R5178 Vss.n1452 Vss.n1451 1.3005
R5179 Vss.n1453 Vss.n1452 1.3005
R5180 Vss.n179 Vss.n178 1.3005
R5181 Vss.n181 Vss.n180 1.3005
R5182 Vss.n180 Vss.n85 1.3005
R5183 Vss.n1523 Vss.n1522 1.3005
R5184 Vss.n1521 Vss.n1520 1.3005
R5185 Vss.n1521 Vss.n167 1.3005
R5186 Vss.n1574 Vss.n1573 1.3005
R5187 Vss.n165 Vss.n164 1.3005
R5188 Vss.n1572 Vss.n165 1.3005
R5189 Vss.n1358 Vss.n195 1.3005
R5190 Vss.n1360 Vss.n1359 1.3005
R5191 Vss.n1359 Vss.n169 1.3005
R5192 Vss.n236 Vss.n225 1.3005
R5193 Vss.n1487 Vss.n1486 1.3005
R5194 Vss.n1486 Vss.n1485 1.3005
R5195 Vss.n1483 Vss.n1482 1.3005
R5196 Vss.n1484 Vss.n1483 1.3005
R5197 Vss.n1507 Vss.n1506 1.3005
R5198 Vss.n1508 Vss.n1507 1.3005
R5199 Vss.n1528 Vss.n1527 1.3005
R5200 Vss.n1529 Vss.n1528 1.3005
R5201 Vss.n240 Vss.n197 1.3005
R5202 Vss.n1239 Vss.n345 1.3005
R5203 Vss.n1238 Vss.n1237 1.3005
R5204 Vss.n1238 Vss.n242 1.3005
R5205 Vss.n953 Vss.n556 1.3005
R5206 Vss.n980 Vss.n979 1.3005
R5207 Vss.n979 Vss.n978 1.3005
R5208 Vss.n557 Vss.n460 1.3005
R5209 Vss.n1132 Vss.n1131 1.3005
R5210 Vss.n1133 Vss.n1132 1.3005
R5211 Vss.n1134 Vss.n458 1.3005
R5212 Vss.n1145 Vss.n1144 1.3005
R5213 Vss.n1144 Vss.n1143 1.3005
R5214 Vss.n1142 Vss.n1141 1.3005
R5215 Vss.n1140 Vss.n1135 1.3005
R5216 Vss.n1140 Vss.n1139 1.3005
R5217 Vss.n1137 Vss.n1136 1.3005
R5218 Vss.n1138 Vss.n1137 1.3005
R5219 Vss.n235 Vss.n224 1.3005
R5220 Vss.n974 Vss.n336 1.3005
R5221 Vss.n972 Vss.n337 1.3005
R5222 Vss.n973 Vss.n972 1.3005
R5223 Vss.n347 Vss.n346 1.3005
R5224 Vss.n1244 Vss.n1243 1.3005
R5225 Vss.n1245 Vss.n1244 1.3005
R5226 Vss.n1344 Vss.n1343 1.3005
R5227 Vss.n1341 Vss.n1340 1.3005
R5228 Vss.n1340 Vss.n1339 1.3005
R5229 Vss.n1354 Vss.n1353 1.3005
R5230 Vss.n1356 Vss.n1355 1.3005
R5231 Vss.n1355 Vss.n291 1.3005
R5232 Vss.n293 Vss.n292 1.3005
R5233 Vss.n1382 Vss.n1381 1.3005
R5234 Vss.n1383 Vss.n1382 1.3005
R5235 Vss.n1387 Vss.n1386 1.3005
R5236 Vss.n289 Vss.n288 1.3005
R5237 Vss.n1385 Vss.n289 1.3005
R5238 Vss.n298 Vss.n297 1.3005
R5239 Vss.n300 Vss.n299 1.3005
R5240 Vss.n299 Vss.n243 1.3005
R5241 Vss.n1440 Vss.n1439 1.3005
R5242 Vss.n1442 Vss.n1441 1.3005
R5243 Vss.n1441 Vss.n246 1.3005
R5244 Vss.n1435 Vss.n1434 1.3005
R5245 Vss.n1432 Vss.n258 1.3005
R5246 Vss.n258 Vss.n257 1.3005
R5247 Vss.n1826 Vss.n1825 1.3005
R5248 Vss.n1822 Vss.n69 1.3005
R5249 Vss.n1815 Vss.n69 1.3005
R5250 Vss.n1819 Vss.n1818 1.3005
R5251 Vss.n74 Vss.n73 1.3005
R5252 Vss.n1817 Vss.n74 1.3005
R5253 Vss.n1688 Vss.n1687 1.3005
R5254 Vss.n1690 Vss.n1689 1.3005
R5255 Vss.n1691 Vss.n1690 1.3005
R5256 Vss.n1693 Vss.n1639 1.3005
R5257 Vss.n1697 Vss.n1696 1.3005
R5258 Vss.n1696 Vss.n1695 1.3005
R5259 Vss.n1664 Vss.n1663 1.3005
R5260 Vss.n1667 Vss.n1666 1.3005
R5261 Vss.n1666 Vss.n1665 1.3005
R5262 Vss.n1801 Vss.n1800 1.3005
R5263 Vss.n1797 Vss.n87 1.3005
R5264 Vss.n1618 Vss.n87 1.3005
R5265 Vss.n1717 Vss.n1716 1.3005
R5266 Vss.n1713 Vss.n1619 1.3005
R5267 Vss.n1677 Vss.n1619 1.3005
R5268 Vss.n142 Vss.n141 1.3005
R5269 Vss.n1722 Vss.n1721 1.3005
R5270 Vss.n1721 Vss.n1720 1.3005
R5271 Vss.n1591 Vss.n1590 1.3005
R5272 Vss.n1587 Vss.n158 1.3005
R5273 Vss.n158 Vss.n143 1.3005
R5274 Vss.n1582 Vss.n144 1.3005
R5275 Vss.n1581 Vss.n1580 1.3005
R5276 Vss.n1581 Vss.n123 1.3005
R5277 Vss.n1594 Vss.n145 1.3005
R5278 Vss.n1609 Vss.n1608 1.3005
R5279 Vss.n1610 Vss.n1609 1.3005
R5280 Vss.n1614 Vss.n1613 1.3005
R5281 Vss.n1612 Vss.n1611 1.3005
R5282 Vss.n1612 Vss.n125 1.3005
R5283 Vss.n127 Vss.n126 1.3005
R5284 Vss.n126 Vss.n124 1.3005
R5285 Vss.n1732 Vss.n1731 1.3005
R5286 Vss.n933 Vss.n929 1.3005
R5287 Vss.n936 Vss.n935 1.3005
R5288 Vss.n935 Vss.n934 1.3005
R5289 Vss.n359 Vss.n328 1.3005
R5290 Vss.n1279 Vss.n1278 1.3005
R5291 Vss.n1280 Vss.n1279 1.3005
R5292 Vss.n1203 Vss.n1202 1.3005
R5293 Vss.n1212 Vss.n1211 1.3005
R5294 Vss.n1213 Vss.n1212 1.3005
R5295 Vss.n397 Vss.n363 1.3005
R5296 Vss.n399 Vss.n398 1.3005
R5297 Vss.n400 Vss.n399 1.3005
R5298 Vss.n416 Vss.n415 1.3005
R5299 Vss.n366 Vss.n365 1.3005
R5300 Vss.n365 Vss.n364 1.3005
R5301 Vss.n1190 Vss.n1189 1.3005
R5302 Vss.n422 Vss.n421 1.3005
R5303 Vss.n1188 Vss.n422 1.3005
R5304 Vss.n439 Vss.n438 1.3005
R5305 Vss.n436 Vss.n435 1.3005
R5306 Vss.n435 Vss.n423 1.3005
R5307 Vss.n1186 Vss.n417 1.3005
R5308 Vss.n1199 Vss.n1198 1.3005
R5309 Vss.n1200 Vss.n1199 1.3005
R5310 Vss.n552 Vss.n536 1.3005
R5311 Vss.n959 Vss.n553 1.3005
R5312 Vss.n960 Vss.n959 1.3005
R5313 Vss.n951 Vss.n554 1.3005
R5314 Vss.n951 Vss.n545 1.3005
R5315 Vss.n956 Vss.n555 1.3005
R5316 Vss.n956 Vss.n955 1.3005
R5317 Vss.n997 Vss.n996 1.3005
R5318 Vss.n991 Vss.n990 1.3005
R5319 Vss.n990 Vss.n537 1.3005
R5320 Vss.n1020 Vss.n451 1.3005
R5321 Vss.n1018 Vss.n1017 1.3005
R5322 Vss.n1019 Vss.n1018 1.3005
R5323 Vss.n1016 Vss.n1015 1.3005
R5324 Vss.n546 Vss.n538 1.3005
R5325 Vss.n549 Vss.n538 1.3005
R5326 Vss.n551 Vss.n548 1.3005
R5327 Vss.n551 Vss.n550 1.3005
R5328 Vss.n989 Vss.n988 1.3005
R5329 Vss.n789 Vss.n788 1.3005
R5330 Vss.n788 Vss.n787 1.3005
R5331 Vss.n806 Vss.n805 1.3005
R5332 Vss.n798 Vss.n797 1.3005
R5333 Vss.n795 Vss.n794 1.3005
R5334 Vss.n796 Vss.n795 1.3005
R5335 Vss.n526 Vss.n517 1.3005
R5336 Vss.n1045 Vss.n1044 1.3005
R5337 Vss.n1046 Vss.n1045 1.3005
R5338 Vss.n446 Vss.n445 1.3005
R5339 Vss.n449 Vss.n448 1.3005
R5340 Vss.n448 Vss.n447 1.3005
R5341 Vss.n1183 Vss.n1182 1.3005
R5342 Vss.n1179 Vss.n426 1.3005
R5343 Vss.n930 Vss.n426 1.3005
R5344 Vss.n1166 Vss.n1165 1.3005
R5345 Vss.n1165 Vss.n425 1.3005
R5346 Vss.n1164 Vss.n1163 1.3005
R5347 Vss.n832 Vss.n831 1.3005
R5348 Vss.n831 Vss.n830 1.3005
R5349 Vss.n829 Vss.n785 1.3005
R5350 Vss.n822 Vss.n783 1.3005
R5351 Vss.n821 Vss.n820 1.3005
R5352 Vss.n821 Vss.n786 1.3005
R5353 Vss.n840 Vss.n839 1.3005
R5354 Vss.n814 Vss.n813 1.3005
R5355 Vss.n813 Vss.n812 1.3005
R5356 Vss.n610 Vss.n599 1.3005
R5357 Vss.n608 Vss.n598 1.3005
R5358 Vss.n609 Vss.n608 1.3005
R5359 Vss.n781 Vss.n780 1.3005
R5360 Vss.n782 Vss.n781 1.3005
R5361 Vss.n778 Vss.n777 1.3005
R5362 Vss.n777 Vss.n591 1.3005
R5363 Vss.n646 Vss.n645 1.3005
R5364 Vss.n645 Vss.n644 1.3005
R5365 Vss.n642 Vss.n625 1.3005
R5366 Vss.n627 Vss.n626 1.3005
R5367 Vss.n637 Vss.n636 1.3005
R5368 Vss.n638 Vss.n637 1.3005
R5369 Vss.n639 Vss.n620 1.3005
R5370 Vss.n653 Vss.n652 1.3005
R5371 Vss.n654 Vss.n653 1.3005
R5372 Vss.n9 Vss.n6 1.3005
R5373 Vss.n1913 Vss.n1912 1.3005
R5374 Vss.n1912 Vss.n1911 1.3005
R5375 Vss.n731 Vss.n730 1.3005
R5376 Vss.n733 Vss.n732 1.3005
R5377 Vss.n732 Vss.n7 1.3005
R5378 Vss.n706 Vss.n705 1.3005
R5379 Vss.n700 Vss.n699 1.3005
R5380 Vss.n699 Vss.n695 1.3005
R5381 Vss.n725 Vss.n724 1.3005
R5382 Vss.n721 Vss.n707 1.3005
R5383 Vss.n707 Vss.n696 1.3005
R5384 Vss.n716 Vss.n697 1.3005
R5385 Vss.n715 Vss.n714 1.3005
R5386 Vss.n715 Vss.n8 1.3005
R5387 Vss.n27 Vss.n26 1.3005
R5388 Vss.n24 Vss.n21 1.3005
R5389 Vss.n25 Vss.n24 1.3005
R5390 Vss.n20 Vss.n17 1.3005
R5391 Vss.n1896 Vss.n17 1.3005
R5392 Vss.n1894 Vss.n1893 1.3005
R5393 Vss.n1895 Vss.n1894 1.3005
R5394 Vss.n615 Vss.n613 1.3005
R5395 Vss.n666 Vss.n665 1.3005
R5396 Vss.n667 Vss.n666 1.3005
R5397 Vss.n619 Vss.n617 1.3005
R5398 Vss.n659 Vss.n658 1.3005
R5399 Vss.n658 Vss.n657 1.3005
R5400 Vss.n37 Vss.n36 1.3005
R5401 Vss.n1880 Vss.n1879 1.3005
R5402 Vss.n1879 Vss.n1878 1.3005
R5403 Vss.n1877 Vss.n1876 1.3005
R5404 Vss.n39 Vss.n38 1.3005
R5405 Vss.n684 Vss.n38 1.3005
R5406 Vss.n683 Vss.n682 1.3005
R5407 Vss.n681 Vss.n671 1.3005
R5408 Vss.n681 Vss.n680 1.3005
R5409 Vss.n679 Vss.n678 1.3005
R5410 Vss.n677 Vss.n672 1.3005
R5411 Vss.n677 Vss.n676 1.3005
R5412 Vss.n674 Vss.n673 1.3005
R5413 Vss.n675 Vss.n674 1.3005
R5414 Vss.n851 Vss.n850 1.3005
R5415 Vss.n590 Vss.n589 1.3005
R5416 Vss.n849 Vss.n590 1.3005
R5417 Vss.n848 Vss.n582 1.3005
R5418 Vss.n880 Vss.n879 1.3005
R5419 Vss.n879 Vss.n878 1.3005
R5420 Vss.n877 Vss.n876 1.3005
R5421 Vss.n875 Vss.n564 1.3005
R5422 Vss.n875 Vss.n874 1.3005
R5423 Vss.n873 Vss.n565 1.3005
R5424 Vss.n871 Vss.n870 1.3005
R5425 Vss.n872 Vss.n871 1.3005
R5426 Vss.n868 Vss.n867 1.3005
R5427 Vss.n867 Vss.n583 1.3005
R5428 Vss.n577 Vss.n575 1.3005
R5429 Vss.n894 Vss.n893 1.3005
R5430 Vss.n895 Vss.n894 1.3005
R5431 Vss.n884 Vss.n580 1.3005
R5432 Vss.n887 Vss.n886 1.3005
R5433 Vss.n886 Vss.n885 1.3005
R5434 Vss.n899 Vss.n567 1.3005
R5435 Vss.n901 Vss.n568 1.3005
R5436 Vss.n901 Vss.n900 1.3005
R5437 Vss.n571 Vss.n569 1.3005
R5438 Vss.n571 Vss.n440 1.3005
R5439 Vss.n906 Vss.n905 1.3005
R5440 Vss.n905 Vss.n904 1.3005
R5441 Vss.n758 Vss.n31 1.3005
R5442 Vss.n760 Vss.n32 1.3005
R5443 Vss.n760 Vss.n759 1.3005
R5444 Vss.n687 Vss.n33 1.3005
R5445 Vss.n687 Vss.n16 1.3005
R5446 Vss.n763 Vss.n34 1.3005
R5447 Vss.n764 Vss.n763 1.3005
R5448 Vss.n766 Vss.n603 1.3005
R5449 Vss.n769 Vss.n768 1.3005
R5450 Vss.n768 Vss.n767 1.3005
R5451 Vss.n594 Vss.n593 1.3005
R5452 Vss.n595 Vss.n594 1.3005
R5453 Vss.n856 Vss.n855 1.3005
R5454 Vss.n857 Vss.n856 1.3005
R5455 Vss.n863 Vss.n862 1.3005
R5456 Vss.n860 Vss.n859 1.3005
R5457 Vss.n861 Vss.n860 1.3005
R5458 Vss.n1160 Vss.n1159 1.3005
R5459 Vss.n1161 Vss.n1160 1.3005
R5460 Vss.n690 Vss.n689 1.3005
R5461 Vss.n739 Vss.n738 1.3005
R5462 Vss.n740 Vss.n739 1.3005
R5463 Vss.n756 Vss.n755 1.3005
R5464 Vss.n752 Vss.n751 1.3005
R5465 Vss.n751 Vss.n750 1.3005
R5466 Vss.n749 Vss.n748 1.3005
R5467 Vss.n747 Vss.n741 1.3005
R5468 Vss.n747 Vss.n746 1.3005
R5469 Vss.n744 Vss.n743 1.3005
R5470 Vss.n745 Vss.n744 1.3005
R5471 Vss.n742 Vss.n30 1.3005
R5472 Vss.n49 Vss.n44 1.29323
R5473 Vss.n49 Vss.n48 1.00923
R5474 Vss.n1851 Vss.n1850 0.999917
R5475 Vss.n1833 Vss.n1832 0.999917
R5476 Vss.n1834 Vss.n1833 0.999917
R5477 Vss.n1851 Vss.n58 0.999917
R5478 Vss.n1504 Vss.n146 0.990409
R5479 Vss.n853 Vss.n563 0.990409
R5480 Vss.n1156 Vss.n1155 0.990409
R5481 Vss.n982 Vss.n457 0.990409
R5482 Vss.n1882 Vss.n35 0.990409
R5483 Vss.n50 Vss.n49 0.984484
R5484 Vss.n1849 Vss.n1848 0.949529
R5485 Vss.n737 Vss.n691 0.92075
R5486 Vss.n838 Vss.n815 0.92075
R5487 Vss.n881 Vss.n581 0.92075
R5488 Vss.n889 Vss.n888 0.92075
R5489 Vss.n1181 Vss.n1180 0.92075
R5490 Vss.n1043 Vss.n518 0.92075
R5491 Vss.n923 Vss.n918 0.92075
R5492 Vss.n1197 Vss.n418 0.92075
R5493 Vss.n1277 Vss.n329 0.92075
R5494 Vss.n1583 Vss.n1579 0.92075
R5495 Vss.n1589 Vss.n1588 0.92075
R5496 Vss.n1715 Vss.n1714 0.92075
R5497 Vss.n1799 Vss.n1798 0.92075
R5498 Vss.n1686 Vss.n1638 0.92075
R5499 Vss.n1820 Vss.n72 0.92075
R5500 Vss.n1824 Vss.n1823 0.92075
R5501 Vss.n1443 Vss.n253 0.92075
R5502 Vss.n1388 Vss.n287 0.92075
R5503 Vss.n1380 Vss.n294 0.92075
R5504 Vss.n1357 Vss.n1352 0.92075
R5505 Vss.n945 Vss.n943 0.92075
R5506 Vss.n1392 Vss.n1391 0.92075
R5507 Vss.n1295 Vss.n1291 0.92075
R5508 Vss.n1350 Vss.n304 0.92075
R5509 Vss.n1218 Vss.n354 0.92075
R5510 Vss.n1207 Vss.n352 0.92075
R5511 Vss.n1305 Vss.n1299 0.92075
R5512 Vss.n376 Vss.n371 0.92075
R5513 Vss.n1420 Vss.n264 0.92075
R5514 Vss.n269 Vss.n263 0.92075
R5515 Vss.n406 Vss.n274 0.92075
R5516 Vss.n1287 Vss.n321 0.92075
R5517 Vss.n384 Vss.n383 0.92075
R5518 Vss.n414 Vss.n367 0.92075
R5519 Vss.n394 Vss.n393 0.92075
R5520 Vss.n1333 Vss.n260 0.92075
R5521 Vss.n1403 Vss.n275 0.92075
R5522 Vss.n1320 Vss.n1319 0.92075
R5523 Vss.n1313 Vss.n1308 0.92075
R5524 Vss.n1265 Vss.n1264 0.92075
R5525 Vss.n968 Vss.n966 0.92075
R5526 Vss.n1275 Vss.n1269 0.92075
R5527 Vss.n1242 Vss.n348 0.92075
R5528 Vss.n1258 Vss.n1257 0.92075
R5529 Vss.n1252 Vss.n341 0.92075
R5530 Vss.n1599 Vss.n152 0.92075
R5531 Vss.n1112 Vss.n1082 0.92075
R5532 Vss.n1096 Vss.n1089 0.92075
R5533 Vss.n1069 Vss.n1068 0.92075
R5534 Vss.n1108 Vss.n1085 0.92075
R5535 Vss.n1561 Vss.n1556 0.92075
R5536 Vss.n139 Vss.n134 0.92075
R5537 Vss.n1792 Vss.n94 0.92075
R5538 Vss.n1671 Vss.n1633 0.92075
R5539 Vss.n1658 Vss.n1653 0.92075
R5540 Vss.n1703 Vss.n1631 0.92075
R5541 Vss.n1699 Vss.n1698 0.92075
R5542 Vss.n1647 Vss.n1646 0.92075
R5543 Vss.n1711 Vss.n1623 0.92075
R5544 Vss.n1130 Vss.n461 0.92075
R5545 Vss.n498 Vss.n497 0.92075
R5546 Vss.n482 Vss.n477 0.92075
R5547 Vss.n492 Vss.n487 0.92075
R5548 Vss.n1127 Vss.n463 0.92075
R5549 Vss.n995 Vss.n992 0.92075
R5550 Vss.n1038 Vss.n524 0.92075
R5551 Vss.n207 Vss.n202 0.92075
R5552 Vss.n1514 Vss.n211 0.92075
R5553 Vss.n1566 Vss.n1565 0.92075
R5554 Vss.n1543 Vss.n1541 0.92075
R5555 Vss.n1552 Vss.n175 0.92075
R5556 Vss.n1376 Vss.n1372 0.92075
R5557 Vss.n1536 Vss.n188 0.92075
R5558 Vss.n1369 Vss.n1364 0.92075
R5559 Vss.n183 Vss.n182 0.92075
R5560 Vss.n1456 Vss.n1450 0.92075
R5561 Vss.n1808 Vss.n79 0.92075
R5562 Vss.n1429 Vss.n78 0.92075
R5563 Vss.n1460 Vss.n1459 0.92075
R5564 Vss.n1575 Vss.n163 0.92075
R5565 Vss.n1524 Vss.n1519 0.92075
R5566 Vss.n1526 Vss.n198 0.92075
R5567 Vss.n1240 Vss.n1236 0.92075
R5568 Vss.n1730 Vss.n128 0.92075
R5569 Vss.n937 Vss.n928 0.92075
R5570 Vss.n1191 Vss.n420 0.92075
R5571 Vss.n804 Vss.n790 0.92075
R5572 Vss.n799 Vss.n793 0.92075
R5573 Vss.n1167 Vss.n432 0.92075
R5574 Vss.n833 Vss.n828 0.92075
R5575 Vss.n823 Vss.n819 0.92075
R5576 Vss.n651 Vss.n621 0.92075
R5577 Vss.n661 Vss.n660 0.92075
R5578 Vss.n647 Vss.n624 0.92075
R5579 Vss.n635 Vss.n628 0.92075
R5580 Vss.n1914 Vss.n5 0.92075
R5581 Vss.n734 Vss.n694 0.92075
R5582 Vss.n717 Vss.n713 0.92075
R5583 Vss.n723 Vss.n722 0.92075
R5584 Vss.n1848 Vss.n60 0.907842
R5585 Vss.n1843 Vss.n1842 0.867167
R5586 Vss.t2 Vss.n65 0.867167
R5587 Vss.n1845 Vss.n57 0.867167
R5588 SARlogic_0.dffrs_12.d SARlogic_0.dffrs_12.nand3_8.A 0.784786
R5589 SARlogic_0.dffrs_13.d SARlogic_0.dffrs_13.nand3_8.A 0.784786
R5590 Vss.n1555 Vss.n93 0.780467
R5591 Vss.n1010 Vss.n1009 0.771017
R5592 Vss.n907 Vss.n906 0.771017
R5593 Vss.n1496 Vss.n1495 0.771017
R5594 Vss.n779 Vss.n778 0.771017
R5595 Vss.n1893 Vss.n1892 0.771017
R5596 adc_PISO_0.avss Vss.n1781 0.762138
R5597 Vss.n1872 Vss.n1871 0.714636
R5598 Vss.n1781 Vss.n1780 0.679217
R5599 Vss.n1150 Vss.n1147 0.669813
R5600 Vss.n1154 Vss.n1153 0.669683
R5601 Vss.n914 Vss.n913 0.669683
R5602 Vss.n1849 comparator_no_offsetcal_0.no_offsetLatch_0.VSS 0.664071
R5603 Vss.n1873 Vss.n41 0.651683
R5604 SARlogic_0.dffrs_12.clk Vss.n1176 0.611214
R5605 Vss.n754 Vss.n42 0.601415
R5606 Vss.n1606 Vss.n1605 0.600912
R5607 Vss.n1768 Vss.n1767 0.471317
R5608 Vss.n852 Vss.n589 0.463217
R5609 Vss.n671 Vss.n670 0.463217
R5610 Vss.n1608 Vss.n1607 0.463217
R5611 Vss.n1762 Vss.n110 0.463217
R5612 Vss.n1763 Vss.n109 0.463217
R5613 Vss.n1756 Vss.n1755 0.463217
R5614 Vss.n1750 Vss.n103 0.463217
R5615 Vss.n1784 Vss.n1783 0.463217
R5616 Vss.n1773 Vss.n104 0.463217
R5617 Vss.n1503 Vss.n1502 0.463217
R5618 Vss.n1488 Vss.n1487 0.463217
R5619 Vss.n1482 Vss.n215 0.463217
R5620 Vss.n1506 Vss.n1505 0.463217
R5621 Vss.n1010 Vss.n542 0.463217
R5622 Vss.n1011 Vss.n541 0.463217
R5623 Vss.n908 Vss.n568 0.463217
R5624 Vss.n907 Vss.n569 0.463217
R5625 Vss.n912 Vss.n564 0.463217
R5626 Vss.n859 Vss.n443 0.463217
R5627 Vss.n1159 Vss.n1158 0.463217
R5628 Vss.n1157 Vss.n444 0.463217
R5629 Vss.n450 Vss.n449 0.463217
R5630 Vss.n1017 Vss.n452 0.463217
R5631 Vss.n985 Vss.n553 0.463217
R5632 Vss.n984 Vss.n554 0.463217
R5633 Vss.n983 Vss.n555 0.463217
R5634 Vss.n981 Vss.n980 0.463217
R5635 Vss.n1146 Vss.n1145 0.463217
R5636 Vss.n1494 Vss.n220 0.463217
R5637 Vss.n1495 Vss.n219 0.463217
R5638 Vss.n776 Vss.n598 0.463217
R5639 Vss.n780 Vss.n779 0.463217
R5640 Vss.n1881 Vss.n1880 0.463217
R5641 Vss.n1885 Vss.n32 0.463217
R5642 Vss.n1884 Vss.n33 0.463217
R5643 Vss.n1883 Vss.n34 0.463217
R5644 Vss.n753 Vss.n752 0.463217
R5645 Vss.n1891 Vss.n21 0.463217
R5646 Vss.n1892 Vss.n20 0.463217
R5647 Vss.n770 Vss.n769 0.463217
R5648 Vss.n593 Vss.n588 0.463217
R5649 Vss.n855 Vss.n854 0.463217
R5650 Vss.n560 Vss.n454 0.441453
R5651 Vss.n63 comparator_no_offsetcal_0.VSS 0.404079
R5652 Vss.n1872 Vss.n42 0.328611
R5653 Vss.n1763 Vss.n1762 0.3083
R5654 Vss.n1756 Vss.n103 0.3083
R5655 Vss.n1783 Vss.n103 0.3083
R5656 Vss.n1488 Vss.n215 0.3083
R5657 Vss.n1505 Vss.n215 0.3083
R5658 Vss.n1011 Vss.n1010 0.3083
R5659 Vss.n908 Vss.n907 0.3083
R5660 Vss.n1158 Vss.n443 0.3083
R5661 Vss.n1158 Vss.n1157 0.3083
R5662 Vss.n985 Vss.n984 0.3083
R5663 Vss.n984 Vss.n983 0.3083
R5664 Vss.n1495 Vss.n1494 0.3083
R5665 Vss.n779 Vss.n776 0.3083
R5666 Vss.n1885 Vss.n1884 0.3083
R5667 Vss.n1884 Vss.n1883 0.3083
R5668 Vss.n1892 Vss.n1891 0.3083
R5669 Vss.n770 Vss.n588 0.3083
R5670 Vss.n854 Vss.n588 0.3083
R5671 Vss.n1767 Vss.n1763 0.3002
R5672 Vss.n915 Vss.n914 0.284919
R5673 Vss.n1765 Vss.n1764 0.252687
R5674 Vss.n1847 Vss.n63 0.238053
R5675 Vss.n1757 Vss.n1756 0.2165
R5676 Vss.n1489 Vss.n1488 0.2165
R5677 Vss.n864 Vss.n443 0.2165
R5678 Vss.n986 Vss.n985 0.2165
R5679 Vss.n1886 Vss.n1885 0.2165
R5680 Vss.n771 Vss.n770 0.2165
R5681 Vss.n1870 Vss.n43 0.211763
R5682 Vss.n925 Vss.n560 0.195855
R5683 comparator_no_offsetcal_0.x5.avss Vss.n1869 0.188808
R5684 comparator_no_offsetcal_0.x3.avss Vss.n62 0.188808
R5685 Vss.n1505 Vss.n1504 0.1748
R5686 Vss.n1157 Vss.n1156 0.1748
R5687 Vss.n1883 Vss.n1882 0.1748
R5688 Vss.n854 Vss.n853 0.1748
R5689 Vss.n983 Vss.n982 0.17465
R5690 Vss.n1848 Vss.n1847 0.163684
R5691 Vss.n1837 comparator_no_offsetcal_0.no_offsetLatch_0.VSS 0.1605
R5692 Vss.n1783 Vss.n1782 0.1598
R5693 Vss.n1859 Vss.n1858 0.154786
R5694 Vss.n1902 Vss.n1899 0.154786
R5695 Vss.n1782 Vss.n104 0.152487
R5696 Vss.n1758 Vss.n1757 0.148459
R5697 Vss.n1490 Vss.n1489 0.148459
R5698 Vss.n865 Vss.n864 0.148459
R5699 Vss.n987 Vss.n986 0.148459
R5700 Vss.n1887 Vss.n1886 0.148459
R5701 Vss.n772 Vss.n771 0.148459
R5702 Vss.n1152 Vss.n1151 0.145432
R5703 Vss.n1149 Vss.n1148 0.145432
R5704 Vss.n1554 Vss.n131 0.143322
R5705 Vss.n926 Vss.n925 0.140365
R5706 Vss.n982 Vss.n981 0.13865
R5707 Vss.n1504 Vss.n1503 0.1385
R5708 Vss.n1156 Vss.n450 0.1385
R5709 Vss.n1882 Vss.n1881 0.1385
R5710 Vss.n853 Vss.n852 0.1385
R5711 Vss.n1148 Vss.n148 0.136253
R5712 Vss.n1855 Vss.n55 0.1355
R5713 Vss.n1904 Vss.n1903 0.1355
R5714 Vss.n1869 Vss.n1868 0.128901
R5715 Vss.n62 Vss.n61 0.127885
R5716 Vss.n430 Vss.n429 0.122607
R5717 Vss.n369 Vss.n368 0.122607
R5718 Vss.n1092 Vss.n1091 0.122607
R5719 Vss.n485 Vss.n474 0.122607
R5720 Vss.n802 Vss.n801 0.122607
R5721 Vss.n826 Vss.n825 0.122607
R5722 Vss.n632 Vss.n631 0.122607
R5723 Vss.n710 Vss.n709 0.122607
R5724 Vss.n927 Vss.n926 0.118169
R5725 Vss.n1701 Vss.n1635 0.115241
R5726 Vss.n60 Vss.n43 0.112526
R5727 Vss.n1861 Vss.n1860 0.109786
R5728 Vss.n1151 Vss.n1150 0.104592
R5729 Vss.n1661 Vss.n1660 0.10457
R5730 Vss.n494 Vss.n462 0.10457
R5731 Vss.n1041 Vss.n1040 0.10457
R5732 Vss.n1727 Vss.n1726 0.10457
R5733 Vss.n835 Vss.n578 0.10457
R5734 Vss.n649 Vss.n616 0.10457
R5735 Vss.n693 Vss.n3 0.10457
R5736 SARlogic_0.dffrs_14.vss Vss.n92 0.102612
R5737 Vss.n1378 SARlogic_0.dffrs_8.vss 0.102537
R5738 Vss.n1289 SARlogic_0.dffrs_10.vss 0.102537
R5739 Vss.n1538 SARlogic_0.dffrs_7.vss 0.101537
R5740 Vss.n1290 SARlogic_0.dffrs_9.vss 0.101537
R5741 Vss.n1153 Vss.n1152 0.0911096
R5742 Vss.n1917 Vss.n2 0.0796966
R5743 Vss.n1177 Vss.n1173 0.078611
R5744 Vss.n927 Vss.n561 0.0781858
R5745 Vss.n1148 Vss.n210 0.0776599
R5746 Vss.n1149 Vss.n340 0.0776599
R5747 Vss.n1152 Vss.n455 0.0776599
R5748 Vss.n1151 Vss.n339 0.0776599
R5749 Vss.n1759 Vss.n113 0.073981
R5750 Vss.n869 Vss.n566 0.073981
R5751 Vss.n547 Vss.n539 0.073981
R5752 Vss.n1491 Vss.n223 0.073981
R5753 Vss.n1888 Vss.n29 0.073981
R5754 Vss.n773 Vss.n601 0.073981
R5755 Vss.n1110 Vss.n150 0.0685048
R5756 Vss.n890 Vss.n579 0.0679983
R5757 Vss.n1067 Vss.n1066 0.0679983
R5758 Vss.n508 Vss.n507 0.0679983
R5759 Vss.n994 Vss.n993 0.0679983
R5760 Vss.n702 Vss.n701 0.0679983
R5761 Vss.n1150 Vss.n456 0.0673674
R5762 Vss.n1153 Vss.n453 0.0673025
R5763 Vss.n914 Vss.n562 0.0673025
R5764 Vss.n1194 Vss.n353 0.0660086
R5765 Vss.n1220 Vss.n353 0.0655096
R5766 Vss.n407 Vss.n387 0.0645882
R5767 Vss.n1193 Vss.n1192 0.0645882
R5768 Vss.n1762 Vss.n1761 0.0635
R5769 Vss.n1012 Vss.n1011 0.0635
R5770 Vss.n909 Vss.n908 0.0635
R5771 Vss.n1494 Vss.n1493 0.0635
R5772 Vss.n776 Vss.n775 0.0635
R5773 Vss.n1891 Vss.n1890 0.0635
R5774 Vss.n1621 Vss.n1620 0.0625376
R5775 Vss.n711 Vss.n710 0.0622481
R5776 Vss.n825 Vss.n817 0.0622481
R5777 Vss.n410 Vss.n368 0.0622481
R5778 Vss.n1093 Vss.n1092 0.0622481
R5779 Vss.n475 Vss.n474 0.0622481
R5780 Vss.n801 Vss.n521 0.0622481
R5781 Vss.n1170 Vss.n429 0.0622481
R5782 Vss.n631 Vss.n630 0.0622481
R5783 Vss.n1542 Vss.n89 0.0616538
R5784 Vss.n1516 Vss.n1515 0.0616538
R5785 Vss.n1447 Vss.n186 0.0616538
R5786 Vss.n1379 Vss.n252 0.0616538
R5787 Vss.n350 Vss.n349 0.0616538
R5788 Vss.n967 Vss.n333 0.0616538
R5789 Vss.n1307 Vss.n316 0.0616538
R5790 Vss.n1288 Vss.n320 0.0616538
R5791 Vss.n944 Vss.n330 0.0616538
R5792 Vss.n1578 Vss.n160 0.0615256
R5793 Vss.n1873 Vss.n1872 0.0600636
R5794 Vss.n1129 Vss.n1128 0.0568904
R5795 Vss.n1039 Vss.n523 0.0568904
R5796 Vss.n883 Vss.n882 0.0568904
R5797 Vss.n736 Vss.n735 0.0568904
R5798 Vss.n151 Vss.n150 0.0566774
R5799 Vss.n1605 Vss.n1604 0.0561349
R5800 Vss.n916 Vss.n915 0.0551896
R5801 Vss.n925 Vss.n428 0.0551896
R5802 Vss.n1661 Vss.n1635 0.054837
R5803 Vss.n1128 Vss.n462 0.054837
R5804 Vss.n1040 Vss.n1039 0.054837
R5805 Vss.n1726 Vss.n131 0.054837
R5806 Vss.n883 Vss.n578 0.054837
R5807 Vss.n618 Vss.n616 0.054837
R5808 Vss.n735 Vss.n693 0.054837
R5809 Vss.n1153 Vss.n454 0.0521009
R5810 Vss.n618 Vss.n40 0.0502328
R5811 Vss.n1605 Vss.n147 0.0480028
R5812 Vss.n1290 Vss.n315 0.0478478
R5813 Vss.n455 Vss.n332 0.0478478
R5814 Vss.n1254 Vss.n339 0.0478478
R5815 Vss.n1649 Vss.n93 0.0478478
R5816 Vss.n1539 Vss.n1538 0.0478478
R5817 Vss.n200 Vss.n129 0.0478478
R5818 Vss.n1794 Vss.n92 0.0478478
R5819 Vss.n210 Vss.n209 0.0478478
R5820 Vss.n1233 Vss.n340 0.0478478
R5821 Vss.n1378 Vss.n187 0.0478478
R5822 Vss.n1297 Vss.n1289 0.0478478
R5823 Vss.n941 Vss.n560 0.0478478
R5824 Vss.n1874 Vss.n40 0.0467
R5825 Vss.n1660 Vss.n1640 0.0466843
R5826 Vss.n494 Vss.n493 0.0466843
R5827 Vss.n1728 Vss.n1727 0.0466843
R5828 Vss.n1041 Vss.n520 0.0466843
R5829 Vss.n835 Vss.n834 0.0466843
R5830 Vss.n649 Vss.n648 0.0466843
R5831 Vss.n924 Vss.n916 0.0465106
R5832 Vss.n1178 Vss.n428 0.0465106
R5833 Vss.n1173 Vss.n1172 0.0465106
R5834 Vss.n1363 Vss.n296 0.0465022
R5835 Vss.n1371 Vss.n1370 0.0465022
R5836 Vss.n1351 Vss.n286 0.0465022
R5837 Vss.n1222 Vss.n1221 0.0465022
R5838 Vss.n1554 Vss.n1553 0.0464521
R5839 Vss.n1860 Vss.n1859 0.0455
R5840 Vss.n1899 Vss.n2 0.0455
R5841 Vss.n817 Vss.n578 0.0415307
R5842 Vss.n410 Vss.n409 0.0415307
R5843 Vss.n1093 Vss.n150 0.0415307
R5844 Vss.n475 Vss.n462 0.0415307
R5845 Vss.n1040 Vss.n521 0.0415307
R5846 Vss.n1171 Vss.n1170 0.0415307
R5847 Vss.n630 Vss.n616 0.0415307
R5848 Vss.n711 Vss.n693 0.0415307
R5849 Vss.n1150 Vss.n1149 0.0413406
R5850 Vss.n413 Vss.n412 0.0405109
R5851 Vss.n1109 Vss.n1084 0.0405109
R5852 Vss.n1095 Vss.n1090 0.0405109
R5853 Vss.n1111 Vss.n1083 0.0405109
R5854 Vss.n1648 Vss.n1640 0.0405109
R5855 Vss.n1659 Vss.n1652 0.0405109
R5856 Vss.n493 Vss.n486 0.0405109
R5857 Vss.n483 Vss.n476 0.0405109
R5858 Vss.n495 Vss.n473 0.0405109
R5859 Vss.n1729 Vss.n1728 0.0405109
R5860 Vss.n1584 Vss.n130 0.0405109
R5861 Vss.n803 Vss.n520 0.0405109
R5862 Vss.n800 Vss.n792 0.0405109
R5863 Vss.n1042 Vss.n519 0.0405109
R5864 Vss.n1168 Vss.n431 0.0405109
R5865 Vss.n834 Vss.n827 0.0405109
R5866 Vss.n824 Vss.n818 0.0405109
R5867 Vss.n837 Vss.n836 0.0405109
R5868 Vss.n648 Vss.n623 0.0405109
R5869 Vss.n634 Vss.n629 0.0405109
R5870 Vss.n650 Vss.n622 0.0405109
R5871 Vss.n1915 Vss.n4 0.0405109
R5872 Vss.n720 Vss.n708 0.0405109
R5873 Vss.n718 Vss.n712 0.0405109
R5874 Vss.n561 Vss.n351 0.040346
R5875 Vss.n1916 Vss.n3 0.0399832
R5876 Vss.n1759 Vss.n1758 0.0389018
R5877 Vss.n865 Vss.n566 0.0389018
R5878 Vss.n987 Vss.n539 0.0389018
R5879 Vss.n1491 Vss.n1490 0.0389018
R5880 Vss.n1888 Vss.n1887 0.0389018
R5881 Vss.n773 Vss.n772 0.0389018
R5882 Vss.n1702 Vss.n1701 0.0368083
R5883 Vss.n1670 Vss.n1634 0.036505
R5884 Vss.n1809 Vss.n71 0.036505
R5885 Vss.n1430 Vss.n1423 0.036505
R5886 Vss.n1422 Vss.n262 0.036505
R5887 Vss.n1404 Vss.n261 0.036505
R5888 Vss.n1314 Vss.n1307 0.0361576
R5889 Vss.n1268 Vss.n330 0.0361576
R5890 Vss.n1256 Vss.n333 0.0361576
R5891 Vss.n1650 Vss.n1621 0.0361576
R5892 Vss.n1449 Vss.n1447 0.0361576
R5893 Vss.n1235 Vss.n350 0.0361576
R5894 Vss.n1586 Vss.n1578 0.0361576
R5895 Vss.n1796 Vss.n89 0.0361576
R5896 Vss.n1518 Vss.n1516 0.0361576
R5897 Vss.n1444 Vss.n252 0.0361576
R5898 Vss.n320 Vss.n318 0.0361576
R5899 Vss.n938 Vss.n926 0.0361576
R5900 Vss.n507 Vss.n456 0.035635
R5901 Vss.n994 Vss.n453 0.035635
R5902 Vss.n579 Vss.n562 0.035635
R5903 Vss.n701 Vss.n692 0.035635
R5904 Vss.n692 Vss.n42 0.0352182
R5905 Vss.n891 Vss.n578 0.0349747
R5906 Vss.n409 Vss.n408 0.0349747
R5907 Vss.n1065 Vss.n150 0.0349747
R5908 Vss.n509 Vss.n462 0.0349747
R5909 Vss.n1040 Vss.n522 0.0349747
R5910 Vss.n1171 Vss.n419 0.0349747
R5911 Vss.n663 Vss.n616 0.0349747
R5912 Vss.n703 Vss.n693 0.0349747
R5913 Vss.n1066 Vss.n149 0.0346145
R5914 Vss.n1712 Vss.n1621 0.0340549
R5915 Vss.n1209 Vss.n351 0.0339793
R5916 Vss.n89 Vss.n88 0.0335769
R5917 Vss.n201 Vss.n160 0.0335769
R5918 Vss.n1515 Vss.n210 0.0335769
R5919 Vss.n1525 Vss.n1516 0.0335769
R5920 Vss.n1457 Vss.n1447 0.0335769
R5921 Vss.n1316 Vss.n252 0.0335769
R5922 Vss.n349 Vss.n340 0.0335769
R5923 Vss.n1241 Vss.n350 0.0335769
R5924 Vss.n967 Vss.n339 0.0335769
R5925 Vss.n1259 Vss.n333 0.0335769
R5926 Vss.n1307 Vss.n314 0.0335769
R5927 Vss.n377 Vss.n320 0.0335769
R5928 Vss.n944 Vss.n455 0.0335769
R5929 Vss.n1276 Vss.n330 0.0335769
R5930 Vss.n1577 Vss.n159 0.0334487
R5931 Vss.n817 Vss.n816 0.0322085
R5932 Vss.n1169 Vss.n430 0.0322085
R5933 Vss.n1298 Vss.n317 0.0322085
R5934 Vss.n1445 Vss.n251 0.0322085
R5935 Vss.n1795 Vss.n90 0.0322085
R5936 Vss.n1322 Vss.n315 0.0322085
R5937 Vss.n411 Vss.n369 0.0322085
R5938 Vss.n411 Vss.n410 0.0322085
R5939 Vss.n1267 Vss.n332 0.0322085
R5940 Vss.n1267 Vss.n331 0.0322085
R5941 Vss.n1255 Vss.n1254 0.0322085
R5942 Vss.n1094 Vss.n1091 0.0322085
R5943 Vss.n1094 Vss.n1093 0.0322085
R5944 Vss.n1651 Vss.n1649 0.0322085
R5945 Vss.n485 Vss.n484 0.0322085
R5946 Vss.n484 Vss.n475 0.0322085
R5947 Vss.n791 Vss.n521 0.0322085
R5948 Vss.n1539 Vss.n185 0.0322085
R5949 Vss.n1234 Vss.n1233 0.0322085
R5950 Vss.n1234 Vss.n1231 0.0322085
R5951 Vss.n1585 Vss.n129 0.0322085
R5952 Vss.n1585 Vss.n132 0.0322085
R5953 Vss.n1651 Vss.n1622 0.0322085
R5954 Vss.n1795 Vss.n1794 0.0322085
R5955 Vss.n209 Vss.n161 0.0322085
R5956 Vss.n1517 Vss.n161 0.0322085
R5957 Vss.n1448 Vss.n185 0.0322085
R5958 Vss.n1445 Vss.n187 0.0322085
R5959 Vss.n1255 Vss.n335 0.0322085
R5960 Vss.n1323 Vss.n1322 0.0322085
R5961 Vss.n1298 Vss.n1297 0.0322085
R5962 Vss.n941 Vss.n940 0.0322085
R5963 Vss.n940 Vss.n561 0.0322085
R5964 Vss.n802 Vss.n791 0.0322085
R5965 Vss.n1170 Vss.n1169 0.0322085
R5966 Vss.n826 Vss.n816 0.0322085
R5967 Vss.n633 Vss.n630 0.0322085
R5968 Vss.n633 Vss.n632 0.0322085
R5969 Vss.n719 Vss.n709 0.0322085
R5970 Vss.n719 Vss.n711 0.0322085
R5971 Vss.n1604 Vss.n1603 0.0317776
R5972 Vss.n925 Vss.n924 0.0308765
R5973 Vss.n1604 Vss.n148 0.0306923
R5974 Vss.n917 Vss.n916 0.0268641
R5975 Vss.n1378 Vss.n295 0.0268641
R5976 Vss.n1289 Vss.n319 0.0268641
R5977 Vss.n385 Vss.n320 0.0268641
R5978 Vss.n1321 Vss.n252 0.0268641
R5979 Vss.n965 Vss.n339 0.0268641
R5980 Vss.n1266 Vss.n333 0.0268641
R5981 Vss.n350 Vss.n338 0.0268641
R5982 Vss.n1253 Vss.n340 0.0268641
R5983 Vss.n1540 Vss.n92 0.0268641
R5984 Vss.n184 Vss.n89 0.0268641
R5985 Vss.n1516 Vss.n199 0.0268641
R5986 Vss.n1621 Vss.n91 0.0268641
R5987 Vss.n1793 Vss.n93 0.0268641
R5988 Vss.n1577 Vss.n1576 0.0268641
R5989 Vss.n208 Vss.n201 0.0268641
R5990 Vss.n1232 Vss.n210 0.0268641
R5991 Vss.n1447 Vss.n1446 0.0268641
R5992 Vss.n1538 Vss.n1537 0.0268641
R5993 Vss.n1307 Vss.n1306 0.0268641
R5994 Vss.n1296 Vss.n1290 0.0268641
R5995 Vss.n942 Vss.n455 0.0268641
R5996 Vss.n939 Vss.n330 0.0268641
R5997 Vss.n428 Vss.n427 0.0268641
R5998 Vss.n1555 Vss.n1554 0.0263346
R5999 Vss.n1611 Vss.n113 0.0258591
R6000 Vss.n1734 Vss.n113 0.0258591
R6001 Vss.n870 Vss.n869 0.0258591
R6002 Vss.n869 Vss.n868 0.0258591
R6003 Vss.n547 Vss.n546 0.0258591
R6004 Vss.n548 Vss.n547 0.0258591
R6005 Vss.n1135 Vss.n223 0.0258591
R6006 Vss.n1136 Vss.n223 0.0258591
R6007 Vss.n741 Vss.n29 0.0258591
R6008 Vss.n743 Vss.n29 0.0258591
R6009 Vss.n672 Vss.n601 0.0258591
R6010 Vss.n673 Vss.n601 0.0258591
R6011 Vss.n1661 Vss.n1622 0.0237454
R6012 Vss.n1662 Vss.n90 0.0235512
R6013 Vss.n1726 Vss.n132 0.0235512
R6014 Vss.n1517 Vss.n133 0.0235512
R6015 Vss.n1448 Vss.n77 0.0235512
R6016 Vss.n259 Vss.n251 0.0235512
R6017 Vss.n1231 Vss.n1230 0.0235512
R6018 Vss.n1229 Vss.n335 0.0235512
R6019 Vss.n1324 Vss.n1323 0.0235512
R6020 Vss.n317 Vss.n273 0.0235512
R6021 Vss.n1228 Vss.n331 0.0235512
R6022 Vss.n662 Vss.n40 0.0232899
R6023 Vss.n1760 Vss.n1759 0.023066
R6024 Vss.n910 Vss.n566 0.023066
R6025 Vss.n1013 Vss.n539 0.023066
R6026 Vss.n1492 Vss.n1491 0.023066
R6027 Vss.n1889 Vss.n1888 0.023066
R6028 Vss.n774 Vss.n773 0.023066
R6029 Vss.n1712 Vss.n1622 0.0226532
R6030 Vss.n1173 Vss.n1171 0.0225109
R6031 Vss.n1228 Vss.n351 0.0225109
R6032 Vss.n1229 Vss.n1228 0.0225109
R6033 Vss.n1230 Vss.n1229 0.0225109
R6034 Vss.n1230 Vss.n133 0.0225109
R6035 Vss.n1725 Vss.n133 0.0225109
R6036 Vss.n1662 Vss.n1661 0.0225109
R6037 Vss.n1662 Vss.n77 0.0225109
R6038 Vss.n259 Vss.n77 0.0225109
R6039 Vss.n1324 Vss.n259 0.0225109
R6040 Vss.n1324 Vss.n273 0.0225109
R6041 Vss.n409 Vss.n273 0.0225109
R6042 Vss.n1422 Vss.n261 0.0223682
R6043 Vss.n1423 Vss.n1422 0.0223682
R6044 Vss.n1423 Vss.n71 0.0223682
R6045 Vss.n1634 Vss.n71 0.0223682
R6046 Vss.n1701 Vss.n1634 0.0223682
R6047 Vss.n387 Vss.n261 0.0223682
R6048 Vss.n1194 Vss.n1193 0.0223682
R6049 Vss.n90 Vss.n88 0.0223376
R6050 Vss.n1525 Vss.n1517 0.0223376
R6051 Vss.n1457 Vss.n1448 0.0223376
R6052 Vss.n1316 Vss.n251 0.0223376
R6053 Vss.n1241 Vss.n1231 0.0223376
R6054 Vss.n1259 Vss.n335 0.0223376
R6055 Vss.n1323 Vss.n314 0.0223376
R6056 Vss.n377 Vss.n317 0.0223376
R6057 Vss.n1276 Vss.n331 0.0223376
R6058 Vss.n162 Vss.n132 0.0222094
R6059 Vss.n1833 Vss.n1831 0.0215413
R6060 Vss.n1852 Vss.n1851 0.0215413
R6061 Vss.n917 Vss.n430 0.0214837
R6062 Vss.n315 Vss.n295 0.0214837
R6063 Vss.n369 Vss.n319 0.0214837
R6064 Vss.n411 Vss.n385 0.0214837
R6065 Vss.n1322 Vss.n1321 0.0214837
R6066 Vss.n965 Vss.n332 0.0214837
R6067 Vss.n1267 Vss.n1266 0.0214837
R6068 Vss.n1255 Vss.n338 0.0214837
R6069 Vss.n1254 Vss.n1253 0.0214837
R6070 Vss.n1091 Vss.n1084 0.0214837
R6071 Vss.n1094 Vss.n1083 0.0214837
R6072 Vss.n1649 Vss.n1648 0.0214837
R6073 Vss.n1652 Vss.n1651 0.0214837
R6074 Vss.n486 Vss.n485 0.0214837
R6075 Vss.n484 Vss.n473 0.0214837
R6076 Vss.n1540 Vss.n1539 0.0214837
R6077 Vss.n185 Vss.n184 0.0214837
R6078 Vss.n1234 Vss.n199 0.0214837
R6079 Vss.n1729 Vss.n129 0.0214837
R6080 Vss.n1585 Vss.n1584 0.0214837
R6081 Vss.n1795 Vss.n91 0.0214837
R6082 Vss.n1794 Vss.n1793 0.0214837
R6083 Vss.n1576 Vss.n161 0.0214837
R6084 Vss.n209 Vss.n208 0.0214837
R6085 Vss.n1233 Vss.n1232 0.0214837
R6086 Vss.n1446 Vss.n1445 0.0214837
R6087 Vss.n1537 Vss.n187 0.0214837
R6088 Vss.n1306 Vss.n1298 0.0214837
R6089 Vss.n1297 Vss.n1296 0.0214837
R6090 Vss.n942 Vss.n941 0.0214837
R6091 Vss.n940 Vss.n939 0.0214837
R6092 Vss.n803 Vss.n802 0.0214837
R6093 Vss.n791 Vss.n519 0.0214837
R6094 Vss.n1169 Vss.n427 0.0214837
R6095 Vss.n827 Vss.n826 0.0214837
R6096 Vss.n837 Vss.n816 0.0214837
R6097 Vss.n632 Vss.n623 0.0214837
R6098 Vss.n633 Vss.n622 0.0214837
R6099 Vss.n709 Vss.n4 0.0214837
R6100 Vss.n719 Vss.n718 0.0214837
R6101 Vss.n1172 Vss.n353 0.0204141
R6102 Vss.n1661 Vss.n1632 0.0200312
R6103 Vss.n1701 Vss.n1700 0.0199048
R6104 Vss.n1669 Vss.n1662 0.019868
R6105 Vss.n1362 Vss.n133 0.019868
R6106 Vss.n1810 Vss.n77 0.019868
R6107 Vss.n1431 Vss.n259 0.019868
R6108 Vss.n1230 Vss.n302 0.019868
R6109 Vss.n1229 Vss.n303 0.019868
R6110 Vss.n1325 Vss.n1324 0.019868
R6111 Vss.n1405 Vss.n273 0.019868
R6112 Vss.n1228 Vss.n1227 0.019868
R6113 Vss.n1725 Vss.n1724 0.0197929
R6114 Vss.n1858 Vss.n55 0.0197857
R6115 Vss.n1903 Vss.n1902 0.0197857
R6116 Vss.n1685 Vss.n1634 0.0197428
R6117 Vss.n1821 Vss.n71 0.0197428
R6118 Vss.n1423 Vss.n70 0.0197428
R6119 Vss.n1422 Vss.n1421 0.0197428
R6120 Vss.n391 Vss.n261 0.0197428
R6121 Vss.n1606 Vss.n146 0.0196349
R6122 Vss.n913 Vss.n563 0.0196349
R6123 Vss.n1155 Vss.n1154 0.0196349
R6124 Vss.n1147 Vss.n457 0.0196349
R6125 Vss.n41 Vss.n35 0.0196349
R6126 adc_PISO_0.dffrs_4.vss Vss.n1873 0.0170545
R6127 Vss.n1220 Vss.n1219 0.0164817
R6128 Vss.n1760 Vss.n112 0.0163358
R6129 Vss.n911 Vss.n910 0.0163358
R6130 Vss.n1014 Vss.n1013 0.0163358
R6131 Vss.n1492 Vss.n222 0.0163358
R6132 Vss.n1889 Vss.n28 0.0163358
R6133 Vss.n774 Vss.n600 0.0163358
R6134 Vss.n1221 Vss.n1220 0.0157888
R6135 Vss.n1221 Vss.n286 0.0157888
R6136 Vss.n1371 Vss.n286 0.0157888
R6137 Vss.n1371 Vss.n296 0.0157888
R6138 Vss.n296 Vss.n174 0.0157888
R6139 Vss.n1208 Vss.n353 0.0150091
R6140 Vss.n1620 Vss.n93 0.0142428
R6141 Vss.n1542 Vss.n92 0.014047
R6142 Vss.n1538 Vss.n186 0.014047
R6143 Vss.n1379 Vss.n1378 0.014047
R6144 Vss.n1290 Vss.n316 0.014047
R6145 Vss.n1289 Vss.n1288 0.014047
R6146 Vss.n1607 Vss.n112 0.0139604
R6147 Vss.n912 Vss.n911 0.0139604
R6148 Vss.n1014 Vss.n452 0.0139604
R6149 Vss.n1146 Vss.n222 0.0139604
R6150 Vss.n753 Vss.n28 0.0139604
R6151 Vss.n670 Vss.n600 0.0139604
R6152 Vss.n1607 Vss.n1606 0.0130367
R6153 Vss.n913 Vss.n912 0.0130367
R6154 Vss.n1154 Vss.n452 0.0130367
R6155 Vss.n1147 Vss.n1146 0.0130367
R6156 Vss.n754 Vss.n753 0.0130367
R6157 Vss.n670 Vss.n41 0.0130367
R6158 Vss.n412 Vss.n411 0.0121902
R6159 Vss.n1322 Vss.n1314 0.0121902
R6160 Vss.n1268 Vss.n1267 0.0121902
R6161 Vss.n1256 Vss.n1255 0.0121902
R6162 Vss.n1095 Vss.n1094 0.0121902
R6163 Vss.n1651 Vss.n1650 0.0121902
R6164 Vss.n484 Vss.n483 0.0121902
R6165 Vss.n1449 Vss.n185 0.0121902
R6166 Vss.n1235 Vss.n1234 0.0121902
R6167 Vss.n1586 Vss.n1585 0.0121902
R6168 Vss.n1796 Vss.n1795 0.0121902
R6169 Vss.n1518 Vss.n161 0.0121902
R6170 Vss.n1445 Vss.n1444 0.0121902
R6171 Vss.n1298 Vss.n318 0.0121902
R6172 Vss.n940 Vss.n938 0.0121902
R6173 Vss.n792 Vss.n791 0.0121902
R6174 Vss.n1169 Vss.n1168 0.0121902
R6175 Vss.n818 Vss.n816 0.0121902
R6176 Vss.n634 Vss.n633 0.0121902
R6177 Vss.n720 Vss.n719 0.0121902
R6178 Vss.n1782 adc_PISO_0.avss 0.0118245
R6179 Vss.n1601 Vss.n151 0.0110968
R6180 Vss.n1701 Vss.n1637 0.0102582
R6181 Vss.n296 Vss.n173 0.00974555
R6182 Vss.n1377 Vss.n1371 0.00974555
R6183 Vss.n1389 Vss.n286 0.00974555
R6184 Vss.n1221 Vss.n285 0.00974555
R6185 Vss.n148 Vss.n147 0.00967928
R6186 Vss.n1562 Vss.n174 0.00967038
R6187 Vss.n413 Vss.n368 0.00915761
R6188 Vss.n1092 Vss.n1090 0.00915761
R6189 Vss.n476 Vss.n474 0.00915761
R6190 Vss.n801 Vss.n800 0.00915761
R6191 Vss.n431 Vss.n429 0.00915761
R6192 Vss.n825 Vss.n824 0.00915761
R6193 Vss.n631 Vss.n629 0.00915761
R6194 Vss.n710 Vss.n708 0.00915761
R6195 Vss.n1603 Vss.n149 0.00760526
R6196 Vss.n1178 Vss.n1177 0.00745509
R6197 Vss.n1219 SARlogic_0.dffrs_11.vss 0.00734312
R6198 Vss.n1660 Vss.n1659 0.00720109
R6199 Vss.n495 Vss.n494 0.00720109
R6200 Vss.n1727 Vss.n130 0.00720109
R6201 Vss.n1042 Vss.n1041 0.00720109
R6202 Vss.n836 Vss.n835 0.00720109
R6203 Vss.n650 Vss.n649 0.00720109
R6204 Vss.n1916 Vss.n1915 0.00720109
R6205 Vss.n712 Vss.n3 0.00720109
R6206 Vss.n1196 Vss.n1194 0.00638507
R6207 Vss.n1110 Vss.n1109 0.00617391
R6208 Vss.n1111 Vss.n1110 0.00617391
R6209 Vss.n1600 Vss.n149 0.00613715
R6210 Vss.n1601 Vss.n1600 0.00613715
R6211 Vss.n1871 Vss 0.00568182
R6212 Vss.n1129 Vss.n456 0.00511663
R6213 Vss.n523 Vss.n453 0.00511663
R6214 Vss.n882 Vss.n562 0.00511663
R6215 Vss.n736 Vss.n692 0.00511663
R6216 Vss.n1874 adc_PISO_0.dffrs_4.vss 0.00480909
R6217 Vss.n915 Vss.n454 0.00478552
R6218 SARlogic_0.dffrs_7.vss Vss.n173 0.0044588
R6219 SARlogic_0.dffrs_8.vss Vss.n1377 0.0044588
R6220 Vss.n1389 SARlogic_0.dffrs_9.vss 0.0044588
R6221 SARlogic_0.dffrs_10.vss Vss.n285 0.0044588
R6222 Vss.n1563 SARlogic_0.dffrs_14.vss 0.00438363
R6223 Vss.n1861 comparator_no_offsetcal_0.x4.VSS 0.00371429
R6224 osu_sc_buf_4_flat_0.VSS Vss.n1917 0.00249115
R6225 Vss.n1602 Vss.n1601 0.00175057
R6226 Vss.n1578 Vss.n1577 0.000628205
R6227 Vss.n162 Vss.n159 0.000628205
R6228 Vss.n1726 Vss.n1725 0.000575167
R6229 Vss.n1553 Vss.n140 0.000575167
R6230 Vss.n1563 Vss.n1562 0.000575167
R6231 Vss.n1554 Vss.n174 0.000550111
R6232 Vss.n891 Vss.n890 0.000544599
R6233 Vss.n408 Vss.n407 0.000544599
R6234 Vss.n1067 Vss.n1065 0.000544599
R6235 Vss.n509 Vss.n508 0.000544599
R6236 Vss.n993 Vss.n522 0.000544599
R6237 Vss.n1192 Vss.n419 0.000544599
R6238 Vss.n663 Vss.n662 0.000544599
R6239 Vss.n703 Vss.n702 0.000544599
R6240 Vss.n1209 Vss.n1208 0.000543311
R6241 Vss.n201 Vss.n200 0.000542735
R6242 Vss.n1702 Vss.n1632 0.000525267
R6243 Vss.n1670 Vss.n1669 0.000525056
R6244 Vss.n1724 Vss.n140 0.000525056
R6245 Vss.n1363 Vss.n1362 0.000525056
R6246 Vss.n1810 Vss.n1809 0.000525056
R6247 Vss.n1431 Vss.n1430 0.000525056
R6248 Vss.n1370 Vss.n302 0.000525056
R6249 Vss.n1351 Vss.n303 0.000525056
R6250 Vss.n1325 Vss.n262 0.000525056
R6251 Vss.n1405 Vss.n1404 0.000525056
R6252 Vss.n1227 Vss.n1222 0.000525056
R6253 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t4 41.0041
R6254 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t9 40.8177
R6255 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t8 40.6313
R6256 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t7 27.3166
R6257 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t5 27.1302
R6258 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t6 26.9438
R6259 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.t0 10.0473
R6260 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n4 9.90747
R6261 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n2 9.90116
R6262 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.t1 6.51042
R6263 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.n7 6.04952
R6264 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_6.C.n1 5.7305
R6265 SARlogic_0.dffrs_12.nand3_2.B SARlogic_0.dffrs_12.nand3_6.C.n0 5.47979
R6266 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C.n3 5.13907
R6267 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n9 4.72925
R6268 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_6.C.n5 4.5005
R6269 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.n8 0.732092
R6270 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t2 0.7285
R6271 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t3 0.7285
R6272 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n6 0.449758
R6273 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_2.B 0.166901
R6274 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_0.A 0.0455
R6275 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C 0.0455
R6276 inv2_0.out.n30 inv2_0.out.t25 34.2529
R6277 inv2_0.out.n24 inv2_0.out.t8 34.2529
R6278 inv2_0.out.n18 inv2_0.out.t13 34.2529
R6279 inv2_0.out.n12 inv2_0.out.t21 34.2529
R6280 inv2_0.out.n6 inv2_0.out.t15 34.2529
R6281 inv2_0.out.n1 inv2_0.out.t28 34.2529
R6282 inv2_0.out.n32 inv2_0.out.t20 34.1797
R6283 inv2_0.out.n26 inv2_0.out.t22 34.1797
R6284 inv2_0.out.n20 inv2_0.out.t17 34.1797
R6285 inv2_0.out.n14 inv2_0.out.t5 34.1797
R6286 inv2_0.out.n8 inv2_0.out.t24 34.1797
R6287 inv2_0.out.n3 inv2_0.out.t7 34.1797
R6288 inv2_0.out.n29 inv2_0.out.t31 19.673
R6289 inv2_0.out.n23 inv2_0.out.t11 19.673
R6290 inv2_0.out.n17 inv2_0.out.t12 19.673
R6291 inv2_0.out.n11 inv2_0.out.t27 19.673
R6292 inv2_0.out.n5 inv2_0.out.t19 19.673
R6293 inv2_0.out.n0 inv2_0.out.t2 19.673
R6294 inv2_0.out.n32 inv2_0.out.t9 19.5798
R6295 inv2_0.out.n26 inv2_0.out.t14 19.5798
R6296 inv2_0.out.n20 inv2_0.out.t6 19.5798
R6297 inv2_0.out.n14 inv2_0.out.t26 19.5798
R6298 inv2_0.out.n8 inv2_0.out.t16 19.5798
R6299 inv2_0.out.n3 inv2_0.out.t30 19.5798
R6300 inv2_0.out.n29 inv2_0.out.t18 19.4007
R6301 inv2_0.out.n23 inv2_0.out.t29 19.4007
R6302 inv2_0.out.n17 inv2_0.out.t3 19.4007
R6303 inv2_0.out.n11 inv2_0.out.t10 19.4007
R6304 inv2_0.out.n5 inv2_0.out.t4 19.4007
R6305 inv2_0.out.n0 inv2_0.out.t23 19.4007
R6306 inv2_0.out.n10 inv2_0.out.n4 15.5531
R6307 inv2_0.out.n36 inv2_0.out.t0 9.6935
R6308 inv2_0.out.n34 inv2_0.out.n33 8.46371
R6309 inv2_0.out.n22 inv2_0.out.n21 8.37371
R6310 inv2_0.out.n28 inv2_0.out.n27 8.32871
R6311 inv2_0.out.n16 inv2_0.out.n15 8.32871
R6312 inv2_0.out.n10 inv2_0.out.n9 8.32871
R6313 inv2_0.out.n31 inv2_0.out.n30 7.87164
R6314 inv2_0.out.n25 inv2_0.out.n24 7.87164
R6315 inv2_0.out.n19 inv2_0.out.n18 7.87164
R6316 inv2_0.out.n13 inv2_0.out.n12 7.87164
R6317 inv2_0.out.n7 inv2_0.out.n6 7.87164
R6318 inv2_0.out.n2 inv2_0.out.n1 7.87164
R6319 inv2_0.out.n34 inv2_0.out.n28 7.26762
R6320 inv2_0.out.n16 inv2_0.out.n10 7.22491
R6321 inv2_0.out.n22 inv2_0.out.n16 7.22491
R6322 inv2_0.out.n28 inv2_0.out.n22 7.22491
R6323 inv2_0.out.n33 inv2_0.out.n32 5.00771
R6324 inv2_0.out.n21 inv2_0.out.n20 5.00771
R6325 inv2_0.out.n27 inv2_0.out.n26 4.96432
R6326 inv2_0.out.n15 inv2_0.out.n14 4.96432
R6327 inv2_0.out.n9 inv2_0.out.n8 4.96432
R6328 inv2_0.out.n4 inv2_0.out.n3 4.96432
R6329 inv2_0.out inv2_0.out.n35 4.85086
R6330 inv2_0.out.n36 inv2_0.out.t1 4.35383
R6331 inv2_0.out.n27 inv2_0.out.n25 2.11068
R6332 inv2_0.out.n15 inv2_0.out.n13 2.11068
R6333 inv2_0.out.n9 inv2_0.out.n7 2.11068
R6334 inv2_0.out.n4 inv2_0.out.n2 2.11068
R6335 inv2_0.out.n33 inv2_0.out.n31 2.06729
R6336 inv2_0.out.n21 inv2_0.out.n19 2.06729
R6337 inv2_0.out inv2_0.out.n36 0.254429
R6338 inv2_0.out.n31 adc_PISO_0.2inmux_0.Load 0.2255
R6339 inv2_0.out.n25 adc_PISO_0.2inmux_2.Load 0.2255
R6340 inv2_0.out.n19 adc_PISO_0.2inmux_3.Load 0.2255
R6341 inv2_0.out.n13 adc_PISO_0.2inmux_4.Load 0.2255
R6342 inv2_0.out.n7 adc_PISO_0.2inmux_5.Load 0.2255
R6343 inv2_0.out.n2 adc_PISO_0.2inmux_1.Load 0.2255
R6344 inv2_0.out.n35 inv2_0.out.n34 0.182025
R6345 inv2_0.out.n30 inv2_0.out.n29 0.106438
R6346 inv2_0.out.n24 inv2_0.out.n23 0.106438
R6347 inv2_0.out.n18 inv2_0.out.n17 0.106438
R6348 inv2_0.out.n12 inv2_0.out.n11 0.106438
R6349 inv2_0.out.n6 inv2_0.out.n5 0.106438
R6350 inv2_0.out.n1 inv2_0.out.n0 0.106438
R6351 inv2_0.out.n35 adc_PISO_0.load 0.0294831
R6352 a_37499_31160.n0 a_37499_31160.t5 34.1797
R6353 a_37499_31160.n0 a_37499_31160.t4 19.5798
R6354 a_37499_31160.n1 a_37499_31160.t2 18.7717
R6355 a_37499_31160.n1 a_37499_31160.t1 9.2885
R6356 a_37499_31160.n2 a_37499_31160.n0 4.93379
R6357 a_37499_31160.n3 a_37499_31160.t3 4.23346
R6358 a_37499_31160.t0 a_37499_31160.n3 3.85546
R6359 a_37499_31160.n2 a_37499_31160.n1 0.4055
R6360 a_37499_31160.n3 a_37499_31160.n2 0.352625
R6361 a_n9429_n2007.n18 a_n9429_n2007.n17 11.2899
R6362 a_n9429_n2007.n17 a_n9429_n2007.n16 8.49339
R6363 a_n9429_n2007.n10 a_n9429_n2007.n9 4.89725
R6364 a_n9429_n2007.n14 a_n9429_n2007.n2 4.89725
R6365 a_n9429_n2007.n13 a_n9429_n2007.n3 4.89725
R6366 a_n9429_n2007.n12 a_n9429_n2007.n5 4.89725
R6367 a_n9429_n2007.n11 a_n9429_n2007.n7 4.89725
R6368 a_n9429_n2007.n13 a_n9429_n2007.n4 4.88712
R6369 a_n9429_n2007.n12 a_n9429_n2007.n6 4.88712
R6370 a_n9429_n2007.n11 a_n9429_n2007.n8 4.88712
R6371 a_n9429_n2007.n1 a_n9429_n2007.n0 4.4
R6372 a_n9429_n2007.n16 a_n9429_n2007.n15 4.35275
R6373 a_n9429_n2007.n18 a_n9429_n2007.t17 2.048
R6374 a_n9429_n2007.t0 a_n9429_n2007.n18 2.048
R6375 a_n9429_n2007.n17 a_n9429_n2007.n1 1.95895
R6376 a_n9429_n2007.n9 a_n9429_n2007.t19 1.0925
R6377 a_n9429_n2007.n9 a_n9429_n2007.t11 1.0925
R6378 a_n9429_n2007.n0 a_n9429_n2007.t8 1.0925
R6379 a_n9429_n2007.n0 a_n9429_n2007.t5 1.0925
R6380 a_n9429_n2007.n2 a_n9429_n2007.t3 1.0925
R6381 a_n9429_n2007.n2 a_n9429_n2007.t7 1.0925
R6382 a_n9429_n2007.n15 a_n9429_n2007.t15 1.0925
R6383 a_n9429_n2007.n15 a_n9429_n2007.t21 1.0925
R6384 a_n9429_n2007.n3 a_n9429_n2007.t12 1.0925
R6385 a_n9429_n2007.n3 a_n9429_n2007.t20 1.0925
R6386 a_n9429_n2007.n4 a_n9429_n2007.t6 1.0925
R6387 a_n9429_n2007.n4 a_n9429_n2007.t9 1.0925
R6388 a_n9429_n2007.n5 a_n9429_n2007.t2 1.0925
R6389 a_n9429_n2007.n5 a_n9429_n2007.t16 1.0925
R6390 a_n9429_n2007.n6 a_n9429_n2007.t14 1.0925
R6391 a_n9429_n2007.n6 a_n9429_n2007.t18 1.0925
R6392 a_n9429_n2007.n7 a_n9429_n2007.t10 1.0925
R6393 a_n9429_n2007.n7 a_n9429_n2007.t1 1.0925
R6394 a_n9429_n2007.n8 a_n9429_n2007.t4 1.0925
R6395 a_n9429_n2007.n8 a_n9429_n2007.t13 1.0925
R6396 a_n9429_n2007.n14 a_n9429_n2007.n13 0.849071
R6397 a_n9429_n2007.n13 a_n9429_n2007.n12 0.849071
R6398 a_n9429_n2007.n12 a_n9429_n2007.n11 0.849071
R6399 a_n9429_n2007.n11 a_n9429_n2007.n10 0.849071
R6400 a_n9429_n2007.n16 a_n9429_n2007.n14 0.534875
R6401 a_n9429_n2007.n10 a_n9429_n2007.n1 0.487625
R6402 SARlogic_0.d1.n3 SARlogic_0.d1.t9 41.0041
R6403 SARlogic_0.d1.n4 SARlogic_0.d1.t7 40.8177
R6404 SARlogic_0.d1.n7 SARlogic_0.d1.t8 40.6313
R6405 SARlogic_0.d1.n1 SARlogic_0.d1.t4 34.2529
R6406 SARlogic_0.d1.n6 SARlogic_0.dffrs_9.clk 33.8765
R6407 SARlogic_0.d1.n7 SARlogic_0.d1.t5 27.3166
R6408 SARlogic_0.d1.n4 SARlogic_0.d1.t12 27.1302
R6409 SARlogic_0.d1.n3 SARlogic_0.d1.t11 26.9438
R6410 SARlogic_0.d1 adc_PISO_0.B2 26.2596
R6411 SARlogic_0.d1.n0 SARlogic_0.d1.t6 19.673
R6412 SARlogic_0.d1.n0 SARlogic_0.d1.t10 19.4007
R6413 SARlogic_0.d1.n9 SARlogic_0.d1.n8 14.0582
R6414 SARlogic_0.d1.n9 SARlogic_0.d1.n6 11.729
R6415 SARlogic_0.d1.n12 SARlogic_0.d1.t1 10.0473
R6416 SARlogic_0.d1.n2 SARlogic_0.d1.n1 8.05164
R6417 SARlogic_0.d1.n11 SARlogic_0.d1.t0 6.51042
R6418 SARlogic_0.d1.n11 SARlogic_0.d1.n10 6.04952
R6419 SARlogic_0.dffrs_9.nand3_1.A SARlogic_0.d1.n3 5.7755
R6420 SARlogic_0.dffrs_9.nand3_6.B SARlogic_0.d1.n4 5.47979
R6421 SARlogic_0.d1.n8 SARlogic_0.d1.n7 5.13907
R6422 SARlogic_0.dffrs_10.nand3_2.Z SARlogic_0.d1.n12 4.72925
R6423 SARlogic_0.d1.n5 SARlogic_0.dffrs_9.nand3_6.B 2.17818
R6424 adc_PISO_0.B2 SARlogic_0.d1.n2 1.87121
R6425 SARlogic_0.d1.n5 SARlogic_0.dffrs_9.nand3_1.A 1.34729
R6426 SARlogic_0.d1.n6 SARlogic_0.d1 0.985679
R6427 SARlogic_0.d1.n12 SARlogic_0.d1.n11 0.732092
R6428 SARlogic_0.d1.n10 SARlogic_0.d1.t3 0.7285
R6429 SARlogic_0.d1.n10 SARlogic_0.d1.t2 0.7285
R6430 SARlogic_0.dffrs_9.clk SARlogic_0.d1.n5 0.610571
R6431 SARlogic_0.dffrs_10.nand3_2.Z SARlogic_0.d1.n9 0.166901
R6432 SARlogic_0.d1.n1 SARlogic_0.d1.n0 0.106438
R6433 SARlogic_0.d1.n8 SARlogic_0.dffrs_10.nand3_7.C 0.0455
R6434 SARlogic_0.d1.n2 adc_PISO_0.2inmux_5.In 0.0455
R6435 a_28027_28820.n0 a_28027_28820.t5 34.1797
R6436 a_28027_28820.n0 a_28027_28820.t4 19.5798
R6437 a_28027_28820.n1 a_28027_28820.t2 18.7717
R6438 a_28027_28820.n1 a_28027_28820.t1 9.2885
R6439 a_28027_28820.n2 a_28027_28820.n0 4.93379
R6440 a_28027_28820.t0 a_28027_28820.n3 4.23346
R6441 a_28027_28820.n3 a_28027_28820.t3 3.85546
R6442 a_28027_28820.n2 a_28027_28820.n1 0.4055
R6443 a_28027_28820.n3 a_28027_28820.n2 0.352625
R6444 Reset.n80 Reset.t25 41.0041
R6445 Reset.n86 Reset.t52 41.0041
R6446 Reset.n66 Reset.t59 41.0041
R6447 Reset.n72 Reset.t1 41.0041
R6448 Reset.n52 Reset.t39 41.0041
R6449 Reset.n58 Reset.t66 41.0041
R6450 Reset.n38 Reset.t48 41.0041
R6451 Reset.n44 Reset.t72 41.0041
R6452 Reset.n24 Reset.t36 41.0041
R6453 Reset.n30 Reset.t64 41.0041
R6454 Reset.n10 Reset.t65 41.0041
R6455 Reset.n16 Reset.t7 41.0041
R6456 Reset.n4 Reset.t38 41.0041
R6457 Reset.n83 Reset.t10 40.8177
R6458 Reset.n82 Reset.t0 40.8177
R6459 Reset.n89 Reset.t26 40.8177
R6460 Reset.n88 Reset.t29 40.8177
R6461 Reset.n69 Reset.t37 40.8177
R6462 Reset.n68 Reset.t28 40.8177
R6463 Reset.n75 Reset.t54 40.8177
R6464 Reset.n74 Reset.t57 40.8177
R6465 Reset.n55 Reset.t30 40.8177
R6466 Reset.n54 Reset.t20 40.8177
R6467 Reset.n61 Reset.t75 40.8177
R6468 Reset.n60 Reset.t51 40.8177
R6469 Reset.n41 Reset.t58 40.8177
R6470 Reset.n40 Reset.t53 40.8177
R6471 Reset.n47 Reset.t42 40.8177
R6472 Reset.n46 Reset.t77 40.8177
R6473 Reset.n27 Reset.t2 40.8177
R6474 Reset.n26 Reset.t78 40.8177
R6475 Reset.n33 Reset.t34 40.8177
R6476 Reset.n32 Reset.t24 40.8177
R6477 Reset.n13 Reset.t76 40.8177
R6478 Reset.n12 Reset.t68 40.8177
R6479 Reset.n19 Reset.t73 40.8177
R6480 Reset.n18 Reset.t13 40.8177
R6481 Reset.n7 Reset.t21 40.8177
R6482 Reset.n6 Reset.t14 40.8177
R6483 Reset.n2 Reset.t63 40.6313
R6484 Reset.n0 Reset.t62 40.6313
R6485 Reset.n2 Reset.t23 27.3166
R6486 Reset.n0 Reset.t79 27.3166
R6487 Reset.n83 Reset.t35 27.1302
R6488 Reset.n82 Reset.t22 27.1302
R6489 Reset.n89 Reset.t45 27.1302
R6490 Reset.n88 Reset.t50 27.1302
R6491 Reset.n69 Reset.t61 27.1302
R6492 Reset.n68 Reset.t49 27.1302
R6493 Reset.n75 Reset.t70 27.1302
R6494 Reset.n74 Reset.t74 27.1302
R6495 Reset.n55 Reset.t55 27.1302
R6496 Reset.n54 Reset.t43 27.1302
R6497 Reset.n61 Reset.t11 27.1302
R6498 Reset.n60 Reset.t67 27.1302
R6499 Reset.n41 Reset.t80 27.1302
R6500 Reset.n40 Reset.t69 27.1302
R6501 Reset.n47 Reset.t60 27.1302
R6502 Reset.n46 Reset.t16 27.1302
R6503 Reset.n27 Reset.t27 27.1302
R6504 Reset.n26 Reset.t17 27.1302
R6505 Reset.n33 Reset.t56 27.1302
R6506 Reset.n32 Reset.t44 27.1302
R6507 Reset.n13 Reset.t18 27.1302
R6508 Reset.n12 Reset.t3 27.1302
R6509 Reset.n19 Reset.t8 27.1302
R6510 Reset.n18 Reset.t31 27.1302
R6511 Reset.n7 Reset.t47 27.1302
R6512 Reset.n6 Reset.t32 27.1302
R6513 Reset.n80 Reset.t81 26.9438
R6514 Reset.n86 Reset.t6 26.9438
R6515 Reset.n66 Reset.t33 26.9438
R6516 Reset.n72 Reset.t5 26.9438
R6517 Reset.n52 Reset.t15 26.9438
R6518 Reset.n58 Reset.t71 26.9438
R6519 Reset.n38 Reset.t19 26.9438
R6520 Reset.n44 Reset.t4 26.9438
R6521 Reset.n24 Reset.t9 26.9438
R6522 Reset.n30 Reset.t46 26.9438
R6523 Reset.n10 Reset.t41 26.9438
R6524 Reset.n16 Reset.t40 26.9438
R6525 Reset.n4 Reset.t12 26.9438
R6526 Reset.n78 SARlogic_0.dffrs_1.resetb 19.0901
R6527 Reset.n64 SARlogic_0.dffrs_2.resetb 19.0901
R6528 Reset.n50 SARlogic_0.dffrs_3.resetb 19.0901
R6529 Reset.n36 SARlogic_0.dffrs_4.resetb 19.0901
R6530 Reset.n22 SARlogic_0.dffrs_5.resetb 19.0901
R6531 Reset.n92 SARlogic_0.dffrs_0.resetb 19.0467
R6532 Reset.n23 SARlogic_0.dffrs_12.resetb 14.0622
R6533 Reset.n84 SARlogic_0.dffrs_14.nand3_1.B 12.1571
R6534 Reset.n90 SARlogic_0.dffrs_0.nand3_1.B 12.1571
R6535 Reset.n70 SARlogic_0.dffrs_7.nand3_1.B 12.1571
R6536 Reset.n76 SARlogic_0.dffrs_1.nand3_1.B 12.1571
R6537 Reset.n56 SARlogic_0.dffrs_8.nand3_1.B 12.1571
R6538 Reset.n62 SARlogic_0.dffrs_2.nand3_1.B 12.1571
R6539 Reset.n42 SARlogic_0.dffrs_9.nand3_1.B 12.1571
R6540 Reset.n48 SARlogic_0.dffrs_3.nand3_1.B 12.1571
R6541 Reset.n28 SARlogic_0.dffrs_10.nand3_1.B 12.1571
R6542 Reset.n34 SARlogic_0.dffrs_4.nand3_1.B 12.1571
R6543 Reset.n14 SARlogic_0.dffrs_11.nand3_1.B 12.1571
R6544 Reset.n20 SARlogic_0.dffrs_5.nand3_1.B 12.1571
R6545 Reset.n8 SARlogic_0.dffrs_12.nand3_1.B 12.1571
R6546 Reset.n3 Reset.n1 9.22229
R6547 Reset.n94 Reset.n93 7.9889
R6548 Reset.n85 Reset.n81 7.75389
R6549 Reset.n91 Reset.n87 7.75389
R6550 Reset.n71 Reset.n67 7.75389
R6551 Reset.n77 Reset.n73 7.75389
R6552 Reset.n57 Reset.n53 7.75389
R6553 Reset.n63 Reset.n59 7.75389
R6554 Reset.n43 Reset.n39 7.75389
R6555 Reset.n49 Reset.n45 7.75389
R6556 Reset.n29 Reset.n25 7.75389
R6557 Reset.n35 Reset.n31 7.75389
R6558 Reset.n15 Reset.n11 7.75389
R6559 Reset.n21 Reset.n17 7.75389
R6560 Reset.n9 Reset.n5 7.75389
R6561 Reset.n94 SARlogic_0.dffrs_13.setb 6.43164
R6562 Reset.n85 Reset.n84 5.93546
R6563 Reset.n91 Reset.n90 5.93546
R6564 Reset.n71 Reset.n70 5.93546
R6565 Reset.n77 Reset.n76 5.93546
R6566 Reset.n57 Reset.n56 5.93546
R6567 Reset.n63 Reset.n62 5.93546
R6568 Reset.n43 Reset.n42 5.93546
R6569 Reset.n49 Reset.n48 5.93546
R6570 Reset.n29 Reset.n28 5.93546
R6571 Reset.n35 Reset.n34 5.93546
R6572 Reset.n15 Reset.n14 5.93546
R6573 Reset.n21 Reset.n20 5.93546
R6574 Reset.n9 Reset.n8 5.93546
R6575 Reset.n78 SARlogic_0.dffrs_7.resetb 5.93246
R6576 Reset.n64 SARlogic_0.dffrs_8.resetb 5.93246
R6577 Reset.n50 SARlogic_0.dffrs_9.resetb 5.93246
R6578 Reset.n36 SARlogic_0.dffrs_10.resetb 5.93246
R6579 Reset.n22 SARlogic_0.dffrs_11.resetb 5.93246
R6580 Reset.n92 SARlogic_0.dffrs_14.resetb 5.88425
R6581 Reset.n81 Reset.n80 5.7305
R6582 Reset.n87 Reset.n86 5.7305
R6583 Reset.n67 Reset.n66 5.7305
R6584 Reset.n73 Reset.n72 5.7305
R6585 Reset.n53 Reset.n52 5.7305
R6586 Reset.n59 Reset.n58 5.7305
R6587 Reset.n39 Reset.n38 5.7305
R6588 Reset.n45 Reset.n44 5.7305
R6589 Reset.n25 Reset.n24 5.7305
R6590 Reset.n31 Reset.n30 5.7305
R6591 Reset.n11 Reset.n10 5.7305
R6592 Reset.n17 Reset.n16 5.7305
R6593 Reset.n5 Reset.n4 5.7305
R6594 SARlogic_0.dffrs_14.nand3_8.B Reset.n83 5.47979
R6595 SARlogic_0.dffrs_14.nand3_1.B Reset.n82 5.47979
R6596 SARlogic_0.dffrs_0.nand3_8.B Reset.n89 5.47979
R6597 SARlogic_0.dffrs_0.nand3_1.B Reset.n88 5.47979
R6598 SARlogic_0.dffrs_7.nand3_8.B Reset.n69 5.47979
R6599 SARlogic_0.dffrs_7.nand3_1.B Reset.n68 5.47979
R6600 SARlogic_0.dffrs_1.nand3_8.B Reset.n75 5.47979
R6601 SARlogic_0.dffrs_1.nand3_1.B Reset.n74 5.47979
R6602 SARlogic_0.dffrs_8.nand3_8.B Reset.n55 5.47979
R6603 SARlogic_0.dffrs_8.nand3_1.B Reset.n54 5.47979
R6604 SARlogic_0.dffrs_2.nand3_8.B Reset.n61 5.47979
R6605 SARlogic_0.dffrs_2.nand3_1.B Reset.n60 5.47979
R6606 SARlogic_0.dffrs_9.nand3_8.B Reset.n41 5.47979
R6607 SARlogic_0.dffrs_9.nand3_1.B Reset.n40 5.47979
R6608 SARlogic_0.dffrs_3.nand3_8.B Reset.n47 5.47979
R6609 SARlogic_0.dffrs_3.nand3_1.B Reset.n46 5.47979
R6610 SARlogic_0.dffrs_10.nand3_8.B Reset.n27 5.47979
R6611 SARlogic_0.dffrs_10.nand3_1.B Reset.n26 5.47979
R6612 SARlogic_0.dffrs_4.nand3_8.B Reset.n33 5.47979
R6613 SARlogic_0.dffrs_4.nand3_1.B Reset.n32 5.47979
R6614 SARlogic_0.dffrs_11.nand3_8.B Reset.n13 5.47979
R6615 SARlogic_0.dffrs_11.nand3_1.B Reset.n12 5.47979
R6616 SARlogic_0.dffrs_5.nand3_8.B Reset.n19 5.47979
R6617 SARlogic_0.dffrs_5.nand3_1.B Reset.n18 5.47979
R6618 SARlogic_0.dffrs_12.nand3_8.B Reset.n7 5.47979
R6619 SARlogic_0.dffrs_12.nand3_1.B Reset.n6 5.47979
R6620 Reset.n3 Reset.n2 5.14711
R6621 Reset.n1 Reset.n0 5.13907
R6622 Reset.n84 SARlogic_0.dffrs_14.nand3_8.B 5.09593
R6623 Reset.n90 SARlogic_0.dffrs_0.nand3_8.B 5.09593
R6624 Reset.n70 SARlogic_0.dffrs_7.nand3_8.B 5.09593
R6625 Reset.n76 SARlogic_0.dffrs_1.nand3_8.B 5.09593
R6626 Reset.n56 SARlogic_0.dffrs_8.nand3_8.B 5.09593
R6627 Reset.n62 SARlogic_0.dffrs_2.nand3_8.B 5.09593
R6628 Reset.n42 SARlogic_0.dffrs_9.nand3_8.B 5.09593
R6629 Reset.n48 SARlogic_0.dffrs_3.nand3_8.B 5.09593
R6630 Reset.n28 SARlogic_0.dffrs_10.nand3_8.B 5.09593
R6631 Reset.n34 SARlogic_0.dffrs_4.nand3_8.B 5.09593
R6632 Reset.n14 SARlogic_0.dffrs_11.nand3_8.B 5.09593
R6633 Reset.n20 SARlogic_0.dffrs_5.nand3_8.B 5.09593
R6634 Reset.n8 SARlogic_0.dffrs_12.nand3_8.B 5.09593
R6635 Reset.n23 Reset.n22 4.5005
R6636 Reset.n37 Reset.n36 4.5005
R6637 Reset.n51 Reset.n50 4.5005
R6638 Reset.n65 Reset.n64 4.5005
R6639 Reset.n79 Reset.n78 4.5005
R6640 Reset.n93 Reset.n92 4.5005
R6641 Reset.n37 Reset.n23 3.6383
R6642 Reset.n51 Reset.n37 3.6383
R6643 Reset.n65 Reset.n51 3.6383
R6644 Reset.n79 Reset.n65 3.6383
R6645 Reset.n93 Reset.n79 3.6113
R6646 SARlogic_0.dffrs_13.setb SARlogic_0.dffrs_13.nand3_0.C 0.783821
R6647 SARlogic_0.reset Reset 0.18425
R6648 SARlogic_0.reset Reset.n94 0.13775
R6649 SARlogic_0.dffrs_14.resetb Reset.n85 0.136036
R6650 SARlogic_0.dffrs_0.resetb Reset.n91 0.136036
R6651 SARlogic_0.dffrs_7.resetb Reset.n71 0.136036
R6652 SARlogic_0.dffrs_1.resetb Reset.n77 0.136036
R6653 SARlogic_0.dffrs_8.resetb Reset.n57 0.136036
R6654 SARlogic_0.dffrs_2.resetb Reset.n63 0.136036
R6655 SARlogic_0.dffrs_9.resetb Reset.n43 0.136036
R6656 SARlogic_0.dffrs_3.resetb Reset.n49 0.136036
R6657 SARlogic_0.dffrs_10.resetb Reset.n29 0.136036
R6658 SARlogic_0.dffrs_4.resetb Reset.n35 0.136036
R6659 SARlogic_0.dffrs_11.resetb Reset.n15 0.136036
R6660 SARlogic_0.dffrs_5.resetb Reset.n21 0.136036
R6661 SARlogic_0.dffrs_12.resetb Reset.n9 0.136036
R6662 Reset.n1 SARlogic_0.dffrs_13.nand3_2.C 0.0455
R6663 Reset.n81 SARlogic_0.dffrs_14.nand3_7.A 0.0455
R6664 Reset.n87 SARlogic_0.dffrs_0.nand3_7.A 0.0455
R6665 Reset.n67 SARlogic_0.dffrs_7.nand3_7.A 0.0455
R6666 Reset.n73 SARlogic_0.dffrs_1.nand3_7.A 0.0455
R6667 Reset.n53 SARlogic_0.dffrs_8.nand3_7.A 0.0455
R6668 Reset.n59 SARlogic_0.dffrs_2.nand3_7.A 0.0455
R6669 Reset.n39 SARlogic_0.dffrs_9.nand3_7.A 0.0455
R6670 Reset.n45 SARlogic_0.dffrs_3.nand3_7.A 0.0455
R6671 Reset.n25 SARlogic_0.dffrs_10.nand3_7.A 0.0455
R6672 Reset.n31 SARlogic_0.dffrs_4.nand3_7.A 0.0455
R6673 Reset.n11 SARlogic_0.dffrs_11.nand3_7.A 0.0455
R6674 Reset.n17 SARlogic_0.dffrs_5.nand3_7.A 0.0455
R6675 Reset.n5 SARlogic_0.dffrs_12.nand3_7.A 0.0455
R6676 SARlogic_0.dffrs_13.nand3_0.C Reset.n3 0.0374643
R6677 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t5 41.0041
R6678 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t4 40.8177
R6679 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t9 40.6313
R6680 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t8 27.3166
R6681 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t6 27.1302
R6682 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t7 26.9438
R6683 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.t3 10.0473
R6684 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n4 9.90747
R6685 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n2 9.90116
R6686 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.t0 6.51042
R6687 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.n7 6.04952
R6688 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_6.C.n1 5.7305
R6689 SARlogic_0.dffrs_14.nand3_2.B SARlogic_0.dffrs_14.nand3_6.C.n0 5.47979
R6690 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C.n3 5.13907
R6691 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n9 4.72925
R6692 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_6.C.n5 4.5005
R6693 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.n8 0.732092
R6694 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t1 0.7285
R6695 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t2 0.7285
R6696 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n6 0.449758
R6697 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_2.B 0.166901
R6698 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_0.A 0.0455
R6699 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C 0.0455
R6700 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t8 41.0041
R6701 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t7 40.8177
R6702 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t6 40.6313
R6703 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t5 27.3166
R6704 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t9 27.1302
R6705 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t4 26.9438
R6706 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.t1 10.0473
R6707 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n4 9.90747
R6708 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n2 9.90116
R6709 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.t0 6.51042
R6710 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.n7 6.04952
R6711 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_6.C.n1 5.7305
R6712 SARlogic_0.dffrs_2.nand3_2.B SARlogic_0.dffrs_2.nand3_6.C.n0 5.47979
R6713 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C.n3 5.13907
R6714 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n9 4.72925
R6715 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_6.C.n5 4.5005
R6716 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.n8 0.732092
R6717 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t3 0.7285
R6718 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t2 0.7285
R6719 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n6 0.449758
R6720 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_2.B 0.166901
R6721 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_0.A 0.0455
R6722 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C 0.0455
R6723 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t4 40.6313
R6724 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t5 27.3166
R6725 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n1 14.2854
R6726 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.t1 10.0473
R6727 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.t2 6.51042
R6728 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.n2 6.04952
R6729 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C.n0 5.13907
R6730 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n4 4.72925
R6731 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.n3 0.732092
R6732 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t0 0.7285
R6733 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t3 0.7285
R6734 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C 0.0455
R6735 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t8 41.0041
R6736 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t5 40.6313
R6737 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t4 40.6313
R6738 SARlogic_0.dffrs_1.Qb SARlogic_0.dffrs_8.setb 28.021
R6739 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t7 27.3166
R6740 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t6 27.3166
R6741 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t9 26.9438
R6742 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.t1 10.0473
R6743 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb.n1 9.84255
R6744 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n3 9.22229
R6745 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.t2 6.51042
R6746 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.n7 6.04952
R6747 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.Qb.n0 5.7305
R6748 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n4 5.14711
R6749 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_1.Qb.n2 5.13907
R6750 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n6 4.94976
R6751 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n9 4.72925
R6752 SARlogic_0.dffrs_8.setb SARlogic_0.dffrs_8.nand3_0.C 0.784786
R6753 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.n8 0.732092
R6754 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t3 0.7285
R6755 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t0 0.7285
R6756 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb 0.175225
R6757 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.nand3_2.A 0.0455
R6758 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_8.nand3_2.C 0.0455
R6759 SARlogic_0.dffrs_8.nand3_0.C SARlogic_0.dffrs_1.Qb.n5 0.0374643
R6760 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t6 41.0041
R6761 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t5 40.8177
R6762 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t7 27.1302
R6763 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t4 26.9438
R6764 SARlogic_0.dffrs_4.nand3_6.A SARlogic_0.dffrs_4.nand3_0.B 17.0041
R6765 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n2 14.8493
R6766 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.t2 10.0473
R6767 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.t3 6.51042
R6768 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.n3 6.04952
R6769 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_8.Z.n0 5.7305
R6770 SARlogic_0.dffrs_4.nand3_0.B SARlogic_0.dffrs_4.nand3_8.Z.n1 5.47979
R6771 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n5 4.72925
R6772 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.n4 0.732092
R6773 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t0 0.7285
R6774 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t1 0.7285
R6775 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_6.A 0.0455
R6776 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t7 40.8177
R6777 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t5 40.6313
R6778 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t6 27.3166
R6779 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t4 27.1302
R6780 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_8.C.n2 14.119
R6781 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.t2 10.0473
R6782 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.t3 6.51042
R6783 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.n4 6.04952
R6784 SARlogic_0.dffrs_4.nand3_7.B SARlogic_0.dffrs_4.nand3_8.C.n0 5.47979
R6785 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C.n1 5.13907
R6786 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n6 4.72925
R6787 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.n5 0.732092
R6788 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t0 0.7285
R6789 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t1 0.7285
R6790 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_7.B 0.438233
R6791 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n3 0.166901
R6792 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C 0.0455
R6793 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t4 40.8177
R6794 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t6 40.6313
R6795 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t7 27.3166
R6796 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t5 27.1302
R6797 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_8.C.n2 14.119
R6798 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.t0 10.0473
R6799 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.t3 6.51042
R6800 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.n4 6.04952
R6801 SARlogic_0.dffrs_1.nand3_7.B SARlogic_0.dffrs_1.nand3_8.C.n0 5.47979
R6802 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C.n1 5.13907
R6803 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n6 4.72925
R6804 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.n5 0.732092
R6805 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t1 0.7285
R6806 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t2 0.7285
R6807 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_7.B 0.438233
R6808 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n3 0.166901
R6809 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C 0.0455
R6810 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t6 40.8177
R6811 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t7 40.6313
R6812 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t4 27.3166
R6813 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t5 27.1302
R6814 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_8.C.n2 14.119
R6815 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.t1 10.0473
R6816 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.t2 6.51042
R6817 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.n4 6.04952
R6818 SARlogic_0.dffrs_5.nand3_7.B SARlogic_0.dffrs_5.nand3_8.C.n0 5.47979
R6819 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C.n1 5.13907
R6820 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n6 4.72925
R6821 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.n5 0.732092
R6822 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t0 0.7285
R6823 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t3 0.7285
R6824 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_7.B 0.438233
R6825 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n3 0.166901
R6826 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C 0.0455
R6827 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t4 41.0041
R6828 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t7 40.8177
R6829 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t6 27.1302
R6830 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t5 26.9438
R6831 SARlogic_0.dffrs_3.nand3_6.A SARlogic_0.dffrs_3.nand3_0.B 17.0041
R6832 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n2 14.8493
R6833 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.t1 10.0473
R6834 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.t2 6.51042
R6835 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.n3 6.04952
R6836 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_8.Z.n0 5.7305
R6837 SARlogic_0.dffrs_3.nand3_0.B SARlogic_0.dffrs_3.nand3_8.Z.n1 5.47979
R6838 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n5 4.72925
R6839 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.n4 0.732092
R6840 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t0 0.7285
R6841 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t3 0.7285
R6842 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_6.A 0.0455
R6843 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t7 40.8177
R6844 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t5 40.6313
R6845 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t6 27.3166
R6846 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t4 27.1302
R6847 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_8.C.n2 14.119
R6848 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.t3 10.0473
R6849 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.t2 6.51042
R6850 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.n4 6.04952
R6851 SARlogic_0.dffrs_3.nand3_7.B SARlogic_0.dffrs_3.nand3_8.C.n0 5.47979
R6852 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C.n1 5.13907
R6853 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n6 4.72925
R6854 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.n5 0.732092
R6855 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t0 0.7285
R6856 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t1 0.7285
R6857 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_7.B 0.438233
R6858 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n3 0.166901
R6859 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C 0.0455
R6860 a_33257_31423.n3 a_33257_31423.t5 41.0041
R6861 a_33257_31423.n2 a_33257_31423.t6 40.8177
R6862 a_33257_31423.n4 a_33257_31423.t9 40.6313
R6863 a_33257_31423.n4 a_33257_31423.t4 27.3166
R6864 a_33257_31423.n2 a_33257_31423.t8 27.1302
R6865 a_33257_31423.n3 a_33257_31423.t7 26.9438
R6866 a_33257_31423.n5 a_33257_31423.n3 15.6312
R6867 a_33257_31423.n5 a_33257_31423.n4 15.046
R6868 a_33257_31423.t0 a_33257_31423.n7 10.0473
R6869 a_33257_31423.n1 a_33257_31423.t3 6.51042
R6870 a_33257_31423.n1 a_33257_31423.n0 6.04952
R6871 a_33257_31423.n6 a_33257_31423.n2 5.64619
R6872 a_33257_31423.n7 a_33257_31423.n6 5.17851
R6873 a_33257_31423.n6 a_33257_31423.n5 4.5005
R6874 a_33257_31423.n7 a_33257_31423.n1 0.732092
R6875 a_33257_31423.n0 a_33257_31423.t1 0.7285
R6876 a_33257_31423.n0 a_33257_31423.t2 0.7285
R6877 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t8 41.0041
R6878 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t7 40.8177
R6879 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t4 40.6313
R6880 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t5 27.3166
R6881 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t9 27.1302
R6882 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t6 26.9438
R6883 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.t1 10.0473
R6884 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n4 9.90747
R6885 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n2 9.90116
R6886 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.t0 6.51042
R6887 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.n7 6.04952
R6888 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_6.C.n1 5.7305
R6889 SARlogic_0.dffrs_5.nand3_2.B SARlogic_0.dffrs_5.nand3_6.C.n0 5.47979
R6890 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C.n3 5.13907
R6891 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n9 4.72925
R6892 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_6.C.n5 4.5005
R6893 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.n8 0.732092
R6894 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t2 0.7285
R6895 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t3 0.7285
R6896 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n6 0.449758
R6897 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_2.B 0.166901
R6898 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_0.A 0.0455
R6899 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C 0.0455
R6900 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t6 40.8177
R6901 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t5 40.6313
R6902 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t7 27.3166
R6903 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t4 27.1302
R6904 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_8.C.n2 14.119
R6905 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.t0 10.0473
R6906 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.t1 6.51042
R6907 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.n4 6.04952
R6908 SARlogic_0.dffrs_12.nand3_7.B SARlogic_0.dffrs_12.nand3_8.C.n0 5.47979
R6909 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C.n1 5.13907
R6910 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n6 4.72925
R6911 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.n5 0.732092
R6912 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t3 0.7285
R6913 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t2 0.7285
R6914 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_7.B 0.438233
R6915 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n3 0.166901
R6916 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C 0.0455
R6917 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t16 49.7997
R6918 comparator_no_offsetcal_0.x3.in comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t11 31.5367
R6919 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t9 19.735
R6920 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 18.0852
R6921 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t0 16.9998
R6922 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 14.5537
R6923 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 14.2885
R6924 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t17 13.6729
R6925 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t12 13.3844
R6926 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t14 13.3445
R6927 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 11.24
R6928 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 7.16477
R6929 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 6.95627
R6930 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 6.75194
R6931 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 6.32624
R6932 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t10 5.04666
R6933 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t13 4.84137
R6934 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 2.836
R6935 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 2.75432
R6936 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t1 1.8205
R6937 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t2 1.8205
R6938 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t4 1.8205
R6939 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t7 1.8205
R6940 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t6 0.8195
R6941 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t3 0.8195
R6942 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t8 0.8195
R6943 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t5 0.8195
R6944 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 0.733357
R6945 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 0.440894
R6946 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 0.426875
R6947 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 0.289009
R6948 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 0.0607115
R6949 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 comparator_no_offsetcal_0.x3.in 0.014
R6950 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t16 49.7997
R6951 comparator_no_offsetcal_0.x5.in comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t12 31.5367
R6952 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t10 19.735
R6953 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 18.9075
R6954 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t0 16.9998
R6955 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t14 13.6729
R6956 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t11 13.3844
R6957 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t17 13.3445
R6958 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 12.247
R6959 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 11.2403
R6960 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 9.4181
R6961 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 7.4449
R6962 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 6.95074
R6963 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 6.75194
R6964 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 6.32761
R6965 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t15 5.04666
R6966 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 4.94262
R6967 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t13 4.84137
R6968 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 2.836
R6969 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 2.75432
R6970 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t7 1.8205
R6971 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t6 1.8205
R6972 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t8 1.8205
R6973 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t5 1.8205
R6974 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t4 0.8195
R6975 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t1 0.8195
R6976 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t2 0.8195
R6977 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t3 0.8195
R6978 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 0.733357
R6979 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 0.5315
R6980 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 0.289009
R6981 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 0.184462
R6982 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 comparator_no_offsetcal_0.x5.in 0.014
R6983 Clk.n0 Clk.t23 41.0041
R6984 Clk.n22 Clk.t5 41.0041
R6985 Clk.n18 Clk.t24 41.0041
R6986 Clk.n14 Clk.t14 41.0041
R6987 Clk.n10 Clk.t1 41.0041
R6988 Clk.n6 Clk.t10 41.0041
R6989 Clk.n3 Clk.t28 41.0041
R6990 Clk.n1 Clk.t25 40.8177
R6991 Clk.n23 Clk.t8 40.8177
R6992 Clk.n19 Clk.t20 40.8177
R6993 Clk.n15 Clk.t17 40.8177
R6994 Clk.n11 Clk.t29 40.8177
R6995 Clk.n7 Clk.t6 40.8177
R6996 Clk.n4 Clk.t2 40.8177
R6997 Clk.n1 Clk.t19 27.1302
R6998 Clk.n23 Clk.t26 27.1302
R6999 Clk.n19 Clk.t4 27.1302
R7000 Clk.n15 Clk.t15 27.1302
R7001 Clk.n11 Clk.t32 27.1302
R7002 Clk.n7 Clk.t30 27.1302
R7003 Clk.n4 Clk.t13 27.1302
R7004 Clk.n0 Clk.t31 26.9438
R7005 Clk.n22 Clk.t16 26.9438
R7006 Clk.n18 Clk.t0 26.9438
R7007 Clk.n14 Clk.t21 26.9438
R7008 Clk.n10 Clk.t7 26.9438
R7009 Clk.n6 Clk.t18 26.9438
R7010 Clk.n3 Clk.t3 26.9438
R7011 Clk.n31 Clk.t12 21.1483
R7012 Clk.n30 Clk.t11 21.1483
R7013 Clk.n29 Clk.t22 21.1483
R7014 Clk.n28 Clk.t9 21.1483
R7015 Clk.n27 Clk.t27 20.5929
R7016 Clk.n9 SARlogic_0.dffrs_5.clk 20.5278
R7017 Clk.n28 Clk.n27 19.1491
R7018 Clk.n21 SARlogic_0.dffrs_1.clk 16.89
R7019 Clk.n17 SARlogic_0.dffrs_2.clk 16.89
R7020 Clk.n13 SARlogic_0.dffrs_3.clk 16.89
R7021 Clk.n9 SARlogic_0.dffrs_4.clk 16.89
R7022 Clk.n25 SARlogic_0.dffrs_0.clk 16.8417
R7023 Clk.n32 Clk.n31 15.5861
R7024 Clk.n26 SARlogic_0.dffrs_13.clk 12.2453
R7025 SARlogic_0.clk Clk.n33 11.0885
R7026 Clk.n26 Clk.n25 8.1113
R7027 SARlogic_0.dffrs_13.nand3_1.A Clk.n0 5.7755
R7028 SARlogic_0.dffrs_0.nand3_1.A Clk.n22 5.7755
R7029 SARlogic_0.dffrs_1.nand3_1.A Clk.n18 5.7755
R7030 SARlogic_0.dffrs_2.nand3_1.A Clk.n14 5.7755
R7031 SARlogic_0.dffrs_3.nand3_1.A Clk.n10 5.7755
R7032 SARlogic_0.dffrs_4.nand3_1.A Clk.n6 5.7755
R7033 SARlogic_0.dffrs_5.nand3_1.A Clk.n3 5.7755
R7034 SARlogic_0.dffrs_13.nand3_6.B Clk.n1 5.47979
R7035 SARlogic_0.dffrs_0.nand3_6.B Clk.n23 5.47979
R7036 SARlogic_0.dffrs_1.nand3_6.B Clk.n19 5.47979
R7037 SARlogic_0.dffrs_2.nand3_6.B Clk.n15 5.47979
R7038 SARlogic_0.dffrs_3.nand3_6.B Clk.n11 5.47979
R7039 SARlogic_0.dffrs_4.nand3_6.B Clk.n7 5.47979
R7040 SARlogic_0.dffrs_5.nand3_6.B Clk.n4 5.47979
R7041 Clk.n33 comparator_no_offsetcal_0.CLK 5.11456
R7042 Clk.n30 Clk.n29 4.47208
R7043 Clk.n13 Clk.n9 3.6383
R7044 Clk.n17 Clk.n13 3.6383
R7045 Clk.n21 Clk.n17 3.6383
R7046 Clk.n25 Clk.n21 3.6113
R7047 Clk.n32 Clk.n27 3.56405
R7048 Clk.n2 SARlogic_0.dffrs_13.nand3_6.B 2.17818
R7049 Clk.n24 SARlogic_0.dffrs_0.nand3_6.B 2.17818
R7050 Clk.n20 SARlogic_0.dffrs_1.nand3_6.B 2.17818
R7051 Clk.n16 SARlogic_0.dffrs_2.nand3_6.B 2.17818
R7052 Clk.n12 SARlogic_0.dffrs_3.nand3_6.B 2.17818
R7053 Clk.n8 SARlogic_0.dffrs_4.nand3_6.B 2.17818
R7054 Clk.n5 SARlogic_0.dffrs_5.nand3_6.B 2.17818
R7055 comparator_no_offsetcal_0.CLK Clk.n32 1.60543
R7056 Clk.n2 SARlogic_0.dffrs_13.nand3_1.A 1.34729
R7057 Clk.n24 SARlogic_0.dffrs_0.nand3_1.A 1.34729
R7058 Clk.n20 SARlogic_0.dffrs_1.nand3_1.A 1.34729
R7059 Clk.n16 SARlogic_0.dffrs_2.nand3_1.A 1.34729
R7060 Clk.n12 SARlogic_0.dffrs_3.nand3_1.A 1.34729
R7061 Clk.n8 SARlogic_0.dffrs_4.nand3_1.A 1.34729
R7062 Clk.n5 SARlogic_0.dffrs_5.nand3_1.A 1.34729
R7063 Clk.n29 Clk.n28 1.01892
R7064 Clk.n31 Clk.n30 1.01892
R7065 SARlogic_0.dffrs_13.clk Clk.n2 0.611214
R7066 SARlogic_0.dffrs_0.clk Clk.n24 0.611214
R7067 SARlogic_0.dffrs_1.clk Clk.n20 0.611214
R7068 SARlogic_0.dffrs_2.clk Clk.n16 0.611214
R7069 SARlogic_0.dffrs_3.clk Clk.n12 0.611214
R7070 SARlogic_0.dffrs_4.clk Clk.n8 0.611214
R7071 SARlogic_0.dffrs_5.clk Clk.n5 0.611214
R7072 Clk.n33 Clk 0.514034
R7073 SARlogic_0.clk Clk.n26 0.13775
R7074 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t8 41.0041
R7075 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t6 40.8177
R7076 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t7 40.6313
R7077 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t4 27.3166
R7078 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t9 27.1302
R7079 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t5 26.9438
R7080 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.t2 10.0473
R7081 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n4 9.90747
R7082 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n2 9.90116
R7083 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.t1 6.51042
R7084 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.n7 6.04952
R7085 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_6.C.n1 5.7305
R7086 SARlogic_0.dffrs_1.nand3_2.B SARlogic_0.dffrs_1.nand3_6.C.n0 5.47979
R7087 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C.n3 5.13907
R7088 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n9 4.72925
R7089 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_6.C.n5 4.5005
R7090 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.n8 0.732092
R7091 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t0 0.7285
R7092 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t3 0.7285
R7093 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n6 0.449758
R7094 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_2.B 0.166901
R7095 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_0.A 0.0455
R7096 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C 0.0455
R7097 SARlogic_0.d2.n3 SARlogic_0.d2.t5 41.0041
R7098 SARlogic_0.d2.n4 SARlogic_0.d2.t11 40.8177
R7099 SARlogic_0.d2.n7 SARlogic_0.d2.t4 40.6313
R7100 SARlogic_0.d2.n1 SARlogic_0.d2.t6 34.2529
R7101 SARlogic_0.d2.n6 SARlogic_0.dffrs_8.clk 34.1594
R7102 SARlogic_0.d2.n7 SARlogic_0.d2.t10 27.3166
R7103 SARlogic_0.d2.n4 SARlogic_0.d2.t9 27.1302
R7104 SARlogic_0.d2.n3 SARlogic_0.d2.t7 26.9438
R7105 SARlogic_0.d2.n0 SARlogic_0.d2.t8 19.673
R7106 SARlogic_0.d2.n0 SARlogic_0.d2.t12 19.4007
R7107 SARlogic_0.d2 adc_PISO_0.B3 17.5376
R7108 SARlogic_0.d2.n9 SARlogic_0.d2.n8 14.0582
R7109 SARlogic_0.d2.n9 SARlogic_0.d2.n6 12.0118
R7110 SARlogic_0.d2.n12 SARlogic_0.d2.t1 10.0473
R7111 SARlogic_0.d2.n2 SARlogic_0.d2.n1 8.05164
R7112 SARlogic_0.d2.n11 SARlogic_0.d2.t2 6.51042
R7113 SARlogic_0.d2.n11 SARlogic_0.d2.n10 6.04952
R7114 SARlogic_0.dffrs_8.nand3_1.A SARlogic_0.d2.n3 5.7755
R7115 SARlogic_0.dffrs_8.nand3_6.B SARlogic_0.d2.n4 5.47979
R7116 SARlogic_0.d2.n8 SARlogic_0.d2.n7 5.13907
R7117 SARlogic_0.dffrs_9.nand3_2.Z SARlogic_0.d2.n12 4.72925
R7118 SARlogic_0.d2.n5 SARlogic_0.dffrs_8.nand3_6.B 2.17818
R7119 adc_PISO_0.B3 SARlogic_0.d2.n2 1.87121
R7120 SARlogic_0.d2.n5 SARlogic_0.dffrs_8.nand3_1.A 1.34729
R7121 SARlogic_0.d2.n12 SARlogic_0.d2.n11 0.732092
R7122 SARlogic_0.d2.n10 SARlogic_0.d2.t3 0.7285
R7123 SARlogic_0.d2.n10 SARlogic_0.d2.t0 0.7285
R7124 SARlogic_0.d2.n6 SARlogic_0.d2 0.698
R7125 SARlogic_0.dffrs_8.clk SARlogic_0.d2.n5 0.610571
R7126 SARlogic_0.dffrs_9.nand3_2.Z SARlogic_0.d2.n9 0.166901
R7127 SARlogic_0.d2.n1 SARlogic_0.d2.n0 0.106438
R7128 SARlogic_0.d2.n8 SARlogic_0.dffrs_9.nand3_7.C 0.0455
R7129 SARlogic_0.d2.n2 adc_PISO_0.2inmux_4.In 0.0455
R7130 a_4841_31422.n3 a_4841_31422.t4 41.0041
R7131 a_4841_31422.n2 a_4841_31422.t6 40.8177
R7132 a_4841_31422.n4 a_4841_31422.t7 40.6313
R7133 a_4841_31422.n4 a_4841_31422.t9 27.3166
R7134 a_4841_31422.n2 a_4841_31422.t8 27.1302
R7135 a_4841_31422.n3 a_4841_31422.t5 26.9438
R7136 a_4841_31422.n5 a_4841_31422.n3 15.6312
R7137 a_4841_31422.n5 a_4841_31422.n4 15.046
R7138 a_4841_31422.t0 a_4841_31422.n7 10.0473
R7139 a_4841_31422.n1 a_4841_31422.t3 6.51042
R7140 a_4841_31422.n1 a_4841_31422.n0 6.04952
R7141 a_4841_31422.n6 a_4841_31422.n2 5.64619
R7142 a_4841_31422.n7 a_4841_31422.n6 5.17851
R7143 a_4841_31422.n6 a_4841_31422.n5 4.5005
R7144 a_4841_31422.n7 a_4841_31422.n1 0.732092
R7145 a_4841_31422.n0 a_4841_31422.t2 0.7285
R7146 a_4841_31422.n0 a_4841_31422.t1 0.7285
R7147 a_4841_33627.n0 a_4841_33627.t4 40.6313
R7148 a_4841_33627.n0 a_4841_33627.t5 27.3166
R7149 a_4841_33627.n1 a_4841_33627.n0 24.1527
R7150 a_4841_33627.n1 a_4841_33627.t1 10.0473
R7151 a_4841_33627.n2 a_4841_33627.t2 6.51042
R7152 a_4841_33627.n3 a_4841_33627.n2 6.04952
R7153 a_4841_33627.n2 a_4841_33627.n1 0.732092
R7154 a_4841_33627.t0 a_4841_33627.n3 0.7285
R7155 a_4841_33627.n3 a_4841_33627.t3 0.7285
R7156 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t6 40.6313
R7157 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.t4 34.1066
R7158 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t7 27.3166
R7159 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t5 19.673
R7160 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t8 19.4007
R7161 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n3 14.6967
R7162 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.t1 10.0473
R7163 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n6 9.39565
R7164 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit.n1 6.70486
R7165 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.t2 6.51042
R7166 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.n4 6.04952
R7167 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n2 5.81514
R7168 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.n5 0.732092
R7169 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t0 0.7285
R7170 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t3 0.7285
R7171 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n7 0.458082
R7172 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.n0 0.252687
R7173 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit 0.0519286
R7174 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t4 40.6313
R7175 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t5 27.3166
R7176 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n1 14.2854
R7177 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.t0 10.0473
R7178 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.t1 6.51042
R7179 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.n2 6.04952
R7180 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C.n0 5.13907
R7181 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n4 4.72925
R7182 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.n3 0.732092
R7183 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t3 0.7285
R7184 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t2 0.7285
R7185 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C 0.0455
R7186 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t5 41.0041
R7187 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t6 40.8177
R7188 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t4 40.6313
R7189 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t9 27.3166
R7190 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t7 27.1302
R7191 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t8 26.9438
R7192 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.t2 10.0473
R7193 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n4 9.90747
R7194 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n2 9.90116
R7195 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.t3 6.51042
R7196 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.n7 6.04952
R7197 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_6.C.n1 5.7305
R7198 SARlogic_0.dffrs_3.nand3_2.B SARlogic_0.dffrs_3.nand3_6.C.n0 5.47979
R7199 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C.n3 5.13907
R7200 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n9 4.72925
R7201 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_6.C.n5 4.5005
R7202 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.n8 0.732092
R7203 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t1 0.7285
R7204 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t0 0.7285
R7205 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n6 0.449758
R7206 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_2.B 0.166901
R7207 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_0.A 0.0455
R7208 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C 0.0455
R7209 a_33337_30170.n2 a_33337_30170.t7 41.0041
R7210 a_33337_30170.n3 a_33337_30170.t4 40.8177
R7211 a_33337_30170.n3 a_33337_30170.t6 27.1302
R7212 a_33337_30170.n2 a_33337_30170.t5 26.9438
R7213 a_33337_30170.n4 a_33337_30170.n3 22.5284
R7214 a_33337_30170.n5 a_33337_30170.n4 19.5781
R7215 a_33337_30170.t0 a_33337_30170.n5 10.0473
R7216 a_33337_30170.n1 a_33337_30170.t1 6.51042
R7217 a_33337_30170.n1 a_33337_30170.n0 6.04952
R7218 a_33337_30170.n4 a_33337_30170.n2 5.7305
R7219 a_33337_30170.n5 a_33337_30170.n1 0.732092
R7220 a_33337_30170.n0 a_33337_30170.t2 0.7285
R7221 a_33337_30170.n0 a_33337_30170.t3 0.7285
R7222 a_33257_33628.n2 a_33257_33628.t4 40.6313
R7223 a_33257_33628.n2 a_33257_33628.t5 27.3166
R7224 a_33257_33628.n3 a_33257_33628.n2 24.1527
R7225 a_33257_33628.t0 a_33257_33628.n3 10.0473
R7226 a_33257_33628.n1 a_33257_33628.t1 6.51042
R7227 a_33257_33628.n1 a_33257_33628.n0 6.04952
R7228 a_33257_33628.n3 a_33257_33628.n1 0.732092
R7229 a_33257_33628.n0 a_33257_33628.t2 0.7285
R7230 a_33257_33628.n0 a_33257_33628.t3 0.7285
R7231 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t5 41.0041
R7232 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t4 40.6313
R7233 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t6 27.3166
R7234 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t7 26.9438
R7235 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d 17.5022
R7236 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d.n2 14.0582
R7237 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.t2 10.0473
R7238 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.t1 6.51042
R7239 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.n4 6.04952
R7240 SARlogic_0.dffrs_0.nand3_8.A SARlogic_0.dffrs_0.d.n0 5.7755
R7241 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_0.d.n1 5.13907
R7242 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n6 4.72925
R7243 SARlogic_0.dffrs_0.d SARlogic_0.dffrs_0.nand3_8.A 0.783821
R7244 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.n5 0.732092
R7245 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t3 0.7285
R7246 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t0 0.7285
R7247 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n3 0.166901
R7248 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_13.nand3_7.C 0.0455
R7249 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t7 41.0041
R7250 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t4 40.6313
R7251 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t8 40.6313
R7252 SARlogic_0.dffrs_13.Qb SARlogic_0.dffrs_14.setb 27.9776
R7253 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t6 27.3166
R7254 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t5 27.3166
R7255 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t9 26.9438
R7256 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.t1 10.0473
R7257 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb.n1 9.84255
R7258 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n3 9.22229
R7259 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.t2 6.51042
R7260 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.n7 6.04952
R7261 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.Qb.n0 5.7305
R7262 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n4 5.14711
R7263 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_13.Qb.n2 5.13907
R7264 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n6 4.94976
R7265 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n9 4.72925
R7266 SARlogic_0.dffrs_14.setb SARlogic_0.dffrs_14.nand3_0.C 0.784786
R7267 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.n8 0.732092
R7268 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t0 0.7285
R7269 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t3 0.7285
R7270 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb 0.175225
R7271 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.nand3_2.A 0.0455
R7272 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_14.nand3_2.C 0.0455
R7273 SARlogic_0.dffrs_14.nand3_0.C SARlogic_0.dffrs_13.Qb.n5 0.0374643
R7274 Comp_out.n0 Comp_out 11.2807
R7275 Comp_out.n6 Comp_out.n5 6.5435
R7276 Comp_out.n3 Comp_out.n2 6.5435
R7277 comparator_no_offsetcal_0.x4.Y Comp_out.n9 4.5005
R7278 comparator_no_offsetcal_0.x4.Y Comp_out.n0 2.3842
R7279 Comp_out.n7 Comp_out.n4 2.17483
R7280 Comp_out.n5 Comp_out.t1 2.03874
R7281 Comp_out.n5 Comp_out.t2 2.03874
R7282 Comp_out.n2 Comp_out.t0 2.03874
R7283 Comp_out.n2 Comp_out.t3 2.03874
R7284 Comp_out.n9 Comp_out.n1 2.00383
R7285 Comp_out.n1 Comp_out.t7 1.13285
R7286 Comp_out.n1 Comp_out.t6 1.13285
R7287 Comp_out.n4 Comp_out.t4 1.13285
R7288 Comp_out.n4 Comp_out.t5 1.13285
R7289 Comp_out.n6 Comp_out.n3 0.5105
R7290 Comp_out.n8 Comp_out.n7 0.5105
R7291 Comp_out.n0 comparator_no_offsetcal_0.Vout 0.3995
R7292 Comp_out.n8 Comp_out.n3 0.2165
R7293 Comp_out.n7 Comp_out.n6 0.2165
R7294 Comp_out.n9 Comp_out.n8 0.1175
R7295 a_9083_28820.n0 a_9083_28820.t4 34.1797
R7296 a_9083_28820.n0 a_9083_28820.t5 19.5798
R7297 a_9083_28820.t1 a_9083_28820.n3 18.7717
R7298 a_9083_28820.n3 a_9083_28820.t0 9.2885
R7299 a_9083_28820.n2 a_9083_28820.n0 4.93379
R7300 a_9083_28820.n1 a_9083_28820.t3 4.23346
R7301 a_9083_28820.n1 a_9083_28820.t2 3.85546
R7302 a_9083_28820.n3 a_9083_28820.n2 0.4055
R7303 a_9083_28820.n2 a_9083_28820.n1 0.352625
R7304 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t7 41.0041
R7305 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t8 40.8177
R7306 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t6 40.6313
R7307 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t5 27.3166
R7308 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t4 27.1302
R7309 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t9 26.9438
R7310 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.t2 10.0473
R7311 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n4 9.90747
R7312 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n2 9.90116
R7313 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.t3 6.51042
R7314 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.n7 6.04952
R7315 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_6.C.n1 5.7305
R7316 SARlogic_0.dffrs_9.nand3_2.B SARlogic_0.dffrs_9.nand3_6.C.n0 5.47979
R7317 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C.n3 5.13907
R7318 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n9 4.72925
R7319 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_6.C.n5 4.5005
R7320 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.n8 0.732092
R7321 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t0 0.7285
R7322 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t1 0.7285
R7323 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n6 0.449758
R7324 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_2.B 0.166901
R7325 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_0.A 0.0455
R7326 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C 0.0455
R7327 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t6 40.8177
R7328 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t7 40.6313
R7329 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t4 27.3166
R7330 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t5 27.1302
R7331 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_8.C.n2 14.119
R7332 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.t1 10.0473
R7333 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.t0 6.51042
R7334 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.n4 6.04952
R7335 SARlogic_0.dffrs_2.nand3_7.B SARlogic_0.dffrs_2.nand3_8.C.n0 5.47979
R7336 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C.n1 5.13907
R7337 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n6 4.72925
R7338 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.n5 0.732092
R7339 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t3 0.7285
R7340 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t2 0.7285
R7341 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_7.B 0.438233
R7342 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n3 0.166901
R7343 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C 0.0455
R7344 a_30255_29264.n0 a_30255_29264.t5 34.1797
R7345 a_30255_29264.n0 a_30255_29264.t4 19.5798
R7346 a_30255_29264.t0 a_30255_29264.n3 10.3401
R7347 a_30255_29264.n3 a_30255_29264.t1 9.2885
R7348 a_30255_29264.n2 a_30255_29264.n0 4.93379
R7349 a_30255_29264.n1 a_30255_29264.t2 4.09202
R7350 a_30255_29264.n1 a_30255_29264.t3 3.95079
R7351 a_30255_29264.n3 a_30255_29264.n2 0.599711
R7352 a_30255_29264.n2 a_30255_29264.n1 0.296375
R7353 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t3 41.0041
R7354 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t2 26.9438
R7355 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t0 9.6935
R7356 adc_PISO_0.dffrs_4.d adc_PISO_0.2inmux_5.OUT.n0 6.55979
R7357 adc_PISO_0.2inmux_5.OUT adc_PISO_0.dffrs_4.d 4.883
R7358 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t1 4.35383
R7359 adc_PISO_0.2inmux_5.OUT adc_PISO_0.2inmux_5.OUT.n1 0.350857
R7360 SARlogic_0.d0.n3 SARlogic_0.d0.t4 41.0041
R7361 SARlogic_0.d0.n4 SARlogic_0.d0.t10 40.8177
R7362 SARlogic_0.d0.n7 SARlogic_0.d0.t5 40.6313
R7363 SARlogic_0.d0.n6 adc_PISO_0.B1 36.2544
R7364 SARlogic_0.d0.n1 SARlogic_0.d0.t9 34.2529
R7365 SARlogic_0.d0.n6 SARlogic_0.dffrs_10.clk 33.5936
R7366 SARlogic_0.d0.n7 SARlogic_0.d0.t12 27.3166
R7367 SARlogic_0.d0.n4 SARlogic_0.d0.t7 27.1302
R7368 SARlogic_0.d0.n3 SARlogic_0.d0.t6 26.9438
R7369 SARlogic_0.d0.n0 SARlogic_0.d0.t11 19.673
R7370 SARlogic_0.d0.n0 SARlogic_0.d0.t8 19.4007
R7371 SARlogic_0.d0.n9 SARlogic_0.d0.n8 14.0582
R7372 SARlogic_0.d0.n9 SARlogic_0.d0.n6 11.4461
R7373 SARlogic_0.d0.n12 SARlogic_0.d0.t1 10.0473
R7374 SARlogic_0.d0.n2 SARlogic_0.d0.n1 8.05164
R7375 SARlogic_0.d0.n11 SARlogic_0.d0.t2 6.51042
R7376 SARlogic_0.d0.n11 SARlogic_0.d0.n10 6.04952
R7377 SARlogic_0.dffrs_10.nand3_1.A SARlogic_0.d0.n3 5.7755
R7378 SARlogic_0.dffrs_10.nand3_6.B SARlogic_0.d0.n4 5.47979
R7379 SARlogic_0.d0.n8 SARlogic_0.d0.n7 5.13907
R7380 SARlogic_0.dffrs_11.nand3_2.Z SARlogic_0.d0.n12 4.72925
R7381 SARlogic_0.d0.n5 SARlogic_0.dffrs_10.nand3_6.B 2.17818
R7382 adc_PISO_0.B1 SARlogic_0.d0.n2 1.87121
R7383 SARlogic_0.d0.n5 SARlogic_0.dffrs_10.nand3_1.A 1.34729
R7384 SARlogic_0.d0.n12 SARlogic_0.d0.n11 0.732092
R7385 SARlogic_0.d0.n10 SARlogic_0.d0.t0 0.7285
R7386 SARlogic_0.d0.n10 SARlogic_0.d0.t3 0.7285
R7387 SARlogic_0.dffrs_10.clk SARlogic_0.d0.n5 0.610571
R7388 SARlogic_0.dffrs_11.nand3_2.Z SARlogic_0.d0.n9 0.166901
R7389 SARlogic_0.d0.n1 SARlogic_0.d0.n0 0.106438
R7390 SARlogic_0.d0.n8 SARlogic_0.dffrs_11.nand3_7.C 0.0455
R7391 SARlogic_0.d0.n2 adc_PISO_0.2inmux_1.In 0.0455
R7392 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t4 41.0041
R7393 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t5 40.8177
R7394 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t9 40.6313
R7395 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t8 27.3166
R7396 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t7 27.1302
R7397 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t6 26.9438
R7398 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.t2 10.0473
R7399 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n4 9.90747
R7400 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n2 9.90116
R7401 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.t3 6.51042
R7402 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.n7 6.04952
R7403 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_6.C.n1 5.7305
R7404 SARlogic_0.dffrs_10.nand3_2.B SARlogic_0.dffrs_10.nand3_6.C.n0 5.47979
R7405 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C.n3 5.13907
R7406 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n9 4.72925
R7407 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_6.C.n5 4.5005
R7408 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.n8 0.732092
R7409 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t1 0.7285
R7410 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t0 0.7285
R7411 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n6 0.449758
R7412 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_2.B 0.166901
R7413 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_0.A 0.0455
R7414 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C 0.0455
R7415 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t8 41.0041
R7416 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t5 40.6313
R7417 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t4 40.6313
R7418 SARlogic_0.dffrs_3.Qb SARlogic_0.dffrs_10.setb 28.021
R7419 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t7 27.3166
R7420 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t6 27.3166
R7421 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t9 26.9438
R7422 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.t2 10.0473
R7423 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb.n1 9.84255
R7424 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n3 9.22229
R7425 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.t1 6.51042
R7426 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.n7 6.04952
R7427 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.Qb.n0 5.7305
R7428 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n4 5.14711
R7429 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_3.Qb.n2 5.13907
R7430 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n6 4.94976
R7431 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n9 4.72925
R7432 SARlogic_0.dffrs_10.setb SARlogic_0.dffrs_10.nand3_0.C 0.784786
R7433 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.n8 0.732092
R7434 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t0 0.7285
R7435 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t3 0.7285
R7436 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb 0.175225
R7437 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.nand3_2.A 0.0455
R7438 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_10.nand3_2.C 0.0455
R7439 SARlogic_0.dffrs_10.nand3_0.C SARlogic_0.dffrs_3.Qb.n5 0.0374643
R7440 a_14313_33628.n2 a_14313_33628.t5 40.6313
R7441 a_14313_33628.n2 a_14313_33628.t4 27.3166
R7442 a_14313_33628.n3 a_14313_33628.n2 24.1527
R7443 a_14313_33628.t0 a_14313_33628.n3 10.0473
R7444 a_14313_33628.n1 a_14313_33628.t2 6.51042
R7445 a_14313_33628.n1 a_14313_33628.n0 6.04952
R7446 a_14313_33628.n3 a_14313_33628.n1 0.732092
R7447 a_14313_33628.n0 a_14313_33628.t3 0.7285
R7448 a_14313_33628.n0 a_14313_33628.t1 0.7285
R7449 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t8 41.0041
R7450 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t4 40.6313
R7451 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t5 40.6313
R7452 SARlogic_0.dffrs_5.Qb SARlogic_0.dffrs_12.setb 28.013
R7453 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t6 27.3166
R7454 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t7 27.3166
R7455 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t9 26.9438
R7456 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.t0 10.0473
R7457 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb.n1 9.84255
R7458 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n3 9.22229
R7459 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.t1 6.51042
R7460 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.n7 6.04952
R7461 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.Qb.n0 5.7305
R7462 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n4 5.14711
R7463 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_5.Qb.n2 5.13907
R7464 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n6 4.94976
R7465 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n9 4.72925
R7466 SARlogic_0.dffrs_12.setb SARlogic_0.dffrs_12.nand3_0.C 0.784786
R7467 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.n8 0.732092
R7468 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t3 0.7285
R7469 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t2 0.7285
R7470 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb 0.175225
R7471 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.nand3_2.A 0.0455
R7472 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_12.nand3_2.C 0.0455
R7473 SARlogic_0.dffrs_12.nand3_0.C SARlogic_0.dffrs_5.Qb.n5 0.0374643
R7474 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t4 40.6313
R7475 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.t8 34.1066
R7476 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t5 27.3166
R7477 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t6 19.673
R7478 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t7 19.4007
R7479 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n3 14.6967
R7480 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.t0 10.0473
R7481 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n6 9.39565
R7482 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.dffrs_1.Q.n1 6.70486
R7483 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.t1 6.51042
R7484 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.n4 6.04952
R7485 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n2 5.81354
R7486 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.n5 0.732092
R7487 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t2 0.7285
R7488 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t3 0.7285
R7489 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n7 0.458082
R7490 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.n0 0.252687
R7491 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.2inmux_3.Bit 0.0519286
R7492 SARlogic_0.d5.n3 SARlogic_0.d5.t4 40.6313
R7493 SARlogic_0.d5.n1 SARlogic_0.d5.t6 34.2529
R7494 SARlogic_0.d5.n3 SARlogic_0.d5.t8 27.3166
R7495 SARlogic_0.d5.n5 adc_PISO_0.B6 23.5656
R7496 SARlogic_0.d5.n0 SARlogic_0.d5.t7 19.673
R7497 SARlogic_0.d5.n0 SARlogic_0.d5.t5 19.4007
R7498 SARlogic_0.d5.n5 SARlogic_0.d5.n4 14.0582
R7499 SARlogic_0.d5.n8 SARlogic_0.d5.t2 10.0473
R7500 SARlogic_0.d5.n2 SARlogic_0.d5.n1 8.05164
R7501 SARlogic_0.d5.n7 SARlogic_0.d5.t1 6.51042
R7502 SARlogic_0.d5.n7 SARlogic_0.d5.n6 6.04952
R7503 SARlogic_0.d5.n4 SARlogic_0.d5.n3 5.13907
R7504 SARlogic_0.dffrs_14.nand3_2.Z SARlogic_0.d5.n8 4.72925
R7505 adc_PISO_0.B6 SARlogic_0.d5.n2 1.87121
R7506 SARlogic_0.d5.n8 SARlogic_0.d5.n7 0.732092
R7507 SARlogic_0.d5.n6 SARlogic_0.d5.t0 0.7285
R7508 SARlogic_0.d5.n6 SARlogic_0.d5.t3 0.7285
R7509 SARlogic_0.dffrs_14.nand3_2.Z SARlogic_0.d5.n5 0.166901
R7510 SARlogic_0.d5.n1 SARlogic_0.d5.n0 0.106438
R7511 SARlogic_0.d5.n4 SARlogic_0.dffrs_14.nand3_7.C 0.0455
R7512 SARlogic_0.d5.n2 adc_PISO_0.2inmux_0.In 0.0455
R7513 a_33257_29218.n0 a_33257_29218.t4 40.8177
R7514 a_33257_29218.n1 a_33257_29218.t7 40.6313
R7515 a_33257_29218.n1 a_33257_29218.t6 27.3166
R7516 a_33257_29218.n0 a_33257_29218.t5 27.1302
R7517 a_33257_29218.n2 a_33257_29218.n1 19.2576
R7518 a_33257_29218.n3 a_33257_29218.t1 10.0473
R7519 a_33257_29218.n4 a_33257_29218.t2 6.51042
R7520 a_33257_29218.n5 a_33257_29218.n4 6.04952
R7521 a_33257_29218.n2 a_33257_29218.n0 5.91752
R7522 a_33257_29218.n3 a_33257_29218.n2 4.89565
R7523 a_33257_29218.n4 a_33257_29218.n3 0.732092
R7524 a_33257_29218.n5 a_33257_29218.t3 0.7285
R7525 a_33257_29218.t0 a_33257_29218.n5 0.7285
R7526 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t5 41.0041
R7527 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t6 40.6313
R7528 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t4 40.6313
R7529 SARlogic_0.dffrs_0.Qb SARlogic_0.dffrs_7.setb 28.021
R7530 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t9 27.3166
R7531 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t7 27.3166
R7532 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t8 26.9438
R7533 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.t3 10.0473
R7534 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb.n1 9.84255
R7535 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n3 9.22229
R7536 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.t2 6.51042
R7537 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.n7 6.04952
R7538 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.Qb.n0 5.7305
R7539 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n4 5.14711
R7540 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_0.Qb.n2 5.13907
R7541 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n6 4.94976
R7542 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n9 4.72925
R7543 SARlogic_0.dffrs_7.setb SARlogic_0.dffrs_7.nand3_0.C 0.784786
R7544 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.n8 0.732092
R7545 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t0 0.7285
R7546 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t1 0.7285
R7547 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb 0.175225
R7548 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.nand3_2.A 0.0455
R7549 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_7.nand3_2.C 0.0455
R7550 SARlogic_0.dffrs_7.nand3_0.C SARlogic_0.dffrs_0.Qb.n5 0.0374643
R7551 a_9083_31160.n0 a_9083_31160.t5 34.1797
R7552 a_9083_31160.n0 a_9083_31160.t4 19.5798
R7553 a_9083_31160.n3 a_9083_31160.t0 18.7717
R7554 a_9083_31160.t1 a_9083_31160.n3 9.2885
R7555 a_9083_31160.n2 a_9083_31160.n0 4.93379
R7556 a_9083_31160.n1 a_9083_31160.t3 4.23346
R7557 a_9083_31160.n1 a_9083_31160.t2 3.85546
R7558 a_9083_31160.n3 a_9083_31160.n2 0.4055
R7559 a_9083_31160.n2 a_9083_31160.n1 0.352625
R7560 a_23785_29218.n0 a_23785_29218.t5 40.8177
R7561 a_23785_29218.n1 a_23785_29218.t4 40.6313
R7562 a_23785_29218.n1 a_23785_29218.t7 27.3166
R7563 a_23785_29218.n0 a_23785_29218.t6 27.1302
R7564 a_23785_29218.n2 a_23785_29218.n1 19.2576
R7565 a_23785_29218.n3 a_23785_29218.t1 10.0473
R7566 a_23785_29218.n4 a_23785_29218.t2 6.51042
R7567 a_23785_29218.n5 a_23785_29218.n4 6.04952
R7568 a_23785_29218.n2 a_23785_29218.n0 5.91752
R7569 a_23785_29218.n3 a_23785_29218.n2 4.89565
R7570 a_23785_29218.n4 a_23785_29218.n3 0.732092
R7571 a_23785_29218.n5 a_23785_29218.t3 0.7285
R7572 a_23785_29218.t0 a_23785_29218.n5 0.7285
R7573 a_23865_30170.n2 a_23865_30170.t7 41.0041
R7574 a_23865_30170.n3 a_23865_30170.t5 40.8177
R7575 a_23865_30170.n3 a_23865_30170.t6 27.1302
R7576 a_23865_30170.n2 a_23865_30170.t4 26.9438
R7577 a_23865_30170.n4 a_23865_30170.n3 22.5284
R7578 a_23865_30170.n5 a_23865_30170.n4 19.5781
R7579 a_23865_30170.t0 a_23865_30170.n5 10.0473
R7580 a_23865_30170.n1 a_23865_30170.t3 6.51042
R7581 a_23865_30170.n1 a_23865_30170.n0 6.04952
R7582 a_23865_30170.n4 a_23865_30170.n2 5.7305
R7583 a_23865_30170.n5 a_23865_30170.n1 0.732092
R7584 a_23865_30170.n0 a_23865_30170.t2 0.7285
R7585 a_23865_30170.n0 a_23865_30170.t1 0.7285
R7586 Piso_out.n5 Piso_out.n4 6.5435
R7587 Piso_out.n2 Piso_out.n1 6.5435
R7588 osu_sc_buf_4_flat_0.Y Piso_out.n8 4.5005
R7589 osu_sc_buf_4_flat_0.Y Piso_out 2.2685
R7590 Piso_out.n6 Piso_out.n3 2.17483
R7591 Piso_out.n4 Piso_out.t1 2.03874
R7592 Piso_out.n4 Piso_out.t3 2.03874
R7593 Piso_out.n1 Piso_out.t0 2.03874
R7594 Piso_out.n1 Piso_out.t2 2.03874
R7595 Piso_out.n8 Piso_out.n0 2.00383
R7596 Piso_out.n0 Piso_out.t7 1.13285
R7597 Piso_out.n0 Piso_out.t5 1.13285
R7598 Piso_out.n3 Piso_out.t4 1.13285
R7599 Piso_out.n3 Piso_out.t6 1.13285
R7600 Piso_out.n5 Piso_out.n2 0.5105
R7601 Piso_out.n7 Piso_out.n6 0.5105
R7602 Piso_out.n7 Piso_out.n2 0.2165
R7603 Piso_out.n6 Piso_out.n5 0.2165
R7604 Piso_out.n8 Piso_out.n7 0.1175
R7605 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t4 40.6313
R7606 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t5 27.3166
R7607 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n1 14.2854
R7608 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.t1 10.0473
R7609 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.t2 6.51042
R7610 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.n2 6.04952
R7611 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C.n0 5.13907
R7612 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n4 4.72925
R7613 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.n3 0.732092
R7614 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t0 0.7285
R7615 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t3 0.7285
R7616 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C 0.0455
R7617 a_42729_33628.n0 a_42729_33628.t4 40.6313
R7618 a_42729_33628.n0 a_42729_33628.t5 27.3166
R7619 a_42729_33628.n1 a_42729_33628.n0 24.1527
R7620 a_42729_33628.n1 a_42729_33628.t1 10.0473
R7621 a_42729_33628.t0 a_42729_33628.n3 6.51042
R7622 a_42729_33628.n3 a_42729_33628.n2 6.04952
R7623 a_42729_33628.n3 a_42729_33628.n1 0.732092
R7624 a_42729_33628.n2 a_42729_33628.t3 0.7285
R7625 a_42729_33628.n2 a_42729_33628.t2 0.7285
R7626 a_42729_31423.n1 a_42729_31423.t4 41.0041
R7627 a_42729_31423.n0 a_42729_31423.t5 40.8177
R7628 a_42729_31423.n2 a_42729_31423.t6 40.6313
R7629 a_42729_31423.n2 a_42729_31423.t9 27.3166
R7630 a_42729_31423.n0 a_42729_31423.t8 27.1302
R7631 a_42729_31423.n1 a_42729_31423.t7 26.9438
R7632 a_42729_31423.n3 a_42729_31423.n1 15.6312
R7633 a_42729_31423.n3 a_42729_31423.n2 15.046
R7634 a_42729_31423.n5 a_42729_31423.t3 10.0473
R7635 a_42729_31423.n6 a_42729_31423.t2 6.51042
R7636 a_42729_31423.n7 a_42729_31423.n6 6.04952
R7637 a_42729_31423.n4 a_42729_31423.n0 5.64619
R7638 a_42729_31423.n5 a_42729_31423.n4 5.17851
R7639 a_42729_31423.n4 a_42729_31423.n3 4.5005
R7640 a_42729_31423.n6 a_42729_31423.n5 0.732092
R7641 a_42729_31423.n7 a_42729_31423.t1 0.7285
R7642 a_42729_31423.t0 a_42729_31423.n7 0.7285
R7643 a_28027_31160.n0 a_28027_31160.t4 34.1797
R7644 a_28027_31160.n0 a_28027_31160.t5 19.5798
R7645 a_28027_31160.n3 a_28027_31160.t0 18.7717
R7646 a_28027_31160.t1 a_28027_31160.n3 9.2885
R7647 a_28027_31160.n2 a_28027_31160.n0 4.93379
R7648 a_28027_31160.n1 a_28027_31160.t3 4.23346
R7649 a_28027_31160.n1 a_28027_31160.t2 3.85546
R7650 a_28027_31160.n3 a_28027_31160.n2 0.4055
R7651 a_28027_31160.n2 a_28027_31160.n1 0.352625
R7652 a_23785_31423.n1 a_23785_31423.t5 41.0041
R7653 a_23785_31423.n0 a_23785_31423.t7 40.8177
R7654 a_23785_31423.n2 a_23785_31423.t4 40.6313
R7655 a_23785_31423.n2 a_23785_31423.t6 27.3166
R7656 a_23785_31423.n0 a_23785_31423.t9 27.1302
R7657 a_23785_31423.n1 a_23785_31423.t8 26.9438
R7658 a_23785_31423.n3 a_23785_31423.n1 15.6312
R7659 a_23785_31423.n3 a_23785_31423.n2 15.046
R7660 a_23785_31423.n5 a_23785_31423.t1 10.0473
R7661 a_23785_31423.n6 a_23785_31423.t3 6.51042
R7662 a_23785_31423.n7 a_23785_31423.n6 6.04952
R7663 a_23785_31423.n4 a_23785_31423.n0 5.64619
R7664 a_23785_31423.n5 a_23785_31423.n4 5.17851
R7665 a_23785_31423.n4 a_23785_31423.n3 4.5005
R7666 a_23785_31423.n6 a_23785_31423.n5 0.732092
R7667 a_23785_31423.n7 a_23785_31423.t2 0.7285
R7668 a_23785_31423.t0 a_23785_31423.n7 0.7285
R7669 Vin1.n7 Vin1.n6 23.1032
R7670 Vin1.n3 Vin1.n2 23.1032
R7671 Vin1.n0 Vin1.t8 22.5295
R7672 Vin1.n2 Vin1.t2 16.3641
R7673 Vin1.n6 Vin1.t6 16.3626
R7674 Vin1.n2 Vin1.t7 16.0225
R7675 Vin1.n6 Vin1.t1 16.021
R7676 Vin1.n8 Vin1.t4 11.5195
R7677 Vin1.n5 Vin1.t3 11.5195
R7678 Vin1.n4 Vin1.t9 11.5195
R7679 Vin1.n1 Vin1.t5 11.5195
R7680 Vin1.n0 Vin1.t0 11.5195
R7681 comparator_no_offsetcal_0.Vin1 Vin1 5.6843
R7682 Vin1.n1 Vin1.n0 4.00673
R7683 comparator_no_offsetcal_0.Vin1 Vin1.n8 3.9441
R7684 Vin1.n7 Vin1.n5 3.16619
R7685 Vin1.n3 Vin1.n1 0.650658
R7686 Vin1.n8 Vin1.n7 0.280193
R7687 Vin1.n4 Vin1.n3 0.279681
R7688 Vin1.n5 Vin1.n4 0.231705
R7689 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t15 19.5626
R7690 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 11.9065
R7691 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 11.2495
R7692 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 11.243
R7693 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 8.80104
R7694 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 6.60725
R7695 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 6.52262
R7696 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 6.386
R7697 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 5.44213
R7698 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 4.36738
R7699 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 4.36738
R7700 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 4.3505
R7701 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 2.2505
R7702 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 2.14009
R7703 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 1.50001
R7704 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 1.49326
R7705 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t0 1.0925
R7706 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t6 1.0925
R7707 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t5 1.0925
R7708 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t10 1.0925
R7709 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t3 1.0925
R7710 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t8 1.0925
R7711 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t11 1.0925
R7712 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t1 1.0925
R7713 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t7 1.0925
R7714 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t2 1.0925
R7715 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 1.0925
R7716 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t4 1.0925
R7717 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t13 0.8195
R7718 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t16 0.8195
R7719 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t14 0.8195
R7720 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t12 0.8195
R7721 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 0.314375
R7722 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 0.16025
R7723 a_n4631_31422.n1 a_n4631_31422.t9 41.0041
R7724 a_n4631_31422.n0 a_n4631_31422.t6 40.8177
R7725 a_n4631_31422.n2 a_n4631_31422.t5 40.6313
R7726 a_n4631_31422.n2 a_n4631_31422.t7 27.3166
R7727 a_n4631_31422.n0 a_n4631_31422.t8 27.1302
R7728 a_n4631_31422.n1 a_n4631_31422.t4 26.9438
R7729 a_n4631_31422.n3 a_n4631_31422.n1 15.6312
R7730 a_n4631_31422.n3 a_n4631_31422.n2 15.046
R7731 a_n4631_31422.n5 a_n4631_31422.t3 10.0473
R7732 a_n4631_31422.t0 a_n4631_31422.n7 6.51042
R7733 a_n4631_31422.n7 a_n4631_31422.n6 6.04952
R7734 a_n4631_31422.n4 a_n4631_31422.n0 5.64619
R7735 a_n4631_31422.n5 a_n4631_31422.n4 5.17851
R7736 a_n4631_31422.n4 a_n4631_31422.n3 4.5005
R7737 a_n4631_31422.n7 a_n4631_31422.n5 0.732092
R7738 a_n4631_31422.n6 a_n4631_31422.t2 0.7285
R7739 a_n4631_31422.n6 a_n4631_31422.t1 0.7285
R7740 a_n4631_33627.n2 a_n4631_33627.t4 40.6313
R7741 a_n4631_33627.n2 a_n4631_33627.t5 27.3166
R7742 a_n4631_33627.n3 a_n4631_33627.n2 24.1527
R7743 a_n4631_33627.t0 a_n4631_33627.n3 10.0473
R7744 a_n4631_33627.n1 a_n4631_33627.t1 6.51042
R7745 a_n4631_33627.n1 a_n4631_33627.n0 6.04952
R7746 a_n4631_33627.n3 a_n4631_33627.n1 0.732092
R7747 a_n4631_33627.n0 a_n4631_33627.t2 0.7285
R7748 a_n4631_33627.n0 a_n4631_33627.t3 0.7285
R7749 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t6 40.8177
R7750 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t7 40.6313
R7751 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t4 27.3166
R7752 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t5 27.1302
R7753 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_8.C.n2 14.119
R7754 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.t1 10.0473
R7755 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.t2 6.51042
R7756 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.n4 6.04952
R7757 SARlogic_0.dffrs_11.nand3_7.B SARlogic_0.dffrs_11.nand3_8.C.n0 5.47979
R7758 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C.n1 5.13907
R7759 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n6 4.72925
R7760 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.n5 0.732092
R7761 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t3 0.7285
R7762 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t0 0.7285
R7763 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_7.B 0.438233
R7764 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n3 0.166901
R7765 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C 0.0455
R7766 SAR_in.n9 SAR_in.t11 41.0041
R7767 SAR_in.n7 SAR_in.t6 41.0041
R7768 SAR_in.n5 SAR_in.t2 41.0041
R7769 SAR_in.n3 SAR_in.t8 41.0041
R7770 SAR_in.n1 SAR_in.t1 41.0041
R7771 SAR_in.n0 SAR_in.t7 41.0041
R7772 SAR_in.n9 SAR_in.t3 26.9438
R7773 SAR_in.n7 SAR_in.t9 26.9438
R7774 SAR_in.n5 SAR_in.t5 26.9438
R7775 SAR_in.n3 SAR_in.t0 26.9438
R7776 SAR_in.n1 SAR_in.t4 26.9438
R7777 SAR_in.n0 SAR_in.t10 26.9438
R7778 SAR_in.n2 SARlogic_0.dffrs_11.d 15.3544
R7779 SAR_in.n8 SARlogic_0.dffrs_7.d 11.7166
R7780 SAR_in.n6 SARlogic_0.dffrs_8.d 11.7166
R7781 SAR_in.n4 SARlogic_0.dffrs_9.d 11.7166
R7782 SAR_in.n2 SARlogic_0.dffrs_10.d 11.7166
R7783 SAR_in.n10 SARlogic_0.dffrs_14.d 11.6732
R7784 SARlogic_0.comp_in SAR_in.n10 7.63655
R7785 SARlogic_0.dffrs_14.nand3_8.A SAR_in.n9 5.7755
R7786 SARlogic_0.dffrs_7.nand3_8.A SAR_in.n7 5.7755
R7787 SARlogic_0.dffrs_8.nand3_8.A SAR_in.n5 5.7755
R7788 SARlogic_0.dffrs_9.nand3_8.A SAR_in.n3 5.7755
R7789 SARlogic_0.dffrs_10.nand3_8.A SAR_in.n1 5.7755
R7790 SARlogic_0.dffrs_11.nand3_8.A SAR_in.n0 5.7755
R7791 SAR_in.n4 SAR_in.n2 3.6383
R7792 SAR_in.n6 SAR_in.n4 3.6383
R7793 SAR_in.n8 SAR_in.n6 3.6383
R7794 SAR_in.n10 SAR_in.n8 3.6113
R7795 SARlogic_0.dffrs_14.d SARlogic_0.dffrs_14.nand3_8.A 0.784786
R7796 SARlogic_0.dffrs_7.d SARlogic_0.dffrs_7.nand3_8.A 0.784786
R7797 SARlogic_0.dffrs_8.d SARlogic_0.dffrs_8.nand3_8.A 0.784786
R7798 SARlogic_0.dffrs_9.d SARlogic_0.dffrs_9.nand3_8.A 0.784786
R7799 SARlogic_0.dffrs_10.d SARlogic_0.dffrs_10.nand3_8.A 0.784786
R7800 SARlogic_0.dffrs_11.d SARlogic_0.dffrs_11.nand3_8.A 0.784786
R7801 SARlogic_0.comp_in SAR_in 0.1775
R7802 a_n9861_31159.n0 a_n9861_31159.t4 34.1797
R7803 a_n9861_31159.n0 a_n9861_31159.t5 19.5798
R7804 a_n9861_31159.n3 a_n9861_31159.t0 18.7717
R7805 a_n9861_31159.t1 a_n9861_31159.n3 9.2885
R7806 a_n9861_31159.n2 a_n9861_31159.n0 4.93379
R7807 a_n9861_31159.n1 a_n9861_31159.t3 4.23346
R7808 a_n9861_31159.n1 a_n9861_31159.t2 3.85546
R7809 a_n9861_31159.n3 a_n9861_31159.n2 0.4055
R7810 a_n9861_31159.n2 a_n9861_31159.n1 0.352625
R7811 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t6 40.8177
R7812 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t7 40.6313
R7813 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t5 27.3166
R7814 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t4 27.1302
R7815 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_8.C.n2 14.119
R7816 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.t0 10.0473
R7817 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.t1 6.51042
R7818 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.n4 6.04952
R7819 SARlogic_0.dffrs_14.nand3_7.B SARlogic_0.dffrs_14.nand3_8.C.n0 5.47979
R7820 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C.n1 5.13907
R7821 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n6 4.72925
R7822 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.n5 0.732092
R7823 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t2 0.7285
R7824 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t3 0.7285
R7825 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_7.B 0.438233
R7826 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n3 0.166901
R7827 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C 0.0455
R7828 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t6 41.0041
R7829 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t7 40.8177
R7830 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t4 27.1302
R7831 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t5 26.9438
R7832 SARlogic_0.dffrs_13.nand3_6.A SARlogic_0.dffrs_13.nand3_0.B 17.0041
R7833 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n2 14.8493
R7834 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.t1 10.0473
R7835 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.t2 6.51042
R7836 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.n3 6.04952
R7837 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_8.Z.n0 5.7305
R7838 SARlogic_0.dffrs_13.nand3_0.B SARlogic_0.dffrs_13.nand3_8.Z.n1 5.47979
R7839 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n5 4.72925
R7840 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.n4 0.732092
R7841 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t3 0.7285
R7842 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t0 0.7285
R7843 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_6.A 0.0455
R7844 a_n389_31159.n0 a_n389_31159.t4 34.1797
R7845 a_n389_31159.n0 a_n389_31159.t5 19.5798
R7846 a_n389_31159.n1 a_n389_31159.t3 18.7717
R7847 a_n389_31159.n1 a_n389_31159.t2 9.2885
R7848 a_n389_31159.n2 a_n389_31159.n0 4.93379
R7849 a_n389_31159.t0 a_n389_31159.n3 4.23346
R7850 a_n389_31159.n3 a_n389_31159.t1 3.85546
R7851 a_n389_31159.n2 a_n389_31159.n1 0.4055
R7852 a_n389_31159.n3 a_n389_31159.n2 0.352625
R7853 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t5 40.8177
R7854 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t7 40.6313
R7855 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t4 27.3166
R7856 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t6 27.1302
R7857 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_8.C.n2 14.119
R7858 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.t1 10.0473
R7859 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.t0 6.51042
R7860 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.n4 6.04952
R7861 SARlogic_0.dffrs_9.nand3_7.B SARlogic_0.dffrs_9.nand3_8.C.n0 5.47979
R7862 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C.n1 5.13907
R7863 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n6 4.72925
R7864 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.n5 0.732092
R7865 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t2 0.7285
R7866 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t3 0.7285
R7867 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_7.B 0.438233
R7868 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n3 0.166901
R7869 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C 0.0455
R7870 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t6 41.0041
R7871 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t7 40.8177
R7872 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t4 40.6313
R7873 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t5 27.3166
R7874 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t8 27.1302
R7875 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t9 26.9438
R7876 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.t3 10.0473
R7877 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n4 9.90747
R7878 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n2 9.90116
R7879 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.t2 6.51042
R7880 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.n7 6.04952
R7881 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_6.C.n1 5.7305
R7882 SARlogic_0.dffrs_0.nand3_2.B SARlogic_0.dffrs_0.nand3_6.C.n0 5.47979
R7883 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C.n3 5.13907
R7884 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n9 4.72925
R7885 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_6.C.n5 4.5005
R7886 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.n8 0.732092
R7887 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t0 0.7285
R7888 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t1 0.7285
R7889 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n6 0.449758
R7890 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_2.B 0.166901
R7891 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_0.A 0.0455
R7892 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C 0.0455
R7893 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t6 40.8177
R7894 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t5 40.6313
R7895 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t7 27.3166
R7896 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t4 27.1302
R7897 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_8.C.n2 14.119
R7898 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.t0 10.0473
R7899 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.t1 6.51042
R7900 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.n4 6.04952
R7901 SARlogic_0.dffrs_0.nand3_7.B SARlogic_0.dffrs_0.nand3_8.C.n0 5.47979
R7902 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C.n1 5.13907
R7903 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n6 4.72925
R7904 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.n5 0.732092
R7905 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t3 0.7285
R7906 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t2 0.7285
R7907 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_7.B 0.438233
R7908 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n3 0.166901
R7909 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C 0.0455
R7910 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t7 41.0041
R7911 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t6 40.8177
R7912 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t5 40.6313
R7913 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t4 27.3166
R7914 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t8 27.1302
R7915 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t9 26.9438
R7916 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.t3 10.0473
R7917 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n4 9.90747
R7918 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n2 9.90116
R7919 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.t2 6.51042
R7920 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.n7 6.04952
R7921 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_6.C.n1 5.7305
R7922 SARlogic_0.dffrs_11.nand3_2.B SARlogic_0.dffrs_11.nand3_6.C.n0 5.47979
R7923 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C.n3 5.13907
R7924 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n9 4.72925
R7925 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_6.C.n5 4.5005
R7926 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.n8 0.732092
R7927 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t0 0.7285
R7928 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t1 0.7285
R7929 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n6 0.449758
R7930 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_2.B 0.166901
R7931 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_0.A 0.0455
R7932 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C 0.0455
R7933 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t4 41.0041
R7934 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t5 40.8177
R7935 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t9 40.6313
R7936 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t8 27.3166
R7937 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t7 27.1302
R7938 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t6 26.9438
R7939 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.t2 10.0473
R7940 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n4 9.90747
R7941 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n2 9.90116
R7942 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.t3 6.51042
R7943 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.n7 6.04952
R7944 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_6.C.n1 5.7305
R7945 SARlogic_0.dffrs_8.nand3_2.B SARlogic_0.dffrs_8.nand3_6.C.n0 5.47979
R7946 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C.n3 5.13907
R7947 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n9 4.72925
R7948 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_6.C.n5 4.5005
R7949 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.n8 0.732092
R7950 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t1 0.7285
R7951 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t0 0.7285
R7952 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n6 0.449758
R7953 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_2.B 0.166901
R7954 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_0.A 0.0455
R7955 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C 0.0455
R7956 a_n389_28819.n0 a_n389_28819.t5 34.1797
R7957 a_n389_28819.n0 a_n389_28819.t4 19.5798
R7958 a_n389_28819.n3 a_n389_28819.t3 18.7717
R7959 a_n389_28819.t0 a_n389_28819.n3 9.2885
R7960 a_n389_28819.n2 a_n389_28819.n0 4.93379
R7961 a_n389_28819.n1 a_n389_28819.t2 4.23346
R7962 a_n389_28819.n1 a_n389_28819.t1 3.85546
R7963 a_n389_28819.n3 a_n389_28819.n2 0.4055
R7964 a_n389_28819.n2 a_n389_28819.n1 0.352625
R7965 a_1839_29263.n0 a_1839_29263.t5 34.1797
R7966 a_1839_29263.n0 a_1839_29263.t4 19.5798
R7967 a_1839_29263.t0 a_1839_29263.n3 10.3401
R7968 a_1839_29263.n3 a_1839_29263.t1 9.2885
R7969 a_1839_29263.n2 a_1839_29263.n0 4.93379
R7970 a_1839_29263.n1 a_1839_29263.t2 4.09202
R7971 a_1839_29263.n1 a_1839_29263.t3 3.95079
R7972 a_1839_29263.n3 a_1839_29263.n2 0.599711
R7973 a_1839_29263.n2 a_1839_29263.n1 0.296375
R7974 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t4 40.6313
R7975 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t5 27.3166
R7976 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n1 14.2854
R7977 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.t1 10.0473
R7978 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.t2 6.51042
R7979 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.n2 6.04952
R7980 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C.n0 5.13907
R7981 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n4 4.72925
R7982 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.n3 0.732092
R7983 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t0 0.7285
R7984 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t3 0.7285
R7985 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C 0.0455
R7986 a_20783_29264.n0 a_20783_29264.t5 34.1797
R7987 a_20783_29264.n0 a_20783_29264.t4 19.5798
R7988 a_20783_29264.n1 a_20783_29264.t3 10.3401
R7989 a_20783_29264.n1 a_20783_29264.t2 9.2885
R7990 a_20783_29264.n2 a_20783_29264.n0 4.93379
R7991 a_20783_29264.t1 a_20783_29264.n3 4.09202
R7992 a_20783_29264.n3 a_20783_29264.t0 3.95079
R7993 a_20783_29264.n2 a_20783_29264.n1 0.599711
R7994 a_20783_29264.n3 a_20783_29264.n2 0.296375
R7995 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t8 40.6313
R7996 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.t6 34.1066
R7997 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t4 27.3166
R7998 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t7 19.673
R7999 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t5 19.4007
R8000 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n3 14.6967
R8001 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.t0 10.0473
R8002 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n6 9.39565
R8003 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit.n1 6.70486
R8004 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.t1 6.51042
R8005 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.n4 6.04952
R8006 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n2 5.81514
R8007 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.n5 0.732092
R8008 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t2 0.7285
R8009 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t3 0.7285
R8010 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n7 0.458082
R8011 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.n0 0.252687
R8012 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit 0.0519286
R8013 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_11.clk 44.4671
R8014 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t7 41.0041
R8015 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t6 40.8177
R8016 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t8 40.6313
R8017 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t5 27.3166
R8018 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t4 27.1302
R8019 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t9 26.9438
R8020 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_12.Q.n4 14.0582
R8021 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.t2 10.0473
R8022 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.t3 6.51042
R8023 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.n6 6.04952
R8024 SARlogic_0.dffrs_11.nand3_1.A SARlogic_0.dffrs_12.Q.n0 5.7755
R8025 SARlogic_0.dffrs_11.nand3_6.B SARlogic_0.dffrs_12.Q.n1 5.47979
R8026 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.Q.n3 5.13907
R8027 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n8 4.72925
R8028 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_6.B 2.17818
R8029 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_1.A 1.34729
R8030 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.n7 0.732092
R8031 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t0 0.7285
R8032 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t1 0.7285
R8033 SARlogic_0.dffrs_11.clk SARlogic_0.dffrs_12.Q.n2 0.610571
R8034 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n5 0.166901
R8035 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.nand3_7.C 0.0455
R8036 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t3 41.0041
R8037 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t2 26.9438
R8038 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t0 9.6935
R8039 adc_PISO_0.dffrs_1.d adc_PISO_0.2inmux_2.OUT.n0 6.55979
R8040 adc_PISO_0.2inmux_2.OUT adc_PISO_0.dffrs_1.d 4.883
R8041 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t1 4.35383
R8042 adc_PISO_0.2inmux_2.OUT adc_PISO_0.2inmux_2.OUT.n1 0.350857
R8043 a_4921_30169.n0 a_4921_30169.t5 41.0041
R8044 a_4921_30169.n1 a_4921_30169.t6 40.8177
R8045 a_4921_30169.n1 a_4921_30169.t4 27.1302
R8046 a_4921_30169.n0 a_4921_30169.t7 26.9438
R8047 a_4921_30169.n2 a_4921_30169.n1 22.5284
R8048 a_4921_30169.n3 a_4921_30169.n2 19.5781
R8049 a_4921_30169.n3 a_4921_30169.t1 10.0473
R8050 a_4921_30169.t0 a_4921_30169.n5 6.51042
R8051 a_4921_30169.n5 a_4921_30169.n4 6.04952
R8052 a_4921_30169.n2 a_4921_30169.n0 5.7305
R8053 a_4921_30169.n5 a_4921_30169.n3 0.732092
R8054 a_4921_30169.n4 a_4921_30169.t3 0.7285
R8055 a_4921_30169.n4 a_4921_30169.t2 0.7285
R8056 a_n4631_29217.n0 a_n4631_29217.t6 40.8177
R8057 a_n4631_29217.n1 a_n4631_29217.t5 40.6313
R8058 a_n4631_29217.n1 a_n4631_29217.t7 27.3166
R8059 a_n4631_29217.n0 a_n4631_29217.t4 27.1302
R8060 a_n4631_29217.n2 a_n4631_29217.n1 19.2576
R8061 a_n4631_29217.n3 a_n4631_29217.t2 10.0473
R8062 a_n4631_29217.n4 a_n4631_29217.t1 6.51042
R8063 a_n4631_29217.n5 a_n4631_29217.n4 6.04952
R8064 a_n4631_29217.n2 a_n4631_29217.n0 5.91752
R8065 a_n4631_29217.n3 a_n4631_29217.n2 4.89565
R8066 a_n4631_29217.n4 a_n4631_29217.n3 0.732092
R8067 a_n4631_29217.n5 a_n4631_29217.t3 0.7285
R8068 a_n4631_29217.t0 a_n4631_29217.n5 0.7285
R8069 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t6 41.0041
R8070 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t5 40.8177
R8071 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t4 40.6313
R8072 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t9 27.3166
R8073 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t7 27.1302
R8074 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t8 26.9438
R8075 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.t0 10.0473
R8076 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n4 9.90747
R8077 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n2 9.90116
R8078 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.t1 6.51042
R8079 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.n7 6.04952
R8080 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_6.C.n1 5.7305
R8081 SARlogic_0.dffrs_7.nand3_2.B SARlogic_0.dffrs_7.nand3_6.C.n0 5.47979
R8082 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C.n3 5.13907
R8083 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n9 4.72925
R8084 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_6.C.n5 4.5005
R8085 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.n8 0.732092
R8086 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t2 0.7285
R8087 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t3 0.7285
R8088 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n6 0.449758
R8089 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_2.B 0.166901
R8090 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_0.A 0.0455
R8091 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C 0.0455
R8092 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t2 41.0041
R8093 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t3 26.9438
R8094 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t1 9.6935
R8095 adc_PISO_0.dffrs_2.d adc_PISO_0.2inmux_3.OUT.n0 6.55979
R8096 adc_PISO_0.2inmux_3.OUT adc_PISO_0.dffrs_2.d 4.883
R8097 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t0 4.35383
R8098 adc_PISO_0.2inmux_3.OUT adc_PISO_0.2inmux_3.OUT.n1 0.350857
R8099 a_14393_30170.n2 a_14393_30170.t4 41.0041
R8100 a_14393_30170.n3 a_14393_30170.t6 40.8177
R8101 a_14393_30170.n3 a_14393_30170.t7 27.1302
R8102 a_14393_30170.n2 a_14393_30170.t5 26.9438
R8103 a_14393_30170.n4 a_14393_30170.n3 22.5284
R8104 a_14393_30170.n5 a_14393_30170.n4 19.5781
R8105 a_14393_30170.t0 a_14393_30170.n5 10.0473
R8106 a_14393_30170.n1 a_14393_30170.t1 6.51042
R8107 a_14393_30170.n1 a_14393_30170.n0 6.04952
R8108 a_14393_30170.n4 a_14393_30170.n2 5.7305
R8109 a_14393_30170.n5 a_14393_30170.n1 0.732092
R8110 a_14393_30170.n0 a_14393_30170.t3 0.7285
R8111 a_14393_30170.n0 a_14393_30170.t2 0.7285
R8112 Vin2.n7 Vin2.n6 23.1032
R8113 Vin2.n3 Vin2.n2 23.1032
R8114 Vin2.n0 Vin2.t6 22.8502
R8115 Vin2.n2 Vin2.t5 16.3656
R8116 Vin2.n6 Vin2.t1 16.3641
R8117 Vin2.n2 Vin2.t2 16.021
R8118 Vin2.n6 Vin2.t4 16.0195
R8119 Vin2.n8 Vin2.t8 11.5195
R8120 Vin2.n5 Vin2.t7 11.5195
R8121 Vin2.n4 Vin2.t0 11.5195
R8122 Vin2.n1 Vin2.t9 11.5195
R8123 Vin2.n0 Vin2.t3 11.5195
R8124 comparator_no_offsetcal_0.Vin2 Vin2 5.6819
R8125 comparator_no_offsetcal_0.Vin2 Vin2.n8 3.94555
R8126 Vin2.n7 Vin2.n5 2.53166
R8127 Vin2.n1 Vin2.n0 2.48408
R8128 Vin2.n3 Vin2.n1 1.40666
R8129 Vin2.n8 Vin2.n7 0.647658
R8130 Vin2.n4 Vin2.n3 0.647132
R8131 Vin2.n5 Vin2.n4 0.234605
R8132 Clk_piso.n19 Clk_piso.t9 41.0041
R8133 Clk_piso.n15 Clk_piso.t16 41.0041
R8134 Clk_piso.n11 Clk_piso.t6 41.0041
R8135 Clk_piso.n7 Clk_piso.t2 41.0041
R8136 Clk_piso.n3 Clk_piso.t0 41.0041
R8137 Clk_piso.n0 Clk_piso.t10 41.0041
R8138 Clk_piso.n20 Clk_piso.t13 40.8177
R8139 Clk_piso.n16 Clk_piso.t11 40.8177
R8140 Clk_piso.n12 Clk_piso.t3 40.8177
R8141 Clk_piso.n8 Clk_piso.t1 40.8177
R8142 Clk_piso.n4 Clk_piso.t15 40.8177
R8143 Clk_piso.n1 Clk_piso.t12 40.8177
R8144 Clk_piso.n20 Clk_piso.t21 27.1302
R8145 Clk_piso.n16 Clk_piso.t19 27.1302
R8146 Clk_piso.n12 Clk_piso.t8 27.1302
R8147 Clk_piso.n8 Clk_piso.t5 27.1302
R8148 Clk_piso.n4 Clk_piso.t22 27.1302
R8149 Clk_piso.n1 Clk_piso.t20 27.1302
R8150 Clk_piso.n19 Clk_piso.t17 26.9438
R8151 Clk_piso.n15 Clk_piso.t23 26.9438
R8152 Clk_piso.n11 Clk_piso.t14 26.9438
R8153 Clk_piso.n7 Clk_piso.t7 26.9438
R8154 Clk_piso.n3 Clk_piso.t4 26.9438
R8155 Clk_piso.n0 Clk_piso.t18 26.9438
R8156 Clk_piso.n6 adc_PISO_0.dffrs_5.clk 23.2034
R8157 Clk_piso.n22 Clk_piso.n18 13.9468
R8158 Clk_piso.n18 Clk_piso.n14 13.9463
R8159 Clk_piso.n10 Clk_piso.n6 13.9457
R8160 Clk_piso.n14 Clk_piso.n10 13.9457
R8161 Clk_piso.n23 Clk_piso 13.1341
R8162 Clk_piso.n22 adc_PISO_0.dffrs_0.clk 9.25764
R8163 Clk_piso.n18 adc_PISO_0.dffrs_1.clk 9.25764
R8164 Clk_piso.n14 adc_PISO_0.dffrs_2.clk 9.25764
R8165 Clk_piso.n10 adc_PISO_0.dffrs_3.clk 9.25764
R8166 Clk_piso.n6 adc_PISO_0.dffrs_4.clk 9.25764
R8167 Clk_piso.n21 Clk_piso.n20 7.65746
R8168 Clk_piso.n17 Clk_piso.n16 7.65746
R8169 Clk_piso.n13 Clk_piso.n12 7.65746
R8170 Clk_piso.n9 Clk_piso.n8 7.65746
R8171 Clk_piso.n5 Clk_piso.n4 7.65746
R8172 Clk_piso.n2 Clk_piso.n1 7.65746
R8173 Clk_piso.n21 Clk_piso.n19 7.12229
R8174 Clk_piso.n17 Clk_piso.n15 7.12229
R8175 Clk_piso.n13 Clk_piso.n11 7.12229
R8176 Clk_piso.n9 Clk_piso.n7 7.12229
R8177 Clk_piso.n5 Clk_piso.n3 7.12229
R8178 Clk_piso.n2 Clk_piso.n0 7.12229
R8179 Clk_piso.n23 Clk_piso.n22 3.49505
R8180 adc_PISO_0.dffrs_0.clk Clk_piso.n21 0.611214
R8181 adc_PISO_0.dffrs_1.clk Clk_piso.n17 0.611214
R8182 adc_PISO_0.dffrs_2.clk Clk_piso.n13 0.611214
R8183 adc_PISO_0.dffrs_3.clk Clk_piso.n9 0.611214
R8184 adc_PISO_0.dffrs_4.clk Clk_piso.n5 0.611214
R8185 adc_PISO_0.dffrs_5.clk Clk_piso.n2 0.611214
R8186 adc_PISO_0.clk Clk_piso.n23 0.0336579
R8187 a_14313_29218.n2 a_14313_29218.t6 40.8177
R8188 a_14313_29218.n3 a_14313_29218.t5 40.6313
R8189 a_14313_29218.n3 a_14313_29218.t4 27.3166
R8190 a_14313_29218.n2 a_14313_29218.t7 27.1302
R8191 a_14313_29218.n4 a_14313_29218.n3 19.2576
R8192 a_14313_29218.t0 a_14313_29218.n5 10.0473
R8193 a_14313_29218.n1 a_14313_29218.t1 6.51042
R8194 a_14313_29218.n1 a_14313_29218.n0 6.04952
R8195 a_14313_29218.n4 a_14313_29218.n2 5.91752
R8196 a_14313_29218.n5 a_14313_29218.n4 4.89565
R8197 a_14313_29218.n5 a_14313_29218.n1 0.732092
R8198 a_14313_29218.n0 a_14313_29218.t3 0.7285
R8199 a_14313_29218.n0 a_14313_29218.t2 0.7285
R8200 a_4841_29217.n2 a_4841_29217.t6 40.8177
R8201 a_4841_29217.n3 a_4841_29217.t5 40.6313
R8202 a_4841_29217.n3 a_4841_29217.t7 27.3166
R8203 a_4841_29217.n2 a_4841_29217.t4 27.1302
R8204 a_4841_29217.n4 a_4841_29217.n3 19.2576
R8205 a_4841_29217.t0 a_4841_29217.n5 10.0473
R8206 a_4841_29217.n1 a_4841_29217.t1 6.51042
R8207 a_4841_29217.n1 a_4841_29217.n0 6.04952
R8208 a_4841_29217.n4 a_4841_29217.n2 5.91752
R8209 a_4841_29217.n5 a_4841_29217.n4 4.89565
R8210 a_4841_29217.n5 a_4841_29217.n1 0.732092
R8211 a_4841_29217.n0 a_4841_29217.t3 0.7285
R8212 a_4841_29217.n0 a_4841_29217.t2 0.7285
R8213 SARlogic_0.d4.n3 SARlogic_0.d4.t11 41.0041
R8214 SARlogic_0.d4.n4 SARlogic_0.d4.t12 40.8177
R8215 SARlogic_0.d4.n7 SARlogic_0.d4.t7 40.6313
R8216 SARlogic_0.d4.n1 SARlogic_0.d4.t10 34.2529
R8217 SARlogic_0.d4.n6 SARlogic_0.dffrs_14.clk 33.675
R8218 SARlogic_0.d4.n7 SARlogic_0.d4.t5 27.3166
R8219 SARlogic_0.d4.n4 SARlogic_0.d4.t8 27.1302
R8220 SARlogic_0.d4.n3 SARlogic_0.d4.t4 26.9438
R8221 SARlogic_0.d4.n0 SARlogic_0.d4.t6 19.673
R8222 SARlogic_0.d4.n0 SARlogic_0.d4.t9 19.4007
R8223 SARlogic_0.d4.n9 SARlogic_0.d4.n8 14.0582
R8224 SARlogic_0.d4.n9 SARlogic_0.d4.n6 11.3593
R8225 SARlogic_0.d4.n12 SARlogic_0.d4.t0 10.0473
R8226 SARlogic_0.d4.n2 SARlogic_0.d4.n1 8.05164
R8227 SARlogic_0.d4.n11 SARlogic_0.d4.t1 6.51042
R8228 SARlogic_0.d4.n11 SARlogic_0.d4.n10 6.04952
R8229 SARlogic_0.dffrs_14.nand3_1.A SARlogic_0.d4.n3 5.7755
R8230 SARlogic_0.dffrs_14.nand3_6.B SARlogic_0.d4.n4 5.47979
R8231 SARlogic_0.d4.n8 SARlogic_0.d4.n7 5.13907
R8232 SARlogic_0.dffrs_7.nand3_2.Z SARlogic_0.d4.n12 4.72925
R8233 SARlogic_0.d4.n6 adc_PISO_0.B5 3.49604
R8234 SARlogic_0.d4.n5 SARlogic_0.dffrs_14.nand3_6.B 2.17818
R8235 adc_PISO_0.B5 SARlogic_0.d4.n2 1.87121
R8236 SARlogic_0.d4.n5 SARlogic_0.dffrs_14.nand3_1.A 1.34729
R8237 SARlogic_0.d4.n12 SARlogic_0.d4.n11 0.732092
R8238 SARlogic_0.d4.n10 SARlogic_0.d4.t3 0.7285
R8239 SARlogic_0.d4.n10 SARlogic_0.d4.t2 0.7285
R8240 SARlogic_0.dffrs_14.clk SARlogic_0.d4.n5 0.611214
R8241 SARlogic_0.dffrs_7.nand3_2.Z SARlogic_0.d4.n9 0.166901
R8242 SARlogic_0.d4.n1 SARlogic_0.d4.n0 0.106438
R8243 SARlogic_0.d4.n8 SARlogic_0.dffrs_7.nand3_7.C 0.0455
R8244 SARlogic_0.d4.n2 adc_PISO_0.2inmux_2.In 0.0455
R8245 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t5 41.0041
R8246 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t7 40.6313
R8247 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t8 40.6313
R8248 SARlogic_0.dffrs_4.Qb SARlogic_0.dffrs_11.setb 28.021
R8249 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t9 27.3166
R8250 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t4 27.3166
R8251 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t6 26.9438
R8252 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.t1 10.0473
R8253 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb.n1 9.84255
R8254 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n3 9.22229
R8255 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.t2 6.51042
R8256 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.n7 6.04952
R8257 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.Qb.n0 5.7305
R8258 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n4 5.14711
R8259 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_4.Qb.n2 5.13907
R8260 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n6 4.94976
R8261 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n9 4.72925
R8262 SARlogic_0.dffrs_11.setb SARlogic_0.dffrs_11.nand3_0.C 0.784786
R8263 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.n8 0.732092
R8264 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t3 0.7285
R8265 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t0 0.7285
R8266 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb 0.175225
R8267 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.nand3_2.A 0.0455
R8268 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_11.nand3_2.C 0.0455
R8269 SARlogic_0.dffrs_11.nand3_0.C SARlogic_0.dffrs_4.Qb.n5 0.0374643
R8270 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t6 40.8177
R8271 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t5 40.6313
R8272 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t7 27.3166
R8273 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t4 27.1302
R8274 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_8.C.n2 14.119
R8275 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.t1 10.0473
R8276 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.t2 6.51042
R8277 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.n4 6.04952
R8278 SARlogic_0.dffrs_8.nand3_7.B SARlogic_0.dffrs_8.nand3_8.C.n0 5.47979
R8279 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C.n1 5.13907
R8280 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n6 4.72925
R8281 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.n5 0.732092
R8282 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t3 0.7285
R8283 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t0 0.7285
R8284 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_7.B 0.438233
R8285 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n3 0.166901
R8286 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C 0.0455
R8287 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t5 41.0041
R8288 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t6 40.8177
R8289 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t4 27.1302
R8290 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t7 26.9438
R8291 SARlogic_0.dffrs_2.nand3_6.A SARlogic_0.dffrs_2.nand3_0.B 17.0041
R8292 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n2 14.8493
R8293 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.t1 10.0473
R8294 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.t0 6.51042
R8295 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.n3 6.04952
R8296 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_8.Z.n0 5.7305
R8297 SARlogic_0.dffrs_2.nand3_0.B SARlogic_0.dffrs_2.nand3_8.Z.n1 5.47979
R8298 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n5 4.72925
R8299 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.n4 0.732092
R8300 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t2 0.7285
R8301 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t3 0.7285
R8302 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_6.A 0.0455
R8303 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t5 40.6313
R8304 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.t6 34.1066
R8305 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t7 27.3166
R8306 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t8 19.673
R8307 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t4 19.4007
R8308 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n3 14.6967
R8309 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.t1 10.0473
R8310 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n6 9.39565
R8311 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.dffrs_3.Q.n1 6.70486
R8312 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.t2 6.51042
R8313 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.n4 6.04952
R8314 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n2 5.81514
R8315 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.n5 0.732092
R8316 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t0 0.7285
R8317 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t3 0.7285
R8318 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n7 0.458082
R8319 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.n0 0.252687
R8320 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.2inmux_5.Bit 0.0519286
R8321 a_39727_29264.n0 a_39727_29264.t5 34.1797
R8322 a_39727_29264.n0 a_39727_29264.t4 19.5798
R8323 a_39727_29264.n3 a_39727_29264.t3 10.3401
R8324 a_39727_29264.t0 a_39727_29264.n3 9.2885
R8325 a_39727_29264.n2 a_39727_29264.n0 4.93379
R8326 a_39727_29264.n1 a_39727_29264.t1 4.09202
R8327 a_39727_29264.n1 a_39727_29264.t2 3.95079
R8328 a_39727_29264.n3 a_39727_29264.n2 0.599711
R8329 a_39727_29264.n2 a_39727_29264.n1 0.296375
R8330 a_42809_30170.n0 a_42809_30170.t5 41.0041
R8331 a_42809_30170.n1 a_42809_30170.t7 40.8177
R8332 a_42809_30170.n1 a_42809_30170.t4 27.1302
R8333 a_42809_30170.n0 a_42809_30170.t6 26.9438
R8334 a_42809_30170.n2 a_42809_30170.n1 22.5284
R8335 a_42809_30170.n3 a_42809_30170.n2 19.5781
R8336 a_42809_30170.n3 a_42809_30170.t3 10.0473
R8337 a_42809_30170.n4 a_42809_30170.t2 6.51042
R8338 a_42809_30170.n5 a_42809_30170.n4 6.04952
R8339 a_42809_30170.n2 a_42809_30170.n0 5.7305
R8340 a_42809_30170.n4 a_42809_30170.n3 0.732092
R8341 a_42809_30170.n5 a_42809_30170.t1 0.7285
R8342 a_42809_30170.t0 a_42809_30170.n5 0.7285
R8343 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t7 40.8177
R8344 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t5 40.6313
R8345 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t6 27.3166
R8346 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t4 27.1302
R8347 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_8.C.n2 14.119
R8348 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.t0 10.0473
R8349 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.t1 6.51042
R8350 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.n4 6.04952
R8351 SARlogic_0.dffrs_10.nand3_7.B SARlogic_0.dffrs_10.nand3_8.C.n0 5.47979
R8352 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C.n1 5.13907
R8353 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n6 4.72925
R8354 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.n5 0.732092
R8355 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t3 0.7285
R8356 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t2 0.7285
R8357 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_7.B 0.438233
R8358 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n3 0.166901
R8359 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C 0.0455
R8360 adc_PISO_0.serial_out.n0 adc_PISO_0.serial_out.t6 45.6255
R8361 adc_PISO_0.serial_out.n1 adc_PISO_0.serial_out.t7 40.6313
R8362 adc_PISO_0.serial_out.n1 adc_PISO_0.serial_out.t4 27.3166
R8363 adc_PISO_0.serial_out.n0 adc_PISO_0.serial_out.t5 20.6838
R8364 adc_PISO_0.serial_out.n5 adc_PISO_0.serial_out.n1 14.6967
R8365 osu_sc_buf_4_flat_0.A adc_PISO_0.serial_out.n0 12.5005
R8366 adc_PISO_0.serial_out.n4 adc_PISO_0.serial_out.t0 10.0473
R8367 adc_PISO_0.serial_out.n5 adc_PISO_0.serial_out.n4 9.39565
R8368 adc_PISO_0.serial_out osu_sc_buf_4_flat_0.A 9.18361
R8369 adc_PISO_0.serial_out.n3 adc_PISO_0.serial_out.t1 6.51042
R8370 adc_PISO_0.serial_out.n3 adc_PISO_0.serial_out.n2 6.04952
R8371 adc_PISO_0.dffrs_5.Q adc_PISO_0.serial_out 5.90514
R8372 adc_PISO_0.serial_out.n4 adc_PISO_0.serial_out.n3 0.732092
R8373 adc_PISO_0.serial_out.n2 adc_PISO_0.serial_out.t2 0.7285
R8374 adc_PISO_0.serial_out.n2 adc_PISO_0.serial_out.t3 0.7285
R8375 adc_PISO_0.dffrs_5.Q adc_PISO_0.serial_out.n5 0.458082
R8376 a_n4551_30169.n0 a_n4551_30169.t5 41.0041
R8377 a_n4551_30169.n1 a_n4551_30169.t7 40.8177
R8378 a_n4551_30169.n1 a_n4551_30169.t4 27.1302
R8379 a_n4551_30169.n0 a_n4551_30169.t6 26.9438
R8380 a_n4551_30169.n2 a_n4551_30169.n1 22.5284
R8381 a_n4551_30169.n3 a_n4551_30169.n2 19.5781
R8382 a_n4551_30169.n3 a_n4551_30169.t1 10.0473
R8383 a_n4551_30169.t0 a_n4551_30169.n5 6.51042
R8384 a_n4551_30169.n5 a_n4551_30169.n4 6.04952
R8385 a_n4551_30169.n2 a_n4551_30169.n0 5.7305
R8386 a_n4551_30169.n5 a_n4551_30169.n3 0.732092
R8387 a_n4551_30169.n4 a_n4551_30169.t2 0.7285
R8388 a_n4551_30169.n4 a_n4551_30169.t3 0.7285
R8389 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t4 41.0041
R8390 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t5 40.8177
R8391 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t7 27.1302
R8392 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t6 26.9438
R8393 SARlogic_0.dffrs_0.nand3_6.A SARlogic_0.dffrs_0.nand3_0.B 17.0041
R8394 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n2 14.8493
R8395 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.t2 10.0473
R8396 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.t3 6.51042
R8397 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.n3 6.04952
R8398 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_8.Z.n0 5.7305
R8399 SARlogic_0.dffrs_0.nand3_0.B SARlogic_0.dffrs_0.nand3_8.Z.n1 5.47979
R8400 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n5 4.72925
R8401 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.n4 0.732092
R8402 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t1 0.7285
R8403 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t0 0.7285
R8404 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_6.A 0.0455
R8405 a_11311_29264.n0 a_11311_29264.t5 34.1797
R8406 a_11311_29264.n0 a_11311_29264.t4 19.5798
R8407 a_11311_29264.n3 a_11311_29264.t3 10.3401
R8408 a_11311_29264.t0 a_11311_29264.n3 9.2885
R8409 a_11311_29264.n2 a_11311_29264.n0 4.93379
R8410 a_11311_29264.n1 a_11311_29264.t2 4.09202
R8411 a_11311_29264.n1 a_11311_29264.t1 3.95079
R8412 a_11311_29264.n3 a_11311_29264.n2 0.599711
R8413 a_11311_29264.n2 a_11311_29264.n1 0.296375
R8414 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t7 41.0041
R8415 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t4 40.8177
R8416 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t5 27.1302
R8417 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t6 26.9438
R8418 SARlogic_0.dffrs_5.nand3_6.A SARlogic_0.dffrs_5.nand3_0.B 17.0041
R8419 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n2 14.8493
R8420 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.t1 10.0473
R8421 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.t0 6.51042
R8422 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.n3 6.04952
R8423 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_8.Z.n0 5.7305
R8424 SARlogic_0.dffrs_5.nand3_0.B SARlogic_0.dffrs_5.nand3_8.Z.n1 5.47979
R8425 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n5 4.72925
R8426 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.n4 0.732092
R8427 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t2 0.7285
R8428 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t3 0.7285
R8429 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_6.A 0.0455
R8430 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t7 40.8177
R8431 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t5 40.6313
R8432 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t6 27.3166
R8433 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t4 27.1302
R8434 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_8.C.n2 14.119
R8435 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.t1 10.0473
R8436 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.t2 6.51042
R8437 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.n4 6.04952
R8438 SARlogic_0.dffrs_13.nand3_7.B SARlogic_0.dffrs_13.nand3_8.C.n0 5.47979
R8439 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C.n1 5.13907
R8440 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n6 4.72925
R8441 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.n5 0.732092
R8442 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t0 0.7285
R8443 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t3 0.7285
R8444 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_7.B 0.438233
R8445 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n3 0.166901
R8446 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C 0.0455
R8447 a_n7633_29263.n0 a_n7633_29263.t4 34.1797
R8448 a_n7633_29263.n0 a_n7633_29263.t5 19.5798
R8449 a_n7633_29263.t0 a_n7633_29263.n3 10.3401
R8450 a_n7633_29263.n3 a_n7633_29263.t1 9.2885
R8451 a_n7633_29263.n2 a_n7633_29263.n0 4.93379
R8452 a_n7633_29263.n1 a_n7633_29263.t2 4.09202
R8453 a_n7633_29263.n1 a_n7633_29263.t3 3.95079
R8454 a_n7633_29263.n3 a_n7633_29263.n2 0.599711
R8455 a_n7633_29263.n2 a_n7633_29263.n1 0.296375
R8456 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t2 41.0041
R8457 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t3 26.9438
R8458 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t0 9.6935
R8459 adc_PISO_0.dffrs_0.d adc_PISO_0.2inmux_0.OUT.n0 6.55979
R8460 adc_PISO_0.2inmux_0.OUT adc_PISO_0.dffrs_0.d 4.883
R8461 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t1 4.35383
R8462 adc_PISO_0.2inmux_0.OUT adc_PISO_0.2inmux_0.OUT.n1 0.350857
R8463 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t4 41.0041
R8464 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t6 40.6313
R8465 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t7 27.3166
R8466 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t5 26.9438
R8467 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_5.d 17.5382
R8468 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_4.Q.n2 14.0582
R8469 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.t1 10.0473
R8470 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.t2 6.51042
R8471 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.n4 6.04952
R8472 SARlogic_0.dffrs_5.nand3_8.A SARlogic_0.dffrs_4.Q.n0 5.7755
R8473 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.Q.n1 5.13907
R8474 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n6 4.72925
R8475 SARlogic_0.dffrs_5.d SARlogic_0.dffrs_5.nand3_8.A 0.784786
R8476 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.n5 0.732092
R8477 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t0 0.7285
R8478 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t3 0.7285
R8479 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n3 0.166901
R8480 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.nand3_7.C 0.0455
R8481 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t4 41.0041
R8482 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t7 40.6313
R8483 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t6 27.3166
R8484 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t5 26.9438
R8485 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_1.d 17.5382
R8486 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_0.Q.n2 14.0582
R8487 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.t2 10.0473
R8488 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.t3 6.51042
R8489 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.n4 6.04952
R8490 SARlogic_0.dffrs_1.nand3_8.A SARlogic_0.dffrs_0.Q.n0 5.7755
R8491 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.Q.n1 5.13907
R8492 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n6 4.72925
R8493 SARlogic_0.dffrs_1.d SARlogic_0.dffrs_1.nand3_8.A 0.784786
R8494 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.n5 0.732092
R8495 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t0 0.7285
R8496 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t1 0.7285
R8497 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n3 0.166901
R8498 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.nand3_7.C 0.0455
R8499 a_18555_28820.n0 a_18555_28820.t5 34.1797
R8500 a_18555_28820.n0 a_18555_28820.t4 19.5798
R8501 a_18555_28820.n1 a_18555_28820.t2 18.7717
R8502 a_18555_28820.n1 a_18555_28820.t1 9.2885
R8503 a_18555_28820.n2 a_18555_28820.n0 4.93379
R8504 a_18555_28820.t0 a_18555_28820.n3 4.23346
R8505 a_18555_28820.n3 a_18555_28820.t3 3.85546
R8506 a_18555_28820.n2 a_18555_28820.n1 0.4055
R8507 a_18555_28820.n3 a_18555_28820.n2 0.352625
R8508 a_23785_33628.n0 a_23785_33628.t4 40.6313
R8509 a_23785_33628.n0 a_23785_33628.t5 27.3166
R8510 a_23785_33628.n1 a_23785_33628.n0 24.1527
R8511 a_23785_33628.n1 a_23785_33628.t1 10.0473
R8512 a_23785_33628.t0 a_23785_33628.n3 6.51042
R8513 a_23785_33628.n3 a_23785_33628.n2 6.04952
R8514 a_23785_33628.n3 a_23785_33628.n1 0.732092
R8515 a_23785_33628.n2 a_23785_33628.t3 0.7285
R8516 a_23785_33628.n2 a_23785_33628.t2 0.7285
R8517 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t6 41.0041
R8518 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t5 40.8177
R8519 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t4 27.1302
R8520 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t7 26.9438
R8521 SARlogic_0.dffrs_1.nand3_6.A SARlogic_0.dffrs_1.nand3_0.B 17.0041
R8522 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n2 14.8493
R8523 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.t1 10.0473
R8524 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.t2 6.51042
R8525 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.n3 6.04952
R8526 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_8.Z.n0 5.7305
R8527 SARlogic_0.dffrs_1.nand3_0.B SARlogic_0.dffrs_1.nand3_8.Z.n1 5.47979
R8528 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n5 4.72925
R8529 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.n4 0.732092
R8530 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t0 0.7285
R8531 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t3 0.7285
R8532 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_6.A 0.0455
R8533 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t4 41.0041
R8534 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t7 40.6313
R8535 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t6 27.3166
R8536 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t5 26.9438
R8537 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d 17.5382
R8538 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d.n2 14.0582
R8539 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.t2 10.0473
R8540 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.t3 6.51042
R8541 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.n4 6.04952
R8542 SARlogic_0.dffrs_2.nand3_8.A SARlogic_0.dffrs_2.d.n0 5.7755
R8543 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_2.d.n1 5.13907
R8544 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n6 4.72925
R8545 SARlogic_0.dffrs_2.d SARlogic_0.dffrs_2.nand3_8.A 0.784786
R8546 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.n5 0.732092
R8547 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t1 0.7285
R8548 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t0 0.7285
R8549 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n3 0.166901
R8550 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_1.nand3_7.C 0.0455
R8551 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t5 40.6313
R8552 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t4 27.3166
R8553 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n1 14.2246
R8554 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.t0 10.0473
R8555 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.t1 6.51042
R8556 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.n2 6.04952
R8557 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.Q.n0 5.13907
R8558 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n4 4.72925
R8559 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.n3 0.732092
R8560 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t2 0.7285
R8561 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t3 0.7285
R8562 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.nand3_7.C 0.0455
R8563 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t5 41.0041
R8564 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t6 40.8177
R8565 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t4 40.6313
R8566 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t7 27.3166
R8567 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t8 27.1302
R8568 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t9 26.9438
R8569 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.t2 10.0473
R8570 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n4 9.90747
R8571 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n2 9.90116
R8572 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.t3 6.51042
R8573 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.n7 6.04952
R8574 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_6.C.n1 5.7305
R8575 SARlogic_0.dffrs_4.nand3_2.B SARlogic_0.dffrs_4.nand3_6.C.n0 5.47979
R8576 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C.n3 5.13907
R8577 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n9 4.72925
R8578 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_6.C.n5 4.5005
R8579 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.n8 0.732092
R8580 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t0 0.7285
R8581 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t1 0.7285
R8582 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n6 0.449758
R8583 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_2.B 0.166901
R8584 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_0.A 0.0455
R8585 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C 0.0455
R8586 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t2 41.0041
R8587 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t3 26.9438
R8588 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t0 9.6935
R8589 adc_PISO_0.dffrs_5.d adc_PISO_0.2inmux_1.OUT.n0 6.55979
R8590 adc_PISO_0.2inmux_1.OUT adc_PISO_0.dffrs_5.d 4.883
R8591 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t1 4.35383
R8592 adc_PISO_0.2inmux_1.OUT adc_PISO_0.2inmux_1.OUT.n1 0.350857
R8593 Load.n0 Load.t1 34.1797
R8594 Load.n0 Load.t0 19.5798
R8595 inv2_0.in Load.n0 4.87271
R8596 inv2_0.in Load 0.868357
R8597 a_42729_29218.n2 a_42729_29218.t5 40.8177
R8598 a_42729_29218.n3 a_42729_29218.t6 40.6313
R8599 a_42729_29218.n3 a_42729_29218.t4 27.3166
R8600 a_42729_29218.n2 a_42729_29218.t7 27.1302
R8601 a_42729_29218.n4 a_42729_29218.n3 19.2576
R8602 a_42729_29218.t0 a_42729_29218.n5 10.0473
R8603 a_42729_29218.n1 a_42729_29218.t1 6.51042
R8604 a_42729_29218.n1 a_42729_29218.n0 6.04952
R8605 a_42729_29218.n4 a_42729_29218.n2 5.91752
R8606 a_42729_29218.n5 a_42729_29218.n4 4.89565
R8607 a_42729_29218.n5 a_42729_29218.n1 0.732092
R8608 a_42729_29218.n0 a_42729_29218.t3 0.7285
R8609 a_42729_29218.n0 a_42729_29218.t2 0.7285
R8610 a_18555_31160.n0 a_18555_31160.t5 34.1797
R8611 a_18555_31160.n0 a_18555_31160.t4 19.5798
R8612 a_18555_31160.n3 a_18555_31160.t0 18.7717
R8613 a_18555_31160.t1 a_18555_31160.n3 9.2885
R8614 a_18555_31160.n2 a_18555_31160.n0 4.93379
R8615 a_18555_31160.n1 a_18555_31160.t3 4.23346
R8616 a_18555_31160.n1 a_18555_31160.t2 3.85546
R8617 a_18555_31160.n3 a_18555_31160.n2 0.4055
R8618 a_18555_31160.n2 a_18555_31160.n1 0.352625
R8619 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t7 41.0041
R8620 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t5 40.8177
R8621 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t6 40.6313
R8622 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t9 27.3166
R8623 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t8 27.1302
R8624 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t4 26.9438
R8625 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.t2 10.0473
R8626 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n4 9.90747
R8627 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n2 9.90116
R8628 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.t3 6.51042
R8629 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.n7 6.04952
R8630 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_6.C.n1 5.7305
R8631 SARlogic_0.dffrs_13.nand3_2.B SARlogic_0.dffrs_13.nand3_6.C.n0 5.47979
R8632 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C.n3 5.13907
R8633 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n9 4.72925
R8634 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_6.C.n5 4.5005
R8635 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.n8 0.732092
R8636 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t1 0.7285
R8637 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t0 0.7285
R8638 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n6 0.449758
R8639 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_2.B 0.166901
R8640 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_0.A 0.0455
R8641 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C 0.0455
R8642 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t4 40.6313
R8643 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t5 27.3166
R8644 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n1 14.2854
R8645 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.t1 10.0473
R8646 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.t2 6.51042
R8647 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.n2 6.04952
R8648 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C.n0 5.13907
R8649 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n4 4.72925
R8650 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.n3 0.732092
R8651 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t3 0.7285
R8652 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t0 0.7285
R8653 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C 0.0455
R8654 a_n9861_28819.n0 a_n9861_28819.t5 34.1797
R8655 a_n9861_28819.n0 a_n9861_28819.t4 19.5798
R8656 a_n9861_28819.n1 a_n9861_28819.t1 18.7717
R8657 a_n9861_28819.n1 a_n9861_28819.t2 9.2885
R8658 a_n9861_28819.n2 a_n9861_28819.n0 4.93379
R8659 a_n9861_28819.t0 a_n9861_28819.n3 4.23346
R8660 a_n9861_28819.n3 a_n9861_28819.t3 3.85546
R8661 a_n9861_28819.n2 a_n9861_28819.n1 0.4055
R8662 a_n9861_28819.n3 a_n9861_28819.n2 0.352625
R8663 a_37499_28820.n0 a_37499_28820.t5 34.1797
R8664 a_37499_28820.n0 a_37499_28820.t4 19.5798
R8665 a_37499_28820.n1 a_37499_28820.t1 18.7717
R8666 a_37499_28820.n1 a_37499_28820.t2 9.2885
R8667 a_37499_28820.n2 a_37499_28820.n0 4.93379
R8668 a_37499_28820.t0 a_37499_28820.n3 4.23346
R8669 a_37499_28820.n3 a_37499_28820.t3 3.85546
R8670 a_37499_28820.n2 a_37499_28820.n1 0.4055
R8671 a_37499_28820.n3 a_37499_28820.n2 0.352625
R8672 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t4 40.6313
R8673 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t5 27.3166
R8674 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n1 14.2854
R8675 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.t2 10.0473
R8676 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.t3 6.51042
R8677 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.n2 6.04952
R8678 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C.n0 5.13907
R8679 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n4 4.72925
R8680 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.n3 0.732092
R8681 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t1 0.7285
R8682 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t0 0.7285
R8683 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C 0.0455
R8684 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t5 41.0041
R8685 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t6 40.6313
R8686 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t4 27.3166
R8687 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t7 26.9438
R8688 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_3.d 17.5382
R8689 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_2.Q.n2 14.0582
R8690 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.t3 10.0473
R8691 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.t2 6.51042
R8692 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.n4 6.04952
R8693 SARlogic_0.dffrs_3.nand3_8.A SARlogic_0.dffrs_2.Q.n0 5.7755
R8694 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.Q.n1 5.13907
R8695 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n6 4.72925
R8696 SARlogic_0.dffrs_3.d SARlogic_0.dffrs_3.nand3_8.A 0.784786
R8697 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.n5 0.732092
R8698 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t0 0.7285
R8699 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t1 0.7285
R8700 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n3 0.166901
R8701 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.nand3_7.C 0.0455
R8702 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t6 40.6313
R8703 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.t5 34.1066
R8704 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t7 27.3166
R8705 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t8 19.673
R8706 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t4 19.4007
R8707 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n3 14.6967
R8708 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.t0 10.0473
R8709 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n6 9.39565
R8710 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.dffrs_2.Q.n1 6.70486
R8711 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.t1 6.51042
R8712 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.n4 6.04952
R8713 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n2 5.81514
R8714 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.n5 0.732092
R8715 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t3 0.7285
R8716 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t2 0.7285
R8717 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n7 0.458082
R8718 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.n0 0.252687
R8719 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.2inmux_4.Bit 0.0519286
R8720 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t4 40.6313
R8721 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t5 27.3166
R8722 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n1 14.2854
R8723 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.t2 10.0473
R8724 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.t3 6.51042
R8725 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.n2 6.04952
R8726 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C.n0 5.13907
R8727 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n4 4.72925
R8728 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.n3 0.732092
R8729 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t0 0.7285
R8730 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t1 0.7285
R8731 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C 0.0455
R8732 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t3 41.0041
R8733 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t2 26.9438
R8734 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t0 9.6935
R8735 adc_PISO_0.dffrs_3.d adc_PISO_0.2inmux_4.OUT.n0 6.55979
R8736 adc_PISO_0.2inmux_4.OUT adc_PISO_0.dffrs_3.d 4.883
R8737 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t1 4.35383
R8738 adc_PISO_0.2inmux_4.OUT adc_PISO_0.2inmux_4.OUT.n1 0.350857
R8739 a_14313_31423.n1 a_14313_31423.t4 41.0041
R8740 a_14313_31423.n0 a_14313_31423.t6 40.8177
R8741 a_14313_31423.n2 a_14313_31423.t5 40.6313
R8742 a_14313_31423.n2 a_14313_31423.t8 27.3166
R8743 a_14313_31423.n0 a_14313_31423.t9 27.1302
R8744 a_14313_31423.n1 a_14313_31423.t7 26.9438
R8745 a_14313_31423.n3 a_14313_31423.n1 15.6312
R8746 a_14313_31423.n3 a_14313_31423.n2 15.046
R8747 a_14313_31423.n5 a_14313_31423.t2 10.0473
R8748 a_14313_31423.n6 a_14313_31423.t3 6.51042
R8749 a_14313_31423.n7 a_14313_31423.n6 6.04952
R8750 a_14313_31423.n4 a_14313_31423.n0 5.64619
R8751 a_14313_31423.n5 a_14313_31423.n4 5.17851
R8752 a_14313_31423.n4 a_14313_31423.n3 4.5005
R8753 a_14313_31423.n6 a_14313_31423.n5 0.732092
R8754 a_14313_31423.n7 a_14313_31423.t1 0.7285
R8755 a_14313_31423.t0 a_14313_31423.n7 0.7285
R8756 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t4 41.0041
R8757 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t7 40.6313
R8758 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t6 40.6313
R8759 SARlogic_0.dffrs_2.Qb SARlogic_0.dffrs_9.setb 28.021
R8760 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t9 27.3166
R8761 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t8 27.3166
R8762 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t5 26.9438
R8763 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.t0 10.0473
R8764 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb.n1 9.84255
R8765 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n3 9.22229
R8766 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.t1 6.51042
R8767 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.n7 6.04952
R8768 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.Qb.n0 5.7305
R8769 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n4 5.14711
R8770 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_2.Qb.n2 5.13907
R8771 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n6 4.94976
R8772 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n9 4.72925
R8773 SARlogic_0.dffrs_9.setb SARlogic_0.dffrs_9.nand3_0.C 0.784786
R8774 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.n8 0.732092
R8775 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t2 0.7285
R8776 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t3 0.7285
R8777 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb 0.175225
R8778 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.nand3_2.A 0.0455
R8779 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_9.nand3_2.C 0.0455
R8780 SARlogic_0.dffrs_9.nand3_0.C SARlogic_0.dffrs_2.Qb.n5 0.0374643
.ends

