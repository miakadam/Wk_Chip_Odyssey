* SPICE3 file created from adc_PISO.ext - technology: (null)

.option scale=5n

X0 a_44488_8266 avdd.t378 avss.t87 avss.t86 nfet_03v3
X1 a_50206_2781 a_48650_3501.t4 avdd.t5 avdd.t4 pfet_03v3
X2 a_6600_2510.t2 a_6520_1558.t4 avdd.t317 avdd.t316 pfet_03v3
X3 a_6520_1558.t2 a_6520_3763.t4 avdd.t307 avdd.t306 pfet_03v3
X4 avdd.t337 dffrs_1.Q.t4 a_20234_3501.t2 avdd.t336 pfet_03v3
X5 avdd.t309 a_6520_3763.t5 2inmux_2.Bit.t3 avdd.t308 pfet_03v3
X6 a_2846_2780 a_1290_3500.t4 avdd.t141 avdd.t140 pfet_03v3
X7 dffrs_4.Qb avdd.t379 a_46158_3857 avss.t85 nfet_03v3
X8 a_15992_3763.t3 clk.t0 a_16256_6060 avss.t289 nfet_03v3
X9 2inmux_1.Bit.t1 dffrs_4.Qb a_46158_6061 avss.t35 nfet_03v3
X10 a_10950_2780 2inmux_2.Bit.t4 avss.t94 avss.t93 nfet_03v3
X11 a_15992_5968.t1 a_15992_3763.t4 a_16256_8265 avss.t233 nfet_03v3
X12 a_39178_3501.t0 load.t0 avdd.t271 avdd.t270 pfet_03v3
X13 avss.t179 dffrs_2.Q.t4 a_29894_2781 avss.t178 nfet_03v3
X14 a_50206_441 a_48650_1161.t4 avss.t215 avss.t214 nfet_03v3
X15 2inmux_1.OUT.t1 a_50878_1605.t4 avss.t163 avss.t162 nfet_03v3
X16 avdd.t319 a_6520_1558.t5 dffrs_0.Qb avdd.t318 pfet_03v3
X17 avss.t100 a_21790_2781 a_22462_1605.t3 avss.t99 nfet_03v3
X18 a_35016_1651 a_34936_1559.t4 avss.t137 avss.t136 nfet_03v3
X19 a_35016_3856 a_34936_3764.t4 avss.t139 avss.t138 nfet_03v3
X20 2inmux_0.OUT.t1 a_3518_1604.t4 avss.t142 avss.t141 nfet_03v3
X21 a_22462_1605.t1 a_21790_441 a_22650_2325 avdd.t25 pfet_03v3
X22 a_29000_1361 load.t1 avdd.t345 avdd.t344 pfet_03v3
X23 avss.t15 a_47944_1361 a_48838_441 avss.t14 nfet_03v3
X24 avdd.t127 avdd.t125 a_44408_3764.t0 avdd.t126 pfet_03v3
X25 a_21790_441 a_20234_1161.t4 avdd.t245 avdd.t244 pfet_03v3
X26 a_1478_2780 load.t2 a_1290_3500.t3 avss.t272 nfet_03v3
X27 avdd.t27 a_29000_1361 a_29706_1161.t0 avdd.t26 pfet_03v3
X28 a_25464_3764.t3 clk.t1 avdd.t355 avdd.t354 pfet_03v3
X29 avdd.t124 avdd.t122 a_6600_2510.t0 avdd.t123 pfet_03v3
X30 a_1478_440 B6.t0 a_1290_1160.t3 avss.t101 nfet_03v3
X31 avdd.t239 a_25464_3764.t4 dffrs_2.Q.t3 avdd.t238 pfet_03v3
X32 a_35200_6061 avdd.t380 a_35016_6061 avss.t84 nfet_03v3
X33 avdd.t137 2inmux_2.Bit.t5 a_10762_3500.t3 avdd.t136 pfet_03v3
X34 a_1290_1160.t1 B6.t1 avdd.t247 avdd.t246 pfet_03v3
X35 2inmux_2.Bit.t1 dffrs_0.Qb avdd.t301 avdd.t300 pfet_03v3
X36 avdd.t357 clk.t2 a_6520_1558.t3 avdd.t356 pfet_03v3
X37 a_35200_8266 a_35016_2511.t4 a_35016_8266 avss.t271 nfet_03v3
X38 avss.t280 2inmux_1.Bit.t4 a_48838_2781 avss.t279 nfet_03v3
X39 avss.t185 a_40734_2781 a_41406_1605.t0 avss.t184 nfet_03v3
X40 avdd.t187 a_44488_2511.t4 a_44408_5969.t1 avdd.t186 pfet_03v3
X41 avdd.t219 a_25464_1559.t4 dffrs_2.Qb avdd.t218 pfet_03v3
X42 a_31262_2781 a_29706_3501.t4 avss.t96 avss.t95 nfet_03v3
X43 a_47944_1361 load.t3 avdd.t347 avdd.t346 pfet_03v3
X44 a_39366_2781 dffrs_3.Q.t4 avss.t191 avss.t190 nfet_03v3
X45 dffrs_0.Qb avdd.t119 avdd.t121 avdd.t120 pfet_03v3
X46 avdd.t23 a_584_1360 a_1290_1160.t0 avdd.t22 pfet_03v3
X47 2inmux_3.OUT.t1 a_22462_1605.t4 avss.t175 avss.t174 nfet_03v3
X48 a_51066_2325 a_50206_441 a_50878_1605.t1 avdd.t21 pfet_03v3
X49 a_12990_1604.t1 a_12318_440 a_13178_2324 avdd.t9 pfet_03v3
X50 a_25464_5969.t3 a_25464_3764.t5 avdd.t241 avdd.t240 pfet_03v3
X51 a_44488_2511.t3 a_44408_1559.t4 avdd.t285 avdd.t284 pfet_03v3
X52 avdd.t118 avdd.t116 a_15992_3763.t0 avdd.t117 pfet_03v3
X53 a_44408_3764.t3 clk.t3 avdd.t359 avdd.t358 pfet_03v3
X54 a_44408_1559.t3 a_44408_3764.t4 avdd.t259 avdd.t258 pfet_03v3
X55 a_20422_2781 load.t4 a_20234_3501.t1 avss.t176 nfet_03v3
X56 avdd.t261 a_44408_3764.t5 2inmux_1.Bit.t3 avdd.t260 pfet_03v3
X57 a_54144_6061 avdd.t381 a_53960_6061 avss.t83 nfet_03v3
X58 a_55630_3857 a_53880_1559.t4 a_55446_3857 avss.t130 nfet_03v3
X59 a_54144_8266 a_53960_2511.t4 a_53960_8266 avss.t152 nfet_03v3
X60 avdd.t303 a_15992_3763.t5 dffrs_1.Q.t1 avdd.t302 pfet_03v3
X61 a_25544_6061 a_25464_5969.t4 avss.t147 avss.t146 nfet_03v3
X62 a_27030_3857 dffrs_2.Q.t5 avss.t181 avss.t180 nfet_03v3
X63 a_25544_8266 avdd.t382 avss.t82 avss.t81 nfet_03v3
X64 dffrs_2.Q.t0 dffrs_2.Qb avdd.t1 avdd.t0 pfet_03v3
X65 a_55630_6061 a_53880_3764.t4 a_55446_6061 avss.t148 nfet_03v3
X66 a_3518_1604.t2 a_2846_440 avss.t18 avss.t17 nfet_03v3
X67 a_27030_6061 avdd.t383 avss.t80 avss.t79 nfet_03v3
X68 a_34936_3764.t2 clk.t4 a_35200_6061 avss.t273 nfet_03v3
X69 a_31262_2781 a_29706_3501.t5 avdd.t305 avdd.t304 pfet_03v3
X70 avdd.t235 dffrs_3.Q.t5 a_39178_3501.t3 avdd.t234 pfet_03v3
X71 a_16072_2510.t2 2inmux_2.OUT.t2 avdd.t371 avdd.t370 pfet_03v3
X72 a_34936_5969.t2 a_34936_3764.t5 a_35200_8266 avss.t140 nfet_03v3
X73 avdd.t287 a_44408_1559.t5 dffrs_4.Qb avdd.t286 pfet_03v3
X74 a_15992_1558.t1 a_16072_2510.t4 avdd.t231 avdd.t230 pfet_03v3
X75 a_39366_441 a_38472_1361 avss.t112 avss.t111 nfet_03v3
X76 a_21790_441 a_20234_1161.t5 avss.t193 avss.t192 nfet_03v3
X77 a_1290_1160.t2 B6.t2 a_1478_440 avss.t117 nfet_03v3
X78 a_44408_5969.t3 a_44408_3764.t6 avdd.t263 avdd.t262 pfet_03v3
X79 avdd.t253 a_15992_1558.t4 dffrs_1.Qb avdd.t252 pfet_03v3
X80 dffrs_2.Qb avdd.t113 avdd.t115 avdd.t114 pfet_03v3
X81 avss.t41 a_12318_2780 a_12990_1604.t3 avss.t40 nfet_03v3
X82 avdd.t233 a_16072_2510.t5 a_15992_5968.t3 avdd.t232 pfet_03v3
X83 a_53880_3764.t1 a_53880_5969.t4 avdd.t203 avdd.t202 pfet_03v3
X84 a_2846_440 a_1290_1160.t4 avss.t211 avss.t210 nfet_03v3
X85 a_44672_1651 avdd.t384 a_44488_1651 avss.t78 nfet_03v3
X86 2inmux_4.OUT.t1 a_31934_1605.t4 avss.t287 avss.t286 nfet_03v3
X87 a_44672_3856 clk.t5 a_44488_3856 avss.t274 nfet_03v3
X88 dffrs_3.Q.t1 avdd.t110 avdd.t112 avdd.t111 pfet_03v3
X89 a_45974_3857 2inmux_1.Bit.t5 avss.t282 avss.t281 nfet_03v3
X90 a_10950_2780 load.t5 a_10762_3500.t1 avss.t177 nfet_03v3
X91 a_25544_2511.t2 2inmux_3.OUT.t2 a_25728_1651 avss.t194 nfet_03v3
X92 a_1478_440 a_584_1360 avss.t27 avss.t26 nfet_03v3
X93 a_16072_6060 a_15992_5968.t4 avss.t116 avss.t115 nfet_03v3
X94 a_25464_1559.t0 a_25544_2511.t4 a_25728_3856 avss.t134 nfet_03v3
X95 a_25728_6061 avdd.t385 a_25544_6061 avss.t77 nfet_03v3
X96 a_45974_6061 avdd.t386 avss.t76 avss.t75 nfet_03v3
X97 a_53880_3764.t2 clk.t6 a_54144_6061 avss.t275 nfet_03v3
X98 dffrs_5.Qb avdd.t387 a_55630_3857 avss.t74 nfet_03v3
X99 a_10762_1160.t3 B5.t0 avdd.t185 avdd.t184 pfet_03v3
X100 a_19528_1361 load.t6 avss.t167 avss.t166 nfet_03v3
X101 a_39366_2781 load.t7 a_39178_3501.t2 avss.t168 nfet_03v3
X102 avdd.t109 avdd.t107 a_35016_2511.t1 avdd.t108 pfet_03v3
X103 a_16072_8265 avdd.t388 avss.t73 avss.t72 nfet_03v3
X104 a_25728_8266 a_25544_2511.t5 a_25544_8266 avss.t135 nfet_03v3
X105 a_53880_5969.t0 a_53880_3764.t5 a_54144_8266 avss.t149 nfet_03v3
X106 dffrs_1.Q.t2 dffrs_1.Qb avdd.t363 avdd.t362 pfet_03v3
X107 a_6520_3763.t3 clk.t7 a_6784_6060 avss.t212 nfet_03v3
X108 avdd.t269 clk.t8 a_34936_1559.t1 avdd.t268 pfet_03v3
X109 avdd.t37 a_12318_2780 a_13178_2324 avdd.t36 pfet_03v3
X110 a_22462_1605.t2 a_21790_441 avss.t29 avss.t28 nfet_03v3
X111 a_53880_5969.t3 avdd.t104 avdd.t106 avdd.t105 pfet_03v3
X112 a_6520_5968.t3 a_6520_3763.t6 a_6784_8265 avss.t236 nfet_03v3
X113 serial_out.t3 dffrs_5.Qb a_55630_6061 avss.t98 nfet_03v3
X114 dffrs_3.Qb dffrs_3.Q.t6 avdd.t257 avdd.t256 pfet_03v3
X115 avss.t110 a_38472_1361 a_39366_441 avss.t109 nfet_03v3
X116 a_39366_441 B2.t0 a_39178_1161.t2 avss.t23 nfet_03v3
X117 dffrs_1.Qb avdd.t101 avdd.t103 avdd.t102 pfet_03v3
X118 serial_out.t1 avdd.t98 avdd.t100 avdd.t99 pfet_03v3
X119 a_16256_1650 avdd.t389 a_16072_1650 avss.t71 nfet_03v3
X120 a_44488_2511.t1 2inmux_5.OUT.t2 a_44672_1651 avss.t128 nfet_03v3
X121 a_6520_3763.t2 a_6520_5968.t4 avdd.t161 avdd.t160 pfet_03v3
X122 a_16256_3855 clk.t9 a_16072_3855 avss.t213 nfet_03v3
X123 a_44408_1559.t2 a_44488_2511.t5 a_44672_3856 avss.t143 nfet_03v3
X124 avss.t25 a_584_1360 a_1478_440 avss.t24 nfet_03v3
X125 a_17558_3856 dffrs_1.Q.t5 avss.t267 avss.t266 nfet_03v3
X126 avdd.t97 avdd.t95 a_53960_2511.t3 avdd.t96 pfet_03v3
X127 a_48650_3501.t2 load.t8 a_48838_2781 avss.t278 nfet_03v3
X128 a_41406_1605.t1 a_40734_441 avss.t240 avss.t239 nfet_03v3
X129 avdd.t181 a_34936_3764.t6 dffrs_3.Q.t0 avdd.t180 pfet_03v3
X130 avdd.t273 clk.t10 a_53880_1559.t3 avdd.t272 pfet_03v3
X131 a_25544_2511.t0 a_25464_1559.t5 avdd.t221 avdd.t220 pfet_03v3
X132 a_25464_1559.t2 a_25464_3764.t6 avdd.t243 avdd.t242 pfet_03v3
X133 dffrs_5.Qb serial_out.t4 avdd.t167 avdd.t166 pfet_03v3
X134 a_12990_1604.t2 a_12318_440 avss.t11 avss.t10 nfet_03v3
X135 2inmux_1.OUT.t0 a_50878_1605.t5 avdd.t213 avdd.t212 pfet_03v3
X136 a_17558_6060 avdd.t390 avss.t70 avss.t69 nfet_03v3
X137 avss.t247 avss.t245 a_1478_2780 avss.t246 nfet_03v3
X138 a_22650_2325 a_21790_2781 avdd.t145 avdd.t144 pfet_03v3
X139 a_35016_2511.t2 2inmux_4.OUT.t2 avdd.t205 avdd.t204 pfet_03v3
X140 a_34936_1559.t3 a_35016_2511.t5 avdd.t343 avdd.t342 pfet_03v3
X141 2inmux_0.OUT.t0 a_3518_1604.t5 avdd.t183 avdd.t182 pfet_03v3
X142 avss.t161 a_50206_2781 a_50878_1605.t3 avss.t160 nfet_03v3
X143 a_40734_2781 a_39178_3501.t4 avss.t165 avss.t164 nfet_03v3
X144 avdd.t375 a_34936_1559.t5 dffrs_3.Qb avdd.t374 pfet_03v3
X145 a_20422_441 B4.t0 a_20234_1161.t3 avss.t16 nfet_03v3
X146 a_48838_2781 2inmux_1.Bit.t6 avss.t252 avss.t251 nfet_03v3
X147 a_6520_5968.t0 avdd.t92 avdd.t94 avdd.t93 pfet_03v3
X148 a_53960_1651 a_53880_1559.t5 avss.t132 avss.t131 nfet_03v3
X149 a_53960_3856 a_53880_3764.t6 avss.t151 avss.t150 nfet_03v3
X150 a_12318_440 a_10762_1160.t4 avss.t114 avss.t113 nfet_03v3
X151 a_41406_1605.t3 a_40734_441 a_41594_2325 avdd.t311 pfet_03v3
X152 a_48650_3501.t3 load.t9 avdd.t353 avdd.t352 pfet_03v3
X153 a_29706_3501.t1 load.t10 a_29894_2781 avss.t217 nfet_03v3
X154 avdd.t91 avdd.t89 a_6520_3763.t0 avdd.t90 pfet_03v3
X155 a_35016_6061 a_34936_5969.t4 avss.t198 avss.t197 nfet_03v3
X156 2inmux_2.Bit.t0 avdd.t86 avdd.t88 avdd.t87 pfet_03v3
X157 a_16072_2510.t3 a_15992_1558.t5 avdd.t255 avdd.t254 pfet_03v3
X158 a_10056_1360 load.t11 avss.t219 avss.t218 nfet_03v3
X159 a_53960_2511.t2 2inmux_1.OUT.t2 avdd.t149 avdd.t148 pfet_03v3
X160 a_35016_8266 avdd.t391 avss.t68 avss.t67 nfet_03v3
X161 a_15992_1558.t0 a_15992_3763.t6 avdd.t281 avdd.t280 pfet_03v3
X162 a_40734_2781 a_39178_3501.t5 avdd.t237 avdd.t236 pfet_03v3
X163 avdd.t85 avdd.t83 a_25544_2511.t3 avdd.t84 pfet_03v3
X164 a_41594_2325 a_40734_2781 avdd.t227 avdd.t226 pfet_03v3
X165 avdd.t299 a_31262_2781 a_32122_2325 avdd.t298 pfet_03v3
X166 avdd.t275 clk.t11 a_25464_1559.t3 avdd.t274 pfet_03v3
X167 a_53880_1559.t2 a_53960_2511.t5 avdd.t197 avdd.t196 pfet_03v3
X168 avdd.t321 2inmux_1.Bit.t7 a_48650_3501.t1 avdd.t320 pfet_03v3
X169 a_6600_2510.t3 2inmux_0.OUT.t2 avdd.t201 avdd.t200 pfet_03v3
X170 a_584_1360 load.t12 avss.t228 avss.t227 nfet_03v3
X171 a_6520_1558.t1 a_6600_2510.t4 avdd.t13 avdd.t12 pfet_03v3
X172 dffrs_3.Qb avdd.t392 a_36686_3857 avss.t66 nfet_03v3
X173 avss.t263 dffrs_1.Q.t6 a_20422_2781 avss.t262 nfet_03v3
X174 2inmux_3.OUT.t0 a_22462_1605.t5 avdd.t223 avdd.t222 pfet_03v3
X175 a_20234_1161.t1 B4.t1 avdd.t7 avdd.t6 pfet_03v3
X176 dffrs_0.Qb 2inmux_2.Bit.t6 avdd.t147 avdd.t146 pfet_03v3
X177 a_20234_1161.t2 B4.t2 a_20422_441 avss.t9 nfet_03v3
X178 dffrs_3.Q.t3 dffrs_3.Qb a_36686_6061 avss.t241 nfet_03v3
X179 a_12318_2780 a_10762_3500.t4 avss.t269 avss.t268 nfet_03v3
X180 avdd.t15 a_6600_2510.t5 a_6520_5968.t1 avdd.t14 pfet_03v3
X181 a_29706_3501.t2 load.t13 avdd.t293 avdd.t292 pfet_03v3
X182 avss.t285 a_2846_2780 a_3518_1604.t3 avss.t284 nfet_03v3
X183 2inmux_5.OUT.t1 a_41406_1605.t4 avss.t235 avss.t234 nfet_03v3
X184 a_44408_3764.t1 a_44408_5969.t4 avdd.t159 avdd.t158 pfet_03v3
X185 a_6600_1650 a_6520_1558.t6 avss.t249 avss.t248 nfet_03v3
X186 a_50206_441 a_48650_1161.t5 avdd.t279 avdd.t278 pfet_03v3
X187 a_2846_440 a_1290_1160.t5 avdd.t267 avdd.t266 pfet_03v3
X188 avdd.t3 a_19528_1361 a_20234_1161.t0 avdd.t2 pfet_03v3
X189 a_6600_3855 a_6520_3763.t7 avss.t238 avss.t237 nfet_03v3
X190 a_3706_2324 a_2846_440 a_3518_1604.t1 avdd.t17 pfet_03v3
X191 avss.t39 a_10056_1360 a_10950_440 avss.t38 nfet_03v3
X192 a_39178_1161.t1 B2.t1 a_39366_441 avss.t260 nfet_03v3
X193 a_20422_441 a_19528_1361 avss.t6 avss.t5 nfet_03v3
X194 a_10950_440 B5.t1 a_10762_1160.t2 avss.t253 nfet_03v3
X195 a_31934_1605.t2 a_31262_441 avss.t89 avss.t88 nfet_03v3
X196 a_15992_3763.t2 clk.t12 avdd.t277 avdd.t276 pfet_03v3
X197 2inmux_1.Bit.t0 dffrs_4.Qb avdd.t31 avdd.t30 pfet_03v3
X198 avdd.t367 a_2846_2780 a_3706_2324 avdd.t366 pfet_03v3
X199 a_40734_441 a_39178_1161.t4 avss.t121 avss.t120 nfet_03v3
X200 a_39178_1161.t0 B2.t2 avdd.t165 avdd.t164 pfet_03v3
X201 a_8270_3856 a_6520_1558.t7 a_8086_3856 avss.t250 nfet_03v3
X202 a_12318_2780 a_10762_3500.t5 avdd.t339 avdd.t338 pfet_03v3
X203 a_13178_2324 a_12318_2780 avdd.t35 avdd.t34 pfet_03v3
X204 a_44408_5969.t0 avdd.t80 avdd.t82 avdd.t81 pfet_03v3
X205 a_8270_6060 a_6520_3763.t8 a_8086_6060 avss.t34 nfet_03v3
X206 2inmux_4.OUT.t0 a_31934_1605.t5 avdd.t373 avdd.t372 pfet_03v3
X207 dffrs_4.Qb avdd.t77 avdd.t79 avdd.t78 pfet_03v3
X208 a_21790_2781 a_20234_3501.t4 avss.t43 avss.t42 nfet_03v3
X209 a_29894_2781 dffrs_2.Q.t6 avss.t183 avss.t182 nfet_03v3
X210 avdd.t33 a_10056_1360 a_10762_1160.t0 avdd.t32 pfet_03v3
X211 2inmux_2.OUT.t1 a_12990_1604.t4 avss.t196 avss.t195 nfet_03v3
X212 a_31934_1605.t1 a_31262_441 a_32122_2325 avdd.t129 pfet_03v3
X213 a_15992_5968.t0 a_15992_3763.t7 avdd.t283 avdd.t282 pfet_03v3
X214 a_6784_1650 avdd.t393 a_6600_1650 avss.t65 nfet_03v3
X215 a_19528_1361 load.t14 avdd.t215 avdd.t214 pfet_03v3
X216 a_22650_2325 a_21790_441 a_22462_1605.t0 avdd.t24 pfet_03v3
X217 a_6784_3855 clk.t13 a_6600_3855 avss.t19 nfet_03v3
X218 a_1290_3500.t0 load.t15 a_1478_2780 avss.t169 nfet_03v3
X219 a_35016_2511.t0 a_34936_1559.t6 avdd.t377 avdd.t376 pfet_03v3
X220 avdd.t76 avdd.t74 a_34936_3764.t0 avdd.t75 pfet_03v3
X221 a_34936_1559.t0 a_34936_3764.t7 avdd.t289 avdd.t288 pfet_03v3
X222 a_44672_6061 avdd.t394 a_44488_6061 avss.t64 nfet_03v3
X223 a_38472_1361 load.t16 avss.t255 avss.t254 nfet_03v3
X224 a_44672_8266 a_44488_2511.t6 a_44488_8266 avss.t144 nfet_03v3
X225 dffrs_0.Qb avdd.t395 a_8270_3856 avss.t63 nfet_03v3
X226 a_27214_3857 a_25464_1559.t6 a_27030_3857 avss.t125 nfet_03v3
X227 a_1478_2780 avss.t242 avss.t244 avss.t243 nfet_03v3
X228 avss.t4 a_19528_1361 a_20422_441 avss.t3 nfet_03v3
X229 a_25464_3764.t2 clk.t14 a_25728_6061 avss.t20 nfet_03v3
X230 a_21790_2781 a_20234_3501.t5 avdd.t369 avdd.t368 pfet_03v3
X231 avdd.t151 dffrs_2.Q.t7 a_29706_3501.t3 avdd.t150 pfet_03v3
X232 a_25464_5969.t2 a_25464_3764.t7 a_25728_8266 avss.t222 nfet_03v3
X233 a_27214_6061 a_25464_3764.t8 a_27030_6061 avss.t223 nfet_03v3
X234 a_10762_1160.t1 B5.t2 a_10950_440 avss.t44 nfet_03v3
X235 a_10950_440 a_10056_1360 avss.t37 avss.t36 nfet_03v3
X236 2inmux_2.Bit.t2 dffrs_0.Qb a_8270_6060 avss.t232 nfet_03v3
X237 a_50878_1605.t0 a_50206_441 a_51066_2325 avdd.t20 pfet_03v3
X238 a_44488_1651 a_44408_1559.t6 avss.t221 avss.t220 nfet_03v3
X239 avss.t231 a_31262_2781 a_31934_1605.t3 avss.t230 nfet_03v3
X240 avdd.t341 a_35016_2511.t6 a_34936_5969.t0 avdd.t340 pfet_03v3
X241 a_1290_3500.t2 load.t17 avdd.t327 avdd.t326 pfet_03v3
X242 a_44488_3856 a_44408_3764.t7 avss.t207 avss.t206 nfet_03v3
X243 a_41594_2325 a_40734_441 a_41406_1605.t2 avdd.t310 pfet_03v3
X244 avdd.t73 avdd.t71 a_53880_3764.t0 avdd.t72 pfet_03v3
X245 a_25464_3764.t1 a_25464_5969.t5 avdd.t207 avdd.t206 pfet_03v3
X246 a_13178_2324 a_12318_440 a_12990_1604.t0 avdd.t8 pfet_03v3
X247 a_29894_2781 load.t18 a_29706_3501.t0 avss.t256 nfet_03v3
X248 a_31262_441 a_29706_1161.t4 avdd.t313 avdd.t312 pfet_03v3
X249 avdd.t155 a_38472_1361 a_39178_1161.t3 avdd.t154 pfet_03v3
X250 dffrs_2.Q.t2 avdd.t68 avdd.t70 avdd.t69 pfet_03v3
X251 a_34936_3764.t3 clk.t15 avdd.t19 avdd.t18 pfet_03v3
X252 avdd.t191 a_53880_3764.t7 serial_out.t0 avdd.t190 pfet_03v3
X253 a_46158_3857 a_44408_1559.t7 a_45974_3857 avss.t159 nfet_03v3
X254 a_16072_2510.t1 2inmux_2.OUT.t3 a_16256_1650 avss.t124 nfet_03v3
X255 a_51066_2325 a_50206_2781 avdd.t211 avdd.t210 pfet_03v3
X256 avdd.t325 avss.t290 a_1290_3500.t1 avdd.t324 pfet_03v3
X257 a_15992_1558.t2 a_16072_2510.t6 a_16256_3855 avss.t188 nfet_03v3
X258 a_29894_441 a_29000_1361 avss.t33 avss.t32 nfet_03v3
X259 a_16256_6060 avdd.t396 a_16072_6060 avss.t62 nfet_03v3
X260 a_44408_3764.t2 clk.t16 a_44672_6061 avss.t90 nfet_03v3
X261 a_17742_3856 a_15992_1558.t6 a_17558_3856 avss.t201 nfet_03v3
X262 a_16256_8265 a_16072_2510.t7 a_16072_8265 avss.t189 nfet_03v3
X263 a_44408_5969.t2 a_44408_3764.t8 a_44672_8266 avss.t208 nfet_03v3
X264 a_46158_6061 a_44408_3764.t9 a_45974_6061 avss.t209 nfet_03v3
X265 dffrs_2.Qb avdd.t397 a_27214_3857 avss.t61 nfet_03v3
X266 a_17742_6060 a_15992_3763.t8 a_17558_6060 avss.t216 nfet_03v3
X267 dffrs_2.Qb dffrs_2.Q.t8 avdd.t153 avdd.t152 pfet_03v3
X268 avdd.t173 a_53880_1559.t6 dffrs_5.Qb avdd.t172 pfet_03v3
X269 avdd.t189 a_53960_2511.t6 a_53880_5969.t2 avdd.t188 pfet_03v3
X270 dffrs_2.Q.t1 dffrs_2.Qb a_27214_6061 avss.t0 nfet_03v3
X271 a_25464_5969.t0 avdd.t65 avdd.t67 avdd.t66 pfet_03v3
X272 a_10056_1360 load.t19 avdd.t329 avdd.t328 pfet_03v3
X273 a_34936_5969.t1 a_34936_3764.t8 avdd.t291 avdd.t290 pfet_03v3
X274 a_31262_441 a_29706_1161.t5 avss.t173 avss.t172 nfet_03v3
X275 a_15992_3763.t1 a_15992_5968.t5 avdd.t265 avdd.t264 pfet_03v3
X276 a_35200_1651 avdd.t398 a_35016_1651 avss.t60 nfet_03v3
X277 a_10762_3500.t0 load.t21 a_10950_2780 avss.t276 nfet_03v3
X278 a_584_1360 load.t20 avdd.t349 avdd.t348 pfet_03v3
X279 a_53880_3764.t3 clk.t17 avdd.t131 avdd.t130 pfet_03v3
X280 2inmux_1.Bit.t2 avdd.t41 avdd.t43 avdd.t42 pfet_03v3
X281 avdd.t64 avdd.t62 a_25464_3764.t0 avdd.t63 pfet_03v3
X282 a_35200_3856 clk.t19 a_35016_3856 avss.t91 nfet_03v3
X283 a_53960_6061 a_53880_5969.t5 avss.t154 avss.t153 nfet_03v3
X284 a_6520_3763.t1 clk.t18 avdd.t133 avdd.t132 pfet_03v3
X285 a_29000_1361 load.t22 avss.t171 avss.t170 nfet_03v3
X286 avdd.t61 avdd.t59 a_44488_2511.t0 avdd.t60 pfet_03v3
X287 avdd.t209 a_50206_2781 a_51066_2325 avdd.t208 pfet_03v3
X288 a_36502_3857 dffrs_3.Q.t7 avss.t203 avss.t202 nfet_03v3
X289 serial_out.t2 dffrs_5.Qb avdd.t139 avdd.t138 pfet_03v3
X290 a_53960_8266 avdd.t399 avss.t59 avss.t58 nfet_03v3
X291 a_3706_2324 a_2846_2780 avdd.t365 avdd.t364 pfet_03v3
X292 avdd.t135 clk.t20 a_44408_1559.t0 avdd.t134 pfet_03v3
X293 2inmux_5.OUT.t0 a_41406_1605.t5 avdd.t169 avdd.t168 pfet_03v3
X294 a_25544_2511.t1 2inmux_3.OUT.t3 avdd.t249 avdd.t248 pfet_03v3
X295 dffrs_1.Qb avdd.t401 a_17742_3856 avss.t55 nfet_03v3
X296 dffrs_4.Qb 2inmux_1.Bit.t8 avdd.t323 avdd.t322 pfet_03v3
X297 a_36502_6061 avdd.t400 avss.t57 avss.t56 nfet_03v3
X298 dffrs_5.Qb avdd.t56 avdd.t58 avdd.t57 pfet_03v3
X299 a_25464_1559.t1 a_25544_2511.t6 avdd.t179 avdd.t178 pfet_03v3
X300 avss.t31 a_29000_1361 a_29894_441 avss.t30 nfet_03v3
X301 dffrs_1.Q.t3 dffrs_1.Qb a_17742_6060 avss.t283 nfet_03v3
X302 a_53880_5969.t1 a_53880_3764.t8 avdd.t193 avdd.t192 pfet_03v3
X303 a_15992_5968.t2 avdd.t53 avdd.t55 avdd.t54 pfet_03v3
X304 a_54144_1651 avdd.t402 a_53960_1651 avss.t54 nfet_03v3
X305 a_10762_3500.t2 load.t23 avdd.t217 avdd.t216 pfet_03v3
X306 avdd.t177 a_25544_2511.t7 a_25464_5969.t1 avdd.t176 pfet_03v3
X307 a_32122_2325 a_31262_441 a_31934_1605.t0 avdd.t128 pfet_03v3
X308 a_25544_1651 a_25464_1559.t7 avss.t127 avss.t126 nfet_03v3
X309 a_6520_5968.t2 a_6520_3763.t9 avdd.t29 avdd.t28 pfet_03v3
X310 a_54144_3856 clk.t21 a_53960_3856 avss.t92 nfet_03v3
X311 a_25544_3856 a_25464_3764.t9 avss.t225 avss.t224 nfet_03v3
X312 a_35016_2511.t3 2inmux_4.OUT.t3 a_35200_1651 avss.t155 nfet_03v3
X313 a_47944_1361 load.t24 avss.t157 avss.t156 nfet_03v3
X314 a_48838_441 B1.t0 a_48650_1161.t1 avss.t45 nfet_03v3
X315 a_55446_3857 serial_out.t5 avss.t123 avss.t122 nfet_03v3
X316 a_50878_1605.t2 a_50206_441 avss.t22 avss.t21 nfet_03v3
X317 a_34936_1559.t2 a_35016_2511.t7 a_35200_3856 avss.t270 nfet_03v3
X318 dffrs_1.Q.t0 avdd.t50 avdd.t52 avdd.t51 pfet_03v3
X319 a_44488_2511.t2 2inmux_5.OUT.t3 avdd.t199 avdd.t198 pfet_03v3
X320 a_48838_2781 load.t25 a_48650_3501.t0 avss.t158 nfet_03v3
X321 a_36686_3857 a_34936_1559.t7 a_36502_3857 avss.t288 nfet_03v3
X322 a_55446_6061 avdd.t403 avss.t53 avss.t52 nfet_03v3
X323 a_6600_6060 a_6520_5968.t5 avss.t119 avss.t118 nfet_03v3
X324 avdd.t143 a_21790_2781 a_22650_2325 avdd.t142 pfet_03v3
X325 avdd.t49 avdd.t47 a_16072_2510.t0 avdd.t48 pfet_03v3
X326 a_44408_1559.t1 a_44488_2511.t7 avdd.t361 avdd.t360 pfet_03v3
X327 avdd.t331 clk.t22 a_15992_1558.t3 avdd.t330 pfet_03v3
X328 a_36686_6061 a_34936_3764.t9 a_36502_6061 avss.t226 nfet_03v3
X329 a_6600_8265 avdd.t404 avss.t51 avss.t50 nfet_03v3
X330 a_48650_1161.t2 B1.t1 avdd.t295 avdd.t294 pfet_03v3
X331 2inmux_2.OUT.t0 a_12990_1604.t5 avdd.t229 avdd.t228 pfet_03v3
X332 avss.t103 2inmux_2.Bit.t7 a_10950_2780 avss.t102 nfet_03v3
X333 dffrs_1.Qb dffrs_1.Q.t7 avdd.t335 avdd.t334 pfet_03v3
X334 avss.t205 dffrs_3.Q.t8 a_39366_2781 avss.t204 nfet_03v3
X335 a_16072_1650 a_15992_1558.t7 avss.t200 avss.t199 nfet_03v3
X336 a_38472_1361 load.t26 avdd.t175 avdd.t174 pfet_03v3
X337 a_40734_441 a_39178_1161.t5 avdd.t163 avdd.t162 pfet_03v3
X338 a_53960_2511.t1 2inmux_1.OUT.t3 a_54144_1651 avss.t106 nfet_03v3
X339 a_29894_441 B3.t0 a_29706_1161.t2 avss.t261 nfet_03v3
X340 a_25728_1651 avdd.t405 a_25544_1651 avss.t49 nfet_03v3
X341 a_34936_3764.t1 a_34936_5969.t5 avdd.t251 avdd.t250 pfet_03v3
X342 a_53960_2511.t0 a_53880_1559.t7 avdd.t171 avdd.t170 pfet_03v3
X343 avdd.t11 a_47944_1361 a_48650_1161.t0 avdd.t10 pfet_03v3
X344 a_6600_2510.t1 2inmux_0.OUT.t3 a_6784_1650 avss.t97 nfet_03v3
X345 a_53880_1559.t0 a_53960_2511.t7 a_54144_3856 avss.t145 nfet_03v3
X346 a_16072_3855 a_15992_3763.t9 avss.t259 avss.t258 nfet_03v3
X347 a_20234_3501.t0 load.t27 a_20422_2781 avss.t133 nfet_03v3
X348 a_25728_3856 clk.t23 a_25544_3856 avss.t257 nfet_03v3
X349 a_53880_1559.t1 a_53880_3764.t9 avdd.t195 avdd.t194 pfet_03v3
X350 avdd.t225 a_40734_2781 a_41594_2325 avdd.t224 pfet_03v3
X351 a_8086_3856 2inmux_2.Bit.t8 avss.t105 avss.t104 nfet_03v3
X352 a_6520_1558.t0 a_6600_2510.t6 a_6784_3855 avss.t1 nfet_03v3
X353 a_32122_2325 a_31262_2781 avdd.t297 avdd.t296 pfet_03v3
X354 a_29706_1161.t3 B3.t1 avdd.t333 avdd.t332 pfet_03v3
X355 a_6784_6060 avdd.t406 a_6600_6060 avss.t48 nfet_03v3
X356 dffrs_3.Q.t2 dffrs_3.Qb avdd.t315 avdd.t314 pfet_03v3
X357 a_50206_2781 a_48650_3501.t5 avss.t8 avss.t7 nfet_03v3
X358 a_48650_1161.t3 B1.t2 a_48838_441 avss.t229 nfet_03v3
X359 a_8086_6060 avdd.t407 avss.t47 avss.t46 nfet_03v3
X360 a_6784_8265 a_6600_2510.t7 a_6600_8265 avss.t2 nfet_03v3
X361 a_20422_2781 dffrs_1.Q.t8 avss.t265 avss.t264 nfet_03v3
X362 a_34936_5969.t3 avdd.t44 avdd.t46 avdd.t45 pfet_03v3
X363 a_2846_2780 a_1290_3500.t5 avss.t108 avss.t107 nfet_03v3
X364 a_29706_1161.t1 B3.t2 a_29894_441 avss.t129 nfet_03v3
X365 dffrs_3.Qb avdd.t38 avdd.t40 avdd.t39 pfet_03v3
X366 a_20234_3501.t3 load.t28 avdd.t351 avdd.t350 pfet_03v3
X367 a_39178_3501.t1 load.t29 a_39366_2781 avss.t277 nfet_03v3
X368 a_48838_441 a_47944_1361 avss.t13 avss.t12 nfet_03v3
X369 a_3518_1604.t0 a_2846_440 a_3706_2324 avdd.t16 pfet_03v3
X370 a_12318_440 a_10762_1160.t5 avdd.t157 avdd.t156 pfet_03v3
X371 a_44488_6061 a_44408_5969.t5 avss.t187 avss.t186 nfet_03v3
R0 avdd.t282 avdd.n390 250.9
R1 avdd.n391 avdd.t54 250.9
R2 avdd.t276 avdd.n401 250.9
R3 avdd.n402 avdd.t264 250.9
R4 avdd.t362 avdd.n396 250.9
R5 avdd.n397 avdd.t51 250.9
R6 avdd.t230 avdd.n413 250.9
R7 avdd.n414 avdd.t280 250.9
R8 avdd.t102 avdd.n407 250.9
R9 avdd.n408 avdd.t334 250.9
R10 avdd.t370 avdd.n425 250.9
R11 avdd.n426 avdd.t254 250.9
R12 avdd.t192 avdd.n98 250.9
R13 avdd.n99 avdd.t105 250.9
R14 avdd.t130 avdd.n109 250.9
R15 avdd.n110 avdd.t202 250.9
R16 avdd.t138 avdd.n104 250.9
R17 avdd.n105 avdd.t99 250.9
R18 avdd.t196 avdd.n121 250.9
R19 avdd.n122 avdd.t194 250.9
R20 avdd.t57 avdd.n115 250.9
R21 avdd.n116 avdd.t166 250.9
R22 avdd.t148 avdd.n132 250.9
R23 avdd.n133 avdd.t170 250.9
R24 avdd.t262 avdd.n171 250.9
R25 avdd.n172 avdd.t81 250.9
R26 avdd.t358 avdd.n182 250.9
R27 avdd.n183 avdd.t158 250.9
R28 avdd.t30 avdd.n177 250.9
R29 avdd.n178 avdd.t42 250.9
R30 avdd.t360 avdd.n194 250.9
R31 avdd.n195 avdd.t258 250.9
R32 avdd.t78 avdd.n188 250.9
R33 avdd.n189 avdd.t322 250.9
R34 avdd.t198 avdd.n205 250.9
R35 avdd.n206 avdd.t284 250.9
R36 avdd.t290 avdd.n244 250.9
R37 avdd.n245 avdd.t45 250.9
R38 avdd.t18 avdd.n255 250.9
R39 avdd.n256 avdd.t250 250.9
R40 avdd.t314 avdd.n250 250.9
R41 avdd.n251 avdd.t111 250.9
R42 avdd.t342 avdd.n267 250.9
R43 avdd.n268 avdd.t288 250.9
R44 avdd.t39 avdd.n261 250.9
R45 avdd.n262 avdd.t256 250.9
R46 avdd.t204 avdd.n278 250.9
R47 avdd.n279 avdd.t376 250.9
R48 avdd.t240 avdd.n317 250.9
R49 avdd.n318 avdd.t66 250.9
R50 avdd.t354 avdd.n328 250.9
R51 avdd.n329 avdd.t206 250.9
R52 avdd.t0 avdd.n323 250.9
R53 avdd.n324 avdd.t69 250.9
R54 avdd.t178 avdd.n340 250.9
R55 avdd.n341 avdd.t242 250.9
R56 avdd.t114 avdd.n334 250.9
R57 avdd.n335 avdd.t152 250.9
R58 avdd.t248 avdd.n351 250.9
R59 avdd.n352 avdd.t220 250.9
R60 avdd.t28 avdd.n4 250.9
R61 avdd.n5 avdd.t93 250.9
R62 avdd.t132 avdd.n528 250.9
R63 avdd.n529 avdd.t160 250.9
R64 avdd.t300 avdd.n9 250.9
R65 avdd.n10 avdd.t87 250.9
R66 avdd.t12 avdd.n516 250.9
R67 avdd.n517 avdd.t306 250.9
R68 avdd.t120 avdd.n522 250.9
R69 avdd.n523 avdd.t146 250.9
R70 avdd.t200 avdd.n465 250.9
R71 avdd.n466 avdd.t316 250.9
R72 avdd.n495 avdd.t140 236.083
R73 avdd.t326 avdd.n491 236.083
R74 avdd.t266 avdd.n499 236.083
R75 avdd.n505 avdd.t246 236.083
R76 avdd.n453 avdd.t338 236.083
R77 avdd.t216 avdd.n450 236.083
R78 avdd.t156 avdd.n433 236.083
R79 avdd.n439 avdd.t184 236.083
R80 avdd.n379 avdd.t368 236.083
R81 avdd.t350 avdd.n376 236.083
R82 avdd.t244 avdd.n359 236.083
R83 avdd.n365 avdd.t6 236.083
R84 avdd.n306 avdd.t304 236.083
R85 avdd.t292 avdd.n303 236.083
R86 avdd.t312 avdd.n286 236.083
R87 avdd.n292 avdd.t332 236.083
R88 avdd.n233 avdd.t236 236.083
R89 avdd.t270 avdd.n230 236.083
R90 avdd.t162 avdd.n213 236.083
R91 avdd.n219 avdd.t164 236.083
R92 avdd.n160 avdd.t4 236.083
R93 avdd.t352 avdd.n157 236.083
R94 avdd.t278 avdd.n140 236.083
R95 avdd.n146 avdd.t294 236.083
R96 avdd.n92 avdd.t212 236.083
R97 avdd.n86 avdd.t210 236.083
R98 avdd.n76 avdd.t168 236.083
R99 avdd.n70 avdd.t226 236.083
R100 avdd.n60 avdd.t372 236.083
R101 avdd.n54 avdd.t296 236.083
R102 avdd.n44 avdd.t222 236.083
R103 avdd.n38 avdd.t144 236.083
R104 avdd.n28 avdd.t228 236.083
R105 avdd.n22 avdd.t34 236.083
R106 avdd.t182 avdd.n470 236.083
R107 avdd.n481 avdd.t364 236.083
R108 avdd.t140 avdd.n494 235.294
R109 avdd.n494 avdd.t326 235.294
R110 avdd.n504 avdd.t266 235.294
R111 avdd.t246 avdd.n504 235.294
R112 avdd.t338 avdd.n452 235.294
R113 avdd.n452 avdd.t216 235.294
R114 avdd.n438 avdd.t156 235.294
R115 avdd.t184 avdd.n438 235.294
R116 avdd.t368 avdd.n378 235.294
R117 avdd.n378 avdd.t350 235.294
R118 avdd.n364 avdd.t244 235.294
R119 avdd.t6 avdd.n364 235.294
R120 avdd.t304 avdd.n305 235.294
R121 avdd.n305 avdd.t292 235.294
R122 avdd.n291 avdd.t312 235.294
R123 avdd.t332 avdd.n291 235.294
R124 avdd.t236 avdd.n232 235.294
R125 avdd.n232 avdd.t270 235.294
R126 avdd.n218 avdd.t162 235.294
R127 avdd.t164 avdd.n218 235.294
R128 avdd.t4 avdd.n159 235.294
R129 avdd.n159 avdd.t352 235.294
R130 avdd.n145 avdd.t278 235.294
R131 avdd.t294 avdd.n145 235.294
R132 avdd.t212 avdd.n91 235.294
R133 avdd.n91 avdd.t20 235.294
R134 avdd.t21 avdd.n89 235.294
R135 avdd.n89 avdd.t208 235.294
R136 avdd.t168 avdd.n75 235.294
R137 avdd.n75 avdd.t311 235.294
R138 avdd.t310 avdd.n73 235.294
R139 avdd.n73 avdd.t224 235.294
R140 avdd.t372 avdd.n59 235.294
R141 avdd.n59 avdd.t129 235.294
R142 avdd.t128 avdd.n57 235.294
R143 avdd.n57 avdd.t298 235.294
R144 avdd.t222 avdd.n43 235.294
R145 avdd.n43 avdd.t25 235.294
R146 avdd.t24 avdd.n41 235.294
R147 avdd.n41 avdd.t142 235.294
R148 avdd.t228 avdd.n27 235.294
R149 avdd.n27 avdd.t9 235.294
R150 avdd.t8 avdd.n25 235.294
R151 avdd.n25 avdd.t36 235.294
R152 avdd.n478 avdd.t182 235.294
R153 avdd.t16 avdd.n478 235.294
R154 avdd.n480 avdd.t17 235.294
R155 avdd.t366 avdd.n480 235.294
R156 avdd.t232 avdd.t282 200
R157 avdd.t54 avdd.t232 200
R158 avdd.t117 avdd.t276 200
R159 avdd.t264 avdd.t117 200
R160 avdd.t302 avdd.t362 200
R161 avdd.t51 avdd.t302 200
R162 avdd.t330 avdd.t230 200
R163 avdd.t280 avdd.t330 200
R164 avdd.t252 avdd.t102 200
R165 avdd.t334 avdd.t252 200
R166 avdd.t48 avdd.t370 200
R167 avdd.t254 avdd.t48 200
R168 avdd.t188 avdd.t192 200
R169 avdd.t105 avdd.t188 200
R170 avdd.t72 avdd.t130 200
R171 avdd.t202 avdd.t72 200
R172 avdd.t190 avdd.t138 200
R173 avdd.t99 avdd.t190 200
R174 avdd.t272 avdd.t196 200
R175 avdd.t194 avdd.t272 200
R176 avdd.t172 avdd.t57 200
R177 avdd.t166 avdd.t172 200
R178 avdd.t96 avdd.t148 200
R179 avdd.t170 avdd.t96 200
R180 avdd.t20 avdd.t21 200
R181 avdd.t210 avdd.t208 200
R182 avdd.t186 avdd.t262 200
R183 avdd.t81 avdd.t186 200
R184 avdd.t126 avdd.t358 200
R185 avdd.t158 avdd.t126 200
R186 avdd.t260 avdd.t30 200
R187 avdd.t42 avdd.t260 200
R188 avdd.t134 avdd.t360 200
R189 avdd.t258 avdd.t134 200
R190 avdd.t286 avdd.t78 200
R191 avdd.t322 avdd.t286 200
R192 avdd.t60 avdd.t198 200
R193 avdd.t284 avdd.t60 200
R194 avdd.t311 avdd.t310 200
R195 avdd.t226 avdd.t224 200
R196 avdd.t340 avdd.t290 200
R197 avdd.t45 avdd.t340 200
R198 avdd.t75 avdd.t18 200
R199 avdd.t250 avdd.t75 200
R200 avdd.t180 avdd.t314 200
R201 avdd.t111 avdd.t180 200
R202 avdd.t268 avdd.t342 200
R203 avdd.t288 avdd.t268 200
R204 avdd.t374 avdd.t39 200
R205 avdd.t256 avdd.t374 200
R206 avdd.t108 avdd.t204 200
R207 avdd.t376 avdd.t108 200
R208 avdd.t129 avdd.t128 200
R209 avdd.t296 avdd.t298 200
R210 avdd.t176 avdd.t240 200
R211 avdd.t66 avdd.t176 200
R212 avdd.t63 avdd.t354 200
R213 avdd.t206 avdd.t63 200
R214 avdd.t238 avdd.t0 200
R215 avdd.t69 avdd.t238 200
R216 avdd.t274 avdd.t178 200
R217 avdd.t242 avdd.t274 200
R218 avdd.t218 avdd.t114 200
R219 avdd.t152 avdd.t218 200
R220 avdd.t84 avdd.t248 200
R221 avdd.t220 avdd.t84 200
R222 avdd.t25 avdd.t24 200
R223 avdd.t144 avdd.t142 200
R224 avdd.t9 avdd.t8 200
R225 avdd.t34 avdd.t36 200
R226 avdd.t14 avdd.t28 200
R227 avdd.t93 avdd.t14 200
R228 avdd.t90 avdd.t132 200
R229 avdd.t160 avdd.t90 200
R230 avdd.t308 avdd.t300 200
R231 avdd.t87 avdd.t308 200
R232 avdd.t356 avdd.t12 200
R233 avdd.t306 avdd.t356 200
R234 avdd.t318 avdd.t120 200
R235 avdd.t146 avdd.t318 200
R236 avdd.t123 avdd.t200 200
R237 avdd.t316 avdd.t123 200
R238 avdd.t17 avdd.t16 200
R239 avdd.t364 avdd.t366 200
R240 avdd.n486 avdd.t324 131.589
R241 avdd.n507 avdd.t22 131.589
R242 avdd.n14 avdd.t136 131.589
R243 avdd.n441 avdd.t32 131.589
R244 avdd.n30 avdd.t336 131.589
R245 avdd.n367 avdd.t2 131.589
R246 avdd.n46 avdd.t150 131.589
R247 avdd.n294 avdd.t26 131.589
R248 avdd.n62 avdd.t234 131.589
R249 avdd.n221 avdd.t154 131.589
R250 avdd.n78 avdd.t320 131.589
R251 avdd.n148 avdd.t10 131.589
R252 avdd.n164 avdd.t346 118.543
R253 avdd.n237 avdd.t174 118.543
R254 avdd.n310 avdd.t344 118.543
R255 avdd.n383 avdd.t214 118.543
R256 avdd.n457 avdd.t328 118.543
R257 avdd.n487 avdd.t348 118.543
R258 avdd.n86 avdd.n85 96.0755
R259 avdd.n87 avdd.n86 96.0755
R260 avdd.n70 avdd.n69 96.0755
R261 avdd.n71 avdd.n70 96.0755
R262 avdd.n54 avdd.n53 96.0755
R263 avdd.n55 avdd.n54 96.0755
R264 avdd.n38 avdd.n37 96.0755
R265 avdd.n39 avdd.n38 96.0755
R266 avdd.n22 avdd.n21 96.0755
R267 avdd.n23 avdd.n22 96.0755
R268 avdd.n481 avdd.n473 96.0755
R269 avdd.n481 avdd.n474 96.0755
R270 avdd.n501 avdd.n499 78.2255
R271 avdd.n505 avdd.n501 78.2255
R272 avdd.n505 avdd.n502 78.2255
R273 avdd.n502 avdd.n499 78.2255
R274 avdd.n435 avdd.n433 78.2255
R275 avdd.n439 avdd.n435 78.2255
R276 avdd.n439 avdd.n436 78.2255
R277 avdd.n436 avdd.n433 78.2255
R278 avdd.n361 avdd.n359 78.2255
R279 avdd.n365 avdd.n361 78.2255
R280 avdd.n365 avdd.n362 78.2255
R281 avdd.n362 avdd.n359 78.2255
R282 avdd.n288 avdd.n286 78.2255
R283 avdd.n292 avdd.n288 78.2255
R284 avdd.n292 avdd.n289 78.2255
R285 avdd.n289 avdd.n286 78.2255
R286 avdd.n215 avdd.n213 78.2255
R287 avdd.n219 avdd.n215 78.2255
R288 avdd.n219 avdd.n216 78.2255
R289 avdd.n216 avdd.n213 78.2255
R290 avdd.n142 avdd.n140 78.2255
R291 avdd.n146 avdd.n142 78.2255
R292 avdd.n146 avdd.n143 78.2255
R293 avdd.n143 avdd.n140 78.2255
R294 avdd.n92 avdd.n83 78.2255
R295 avdd.n92 avdd.n84 78.2255
R296 avdd.n160 avdd.n155 78.2255
R297 avdd.n160 avdd.n156 78.2255
R298 avdd.n157 avdd.n155 78.2255
R299 avdd.n157 avdd.n156 78.2255
R300 avdd.n76 avdd.n67 78.2255
R301 avdd.n76 avdd.n68 78.2255
R302 avdd.n233 avdd.n228 78.2255
R303 avdd.n233 avdd.n229 78.2255
R304 avdd.n230 avdd.n228 78.2255
R305 avdd.n230 avdd.n229 78.2255
R306 avdd.n60 avdd.n51 78.2255
R307 avdd.n60 avdd.n52 78.2255
R308 avdd.n306 avdd.n301 78.2255
R309 avdd.n306 avdd.n302 78.2255
R310 avdd.n303 avdd.n301 78.2255
R311 avdd.n303 avdd.n302 78.2255
R312 avdd.n44 avdd.n35 78.2255
R313 avdd.n44 avdd.n36 78.2255
R314 avdd.n379 avdd.n374 78.2255
R315 avdd.n379 avdd.n375 78.2255
R316 avdd.n376 avdd.n374 78.2255
R317 avdd.n376 avdd.n375 78.2255
R318 avdd.n28 avdd.n19 78.2255
R319 avdd.n28 avdd.n20 78.2255
R320 avdd.n453 avdd.n448 78.2255
R321 avdd.n453 avdd.n449 78.2255
R322 avdd.n450 avdd.n448 78.2255
R323 avdd.n450 avdd.n449 78.2255
R324 avdd.n475 avdd.n470 78.2255
R325 avdd.n476 avdd.n470 78.2255
R326 avdd.n495 avdd.n484 78.2255
R327 avdd.n495 avdd.n485 78.2255
R328 avdd.n491 avdd.n484 78.2255
R329 avdd.n491 avdd.n485 78.2255
R330 avdd.n391 avdd.n390 68.0765
R331 avdd.n402 avdd.n401 68.0765
R332 avdd.n397 avdd.n396 68.0765
R333 avdd.n414 avdd.n413 68.0765
R334 avdd.n408 avdd.n407 68.0765
R335 avdd.n426 avdd.n425 68.0765
R336 avdd.n99 avdd.n98 68.0765
R337 avdd.n110 avdd.n109 68.0765
R338 avdd.n105 avdd.n104 68.0765
R339 avdd.n122 avdd.n121 68.0765
R340 avdd.n116 avdd.n115 68.0765
R341 avdd.n133 avdd.n132 68.0765
R342 avdd.n172 avdd.n171 68.0765
R343 avdd.n183 avdd.n182 68.0765
R344 avdd.n178 avdd.n177 68.0765
R345 avdd.n195 avdd.n194 68.0765
R346 avdd.n189 avdd.n188 68.0765
R347 avdd.n206 avdd.n205 68.0765
R348 avdd.n245 avdd.n244 68.0765
R349 avdd.n256 avdd.n255 68.0765
R350 avdd.n251 avdd.n250 68.0765
R351 avdd.n268 avdd.n267 68.0765
R352 avdd.n262 avdd.n261 68.0765
R353 avdd.n279 avdd.n278 68.0765
R354 avdd.n318 avdd.n317 68.0765
R355 avdd.n329 avdd.n328 68.0765
R356 avdd.n324 avdd.n323 68.0765
R357 avdd.n341 avdd.n340 68.0765
R358 avdd.n335 avdd.n334 68.0765
R359 avdd.n352 avdd.n351 68.0765
R360 avdd.n5 avdd.n4 68.0765
R361 avdd.n529 avdd.n528 68.0765
R362 avdd.n10 avdd.n9 68.0765
R363 avdd.n517 avdd.n516 68.0765
R364 avdd.n523 avdd.n522 68.0765
R365 avdd.n466 avdd.n465 68.0765
R366 avdd.n85 avdd.n83 59.8505
R367 avdd.n87 avdd.n84 59.8505
R368 avdd.n69 avdd.n67 59.8505
R369 avdd.n71 avdd.n68 59.8505
R370 avdd.n53 avdd.n51 59.8505
R371 avdd.n55 avdd.n52 59.8505
R372 avdd.n37 avdd.n35 59.8505
R373 avdd.n39 avdd.n36 59.8505
R374 avdd.n21 avdd.n19 59.8505
R375 avdd.n23 avdd.n20 59.8505
R376 avdd.n475 avdd.n473 59.8505
R377 avdd.n476 avdd.n474 59.8505
R378 avdd.n419 avdd.t101 41.0041
R379 avdd.n126 avdd.t56 41.0041
R380 avdd.n199 avdd.t77 41.0041
R381 avdd.n272 avdd.t38 41.0041
R382 avdd.n345 avdd.t113 41.0041
R383 avdd.n459 avdd.t119 41.0041
R384 avdd.n421 avdd.t47 40.8177
R385 avdd.n420 avdd.t116 40.8177
R386 avdd.n128 avdd.t95 40.8177
R387 avdd.n127 avdd.t71 40.8177
R388 avdd.n201 avdd.t59 40.8177
R389 avdd.n200 avdd.t125 40.8177
R390 avdd.n274 avdd.t107 40.8177
R391 avdd.n273 avdd.t74 40.8177
R392 avdd.n347 avdd.t83 40.8177
R393 avdd.n346 avdd.t62 40.8177
R394 avdd.n461 avdd.t122 40.8177
R395 avdd.n460 avdd.t89 40.8177
R396 avdd.n386 avdd.t53 40.6313
R397 avdd.n385 avdd.t50 40.6313
R398 avdd.n94 avdd.t104 40.6313
R399 avdd.n93 avdd.t98 40.6313
R400 avdd.n167 avdd.t80 40.6313
R401 avdd.n166 avdd.t41 40.6313
R402 avdd.n240 avdd.t44 40.6313
R403 avdd.n239 avdd.t110 40.6313
R404 avdd.n313 avdd.t65 40.6313
R405 avdd.n312 avdd.t68 40.6313
R406 avdd.n1 avdd.t92 40.6313
R407 avdd.n0 avdd.t86 40.6313
R408 avdd.n503 avdd.n501 36.2255
R409 avdd.n503 avdd.n502 36.2255
R410 avdd.n437 avdd.n435 36.2255
R411 avdd.n437 avdd.n436 36.2255
R412 avdd.n363 avdd.n361 36.2255
R413 avdd.n363 avdd.n362 36.2255
R414 avdd.n290 avdd.n288 36.2255
R415 avdd.n290 avdd.n289 36.2255
R416 avdd.n217 avdd.n215 36.2255
R417 avdd.n217 avdd.n216 36.2255
R418 avdd.n144 avdd.n142 36.2255
R419 avdd.n144 avdd.n143 36.2255
R420 avdd.n88 avdd.n85 36.2255
R421 avdd.n88 avdd.n87 36.2255
R422 avdd.n90 avdd.n83 36.2255
R423 avdd.n90 avdd.n84 36.2255
R424 avdd.n158 avdd.n155 36.2255
R425 avdd.n158 avdd.n156 36.2255
R426 avdd.n72 avdd.n69 36.2255
R427 avdd.n72 avdd.n71 36.2255
R428 avdd.n74 avdd.n67 36.2255
R429 avdd.n74 avdd.n68 36.2255
R430 avdd.n231 avdd.n228 36.2255
R431 avdd.n231 avdd.n229 36.2255
R432 avdd.n56 avdd.n53 36.2255
R433 avdd.n56 avdd.n55 36.2255
R434 avdd.n58 avdd.n51 36.2255
R435 avdd.n58 avdd.n52 36.2255
R436 avdd.n304 avdd.n301 36.2255
R437 avdd.n304 avdd.n302 36.2255
R438 avdd.n40 avdd.n37 36.2255
R439 avdd.n40 avdd.n39 36.2255
R440 avdd.n42 avdd.n35 36.2255
R441 avdd.n42 avdd.n36 36.2255
R442 avdd.n377 avdd.n374 36.2255
R443 avdd.n377 avdd.n375 36.2255
R444 avdd.n24 avdd.n21 36.2255
R445 avdd.n24 avdd.n23 36.2255
R446 avdd.n26 avdd.n19 36.2255
R447 avdd.n26 avdd.n20 36.2255
R448 avdd.n451 avdd.n448 36.2255
R449 avdd.n451 avdd.n449 36.2255
R450 avdd.n479 avdd.n473 36.2255
R451 avdd.n479 avdd.n474 36.2255
R452 avdd.n477 avdd.n475 36.2255
R453 avdd.n477 avdd.n476 36.2255
R454 avdd.n493 avdd.n484 36.2255
R455 avdd.n493 avdd.n485 36.2255
R456 avdd.n386 avdd.t388 27.3166
R457 avdd.n385 avdd.t390 27.3166
R458 avdd.n94 avdd.t399 27.3166
R459 avdd.n93 avdd.t403 27.3166
R460 avdd.n167 avdd.t378 27.3166
R461 avdd.n166 avdd.t386 27.3166
R462 avdd.n240 avdd.t391 27.3166
R463 avdd.n239 avdd.t400 27.3166
R464 avdd.n313 avdd.t382 27.3166
R465 avdd.n312 avdd.t383 27.3166
R466 avdd.n1 avdd.t404 27.3166
R467 avdd.n0 avdd.t407 27.3166
R468 avdd.n421 avdd.t389 27.1302
R469 avdd.n420 avdd.t396 27.1302
R470 avdd.n128 avdd.t402 27.1302
R471 avdd.n127 avdd.t381 27.1302
R472 avdd.n201 avdd.t384 27.1302
R473 avdd.n200 avdd.t394 27.1302
R474 avdd.n274 avdd.t398 27.1302
R475 avdd.n273 avdd.t380 27.1302
R476 avdd.n347 avdd.t405 27.1302
R477 avdd.n346 avdd.t385 27.1302
R478 avdd.n461 avdd.t393 27.1302
R479 avdd.n460 avdd.t406 27.1302
R480 avdd.n419 avdd.t401 26.9438
R481 avdd.n126 avdd.t387 26.9438
R482 avdd.n199 avdd.t379 26.9438
R483 avdd.n272 avdd.t392 26.9438
R484 avdd.n345 avdd.t397 26.9438
R485 avdd.n459 avdd.t395 26.9438
R486 avdd.n429 dffrs_1.resetb 18.2415
R487 avdd.n136 dffrs_5.resetb 18.2415
R488 avdd.n209 dffrs_4.resetb 18.2415
R489 avdd.n282 dffrs_3.resetb 18.2415
R490 avdd.n355 dffrs_2.resetb 18.2415
R491 avdd.n469 dffrs_0.resetb 18.2415
R492 avdd.n394 avdd.n388 18.0418
R493 avdd.n102 avdd.n96 18.0418
R494 avdd.n175 avdd.n169 18.0418
R495 avdd.n248 avdd.n242 18.0418
R496 avdd.n321 avdd.n315 18.0418
R497 avdd.n534 avdd.n533 18.0418
R498 avdd.n422 avdd.n420 17.6364
R499 avdd.n129 avdd.n127 17.6364
R500 avdd.n202 avdd.n200 17.6364
R501 avdd.n275 avdd.n273 17.6364
R502 avdd.n348 avdd.n346 17.6364
R503 avdd.n462 avdd.n460 17.6364
R504 avdd.n387 avdd.n385 14.3609
R505 avdd.n95 avdd.n93 14.3609
R506 avdd.n168 avdd.n166 14.3609
R507 avdd.n241 avdd.n239 14.3609
R508 avdd.n314 avdd.n312 14.3609
R509 avdd.n2 avdd.n0 14.3609
R510 avdd.n394 avdd.n393 13.5174
R511 avdd.n102 avdd.n101 13.5174
R512 avdd.n175 avdd.n174 13.5174
R513 avdd.n248 avdd.n247 13.5174
R514 avdd.n321 avdd.n320 13.5174
R515 avdd.n533 avdd.n7 13.5174
R516 avdd.n405 avdd.n404 13.5005
R517 avdd.n405 avdd.n399 13.5005
R518 avdd.n417 avdd.n416 13.5005
R519 avdd.n411 avdd.n410 13.5005
R520 avdd.n429 avdd.n428 13.5005
R521 avdd.n113 avdd.n112 13.5005
R522 avdd.n113 avdd.n107 13.5005
R523 avdd.n125 avdd.n124 13.5005
R524 avdd.n119 avdd.n118 13.5005
R525 avdd.n136 avdd.n135 13.5005
R526 avdd.n186 avdd.n185 13.5005
R527 avdd.n186 avdd.n180 13.5005
R528 avdd.n198 avdd.n197 13.5005
R529 avdd.n192 avdd.n191 13.5005
R530 avdd.n209 avdd.n208 13.5005
R531 avdd.n259 avdd.n258 13.5005
R532 avdd.n259 avdd.n253 13.5005
R533 avdd.n271 avdd.n270 13.5005
R534 avdd.n265 avdd.n264 13.5005
R535 avdd.n282 avdd.n281 13.5005
R536 avdd.n332 avdd.n331 13.5005
R537 avdd.n332 avdd.n326 13.5005
R538 avdd.n344 avdd.n343 13.5005
R539 avdd.n338 avdd.n337 13.5005
R540 avdd.n355 avdd.n354 13.5005
R541 avdd.n532 avdd.n531 13.5005
R542 avdd.n532 avdd.n12 13.5005
R543 avdd.n520 avdd.n519 13.5005
R544 avdd.n526 avdd.n525 13.5005
R545 avdd.n469 avdd.n468 13.5005
R546 avdd.n423 avdd.n419 13.4839
R547 avdd.n130 avdd.n126 13.4839
R548 avdd.n203 avdd.n199 13.4839
R549 avdd.n276 avdd.n272 13.4839
R550 avdd.n349 avdd.n345 13.4839
R551 avdd.n463 avdd.n459 13.4839
R552 avdd.n422 avdd.n421 10.5752
R553 avdd.n129 avdd.n128 10.5752
R554 avdd.n202 avdd.n201 10.5752
R555 avdd.n275 avdd.n274 10.5752
R556 avdd.n348 avdd.n347 10.5752
R557 avdd.n462 avdd.n461 10.5752
R558 avdd.n393 avdd.n390 6.4802
R559 avdd.n404 avdd.n401 6.4802
R560 avdd.n399 avdd.n396 6.4802
R561 avdd.n416 avdd.n413 6.4802
R562 avdd.n410 avdd.n407 6.4802
R563 avdd.n428 avdd.n425 6.4802
R564 avdd.n101 avdd.n98 6.4802
R565 avdd.n112 avdd.n109 6.4802
R566 avdd.n107 avdd.n104 6.4802
R567 avdd.n124 avdd.n121 6.4802
R568 avdd.n118 avdd.n115 6.4802
R569 avdd.n135 avdd.n132 6.4802
R570 avdd.n174 avdd.n171 6.4802
R571 avdd.n185 avdd.n182 6.4802
R572 avdd.n180 avdd.n177 6.4802
R573 avdd.n197 avdd.n194 6.4802
R574 avdd.n191 avdd.n188 6.4802
R575 avdd.n208 avdd.n205 6.4802
R576 avdd.n247 avdd.n244 6.4802
R577 avdd.n258 avdd.n255 6.4802
R578 avdd.n253 avdd.n250 6.4802
R579 avdd.n270 avdd.n267 6.4802
R580 avdd.n264 avdd.n261 6.4802
R581 avdd.n281 avdd.n278 6.4802
R582 avdd.n320 avdd.n317 6.4802
R583 avdd.n331 avdd.n328 6.4802
R584 avdd.n326 avdd.n323 6.4802
R585 avdd.n343 avdd.n340 6.4802
R586 avdd.n337 avdd.n334 6.4802
R587 avdd.n354 avdd.n351 6.4802
R588 avdd.n7 avdd.n4 6.4802
R589 avdd.n531 avdd.n528 6.4802
R590 avdd.n12 avdd.n9 6.4802
R591 avdd.n519 avdd.n516 6.4802
R592 avdd.n525 avdd.n522 6.4802
R593 avdd.n468 avdd.n465 6.4802
R594 avdd.n393 avdd.n389 6.25878
R595 avdd.n404 avdd.n400 6.25878
R596 avdd.n399 avdd.n395 6.25878
R597 avdd.n416 avdd.n412 6.25878
R598 avdd.n410 avdd.n406 6.25878
R599 avdd.n428 avdd.n424 6.25878
R600 avdd.n101 avdd.n97 6.25878
R601 avdd.n112 avdd.n108 6.25878
R602 avdd.n107 avdd.n103 6.25878
R603 avdd.n124 avdd.n120 6.25878
R604 avdd.n118 avdd.n114 6.25878
R605 avdd.n135 avdd.n131 6.25878
R606 avdd.n174 avdd.n170 6.25878
R607 avdd.n185 avdd.n181 6.25878
R608 avdd.n180 avdd.n176 6.25878
R609 avdd.n197 avdd.n193 6.25878
R610 avdd.n191 avdd.n187 6.25878
R611 avdd.n208 avdd.n204 6.25878
R612 avdd.n247 avdd.n243 6.25878
R613 avdd.n258 avdd.n254 6.25878
R614 avdd.n253 avdd.n249 6.25878
R615 avdd.n270 avdd.n266 6.25878
R616 avdd.n264 avdd.n260 6.25878
R617 avdd.n281 avdd.n277 6.25878
R618 avdd.n320 avdd.n316 6.25878
R619 avdd.n331 avdd.n327 6.25878
R620 avdd.n326 avdd.n322 6.25878
R621 avdd.n343 avdd.n339 6.25878
R622 avdd.n337 avdd.n333 6.25878
R623 avdd.n354 avdd.n350 6.25878
R624 avdd.n7 avdd.n3 6.25878
R625 avdd.n531 avdd.n527 6.25878
R626 avdd.n12 avdd.n8 6.25878
R627 avdd.n519 avdd.n515 6.25878
R628 avdd.n525 avdd.n521 6.25878
R629 avdd.n468 avdd.n464 6.25878
R630 avdd.n423 avdd.n422 5.93546
R631 avdd.n130 avdd.n129 5.93546
R632 avdd.n203 avdd.n202 5.93546
R633 avdd.n276 avdd.n275 5.93546
R634 avdd.n349 avdd.n348 5.93546
R635 avdd.n463 avdd.n462 5.93546
R636 avdd.n393 avdd.n392 5.44497
R637 avdd.n404 avdd.n403 5.44497
R638 avdd.n399 avdd.n398 5.44497
R639 avdd.n416 avdd.n415 5.44497
R640 avdd.n410 avdd.n409 5.44497
R641 avdd.n428 avdd.n427 5.44497
R642 avdd.n101 avdd.n100 5.44497
R643 avdd.n112 avdd.n111 5.44497
R644 avdd.n107 avdd.n106 5.44497
R645 avdd.n124 avdd.n123 5.44497
R646 avdd.n118 avdd.n117 5.44497
R647 avdd.n135 avdd.n134 5.44497
R648 avdd.n174 avdd.n173 5.44497
R649 avdd.n185 avdd.n184 5.44497
R650 avdd.n180 avdd.n179 5.44497
R651 avdd.n197 avdd.n196 5.44497
R652 avdd.n191 avdd.n190 5.44497
R653 avdd.n208 avdd.n207 5.44497
R654 avdd.n247 avdd.n246 5.44497
R655 avdd.n258 avdd.n257 5.44497
R656 avdd.n253 avdd.n252 5.44497
R657 avdd.n270 avdd.n269 5.44497
R658 avdd.n264 avdd.n263 5.44497
R659 avdd.n281 avdd.n280 5.44497
R660 avdd.n320 avdd.n319 5.44497
R661 avdd.n331 avdd.n330 5.44497
R662 avdd.n326 avdd.n325 5.44497
R663 avdd.n343 avdd.n342 5.44497
R664 avdd.n337 avdd.n336 5.44497
R665 avdd.n354 avdd.n353 5.44497
R666 avdd.n7 avdd.n6 5.44497
R667 avdd.n531 avdd.n530 5.44497
R668 avdd.n12 avdd.n11 5.44497
R669 avdd.n519 avdd.n518 5.44497
R670 avdd.n525 avdd.n524 5.44497
R671 avdd.n468 avdd.n467 5.44497
R672 avdd.n387 avdd.n386 5.14711
R673 avdd.n95 avdd.n94 5.14711
R674 avdd.n168 avdd.n167 5.14711
R675 avdd.n241 avdd.n240 5.14711
R676 avdd.n314 avdd.n313 5.14711
R677 avdd.n2 avdd.n1 5.14711
R678 avdd.n511 avdd.n510 2.49936
R679 avdd.n445 avdd.n444 2.49936
R680 avdd.n371 avdd.n370 2.49936
R681 avdd.n298 avdd.n297 2.49936
R682 avdd.n225 avdd.n224 2.49936
R683 avdd.n152 avdd.n151 2.49936
R684 avdd.n510 avdd.n499 1.93883
R685 avdd.n444 avdd.n433 1.93883
R686 avdd.n370 avdd.n359 1.93883
R687 avdd.n297 avdd.n286 1.93883
R688 avdd.n224 avdd.n213 1.93883
R689 avdd.n151 avdd.n140 1.93883
R690 avdd.n392 avdd.t55 1.85637
R691 avdd.n403 avdd.t265 1.85637
R692 avdd.n398 avdd.t52 1.85637
R693 avdd.n415 avdd.t281 1.85637
R694 avdd.n409 avdd.t335 1.85637
R695 avdd.n427 avdd.t255 1.85637
R696 avdd.n100 avdd.t106 1.85637
R697 avdd.n111 avdd.t203 1.85637
R698 avdd.n106 avdd.t100 1.85637
R699 avdd.n123 avdd.t195 1.85637
R700 avdd.n117 avdd.t167 1.85637
R701 avdd.n134 avdd.t171 1.85637
R702 avdd.n173 avdd.t82 1.85637
R703 avdd.n184 avdd.t159 1.85637
R704 avdd.n179 avdd.t43 1.85637
R705 avdd.n196 avdd.t259 1.85637
R706 avdd.n190 avdd.t323 1.85637
R707 avdd.n207 avdd.t285 1.85637
R708 avdd.n246 avdd.t46 1.85637
R709 avdd.n257 avdd.t251 1.85637
R710 avdd.n252 avdd.t112 1.85637
R711 avdd.n269 avdd.t289 1.85637
R712 avdd.n263 avdd.t257 1.85637
R713 avdd.n280 avdd.t377 1.85637
R714 avdd.n319 avdd.t67 1.85637
R715 avdd.n330 avdd.t207 1.85637
R716 avdd.n325 avdd.t70 1.85637
R717 avdd.n342 avdd.t243 1.85637
R718 avdd.n336 avdd.t153 1.85637
R719 avdd.n353 avdd.t221 1.85637
R720 avdd.n6 avdd.t94 1.85637
R721 avdd.n530 avdd.t161 1.85637
R722 avdd.n11 avdd.t88 1.85637
R723 avdd.n518 avdd.t307 1.85637
R724 avdd.n524 avdd.t147 1.85637
R725 avdd.n467 avdd.t317 1.85637
R726 avdd.n138 avdd.n92 1.80479
R727 avdd.n211 avdd.n76 1.80479
R728 avdd.n284 avdd.n60 1.80479
R729 avdd.n357 avdd.n44 1.80479
R730 avdd.n431 avdd.n28 1.80479
R731 avdd.n513 avdd.n470 1.80479
R732 avdd.n161 avdd.n160 1.78583
R733 avdd.n234 avdd.n233 1.78583
R734 avdd.n307 avdd.n306 1.78583
R735 avdd.n380 avdd.n379 1.78583
R736 avdd.n454 avdd.n453 1.78583
R737 avdd.n496 avdd.n495 1.78583
R738 avdd.n164 avdd.t347 1.74654
R739 avdd.n237 avdd.t175 1.74654
R740 avdd.n310 avdd.t345 1.74654
R741 avdd.n383 avdd.t215 1.74654
R742 avdd.n457 avdd.t329 1.74654
R743 avdd.n487 avdd.t349 1.74654
R744 avdd.n486 avdd.t325 1.49467
R745 avdd.n507 avdd.t23 1.49467
R746 avdd.n506 avdd.t247 1.49467
R747 avdd.n14 avdd.t137 1.49467
R748 avdd.n441 avdd.t33 1.49467
R749 avdd.n440 avdd.t185 1.49467
R750 avdd.n30 avdd.t337 1.49467
R751 avdd.n367 avdd.t3 1.49467
R752 avdd.n366 avdd.t7 1.49467
R753 avdd.n46 avdd.t151 1.49467
R754 avdd.n294 avdd.t27 1.49467
R755 avdd.n293 avdd.t333 1.49467
R756 avdd.n62 avdd.t235 1.49467
R757 avdd.n221 avdd.t155 1.49467
R758 avdd.n220 avdd.t165 1.49467
R759 avdd.n78 avdd.t321 1.49467
R760 avdd.n148 avdd.t11 1.49467
R761 avdd.n147 avdd.t295 1.49467
R762 avdd.n77 avdd.t353 1.49467
R763 avdd.n61 avdd.t271 1.49467
R764 avdd.n45 avdd.t293 1.49467
R765 avdd.n29 avdd.t351 1.49467
R766 avdd.n13 avdd.t217 1.49467
R767 avdd.n490 avdd.t327 1.49467
R768 avdd.n500 avdd.t267 1.47383
R769 avdd.n434 avdd.t157 1.47383
R770 avdd.n360 avdd.t245 1.47383
R771 avdd.n287 avdd.t313 1.47383
R772 avdd.n214 avdd.t163 1.47383
R773 avdd.n141 avdd.t279 1.47383
R774 avdd.n80 avdd.t211 1.47383
R775 avdd.n81 avdd.t209 1.47383
R776 avdd.n82 avdd.t213 1.47383
R777 avdd.n79 avdd.t5 1.47383
R778 avdd.n64 avdd.t227 1.47383
R779 avdd.n65 avdd.t225 1.47383
R780 avdd.n66 avdd.t169 1.47383
R781 avdd.n63 avdd.t237 1.47383
R782 avdd.n48 avdd.t297 1.47383
R783 avdd.n49 avdd.t299 1.47383
R784 avdd.n50 avdd.t373 1.47383
R785 avdd.n47 avdd.t305 1.47383
R786 avdd.n32 avdd.t145 1.47383
R787 avdd.n33 avdd.t143 1.47383
R788 avdd.n34 avdd.t223 1.47383
R789 avdd.n31 avdd.t369 1.47383
R790 avdd.n16 avdd.t35 1.47383
R791 avdd.n17 avdd.t37 1.47383
R792 avdd.n18 avdd.t229 1.47383
R793 avdd.n15 avdd.t339 1.47383
R794 avdd.n482 avdd.t365 1.47383
R795 avdd.n472 avdd.t367 1.47383
R796 avdd.n471 avdd.t183 1.47383
R797 avdd.n492 avdd.t141 1.47383
R798 avdd.n210 avdd.n165 1.19311
R799 avdd.n283 avdd.n238 1.19311
R800 avdd.n356 avdd.n311 1.19311
R801 avdd.n418 avdd.n384 1.19311
R802 avdd.n514 avdd.n458 1.19311
R803 avdd.n392 avdd.n391 1.04105
R804 avdd.n403 avdd.n402 1.04105
R805 avdd.n398 avdd.n397 1.04105
R806 avdd.n415 avdd.n414 1.04105
R807 avdd.n409 avdd.n408 1.04105
R808 avdd.n427 avdd.n426 1.04105
R809 avdd.n100 avdd.n99 1.04105
R810 avdd.n111 avdd.n110 1.04105
R811 avdd.n106 avdd.n105 1.04105
R812 avdd.n123 avdd.n122 1.04105
R813 avdd.n117 avdd.n116 1.04105
R814 avdd.n134 avdd.n133 1.04105
R815 avdd.n173 avdd.n172 1.04105
R816 avdd.n184 avdd.n183 1.04105
R817 avdd.n179 avdd.n178 1.04105
R818 avdd.n196 avdd.n195 1.04105
R819 avdd.n190 avdd.n189 1.04105
R820 avdd.n207 avdd.n206 1.04105
R821 avdd.n246 avdd.n245 1.04105
R822 avdd.n257 avdd.n256 1.04105
R823 avdd.n252 avdd.n251 1.04105
R824 avdd.n269 avdd.n268 1.04105
R825 avdd.n263 avdd.n262 1.04105
R826 avdd.n280 avdd.n279 1.04105
R827 avdd.n319 avdd.n318 1.04105
R828 avdd.n330 avdd.n329 1.04105
R829 avdd.n325 avdd.n324 1.04105
R830 avdd.n342 avdd.n341 1.04105
R831 avdd.n336 avdd.n335 1.04105
R832 avdd.n353 avdd.n352 1.04105
R833 avdd.n6 avdd.n5 1.04105
R834 avdd.n530 avdd.n529 1.04105
R835 avdd.n11 avdd.n10 1.04105
R836 avdd.n518 avdd.n517 1.04105
R837 avdd.n524 avdd.n523 1.04105
R838 avdd.n467 avdd.n466 1.04105
R839 avdd.n138 avdd.n137 0.809622
R840 avdd.n211 avdd.n210 0.809622
R841 avdd.n284 avdd.n283 0.809622
R842 avdd.n357 avdd.n356 0.809622
R843 avdd.n431 avdd.n430 0.809622
R844 avdd.n514 avdd.n513 0.809622
R845 avdd.n503 avdd.n500 0.788
R846 avdd.n504 avdd.n503 0.788
R847 avdd.n506 avdd.n505 0.788
R848 avdd.n437 avdd.n434 0.788
R849 avdd.n438 avdd.n437 0.788
R850 avdd.n440 avdd.n439 0.788
R851 avdd.n363 avdd.n360 0.788
R852 avdd.n364 avdd.n363 0.788
R853 avdd.n366 avdd.n365 0.788
R854 avdd.n290 avdd.n287 0.788
R855 avdd.n291 avdd.n290 0.788
R856 avdd.n293 avdd.n292 0.788
R857 avdd.n217 avdd.n214 0.788
R858 avdd.n218 avdd.n217 0.788
R859 avdd.n220 avdd.n219 0.788
R860 avdd.n144 avdd.n141 0.788
R861 avdd.n145 avdd.n144 0.788
R862 avdd.n147 avdd.n146 0.788
R863 avdd.n88 avdd.n81 0.788
R864 avdd.n89 avdd.n88 0.788
R865 avdd.n90 avdd.n82 0.788
R866 avdd.n91 avdd.n90 0.788
R867 avdd.n86 avdd.n80 0.788
R868 avdd.n158 avdd.n79 0.788
R869 avdd.n159 avdd.n158 0.788
R870 avdd.n157 avdd.n77 0.788
R871 avdd.n72 avdd.n65 0.788
R872 avdd.n73 avdd.n72 0.788
R873 avdd.n74 avdd.n66 0.788
R874 avdd.n75 avdd.n74 0.788
R875 avdd.n70 avdd.n64 0.788
R876 avdd.n231 avdd.n63 0.788
R877 avdd.n232 avdd.n231 0.788
R878 avdd.n230 avdd.n61 0.788
R879 avdd.n56 avdd.n49 0.788
R880 avdd.n57 avdd.n56 0.788
R881 avdd.n58 avdd.n50 0.788
R882 avdd.n59 avdd.n58 0.788
R883 avdd.n54 avdd.n48 0.788
R884 avdd.n304 avdd.n47 0.788
R885 avdd.n305 avdd.n304 0.788
R886 avdd.n303 avdd.n45 0.788
R887 avdd.n40 avdd.n33 0.788
R888 avdd.n41 avdd.n40 0.788
R889 avdd.n42 avdd.n34 0.788
R890 avdd.n43 avdd.n42 0.788
R891 avdd.n38 avdd.n32 0.788
R892 avdd.n377 avdd.n31 0.788
R893 avdd.n378 avdd.n377 0.788
R894 avdd.n376 avdd.n29 0.788
R895 avdd.n24 avdd.n17 0.788
R896 avdd.n25 avdd.n24 0.788
R897 avdd.n26 avdd.n18 0.788
R898 avdd.n27 avdd.n26 0.788
R899 avdd.n22 avdd.n16 0.788
R900 avdd.n451 avdd.n15 0.788
R901 avdd.n452 avdd.n451 0.788
R902 avdd.n450 avdd.n13 0.788
R903 avdd.n479 avdd.n472 0.788
R904 avdd.n480 avdd.n479 0.788
R905 avdd.n477 avdd.n471 0.788
R906 avdd.n478 avdd.n477 0.788
R907 avdd.n482 avdd.n481 0.788
R908 avdd.n493 avdd.n492 0.788
R909 avdd.n494 avdd.n493 0.788
R910 avdd.n491 avdd.n490 0.788
R911 avdd.n388 avdd.n387 0.754571
R912 avdd.n96 avdd.n95 0.754571
R913 avdd.n169 avdd.n168 0.754571
R914 avdd.n242 avdd.n241 0.754571
R915 avdd.n315 avdd.n314 0.754571
R916 avdd.n534 avdd.n2 0.754571
R917 avdd.n389 avdd.t283 0.7285
R918 avdd.n389 avdd.t233 0.7285
R919 avdd.n400 avdd.t277 0.7285
R920 avdd.n400 avdd.t118 0.7285
R921 avdd.n395 avdd.t363 0.7285
R922 avdd.n395 avdd.t303 0.7285
R923 avdd.n412 avdd.t231 0.7285
R924 avdd.n412 avdd.t331 0.7285
R925 avdd.n406 avdd.t103 0.7285
R926 avdd.n406 avdd.t253 0.7285
R927 avdd.n424 avdd.t371 0.7285
R928 avdd.n424 avdd.t49 0.7285
R929 avdd.n97 avdd.t193 0.7285
R930 avdd.n97 avdd.t189 0.7285
R931 avdd.n108 avdd.t131 0.7285
R932 avdd.n108 avdd.t73 0.7285
R933 avdd.n103 avdd.t139 0.7285
R934 avdd.n103 avdd.t191 0.7285
R935 avdd.n120 avdd.t197 0.7285
R936 avdd.n120 avdd.t273 0.7285
R937 avdd.n114 avdd.t58 0.7285
R938 avdd.n114 avdd.t173 0.7285
R939 avdd.n131 avdd.t149 0.7285
R940 avdd.n131 avdd.t97 0.7285
R941 avdd.n170 avdd.t263 0.7285
R942 avdd.n170 avdd.t187 0.7285
R943 avdd.n181 avdd.t359 0.7285
R944 avdd.n181 avdd.t127 0.7285
R945 avdd.n176 avdd.t31 0.7285
R946 avdd.n176 avdd.t261 0.7285
R947 avdd.n193 avdd.t361 0.7285
R948 avdd.n193 avdd.t135 0.7285
R949 avdd.n187 avdd.t79 0.7285
R950 avdd.n187 avdd.t287 0.7285
R951 avdd.n204 avdd.t199 0.7285
R952 avdd.n204 avdd.t61 0.7285
R953 avdd.n243 avdd.t291 0.7285
R954 avdd.n243 avdd.t341 0.7285
R955 avdd.n254 avdd.t19 0.7285
R956 avdd.n254 avdd.t76 0.7285
R957 avdd.n249 avdd.t315 0.7285
R958 avdd.n249 avdd.t181 0.7285
R959 avdd.n266 avdd.t343 0.7285
R960 avdd.n266 avdd.t269 0.7285
R961 avdd.n260 avdd.t40 0.7285
R962 avdd.n260 avdd.t375 0.7285
R963 avdd.n277 avdd.t205 0.7285
R964 avdd.n277 avdd.t109 0.7285
R965 avdd.n316 avdd.t241 0.7285
R966 avdd.n316 avdd.t177 0.7285
R967 avdd.n327 avdd.t355 0.7285
R968 avdd.n327 avdd.t64 0.7285
R969 avdd.n322 avdd.t1 0.7285
R970 avdd.n322 avdd.t239 0.7285
R971 avdd.n339 avdd.t179 0.7285
R972 avdd.n339 avdd.t275 0.7285
R973 avdd.n333 avdd.t115 0.7285
R974 avdd.n333 avdd.t219 0.7285
R975 avdd.n350 avdd.t249 0.7285
R976 avdd.n350 avdd.t85 0.7285
R977 avdd.n3 avdd.t29 0.7285
R978 avdd.n3 avdd.t15 0.7285
R979 avdd.n527 avdd.t133 0.7285
R980 avdd.n527 avdd.t91 0.7285
R981 avdd.n8 avdd.t301 0.7285
R982 avdd.n8 avdd.t309 0.7285
R983 avdd.n515 avdd.t13 0.7285
R984 avdd.n515 avdd.t357 0.7285
R985 avdd.n521 avdd.t121 0.7285
R986 avdd.n521 avdd.t319 0.7285
R987 avdd.n464 avdd.t201 0.7285
R988 avdd.n464 avdd.t124 0.7285
R989 avdd.n509 avdd.n500 0.561043
R990 avdd.n443 avdd.n434 0.561043
R991 avdd.n369 avdd.n360 0.561043
R992 avdd.n296 avdd.n287 0.561043
R993 avdd.n223 avdd.n214 0.561043
R994 avdd.n150 avdd.n141 0.561043
R995 avdd.n154 avdd.n80 0.561043
R996 avdd.n153 avdd.n81 0.561043
R997 avdd.n139 avdd.n82 0.561043
R998 avdd.n162 avdd.n79 0.561043
R999 avdd.n227 avdd.n64 0.561043
R1000 avdd.n226 avdd.n65 0.561043
R1001 avdd.n212 avdd.n66 0.561043
R1002 avdd.n235 avdd.n63 0.561043
R1003 avdd.n300 avdd.n48 0.561043
R1004 avdd.n299 avdd.n49 0.561043
R1005 avdd.n285 avdd.n50 0.561043
R1006 avdd.n308 avdd.n47 0.561043
R1007 avdd.n373 avdd.n32 0.561043
R1008 avdd.n372 avdd.n33 0.561043
R1009 avdd.n358 avdd.n34 0.561043
R1010 avdd.n381 avdd.n31 0.561043
R1011 avdd.n447 avdd.n16 0.561043
R1012 avdd.n446 avdd.n17 0.561043
R1013 avdd.n432 avdd.n18 0.561043
R1014 avdd.n455 avdd.n15 0.561043
R1015 avdd.n497 avdd.n482 0.561043
R1016 avdd.n498 avdd.n472 0.561043
R1017 avdd.n512 avdd.n471 0.561043
R1018 avdd.n492 avdd.n483 0.561043
R1019 avdd.n488 avdd.n487 0.510024
R1020 avdd.n165 avdd.n163 0.490037
R1021 avdd.n238 avdd.n236 0.490037
R1022 avdd.n311 avdd.n309 0.490037
R1023 avdd.n384 avdd.n382 0.490037
R1024 avdd.n458 avdd.n456 0.490037
R1025 avdd.n165 avdd.n164 0.436534
R1026 avdd.n238 avdd.n237 0.436534
R1027 avdd.n311 avdd.n310 0.436534
R1028 avdd.n384 avdd.n383 0.436534
R1029 avdd.n458 avdd.n457 0.436534
R1030 avdd.n489 avdd.n488 0.415037
R1031 avdd.n509 avdd.n508 0.255737
R1032 avdd.n443 avdd.n442 0.255737
R1033 avdd.n369 avdd.n368 0.255737
R1034 avdd.n296 avdd.n295 0.255737
R1035 avdd.n223 avdd.n222 0.255737
R1036 avdd.n150 avdd.n149 0.255737
R1037 avdd.n163 avdd.n162 0.255737
R1038 avdd.n236 avdd.n235 0.255737
R1039 avdd.n309 avdd.n308 0.255737
R1040 avdd.n382 avdd.n381 0.255737
R1041 avdd.n456 avdd.n455 0.255737
R1042 avdd.n489 avdd.n483 0.255737
R1043 avdd.n162 avdd.n161 0.2165
R1044 avdd.n235 avdd.n234 0.2165
R1045 avdd.n308 avdd.n307 0.2165
R1046 avdd.n381 avdd.n380 0.2165
R1047 avdd.n455 avdd.n454 0.2165
R1048 avdd.n496 avdd.n483 0.2165
R1049 avdd.n161 avdd.n154 0.148424
R1050 avdd.n234 avdd.n227 0.148424
R1051 avdd.n307 avdd.n300 0.148424
R1052 avdd.n380 avdd.n373 0.148424
R1053 avdd.n454 avdd.n447 0.148424
R1054 avdd.n497 avdd.n496 0.148424
R1055 dffrs_1.resetb avdd.n423 0.136036
R1056 dffrs_5.resetb avdd.n130 0.136036
R1057 dffrs_4.resetb avdd.n203 0.136036
R1058 dffrs_3.resetb avdd.n276 0.136036
R1059 dffrs_2.resetb avdd.n349 0.136036
R1060 dffrs_0.resetb avdd.n463 0.136036
R1061 avdd.n510 avdd.n509 0.0635
R1062 avdd.n444 avdd.n443 0.0635
R1063 avdd.n370 avdd.n369 0.0635
R1064 avdd.n297 avdd.n296 0.0635
R1065 avdd.n224 avdd.n223 0.0635
R1066 avdd.n151 avdd.n150 0.0635
R1067 avdd.n154 avdd.n153 0.0452384
R1068 avdd.n227 avdd.n226 0.0452384
R1069 avdd.n300 avdd.n299 0.0452384
R1070 avdd.n373 avdd.n372 0.0452384
R1071 avdd.n447 avdd.n446 0.0452384
R1072 avdd.n498 avdd.n497 0.0452384
R1073 avdd.n119 avdd.n113 0.0405727
R1074 avdd.n192 avdd.n186 0.0405727
R1075 avdd.n265 avdd.n259 0.0405727
R1076 avdd.n338 avdd.n332 0.0405727
R1077 avdd.n411 avdd.n405 0.0405727
R1078 avdd.n532 avdd.n526 0.0405727
R1079 avdd.n388 dffrs_1.setb 0.032
R1080 avdd.n96 dffrs_5.setb 0.032
R1081 avdd.n169 dffrs_4.setb 0.032
R1082 avdd.n242 dffrs_3.setb 0.032
R1083 avdd.n315 dffrs_2.setb 0.032
R1084 dffrs_0.setb avdd.n534 0.032
R1085 avdd.n508 avdd.n506 0.0313054
R1086 avdd.n508 avdd.n507 0.0313054
R1087 avdd.n442 avdd.n440 0.0313054
R1088 avdd.n442 avdd.n441 0.0313054
R1089 avdd.n368 avdd.n366 0.0313054
R1090 avdd.n368 avdd.n367 0.0313054
R1091 avdd.n295 avdd.n293 0.0313054
R1092 avdd.n295 avdd.n294 0.0313054
R1093 avdd.n222 avdd.n220 0.0313054
R1094 avdd.n222 avdd.n221 0.0313054
R1095 avdd.n149 avdd.n147 0.0313054
R1096 avdd.n149 avdd.n148 0.0313054
R1097 avdd.n163 avdd.n77 0.0313054
R1098 avdd.n163 avdd.n78 0.0313054
R1099 avdd.n236 avdd.n61 0.0313054
R1100 avdd.n236 avdd.n62 0.0313054
R1101 avdd.n309 avdd.n45 0.0313054
R1102 avdd.n309 avdd.n46 0.0313054
R1103 avdd.n382 avdd.n29 0.0313054
R1104 avdd.n382 avdd.n30 0.0313054
R1105 avdd.n456 avdd.n13 0.0313054
R1106 avdd.n456 avdd.n14 0.0313054
R1107 avdd.n490 avdd.n489 0.0313054
R1108 avdd.n489 avdd.n486 0.0313054
R1109 avdd.n152 avdd.n139 0.0295407
R1110 avdd.n225 avdd.n212 0.0295407
R1111 avdd.n298 avdd.n285 0.0295407
R1112 avdd.n371 avdd.n358 0.0295407
R1113 avdd.n445 avdd.n432 0.0295407
R1114 avdd.n512 avdd.n511 0.0295407
R1115 avdd.n137 avdd.n125 0.0288636
R1116 avdd.n210 avdd.n198 0.0288636
R1117 avdd.n283 avdd.n271 0.0288636
R1118 avdd.n356 avdd.n344 0.0288636
R1119 avdd.n520 avdd.n514 0.0288636
R1120 avdd.n418 avdd.n417 0.0288455
R1121 avdd.n113 avdd.n102 0.0237
R1122 avdd.n186 avdd.n175 0.0237
R1123 avdd.n259 avdd.n248 0.0237
R1124 avdd.n332 avdd.n321 0.0237
R1125 avdd.n405 avdd.n394 0.0237
R1126 avdd.n533 avdd.n532 0.0237
R1127 avdd.n153 avdd.n152 0.0161977
R1128 avdd.n226 avdd.n225 0.0161977
R1129 avdd.n299 avdd.n298 0.0161977
R1130 avdd.n372 avdd.n371 0.0161977
R1131 avdd.n446 avdd.n445 0.0161977
R1132 avdd.n511 avdd.n498 0.0161977
R1133 avdd.n139 avdd.n138 0.0129273
R1134 avdd.n212 avdd.n211 0.0129273
R1135 avdd.n285 avdd.n284 0.0129273
R1136 avdd.n358 avdd.n357 0.0129273
R1137 avdd.n432 avdd.n431 0.0129273
R1138 avdd.n513 avdd.n512 0.0129273
R1139 avdd.n488 avdd 0.0128676
R1140 avdd.n137 avdd.n136 0.0122273
R1141 avdd.n210 avdd.n209 0.0122273
R1142 avdd.n283 avdd.n282 0.0122273
R1143 avdd.n356 avdd.n355 0.0122273
R1144 avdd.n430 avdd.n429 0.0122273
R1145 avdd.n514 avdd.n469 0.0122273
R1146 avdd.n125 avdd.n119 0.000518182
R1147 avdd.n198 avdd.n192 0.000518182
R1148 avdd.n271 avdd.n265 0.000518182
R1149 avdd.n344 avdd.n338 0.000518182
R1150 avdd.n417 avdd.n411 0.000518182
R1151 avdd.n430 avdd.n418 0.000518182
R1152 avdd.n526 avdd.n520 0.000518182
R1153 avss.n259 avss.n258 21124.8
R1154 avss.n216 avss.n215 21124.8
R1155 avss.n173 avss.n172 21124.8
R1156 avss.n124 avss.n51 21034.5
R1157 avss.n787 avss.n786 21034.5
R1158 avss.n321 avss.n301 21026.3
R1159 avss.n374 avss.n373 21012.5
R1160 avss.n474 avss.n473 21012.5
R1161 avss.n574 avss.n573 21012.5
R1162 avss.n674 avss.n673 21012.5
R1163 avss.n757 avss.n756 21000
R1164 avss.n825 avss.n824 21000
R1165 avss.n381 avss.n267 16221.9
R1166 avss.n481 avss.n224 16221.9
R1167 avss.n581 avss.n181 16221.9
R1168 avss.n681 avss.n132 16221.9
R1169 avss.n785 avss.n53 16221.9
R1170 avss.n836 avss.n833 11510.4
R1171 avss.n382 avss.n381 11510.4
R1172 avss.n482 avss.n481 11510.4
R1173 avss.n582 avss.n581 11510.4
R1174 avss.n682 avss.n681 11510.4
R1175 avss.n764 avss.n53 11510.4
R1176 avss.n836 avss.n6 11510.4
R1177 avss.n826 avss.n825 7422.73
R1178 avss.n758 avss.n757 7422.73
R1179 avss.n373 avss.n372 7422.62
R1180 avss.n473 avss.n472 7422.62
R1181 avss.n573 avss.n572 7422.62
R1182 avss.n673 avss.n672 7422.62
R1183 avss.n423 avss.n422 6961.73
R1184 avss.n523 avss.n522 6961.73
R1185 avss.n623 avss.n622 6961.73
R1186 avss.n716 avss.n715 6961.73
R1187 avss.n55 avss.n50 6961.73
R1188 avss.n854 avss.n5 6190.48
R1189 avss.n781 avss.n81 6190.48
R1190 avss.n699 avss.n139 6190.48
R1191 avss.n606 avss.n182 6190.48
R1192 avss.n506 avss.n225 6190.48
R1193 avss.n406 avss.n268 6190.48
R1194 avss.n323 avss.n322 5557.62
R1195 avss.n323 avss.n291 5551.58
R1196 avss.n423 avss.n250 5551.58
R1197 avss.n523 avss.n207 5551.58
R1198 avss.n623 avss.n164 5551.58
R1199 avss.n716 avss.n116 5551.58
R1200 avss.n55 avss.n42 5551.58
R1201 avss.n408 avss.n249 5290.17
R1202 avss.n508 avss.n206 5290.17
R1203 avss.n608 avss.n163 5290.17
R1204 avss.n701 avss.n115 5286.93
R1205 avss.n783 avss.n41 5286.93
R1206 avss.n854 avss.n853 4683.14
R1207 avss.n300 avss.n299 4273.71
R1208 avss.n409 avss.n408 4062.5
R1209 avss.n509 avss.n508 4062.5
R1210 avss.n609 avss.n608 4062.5
R1211 avss.n702 avss.n701 4062.5
R1212 avss.n784 avss.n783 4062.5
R1213 avss.n322 avss.n300 3568.02
R1214 avss.n854 avss.n6 3123.51
R1215 avss.n374 avss.n284 2944.22
R1216 avss.n474 avss.n241 2944.22
R1217 avss.n574 avss.n198 2944.22
R1218 avss.n674 avss.n155 2944.22
R1219 avss.n756 avss.n750 2944.22
R1220 avss.n824 avss.n822 2944.22
R1221 avss.n267 avss.n258 2845.46
R1222 avss.n224 avss.n215 2845.46
R1223 avss.n181 avss.n172 2845.46
R1224 avss.n786 avss.n785 2845.46
R1225 avss.n132 avss.n124 2843.75
R1226 avss.n325 avss.n283 2257.8
R1227 avss.n425 avss.n240 2257.8
R1228 avss.n525 avss.n197 2257.8
R1229 avss.n625 avss.n154 2257.8
R1230 avss.n97 avss.n52 2257.8
R1231 avss.n789 avss.n23 2257.8
R1232 avss.n702 avss.n132 1878.69
R1233 avss.n409 avss.n267 1876.98
R1234 avss.n509 avss.n224 1876.98
R1235 avss.n609 avss.n181 1876.98
R1236 avss.n785 avss.n784 1876.98
R1237 avss.n347 avss.n346 1486.9
R1238 avss.n309 avss.n300 1212.42
R1239 avss.n422 avss.n258 1205.08
R1240 avss.n522 avss.n215 1205.08
R1241 avss.n622 avss.n172 1205.08
R1242 avss.n715 avss.n124 1205.08
R1243 avss.n786 avss.n50 1205.08
R1244 avss.n301 avss.n267 1135.55
R1245 avss.n259 avss.n224 1135.55
R1246 avss.n216 avss.n181 1135.55
R1247 avss.n173 avss.n132 1135.55
R1248 avss.n785 avss.n51 1135.55
R1249 avss.n788 avss.n787 1135.55
R1250 avss.n325 avss.n267 1122.24
R1251 avss.n425 avss.n224 1122.24
R1252 avss.n525 avss.n181 1122.24
R1253 avss.n625 avss.n132 1122.24
R1254 avss.n785 avss.n52 1122.24
R1255 avss.n789 avss.n788 1122.24
R1256 avss.n739 avss.n738 977.434
R1257 avss.n811 avss.n810 977.434
R1258 avss.n447 avss.n446 977.068
R1259 avss.n547 avss.n546 977.068
R1260 avss.n647 avss.n646 977.068
R1261 avss.n738 avss.n115 904.402
R1262 avss.n810 avss.n41 904.402
R1263 avss.n446 avss.n249 904.062
R1264 avss.n546 avss.n206 904.062
R1265 avss.n646 avss.n163 904.062
R1266 avss.n322 avss.n321 897.806
R1267 avss.n323 avss.n298 832.22
R1268 avss.n423 avss.n257 832.22
R1269 avss.n523 avss.n214 832.22
R1270 avss.n623 avss.n171 832.22
R1271 avss.n716 avss.n123 832.22
R1272 avss.n56 avss.n55 832.22
R1273 avss.n324 avss.n323 832.101
R1274 avss.n424 avss.n423 832.101
R1275 avss.n524 avss.n523 832.101
R1276 avss.n624 avss.n623 832.101
R1277 avss.n717 avss.n716 832.101
R1278 avss.n55 avss.n54 832.101
R1279 avss.n75 avss.n41 784.409
R1280 avss.n133 avss.n115 784.37
R1281 avss.n588 avss.n163 784.37
R1282 avss.n488 avss.n206 784.37
R1283 avss.n388 avss.n249 784.37
R1284 avss.n788 avss.n6 697.039
R1285 avss.n374 avss.n283 665.564
R1286 avss.n474 avss.n240 665.564
R1287 avss.n574 avss.n197 665.564
R1288 avss.n674 avss.n154 665.564
R1289 avss.n756 avss.n97 665.564
R1290 avss.n824 avss.n23 665.564
R1291 avss.n822 avss.n821 654.253
R1292 avss.n750 avss.n749 654.253
R1293 avss.n156 avss.n155 654.005
R1294 avss.n199 avss.n198 654.005
R1295 avss.n242 avss.n241 654.005
R1296 avss.n285 avss.n284 654.005
R1297 avss.n750 avss.n98 648.784
R1298 avss.n822 avss.n24 648.784
R1299 avss.n348 avss.n284 648.54
R1300 avss.n448 avss.n241 648.54
R1301 avss.n548 avss.n198 648.54
R1302 avss.n648 avss.n155 648.54
R1303 avss.t210 avss.n826 590.909
R1304 avss.n827 avss.t210 590.909
R1305 avss.n827 avss.t117 590.909
R1306 avss.n833 avss.t101 590.909
R1307 avss.n833 avss.t24 590.909
R1308 avss.t26 avss.n832 590.909
R1309 avss.t7 avss.n375 590.909
R1310 avss.n379 avss.t7 590.909
R1311 avss.t278 avss.n379 590.909
R1312 avss.n381 avss.t158 590.909
R1313 avss.n381 avss.t279 590.909
R1314 avss.n405 avss.t251 590.909
R1315 avss.t164 avss.n475 590.909
R1316 avss.n479 avss.t164 590.909
R1317 avss.t277 avss.n479 590.909
R1318 avss.n481 avss.t168 590.909
R1319 avss.n481 avss.t204 590.909
R1320 avss.n505 avss.t190 590.909
R1321 avss.t95 avss.n575 590.909
R1322 avss.n579 avss.t95 590.909
R1323 avss.t217 avss.n579 590.909
R1324 avss.n581 avss.t256 590.909
R1325 avss.n581 avss.t178 590.909
R1326 avss.n605 avss.t182 590.909
R1327 avss.t42 avss.n675 590.909
R1328 avss.n679 avss.t42 590.909
R1329 avss.t133 avss.n679 590.909
R1330 avss.n681 avss.t176 590.909
R1331 avss.n681 avss.t262 590.909
R1332 avss.n698 avss.t264 590.909
R1333 avss.t113 avss.n758 590.909
R1334 avss.n762 avss.t113 590.909
R1335 avss.t44 avss.n762 590.909
R1336 avss.n764 avss.t253 590.909
R1337 avss.t38 avss.n764 590.909
R1338 avss.n765 avss.t36 590.909
R1339 avss.n755 avss.t268 590.909
R1340 avss.t268 avss.n754 590.909
R1341 avss.n754 avss.t276 590.909
R1342 avss.t177 avss.n53 590.909
R1343 avss.t102 avss.n53 590.909
R1344 avss.n780 avss.t93 590.909
R1345 avss.n823 avss.t107 590.909
R1346 avss.n837 avss.t107 590.909
R1347 avss.n837 avss.t169 590.909
R1348 avss.t272 avss.n836 590.909
R1349 avss.n836 avss.t246 590.909
R1350 avss.n855 avss.t243 590.909
R1351 avss.n372 avss.t214 590.462
R1352 avss.t214 avss.n371 590.462
R1353 avss.n371 avss.t229 590.462
R1354 avss.n382 avss.t45 590.462
R1355 avss.t14 avss.n382 590.462
R1356 avss.n383 avss.t12 590.462
R1357 avss.n472 avss.t120 590.462
R1358 avss.t120 avss.n471 590.462
R1359 avss.n471 avss.t260 590.462
R1360 avss.n482 avss.t23 590.462
R1361 avss.t109 avss.n482 590.462
R1362 avss.n483 avss.t111 590.462
R1363 avss.n572 avss.t172 590.462
R1364 avss.t172 avss.n571 590.462
R1365 avss.n571 avss.t129 590.462
R1366 avss.n582 avss.t261 590.462
R1367 avss.t30 avss.n582 590.462
R1368 avss.n583 avss.t32 590.462
R1369 avss.n672 avss.t192 590.462
R1370 avss.t192 avss.n671 590.462
R1371 avss.n671 avss.t9 590.462
R1372 avss.n682 avss.t16 590.462
R1373 avss.t3 avss.n682 590.462
R1374 avss.n683 avss.t5 590.462
R1375 avss.n309 avss.t98 582.165
R1376 avss.t52 avss.n298 582.165
R1377 avss.n410 avss.t35 582.165
R1378 avss.t75 avss.n257 582.165
R1379 avss.n510 avss.t241 582.165
R1380 avss.t56 avss.n214 582.165
R1381 avss.n610 avss.t0 582.165
R1382 avss.t79 avss.n171 582.165
R1383 avss.n703 avss.t283 582.165
R1384 avss.t69 avss.n123 582.165
R1385 avss.n74 avss.t232 582.165
R1386 avss.n56 avss.t46 582.165
R1387 avss.t275 avss.n324 581.712
R1388 avss.n326 avss.t153 581.712
R1389 avss.n320 avss.t149 581.712
R1390 avss.n302 avss.t58 581.712
R1391 avss.t90 avss.n424 581.712
R1392 avss.n426 avss.t186 581.712
R1393 avss.n421 avss.t208 581.712
R1394 avss.n260 avss.t86 581.712
R1395 avss.t273 avss.n524 581.712
R1396 avss.n526 avss.t197 581.712
R1397 avss.n521 avss.t140 581.712
R1398 avss.n217 avss.t67 581.712
R1399 avss.t20 avss.n624 581.712
R1400 avss.n626 avss.t146 581.712
R1401 avss.n621 avss.t222 581.712
R1402 avss.n174 avss.t81 581.712
R1403 avss.t289 avss.n717 581.712
R1404 avss.n718 avss.t115 581.712
R1405 avss.n714 avss.t233 581.712
R1406 avss.n125 avss.t72 581.712
R1407 avss.n54 avss.t212 581.712
R1408 avss.n790 avss.t118 581.712
R1409 avss.n60 avss.t236 581.712
R1410 avss.t50 avss.n49 581.712
R1411 avss.t145 avss.n334 581.712
R1412 avss.n335 avss.t150 581.712
R1413 avss.t143 avss.n434 581.712
R1414 avss.n435 avss.t206 581.712
R1415 avss.t270 avss.n534 581.712
R1416 avss.n535 avss.t138 581.712
R1417 avss.t134 avss.n634 581.712
R1418 avss.n635 avss.t224 581.712
R1419 avss.t188 avss.n726 581.712
R1420 avss.n727 avss.t258 581.712
R1421 avss.t1 avss.n798 581.712
R1422 avss.n799 avss.t237 581.712
R1423 avss.n701 avss.n699 574.192
R1424 avss.n408 avss.n406 574.061
R1425 avss.n508 avss.n506 574.061
R1426 avss.n608 avss.n606 574.061
R1427 avss.n783 avss.n781 574.061
R1428 avss.n334 avss.n291 548.058
R1429 avss.n434 avss.n250 548.058
R1430 avss.n534 avss.n207 548.058
R1431 avss.n634 avss.n164 548.058
R1432 avss.n726 avss.n116 548.058
R1433 avss.n798 avss.n42 548.058
R1434 avss.t117 avss.t101 502.274
R1435 avss.t24 avss.t26 502.274
R1436 avss.t158 avss.t278 502.274
R1437 avss.t279 avss.t251 502.274
R1438 avss.t168 avss.t277 502.274
R1439 avss.t204 avss.t190 502.274
R1440 avss.t256 avss.t217 502.274
R1441 avss.t178 avss.t182 502.274
R1442 avss.t176 avss.t133 502.274
R1443 avss.t262 avss.t264 502.274
R1444 avss.t253 avss.t44 502.274
R1445 avss.t36 avss.t38 502.274
R1446 avss.t276 avss.t177 502.274
R1447 avss.t93 avss.t102 502.274
R1448 avss.t169 avss.t272 502.274
R1449 avss.t246 avss.t243 502.274
R1450 avss.t229 avss.t45 501.892
R1451 avss.t12 avss.t14 501.892
R1452 avss.t260 avss.t23 501.892
R1453 avss.t111 avss.t109 501.892
R1454 avss.t129 avss.t261 501.892
R1455 avss.t32 avss.t30 501.892
R1456 avss.t9 avss.t16 501.892
R1457 avss.t5 avss.t3 501.892
R1458 avss.n345 avss.n291 484.702
R1459 avss.n445 avss.n250 484.702
R1460 avss.n545 avss.n207 484.702
R1461 avss.n645 avss.n164 484.702
R1462 avss.n737 avss.n116 484.702
R1463 avss.n809 avss.n42 484.702
R1464 avss.t98 avss.t148 465.733
R1465 avss.t148 avss.t52 465.733
R1466 avss.t35 avss.t209 465.733
R1467 avss.t209 avss.t75 465.733
R1468 avss.t241 avss.t226 465.733
R1469 avss.t226 avss.t56 465.733
R1470 avss.t0 avss.t223 465.733
R1471 avss.t223 avss.t79 465.733
R1472 avss.t283 avss.t216 465.733
R1473 avss.t216 avss.t69 465.733
R1474 avss.t34 avss.t232 465.733
R1475 avss.t46 avss.t34 465.733
R1476 avss.t83 avss.t275 465.37
R1477 avss.t153 avss.t83 465.37
R1478 avss.t152 avss.t149 465.37
R1479 avss.t58 avss.t152 465.37
R1480 avss.t64 avss.t90 465.37
R1481 avss.t186 avss.t64 465.37
R1482 avss.t144 avss.t208 465.37
R1483 avss.t86 avss.t144 465.37
R1484 avss.t84 avss.t273 465.37
R1485 avss.t197 avss.t84 465.37
R1486 avss.t271 avss.t140 465.37
R1487 avss.t67 avss.t271 465.37
R1488 avss.t77 avss.t20 465.37
R1489 avss.t146 avss.t77 465.37
R1490 avss.t135 avss.t222 465.37
R1491 avss.t81 avss.t135 465.37
R1492 avss.t62 avss.t289 465.37
R1493 avss.t115 avss.t62 465.37
R1494 avss.t189 avss.t233 465.37
R1495 avss.t72 avss.t189 465.37
R1496 avss.t212 avss.t48 465.37
R1497 avss.t48 avss.t118 465.37
R1498 avss.t236 avss.t2 465.37
R1499 avss.t2 avss.t50 465.37
R1500 avss.t92 avss.t145 465.37
R1501 avss.t150 avss.t92 465.37
R1502 avss.t274 avss.t143 465.37
R1503 avss.t206 avss.t274 465.37
R1504 avss.t91 avss.t270 465.37
R1505 avss.t138 avss.t91 465.37
R1506 avss.t257 avss.t134 465.37
R1507 avss.t224 avss.t257 465.37
R1508 avss.t213 avss.t188 465.37
R1509 avss.t258 avss.t213 465.37
R1510 avss.t19 avss.t1 465.37
R1511 avss.t237 avss.t19 465.37
R1512 avss.n832 avss.n5 361.01
R1513 avss.n765 avss.n81 361.01
R1514 avss.n683 avss.n139 360.803
R1515 avss.n583 avss.n182 360.803
R1516 avss.n483 avss.n225 360.803
R1517 avss.n383 avss.n268 360.803
R1518 avss.n80 avss.t218 348.214
R1519 avss.n75 avss.t218 348.214
R1520 avss.n7 avss.t227 348.214
R1521 avss.n853 avss.t227 348.214
R1522 avss.n138 avss.t166 348.06
R1523 avss.n133 avss.t166 348.06
R1524 avss.t170 avss.n587 348.06
R1525 avss.n588 avss.t170 348.06
R1526 avss.t254 avss.n487 348.06
R1527 avss.n488 avss.t254 348.06
R1528 avss.t156 avss.n387 348.06
R1529 avss.n388 avss.t156 348.06
R1530 avss.n299 avss.t74 338.849
R1531 avss.t122 avss.n345 338.849
R1532 avss.n407 avss.t85 338.849
R1533 avss.n507 avss.t66 338.849
R1534 avss.n607 avss.t61 338.849
R1535 avss.n700 avss.t55 338.849
R1536 avss.n782 avss.t63 338.849
R1537 avss.n821 avss.t141 314.01
R1538 avss.n33 avss.t141 314.01
R1539 avss.n32 avss.t17 314.01
R1540 avss.n29 avss.t17 314.01
R1541 avss.n28 avss.t284 314.01
R1542 avss.t284 avss.n22 314.01
R1543 avss.n749 avss.t195 314.01
R1544 avss.n107 avss.t195 314.01
R1545 avss.n106 avss.t10 314.01
R1546 avss.n103 avss.t10 314.01
R1547 avss.n102 avss.t40 314.01
R1548 avss.t40 avss.n96 314.01
R1549 avss.n156 avss.t174 313.884
R1550 avss.n658 avss.t174 313.884
R1551 avss.n659 avss.t28 313.884
R1552 avss.n663 avss.t28 313.884
R1553 avss.t99 avss.n666 313.884
R1554 avss.n667 avss.t99 313.884
R1555 avss.n199 avss.t286 313.884
R1556 avss.n558 avss.t286 313.884
R1557 avss.n559 avss.t88 313.884
R1558 avss.n563 avss.t88 313.884
R1559 avss.t230 avss.n566 313.884
R1560 avss.n567 avss.t230 313.884
R1561 avss.n242 avss.t234 313.884
R1562 avss.n458 avss.t234 313.884
R1563 avss.n459 avss.t239 313.884
R1564 avss.n463 avss.t239 313.884
R1565 avss.t184 avss.n466 313.884
R1566 avss.n467 avss.t184 313.884
R1567 avss.n285 avss.t162 313.884
R1568 avss.n358 avss.t162 313.884
R1569 avss.n359 avss.t21 313.884
R1570 avss.n363 avss.t21 313.884
R1571 avss.t160 avss.n366 313.884
R1572 avss.n367 avss.t160 313.884
R1573 avss.n81 avss.n80 300.336
R1574 avss.n7 avss.n5 300.336
R1575 avss.n139 avss.n138 300.202
R1576 avss.n587 avss.n182 300.202
R1577 avss.n487 avss.n225 300.202
R1578 avss.n387 avss.n268 300.202
R1579 avss.n739 avss.t124 279.964
R1580 avss.t199 avss.n98 279.964
R1581 avss.n811 avss.t97 279.964
R1582 avss.t248 avss.n24 279.964
R1583 avss.t106 avss.n347 279.858
R1584 avss.n348 avss.t131 279.858
R1585 avss.t128 avss.n447 279.858
R1586 avss.n448 avss.t220 279.858
R1587 avss.t155 avss.n547 279.858
R1588 avss.n548 avss.t136 279.858
R1589 avss.t194 avss.n647 279.858
R1590 avss.n648 avss.t126 279.858
R1591 avss.t130 avss.t122 271.079
R1592 avss.t85 avss.t159 271.079
R1593 avss.t159 avss.t281 271.079
R1594 avss.t66 avss.t288 271.079
R1595 avss.t288 avss.t202 271.079
R1596 avss.t61 avss.t125 271.079
R1597 avss.t125 avss.t180 271.079
R1598 avss.t55 avss.t201 271.079
R1599 avss.t201 avss.t266 271.079
R1600 avss.t63 avss.t250 271.079
R1601 avss.t250 avss.t104 271.079
R1602 avss.n33 avss.n32 266.909
R1603 avss.n29 avss.n28 266.909
R1604 avss.n107 avss.n106 266.909
R1605 avss.n103 avss.n102 266.909
R1606 avss.n659 avss.n658 266.801
R1607 avss.n666 avss.n663 266.801
R1608 avss.n559 avss.n558 266.801
R1609 avss.n566 avss.n563 266.801
R1610 avss.n459 avss.n458 266.801
R1611 avss.n466 avss.n463 266.801
R1612 avss.n359 avss.n358 266.801
R1613 avss.n366 avss.n363 266.801
R1614 avss.t124 avss.t71 223.97
R1615 avss.t71 avss.t199 223.97
R1616 avss.t97 avss.t65 223.97
R1617 avss.t65 avss.t248 223.97
R1618 avss.t54 avss.t106 223.887
R1619 avss.t131 avss.t54 223.887
R1620 avss.t78 avss.t128 223.887
R1621 avss.t220 avss.t78 223.887
R1622 avss.t60 avss.t155 223.887
R1623 avss.t136 avss.t60 223.887
R1624 avss.t49 avss.t194 223.887
R1625 avss.t126 avss.t49 223.887
R1626 avss.n346 avss.t130 220.988
R1627 avss.n446 avss.n445 213.623
R1628 avss.n546 avss.n545 213.623
R1629 avss.n646 avss.n645 213.623
R1630 avss.n738 avss.n737 213.623
R1631 avss.n810 avss.n809 213.623
R1632 avss.n410 avss.n409 151.869
R1633 avss.n510 avss.n509 151.869
R1634 avss.n610 avss.n609 151.869
R1635 avss.n703 avss.n702 151.869
R1636 avss.n784 avss.n74 151.869
R1637 avss.n326 avss.n325 151.751
R1638 avss.n321 avss.n320 151.751
R1639 avss.n302 avss.n301 151.751
R1640 avss.n426 avss.n425 151.751
R1641 avss.n422 avss.n421 151.751
R1642 avss.n260 avss.n259 151.751
R1643 avss.n526 avss.n525 151.751
R1644 avss.n522 avss.n521 151.751
R1645 avss.n217 avss.n216 151.751
R1646 avss.n626 avss.n625 151.751
R1647 avss.n622 avss.n621 151.751
R1648 avss.n174 avss.n173 151.751
R1649 avss.n718 avss.n52 151.751
R1650 avss.n715 avss.n714 151.751
R1651 avss.n125 avss.n51 151.751
R1652 avss.n790 avss.n789 151.751
R1653 avss.n60 avss.n50 151.751
R1654 avss.n787 avss.n49 151.751
R1655 avss.n335 avss.n283 151.751
R1656 avss.n435 avss.n240 151.751
R1657 avss.n535 avss.n197 151.751
R1658 avss.n635 avss.n154 151.751
R1659 avss.n727 avss.n97 151.751
R1660 avss.n799 avss.n23 151.751
R1661 avss.n375 avss.n374 147.727
R1662 avss.n406 avss.n405 147.727
R1663 avss.n475 avss.n474 147.727
R1664 avss.n506 avss.n505 147.727
R1665 avss.n575 avss.n574 147.727
R1666 avss.n606 avss.n605 147.727
R1667 avss.n675 avss.n674 147.727
R1668 avss.n699 avss.n698 147.727
R1669 avss.n756 avss.n755 147.727
R1670 avss.n781 avss.n780 147.727
R1671 avss.n824 avss.n823 147.727
R1672 avss.n855 avss.n854 147.727
R1673 avss.n446 avss.t281 125.228
R1674 avss.n546 avss.t202 125.228
R1675 avss.n646 avss.t180 125.228
R1676 avss.n738 avss.t266 125.228
R1677 avss.n810 avss.t104 125.228
R1678 avss.n408 avss.n407 88.3958
R1679 avss.n508 avss.n507 88.3958
R1680 avss.n608 avss.n607 88.3958
R1681 avss.n701 avss.n700 88.3958
R1682 avss.n783 avss.n782 88.3958
R1683 avss.n856 avss.n3 87.3061
R1684 avss.n856 avss.n4 87.3061
R1685 avss.n779 avss.n82 87.3061
R1686 avss.n779 avss.n83 87.3061
R1687 avss.n766 avss.n94 87.3061
R1688 avss.n766 avss.n95 87.3061
R1689 avss.n697 avss.n140 87.3061
R1690 avss.n697 avss.n141 87.3061
R1691 avss.n684 avss.n151 87.3061
R1692 avss.n684 avss.n152 87.3061
R1693 avss.n604 avss.n183 87.3061
R1694 avss.n604 avss.n184 87.3061
R1695 avss.n584 avss.n194 87.3061
R1696 avss.n584 avss.n195 87.3061
R1697 avss.n504 avss.n226 87.3061
R1698 avss.n504 avss.n227 87.3061
R1699 avss.n484 avss.n237 87.3061
R1700 avss.n484 avss.n238 87.3061
R1701 avss.n404 avss.n269 87.3061
R1702 avss.n404 avss.n270 87.3061
R1703 avss.n384 avss.n280 87.3061
R1704 avss.n384 avss.n281 87.3061
R1705 avss.n831 avss.n20 87.3061
R1706 avss.n831 avss.n830 87.3061
R1707 avss.n825 avss.n22 78.5029
R1708 avss.n757 avss.n96 78.5029
R1709 avss.n673 avss.n667 78.4713
R1710 avss.n573 avss.n567 78.4713
R1711 avss.n473 avss.n467 78.4713
R1712 avss.n373 avss.n367 78.4713
R1713 avss.n17 avss.n16 67.4727
R1714 avss.n18 avss.n16 67.4727
R1715 avss.n751 avss.n87 67.4727
R1716 avss.n752 avss.n87 67.4727
R1717 avss.n759 avss.n91 67.4727
R1718 avss.n760 avss.n91 67.4727
R1719 avss.n676 avss.n144 67.4727
R1720 avss.n677 avss.n144 67.4727
R1721 avss.n668 avss.n148 67.4727
R1722 avss.n669 avss.n148 67.4727
R1723 avss.n576 avss.n187 67.4727
R1724 avss.n577 avss.n187 67.4727
R1725 avss.n568 avss.n191 67.4727
R1726 avss.n569 avss.n191 67.4727
R1727 avss.n476 avss.n230 67.4727
R1728 avss.n477 avss.n230 67.4727
R1729 avss.n468 avss.n234 67.4727
R1730 avss.n469 avss.n234 67.4727
R1731 avss.n376 avss.n273 67.4727
R1732 avss.n377 avss.n273 67.4727
R1733 avss.n368 avss.n277 67.4727
R1734 avss.n369 avss.n277 67.4727
R1735 avss.n21 avss.n12 67.4727
R1736 avss.n829 avss.n12 67.4727
R1737 avss.n17 avss.n3 66.5005
R1738 avss.n18 avss.n4 66.5005
R1739 avss.n751 avss.n82 66.5005
R1740 avss.n752 avss.n83 66.5005
R1741 avss.n759 avss.n94 66.5005
R1742 avss.n760 avss.n95 66.5005
R1743 avss.n676 avss.n140 66.5005
R1744 avss.n677 avss.n141 66.5005
R1745 avss.n668 avss.n151 66.5005
R1746 avss.n669 avss.n152 66.5005
R1747 avss.n576 avss.n183 66.5005
R1748 avss.n577 avss.n184 66.5005
R1749 avss.n568 avss.n194 66.5005
R1750 avss.n569 avss.n195 66.5005
R1751 avss.n476 avss.n226 66.5005
R1752 avss.n477 avss.n227 66.5005
R1753 avss.n468 avss.n237 66.5005
R1754 avss.n469 avss.n238 66.5005
R1755 avss.n376 avss.n269 66.5005
R1756 avss.n377 avss.n270 66.5005
R1757 avss.n368 avss.n280 66.5005
R1758 avss.n369 avss.n281 66.5005
R1759 avss.n21 avss.n20 66.5005
R1760 avss.n830 avss.n829 66.5005
R1761 avss.n319 avss.n303 61.0571
R1762 avss.n420 avss.n261 61.0571
R1763 avss.n520 avss.n218 61.0571
R1764 avss.n620 avss.n175 61.0571
R1765 avss.n713 avss.n126 61.0571
R1766 avss.n62 avss.n61 61.0571
R1767 avss.n800 avss.n797 61.0561
R1768 avss.n808 avss.n43 61.0561
R1769 avss.n813 avss.n812 61.0561
R1770 avss.n728 avss.n725 61.0561
R1771 avss.n736 avss.n117 61.0561
R1772 avss.n741 avss.n740 61.0561
R1773 avss.n636 avss.n633 61.0561
R1774 avss.n644 avss.n165 61.0561
R1775 avss.n649 avss.n162 61.0561
R1776 avss.n536 avss.n533 61.0561
R1777 avss.n544 avss.n208 61.0561
R1778 avss.n549 avss.n205 61.0561
R1779 avss.n436 avss.n433 61.0561
R1780 avss.n444 avss.n251 61.0561
R1781 avss.n449 avss.n248 61.0561
R1782 avss.n336 avss.n333 61.0561
R1783 avss.n344 avss.n292 61.0561
R1784 avss.n349 avss.n290 61.0561
R1785 avss.n327 avss.n297 61.0561
R1786 avss.n311 avss.n310 61.0561
R1787 avss.n427 avss.n256 61.0561
R1788 avss.n412 avss.n411 61.0561
R1789 avss.n527 avss.n213 61.0561
R1790 avss.n512 avss.n511 61.0561
R1791 avss.n627 avss.n170 61.0561
R1792 avss.n612 avss.n611 61.0561
R1793 avss.n719 avss.n122 61.0561
R1794 avss.n705 avss.n704 61.0561
R1795 avss.n791 avss.n48 61.0561
R1796 avss.n73 avss.n57 61.0561
R1797 avss.n346 avss.t74 50.0912
R1798 avss.n31 avss.n30 44.1404
R1799 avss.n27 avss.n13 44.1404
R1800 avss.n79 avss.n76 44.1404
R1801 avss.n105 avss.n104 44.1404
R1802 avss.n101 avss.n90 44.1404
R1803 avss.n137 avss.n134 44.1404
R1804 avss.n662 avss.n660 44.1404
R1805 avss.n665 avss.n147 44.1404
R1806 avss.n589 avss.n586 44.1404
R1807 avss.n562 avss.n560 44.1404
R1808 avss.n565 avss.n190 44.1404
R1809 avss.n489 avss.n486 44.1404
R1810 avss.n462 avss.n460 44.1404
R1811 avss.n465 avss.n233 44.1404
R1812 avss.n389 avss.n386 44.1404
R1813 avss.n852 avss.n8 44.1404
R1814 avss.n365 avss.n276 44.1394
R1815 avss.n362 avss.n360 44.1394
R1816 avss.n357 avss.n286 44.1394
R1817 avss.n820 avss.n34 44.1394
R1818 avss.n748 avss.n108 44.1394
R1819 avss.n657 avss.n157 44.1394
R1820 avss.n557 avss.n200 44.1394
R1821 avss.n457 avss.n243 44.1394
R1822 avss.n1 avss.t290 34.1066
R1823 avss.n835 avss.n3 20.8061
R1824 avss.n835 avss.n4 20.8061
R1825 avss.n838 avss.n17 20.8061
R1826 avss.n838 avss.n18 20.8061
R1827 avss.n84 avss.n82 20.8061
R1828 avss.n84 avss.n83 20.8061
R1829 avss.n753 avss.n751 20.8061
R1830 avss.n753 avss.n752 20.8061
R1831 avss.n763 avss.n94 20.8061
R1832 avss.n763 avss.n95 20.8061
R1833 avss.n761 avss.n759 20.8061
R1834 avss.n761 avss.n760 20.8061
R1835 avss.n680 avss.n140 20.8061
R1836 avss.n680 avss.n141 20.8061
R1837 avss.n678 avss.n676 20.8061
R1838 avss.n678 avss.n677 20.8061
R1839 avss.n153 avss.n151 20.8061
R1840 avss.n153 avss.n152 20.8061
R1841 avss.n670 avss.n668 20.8061
R1842 avss.n670 avss.n669 20.8061
R1843 avss.n580 avss.n183 20.8061
R1844 avss.n580 avss.n184 20.8061
R1845 avss.n578 avss.n576 20.8061
R1846 avss.n578 avss.n577 20.8061
R1847 avss.n196 avss.n194 20.8061
R1848 avss.n196 avss.n195 20.8061
R1849 avss.n570 avss.n568 20.8061
R1850 avss.n570 avss.n569 20.8061
R1851 avss.n480 avss.n226 20.8061
R1852 avss.n480 avss.n227 20.8061
R1853 avss.n478 avss.n476 20.8061
R1854 avss.n478 avss.n477 20.8061
R1855 avss.n239 avss.n237 20.8061
R1856 avss.n239 avss.n238 20.8061
R1857 avss.n470 avss.n468 20.8061
R1858 avss.n470 avss.n469 20.8061
R1859 avss.n380 avss.n269 20.8061
R1860 avss.n380 avss.n270 20.8061
R1861 avss.n378 avss.n376 20.8061
R1862 avss.n378 avss.n377 20.8061
R1863 avss.n282 avss.n280 20.8061
R1864 avss.n282 avss.n281 20.8061
R1865 avss.n370 avss.n368 20.8061
R1866 avss.n370 avss.n369 20.8061
R1867 avss.n828 avss.n21 20.8061
R1868 avss.n829 avss.n828 20.8061
R1869 avss.n20 avss.n19 20.8061
R1870 avss.n830 avss.n19 20.8061
R1871 avss.n0 avss.t245 19.673
R1872 avss.n0 avss.t242 19.4007
R1873 avss.n859 avss.n858 14.6135
R1874 avss.n289 avss.n287 9.0005
R1875 avss.n340 avss.n339 9.0005
R1876 avss.n318 avss.n317 9.0005
R1877 avss.n305 avss.n294 9.0005
R1878 avss.n308 avss.n307 9.0005
R1879 avss.n314 avss.n313 9.0005
R1880 avss.n296 avss.n295 9.0005
R1881 avss.n330 avss.n329 9.0005
R1882 avss.n338 avss.n288 9.0005
R1883 avss.n352 avss.n351 9.0005
R1884 avss.n247 avss.n245 9.0005
R1885 avss.n440 avss.n439 9.0005
R1886 avss.n419 avss.n418 9.0005
R1887 avss.n263 avss.n253 9.0005
R1888 avss.n266 avss.n265 9.0005
R1889 avss.n415 avss.n414 9.0005
R1890 avss.n255 avss.n254 9.0005
R1891 avss.n430 avss.n429 9.0005
R1892 avss.n438 avss.n246 9.0005
R1893 avss.n452 avss.n451 9.0005
R1894 avss.n204 avss.n202 9.0005
R1895 avss.n540 avss.n539 9.0005
R1896 avss.n519 avss.n518 9.0005
R1897 avss.n220 avss.n210 9.0005
R1898 avss.n223 avss.n222 9.0005
R1899 avss.n515 avss.n514 9.0005
R1900 avss.n212 avss.n211 9.0005
R1901 avss.n530 avss.n529 9.0005
R1902 avss.n538 avss.n203 9.0005
R1903 avss.n552 avss.n551 9.0005
R1904 avss.n161 avss.n159 9.0005
R1905 avss.n640 avss.n639 9.0005
R1906 avss.n619 avss.n618 9.0005
R1907 avss.n177 avss.n167 9.0005
R1908 avss.n180 avss.n179 9.0005
R1909 avss.n615 avss.n614 9.0005
R1910 avss.n169 avss.n168 9.0005
R1911 avss.n630 avss.n629 9.0005
R1912 avss.n638 avss.n160 9.0005
R1913 avss.n652 avss.n651 9.0005
R1914 avss.n114 avss.n112 9.0005
R1915 avss.n732 avss.n731 9.0005
R1916 avss.n712 avss.n711 9.0005
R1917 avss.n128 avss.n119 9.0005
R1918 avss.n131 avss.n130 9.0005
R1919 avss.n708 avss.n707 9.0005
R1920 avss.n121 avss.n120 9.0005
R1921 avss.n722 avss.n721 9.0005
R1922 avss.n730 avss.n113 9.0005
R1923 avss.n744 avss.n743 9.0005
R1924 avss.n40 avss.n38 9.0005
R1925 avss.n804 avss.n803 9.0005
R1926 avss.n66 avss.n65 9.0005
R1927 avss.n64 avss.n45 9.0005
R1928 avss.n72 avss.n58 9.0005
R1929 avss.n71 avss.n69 9.0005
R1930 avss.n47 avss.n46 9.0005
R1931 avss.n794 avss.n793 9.0005
R1932 avss.n802 avss.n39 9.0005
R1933 avss.n816 avss.n815 9.0005
R1934 avss.n342 avss.n292 6.9012
R1935 avss.n442 avss.n251 6.9012
R1936 avss.n542 avss.n208 6.9012
R1937 avss.n642 avss.n165 6.9012
R1938 avss.n734 avss.n117 6.9012
R1939 avss.n806 avss.n43 6.9012
R1940 avss.n339 avss.n333 6.46296
R1941 avss.n297 avss.n296 6.46296
R1942 avss.n310 avss.n308 6.46296
R1943 avss.n439 avss.n433 6.46296
R1944 avss.n256 avss.n255 6.46296
R1945 avss.n411 avss.n266 6.46296
R1946 avss.n539 avss.n533 6.46296
R1947 avss.n213 avss.n212 6.46296
R1948 avss.n511 avss.n223 6.46296
R1949 avss.n639 avss.n633 6.46296
R1950 avss.n170 avss.n169 6.46296
R1951 avss.n611 avss.n180 6.46296
R1952 avss.n731 avss.n725 6.46296
R1953 avss.n122 avss.n121 6.46296
R1954 avss.n704 avss.n131 6.46296
R1955 avss.n803 avss.n797 6.46296
R1956 avss.n48 avss.n47 6.46296
R1957 avss.n73 avss.n72 6.46296
R1958 avss.n290 avss.n289 6.4618
R1959 avss.n319 avss.n318 6.4618
R1960 avss.n248 avss.n247 6.4618
R1961 avss.n420 avss.n419 6.4618
R1962 avss.n205 avss.n204 6.4618
R1963 avss.n520 avss.n519 6.4618
R1964 avss.n162 avss.n161 6.4618
R1965 avss.n620 avss.n619 6.4618
R1966 avss.n740 avss.n114 6.4618
R1967 avss.n713 avss.n712 6.4618
R1968 avss.n812 avss.n40 6.4618
R1969 avss.n65 avss.n61 6.4618
R1970 avss.n343 avss.n342 5.47239
R1971 avss.n443 avss.n442 5.47239
R1972 avss.n543 avss.n542 5.47239
R1973 avss.n643 avss.n642 5.47239
R1974 avss.n735 avss.n734 5.47239
R1975 avss.n807 avss.n806 5.47239
R1976 avss.n859 avss.n1 5.18044
R1977 avss.n351 avss.n350 5.03414
R1978 avss.n338 avss.n337 5.03414
R1979 avss.n329 avss.n328 5.03414
R1980 avss.n313 avss.n312 5.03414
R1981 avss.n305 avss.n304 5.03414
R1982 avss.n451 avss.n450 5.03414
R1983 avss.n438 avss.n437 5.03414
R1984 avss.n429 avss.n428 5.03414
R1985 avss.n414 avss.n413 5.03414
R1986 avss.n263 avss.n262 5.03414
R1987 avss.n551 avss.n550 5.03414
R1988 avss.n538 avss.n537 5.03414
R1989 avss.n529 avss.n528 5.03414
R1990 avss.n514 avss.n513 5.03414
R1991 avss.n220 avss.n219 5.03414
R1992 avss.n651 avss.n650 5.03414
R1993 avss.n638 avss.n637 5.03414
R1994 avss.n629 avss.n628 5.03414
R1995 avss.n614 avss.n613 5.03414
R1996 avss.n177 avss.n176 5.03414
R1997 avss.n743 avss.n742 5.03414
R1998 avss.n730 avss.n729 5.03414
R1999 avss.n721 avss.n720 5.03414
R2000 avss.n707 avss.n706 5.03414
R2001 avss.n128 avss.n127 5.03414
R2002 avss.n815 avss.n814 5.03414
R2003 avss.n802 avss.n801 5.03414
R2004 avss.n793 avss.n792 5.03414
R2005 avss.n71 avss.n70 5.03414
R2006 avss.n64 avss.n63 5.03414
R2007 avss.n26 avss.t285 4.84702
R2008 avss.n25 avss.t18 4.84702
R2009 avss.n100 avss.t41 4.84702
R2010 avss.n99 avss.t11 4.84702
R2011 avss.n664 avss.t100 4.84702
R2012 avss.n661 avss.t29 4.84702
R2013 avss.n564 avss.t231 4.84702
R2014 avss.n561 avss.t89 4.84702
R2015 avss.n464 avss.t185 4.84702
R2016 avss.n461 avss.t240 4.84702
R2017 avss.n364 avss.t161 4.84702
R2018 avss.n361 avss.t22 4.84702
R2019 avss.n272 avss.t8 4.7885
R2020 avss.n271 avss.t280 4.7885
R2021 avss.n403 avss.t252 4.7885
R2022 avss.n350 avss.t132 4.7885
R2023 avss.n337 avss.t151 4.7885
R2024 avss.n343 avss.t123 4.7885
R2025 avss.n328 avss.t154 4.7885
R2026 avss.n312 avss.t53 4.7885
R2027 avss.n304 avss.t59 4.7885
R2028 avss.n229 avss.t165 4.7885
R2029 avss.n228 avss.t205 4.7885
R2030 avss.n503 avss.t191 4.7885
R2031 avss.n450 avss.t221 4.7885
R2032 avss.n437 avss.t207 4.7885
R2033 avss.n443 avss.t282 4.7885
R2034 avss.n428 avss.t187 4.7885
R2035 avss.n413 avss.t76 4.7885
R2036 avss.n262 avss.t87 4.7885
R2037 avss.n186 avss.t96 4.7885
R2038 avss.n185 avss.t179 4.7885
R2039 avss.n603 avss.t183 4.7885
R2040 avss.n550 avss.t137 4.7885
R2041 avss.n537 avss.t139 4.7885
R2042 avss.n543 avss.t203 4.7885
R2043 avss.n528 avss.t198 4.7885
R2044 avss.n513 avss.t57 4.7885
R2045 avss.n219 avss.t68 4.7885
R2046 avss.n143 avss.t43 4.7885
R2047 avss.n142 avss.t263 4.7885
R2048 avss.n696 avss.t265 4.7885
R2049 avss.n650 avss.t127 4.7885
R2050 avss.n637 avss.t225 4.7885
R2051 avss.n643 avss.t181 4.7885
R2052 avss.n628 avss.t147 4.7885
R2053 avss.n613 avss.t80 4.7885
R2054 avss.n176 avss.t82 4.7885
R2055 avss.n86 avss.t269 4.7885
R2056 avss.n85 avss.t103 4.7885
R2057 avss.n778 avss.t94 4.7885
R2058 avss.n742 avss.t200 4.7885
R2059 avss.n729 avss.t259 4.7885
R2060 avss.n735 avss.t267 4.7885
R2061 avss.n720 avss.t116 4.7885
R2062 avss.n706 avss.t70 4.7885
R2063 avss.n127 avss.t73 4.7885
R2064 avss.n814 avss.t249 4.7885
R2065 avss.n801 avss.t238 4.7885
R2066 avss.n807 avss.t105 4.7885
R2067 avss.n792 avss.t119 4.7885
R2068 avss.n70 avss.t47 4.7885
R2069 avss.n63 avss.t51 4.7885
R2070 avss.n839 avss.t108 4.7885
R2071 avss.n834 avss.t247 4.7885
R2072 avss.n857 avss.t244 4.7885
R2073 avss.n10 avss.t25 4.7885
R2074 avss.n11 avss.t211 4.7885
R2075 avss.n9 avss.t27 4.7885
R2076 avss.n36 avss.t142 4.7885
R2077 avss.n77 avss.t219 4.7885
R2078 avss.n92 avss.t114 4.7885
R2079 avss.n93 avss.t39 4.7885
R2080 avss.n767 avss.t37 4.7885
R2081 avss.n110 avss.t196 4.7885
R2082 avss.n135 avss.t167 4.7885
R2083 avss.n149 avss.t193 4.7885
R2084 avss.n150 avss.t4 4.7885
R2085 avss.n685 avss.t6 4.7885
R2086 avss.n656 avss.t175 4.7885
R2087 avss.n590 avss.t171 4.7885
R2088 avss.n192 avss.t173 4.7885
R2089 avss.n193 avss.t31 4.7885
R2090 avss.n585 avss.t33 4.7885
R2091 avss.n556 avss.t287 4.7885
R2092 avss.n490 avss.t255 4.7885
R2093 avss.n235 avss.t121 4.7885
R2094 avss.n236 avss.t110 4.7885
R2095 avss.n485 avss.t112 4.7885
R2096 avss.n456 avss.t235 4.7885
R2097 avss.n390 avss.t157 4.7885
R2098 avss.n278 avss.t215 4.7885
R2099 avss.n279 avss.t15 4.7885
R2100 avss.n385 avss.t13 4.7885
R2101 avss.n356 avss.t163 4.7885
R2102 avss.n851 avss.t228 4.7885
R2103 avss.n342 avss.n341 4.28213
R2104 avss.n442 avss.n441 4.28213
R2105 avss.n542 avss.n541 4.28213
R2106 avss.n642 avss.n641 4.28213
R2107 avss.n734 avss.n733 4.28213
R2108 avss.n806 avss.n805 4.28213
R2109 avss.n400 avss.n399 3.51467
R2110 avss.n500 avss.n499 3.51467
R2111 avss.n600 avss.n599 3.51467
R2112 avss.n693 avss.n692 3.51467
R2113 avss.n775 avss.n774 3.51467
R2114 avss.n842 avss.n841 3.51467
R2115 avss.n400 avss.n273 2.06002
R2116 avss.n500 avss.n230 2.06002
R2117 avss.n600 avss.n187 2.06002
R2118 avss.n693 avss.n144 2.06002
R2119 avss.n775 avss.n87 2.06002
R2120 avss.n841 avss.n16 2.06002
R2121 avss.n354 avss.n286 1.92616
R2122 avss.n845 avss.n12 1.90702
R2123 avss.n820 avss.n819 1.90702
R2124 avss.n31 avss.n15 1.90702
R2125 avss.n844 avss.n13 1.90702
R2126 avss.n79 avss.n78 1.90702
R2127 avss.n771 avss.n91 1.90702
R2128 avss.n748 avss.n747 1.90702
R2129 avss.n105 avss.n88 1.90702
R2130 avss.n772 avss.n90 1.90702
R2131 avss.n137 avss.n136 1.90702
R2132 avss.n689 avss.n148 1.90702
R2133 avss.n158 avss.n157 1.90702
R2134 avss.n660 avss.n145 1.90702
R2135 avss.n690 avss.n147 1.90702
R2136 avss.n591 avss.n586 1.90702
R2137 avss.n596 avss.n191 1.90702
R2138 avss.n201 avss.n200 1.90702
R2139 avss.n560 avss.n188 1.90702
R2140 avss.n597 avss.n190 1.90702
R2141 avss.n491 avss.n486 1.90702
R2142 avss.n496 avss.n234 1.90702
R2143 avss.n244 avss.n243 1.90702
R2144 avss.n460 avss.n231 1.90702
R2145 avss.n497 avss.n233 1.90702
R2146 avss.n391 avss.n386 1.90702
R2147 avss.n396 avss.n277 1.90702
R2148 avss.n360 avss.n274 1.90702
R2149 avss.n397 avss.n276 1.90702
R2150 avss.n850 avss.n8 1.90702
R2151 2inmux_0.Bit avss.n859 1.54251
R2152 avss.n310 avss.n309 1.3005
R2153 avss.n312 avss.n311 1.3005
R2154 avss.n311 avss.n298 1.3005
R2155 avss.n324 avss.n297 1.3005
R2156 avss.n328 avss.n327 1.3005
R2157 avss.n327 avss.n326 1.3005
R2158 avss.n304 avss.n303 1.3005
R2159 avss.n303 avss.n302 1.3005
R2160 avss.n320 avss.n319 1.3005
R2161 avss.n411 avss.n410 1.3005
R2162 avss.n413 avss.n412 1.3005
R2163 avss.n412 avss.n257 1.3005
R2164 avss.n424 avss.n256 1.3005
R2165 avss.n428 avss.n427 1.3005
R2166 avss.n427 avss.n426 1.3005
R2167 avss.n262 avss.n261 1.3005
R2168 avss.n261 avss.n260 1.3005
R2169 avss.n421 avss.n420 1.3005
R2170 avss.n511 avss.n510 1.3005
R2171 avss.n513 avss.n512 1.3005
R2172 avss.n512 avss.n214 1.3005
R2173 avss.n524 avss.n213 1.3005
R2174 avss.n528 avss.n527 1.3005
R2175 avss.n527 avss.n526 1.3005
R2176 avss.n219 avss.n218 1.3005
R2177 avss.n218 avss.n217 1.3005
R2178 avss.n521 avss.n520 1.3005
R2179 avss.n611 avss.n610 1.3005
R2180 avss.n613 avss.n612 1.3005
R2181 avss.n612 avss.n171 1.3005
R2182 avss.n624 avss.n170 1.3005
R2183 avss.n628 avss.n627 1.3005
R2184 avss.n627 avss.n626 1.3005
R2185 avss.n176 avss.n175 1.3005
R2186 avss.n175 avss.n174 1.3005
R2187 avss.n621 avss.n620 1.3005
R2188 avss.n704 avss.n703 1.3005
R2189 avss.n706 avss.n705 1.3005
R2190 avss.n705 avss.n123 1.3005
R2191 avss.n717 avss.n122 1.3005
R2192 avss.n720 avss.n719 1.3005
R2193 avss.n719 avss.n718 1.3005
R2194 avss.n127 avss.n126 1.3005
R2195 avss.n126 avss.n125 1.3005
R2196 avss.n714 avss.n713 1.3005
R2197 avss.n74 avss.n73 1.3005
R2198 avss.n70 avss.n57 1.3005
R2199 avss.n57 avss.n56 1.3005
R2200 avss.n54 avss.n48 1.3005
R2201 avss.n792 avss.n791 1.3005
R2202 avss.n791 avss.n790 1.3005
R2203 avss.n63 avss.n62 1.3005
R2204 avss.n62 avss.n49 1.3005
R2205 avss.n61 avss.n60 1.3005
R2206 avss.n828 avss.n11 1.3005
R2207 avss.n828 avss.n827 1.3005
R2208 avss.n826 avss.n12 1.3005
R2209 avss.n19 avss.n10 1.3005
R2210 avss.n833 avss.n19 1.3005
R2211 avss.n831 avss.n9 1.3005
R2212 avss.n832 avss.n831 1.3005
R2213 avss.n821 avss.n820 1.3005
R2214 avss.n36 avss.n34 1.3005
R2215 avss.n34 avss.n33 1.3005
R2216 avss.n32 avss.n31 1.3005
R2217 avss.n30 avss.n25 1.3005
R2218 avss.n30 avss.n29 1.3005
R2219 avss.n27 avss.n26 1.3005
R2220 avss.n28 avss.n27 1.3005
R2221 avss.n22 avss.n13 1.3005
R2222 avss.n77 avss.n76 1.3005
R2223 avss.n76 avss.n75 1.3005
R2224 avss.n80 avss.n79 1.3005
R2225 avss.n749 avss.n748 1.3005
R2226 avss.n110 avss.n108 1.3005
R2227 avss.n108 avss.n107 1.3005
R2228 avss.n106 avss.n105 1.3005
R2229 avss.n104 avss.n99 1.3005
R2230 avss.n104 avss.n103 1.3005
R2231 avss.n101 avss.n100 1.3005
R2232 avss.n102 avss.n101 1.3005
R2233 avss.n96 avss.n90 1.3005
R2234 avss.n135 avss.n134 1.3005
R2235 avss.n134 avss.n133 1.3005
R2236 avss.n138 avss.n137 1.3005
R2237 avss.n157 avss.n156 1.3005
R2238 avss.n657 avss.n656 1.3005
R2239 avss.n658 avss.n657 1.3005
R2240 avss.n660 avss.n659 1.3005
R2241 avss.n662 avss.n661 1.3005
R2242 avss.n663 avss.n662 1.3005
R2243 avss.n665 avss.n664 1.3005
R2244 avss.n666 avss.n665 1.3005
R2245 avss.n667 avss.n147 1.3005
R2246 avss.n590 avss.n589 1.3005
R2247 avss.n589 avss.n588 1.3005
R2248 avss.n587 avss.n586 1.3005
R2249 avss.n200 avss.n199 1.3005
R2250 avss.n557 avss.n556 1.3005
R2251 avss.n558 avss.n557 1.3005
R2252 avss.n560 avss.n559 1.3005
R2253 avss.n562 avss.n561 1.3005
R2254 avss.n563 avss.n562 1.3005
R2255 avss.n565 avss.n564 1.3005
R2256 avss.n566 avss.n565 1.3005
R2257 avss.n567 avss.n190 1.3005
R2258 avss.n490 avss.n489 1.3005
R2259 avss.n489 avss.n488 1.3005
R2260 avss.n487 avss.n486 1.3005
R2261 avss.n243 avss.n242 1.3005
R2262 avss.n457 avss.n456 1.3005
R2263 avss.n458 avss.n457 1.3005
R2264 avss.n460 avss.n459 1.3005
R2265 avss.n462 avss.n461 1.3005
R2266 avss.n463 avss.n462 1.3005
R2267 avss.n465 avss.n464 1.3005
R2268 avss.n466 avss.n465 1.3005
R2269 avss.n467 avss.n233 1.3005
R2270 avss.n390 avss.n389 1.3005
R2271 avss.n389 avss.n388 1.3005
R2272 avss.n387 avss.n386 1.3005
R2273 avss.n286 avss.n285 1.3005
R2274 avss.n357 avss.n356 1.3005
R2275 avss.n358 avss.n357 1.3005
R2276 avss.n360 avss.n359 1.3005
R2277 avss.n362 avss.n361 1.3005
R2278 avss.n363 avss.n362 1.3005
R2279 avss.n365 avss.n364 1.3005
R2280 avss.n366 avss.n365 1.3005
R2281 avss.n367 avss.n276 1.3005
R2282 avss.n347 avss.n290 1.3005
R2283 avss.n350 avss.n349 1.3005
R2284 avss.n349 avss.n348 1.3005
R2285 avss.n299 avss.n292 1.3005
R2286 avss.n344 avss.n343 1.3005
R2287 avss.n345 avss.n344 1.3005
R2288 avss.n334 avss.n333 1.3005
R2289 avss.n337 avss.n336 1.3005
R2290 avss.n336 avss.n335 1.3005
R2291 avss.n372 avss.n277 1.3005
R2292 avss.n370 avss.n278 1.3005
R2293 avss.n371 avss.n370 1.3005
R2294 avss.n282 avss.n279 1.3005
R2295 avss.n382 avss.n282 1.3005
R2296 avss.n385 avss.n384 1.3005
R2297 avss.n384 avss.n383 1.3005
R2298 avss.n375 avss.n273 1.3005
R2299 avss.n378 avss.n272 1.3005
R2300 avss.n379 avss.n378 1.3005
R2301 avss.n380 avss.n271 1.3005
R2302 avss.n381 avss.n380 1.3005
R2303 avss.n404 avss.n403 1.3005
R2304 avss.n405 avss.n404 1.3005
R2305 avss.n447 avss.n248 1.3005
R2306 avss.n450 avss.n449 1.3005
R2307 avss.n449 avss.n448 1.3005
R2308 avss.n407 avss.n251 1.3005
R2309 avss.n444 avss.n443 1.3005
R2310 avss.n445 avss.n444 1.3005
R2311 avss.n434 avss.n433 1.3005
R2312 avss.n437 avss.n436 1.3005
R2313 avss.n436 avss.n435 1.3005
R2314 avss.n472 avss.n234 1.3005
R2315 avss.n470 avss.n235 1.3005
R2316 avss.n471 avss.n470 1.3005
R2317 avss.n239 avss.n236 1.3005
R2318 avss.n482 avss.n239 1.3005
R2319 avss.n485 avss.n484 1.3005
R2320 avss.n484 avss.n483 1.3005
R2321 avss.n475 avss.n230 1.3005
R2322 avss.n478 avss.n229 1.3005
R2323 avss.n479 avss.n478 1.3005
R2324 avss.n480 avss.n228 1.3005
R2325 avss.n481 avss.n480 1.3005
R2326 avss.n504 avss.n503 1.3005
R2327 avss.n505 avss.n504 1.3005
R2328 avss.n547 avss.n205 1.3005
R2329 avss.n550 avss.n549 1.3005
R2330 avss.n549 avss.n548 1.3005
R2331 avss.n507 avss.n208 1.3005
R2332 avss.n544 avss.n543 1.3005
R2333 avss.n545 avss.n544 1.3005
R2334 avss.n534 avss.n533 1.3005
R2335 avss.n537 avss.n536 1.3005
R2336 avss.n536 avss.n535 1.3005
R2337 avss.n572 avss.n191 1.3005
R2338 avss.n570 avss.n192 1.3005
R2339 avss.n571 avss.n570 1.3005
R2340 avss.n196 avss.n193 1.3005
R2341 avss.n582 avss.n196 1.3005
R2342 avss.n585 avss.n584 1.3005
R2343 avss.n584 avss.n583 1.3005
R2344 avss.n575 avss.n187 1.3005
R2345 avss.n578 avss.n186 1.3005
R2346 avss.n579 avss.n578 1.3005
R2347 avss.n580 avss.n185 1.3005
R2348 avss.n581 avss.n580 1.3005
R2349 avss.n604 avss.n603 1.3005
R2350 avss.n605 avss.n604 1.3005
R2351 avss.n647 avss.n162 1.3005
R2352 avss.n650 avss.n649 1.3005
R2353 avss.n649 avss.n648 1.3005
R2354 avss.n607 avss.n165 1.3005
R2355 avss.n644 avss.n643 1.3005
R2356 avss.n645 avss.n644 1.3005
R2357 avss.n634 avss.n633 1.3005
R2358 avss.n637 avss.n636 1.3005
R2359 avss.n636 avss.n635 1.3005
R2360 avss.n672 avss.n148 1.3005
R2361 avss.n670 avss.n149 1.3005
R2362 avss.n671 avss.n670 1.3005
R2363 avss.n153 avss.n150 1.3005
R2364 avss.n682 avss.n153 1.3005
R2365 avss.n685 avss.n684 1.3005
R2366 avss.n684 avss.n683 1.3005
R2367 avss.n675 avss.n144 1.3005
R2368 avss.n678 avss.n143 1.3005
R2369 avss.n679 avss.n678 1.3005
R2370 avss.n680 avss.n142 1.3005
R2371 avss.n681 avss.n680 1.3005
R2372 avss.n697 avss.n696 1.3005
R2373 avss.n698 avss.n697 1.3005
R2374 avss.n740 avss.n739 1.3005
R2375 avss.n742 avss.n741 1.3005
R2376 avss.n741 avss.n98 1.3005
R2377 avss.n700 avss.n117 1.3005
R2378 avss.n736 avss.n735 1.3005
R2379 avss.n737 avss.n736 1.3005
R2380 avss.n726 avss.n725 1.3005
R2381 avss.n729 avss.n728 1.3005
R2382 avss.n728 avss.n727 1.3005
R2383 avss.n758 avss.n91 1.3005
R2384 avss.n761 avss.n92 1.3005
R2385 avss.n762 avss.n761 1.3005
R2386 avss.n763 avss.n93 1.3005
R2387 avss.n764 avss.n763 1.3005
R2388 avss.n767 avss.n766 1.3005
R2389 avss.n766 avss.n765 1.3005
R2390 avss.n755 avss.n87 1.3005
R2391 avss.n753 avss.n86 1.3005
R2392 avss.n754 avss.n753 1.3005
R2393 avss.n85 avss.n84 1.3005
R2394 avss.n84 avss.n53 1.3005
R2395 avss.n779 avss.n778 1.3005
R2396 avss.n780 avss.n779 1.3005
R2397 avss.n812 avss.n811 1.3005
R2398 avss.n814 avss.n813 1.3005
R2399 avss.n813 avss.n24 1.3005
R2400 avss.n782 avss.n43 1.3005
R2401 avss.n808 avss.n807 1.3005
R2402 avss.n809 avss.n808 1.3005
R2403 avss.n798 avss.n797 1.3005
R2404 avss.n801 avss.n800 1.3005
R2405 avss.n800 avss.n799 1.3005
R2406 avss.n823 avss.n16 1.3005
R2407 avss.n839 avss.n838 1.3005
R2408 avss.n838 avss.n837 1.3005
R2409 avss.n835 avss.n834 1.3005
R2410 avss.n836 avss.n835 1.3005
R2411 avss.n857 avss.n856 1.3005
R2412 avss.n856 avss.n855 1.3005
R2413 avss.n852 avss.n851 1.3005
R2414 avss.n853 avss.n852 1.3005
R2415 avss.n8 avss.n7 1.3005
R2416 avss.n819 avss.n35 0.990409
R2417 avss.n747 avss.n109 0.990409
R2418 avss.n592 avss.n158 0.990409
R2419 avss.n492 avss.n201 0.990409
R2420 avss.n392 avss.n244 0.990409
R2421 avss.n351 avss.n289 0.92075
R2422 avss.n339 avss.n338 0.92075
R2423 avss.n329 avss.n296 0.92075
R2424 avss.n313 avss.n308 0.92075
R2425 avss.n318 avss.n305 0.92075
R2426 avss.n451 avss.n247 0.92075
R2427 avss.n439 avss.n438 0.92075
R2428 avss.n429 avss.n255 0.92075
R2429 avss.n414 avss.n266 0.92075
R2430 avss.n419 avss.n263 0.92075
R2431 avss.n551 avss.n204 0.92075
R2432 avss.n539 avss.n538 0.92075
R2433 avss.n529 avss.n212 0.92075
R2434 avss.n514 avss.n223 0.92075
R2435 avss.n519 avss.n220 0.92075
R2436 avss.n651 avss.n161 0.92075
R2437 avss.n639 avss.n638 0.92075
R2438 avss.n629 avss.n169 0.92075
R2439 avss.n614 avss.n180 0.92075
R2440 avss.n619 avss.n177 0.92075
R2441 avss.n743 avss.n114 0.92075
R2442 avss.n731 avss.n730 0.92075
R2443 avss.n721 avss.n121 0.92075
R2444 avss.n707 avss.n131 0.92075
R2445 avss.n712 avss.n128 0.92075
R2446 avss.n815 avss.n40 0.92075
R2447 avss.n803 avss.n802 0.92075
R2448 avss.n793 avss.n47 0.92075
R2449 avss.n72 avss.n71 0.92075
R2450 avss.n65 avss.n64 0.92075
R2451 avss.n403 avss.n402 0.771017
R2452 avss.n503 avss.n502 0.771017
R2453 avss.n603 avss.n602 0.771017
R2454 avss.n696 avss.n695 0.771017
R2455 avss.n778 avss.n777 0.771017
R2456 avss.n354 avss.n353 0.709028
R2457 avss.n454 avss.n453 0.709028
R2458 avss.n554 avss.n553 0.709028
R2459 avss.n654 avss.n653 0.709028
R2460 avss.n746 avss.n745 0.709028
R2461 avss.n818 avss.n817 0.709028
R2462 avss.n858 avss.n857 0.471317
R2463 avss.n401 avss.n272 0.463217
R2464 avss.n402 avss.n271 0.463217
R2465 avss.n501 avss.n229 0.463217
R2466 avss.n502 avss.n228 0.463217
R2467 avss.n601 avss.n186 0.463217
R2468 avss.n602 avss.n185 0.463217
R2469 avss.n694 avss.n143 0.463217
R2470 avss.n695 avss.n142 0.463217
R2471 avss.n776 avss.n86 0.463217
R2472 avss.n777 avss.n85 0.463217
R2473 avss.n840 avss.n839 0.463217
R2474 avss.n834 avss.n2 0.463217
R2475 avss.n847 avss.n10 0.463217
R2476 avss.n846 avss.n11 0.463217
R2477 avss.n848 avss.n9 0.463217
R2478 avss.n37 avss.n36 0.463217
R2479 avss.n78 avss.n77 0.463217
R2480 avss.n770 avss.n92 0.463217
R2481 avss.n769 avss.n93 0.463217
R2482 avss.n768 avss.n767 0.463217
R2483 avss.n111 avss.n110 0.463217
R2484 avss.n136 avss.n135 0.463217
R2485 avss.n688 avss.n149 0.463217
R2486 avss.n687 avss.n150 0.463217
R2487 avss.n686 avss.n685 0.463217
R2488 avss.n656 avss.n655 0.463217
R2489 avss.n591 avss.n590 0.463217
R2490 avss.n595 avss.n192 0.463217
R2491 avss.n594 avss.n193 0.463217
R2492 avss.n593 avss.n585 0.463217
R2493 avss.n556 avss.n555 0.463217
R2494 avss.n491 avss.n490 0.463217
R2495 avss.n495 avss.n235 0.463217
R2496 avss.n494 avss.n236 0.463217
R2497 avss.n493 avss.n485 0.463217
R2498 avss.n456 avss.n455 0.463217
R2499 avss.n391 avss.n390 0.463217
R2500 avss.n395 avss.n278 0.463217
R2501 avss.n394 avss.n279 0.463217
R2502 avss.n393 avss.n385 0.463217
R2503 avss.n356 avss.n355 0.463217
R2504 avss.n851 avss.n850 0.463217
R2505 avss.n402 avss.n401 0.3083
R2506 avss.n502 avss.n501 0.3083
R2507 avss.n602 avss.n601 0.3083
R2508 avss.n695 avss.n694 0.3083
R2509 avss.n777 avss.n776 0.3083
R2510 avss.n840 avss.n2 0.3083
R2511 avss.n847 avss.n846 0.3083
R2512 avss.n848 avss.n847 0.3083
R2513 avss.n770 avss.n769 0.3083
R2514 avss.n769 avss.n768 0.3083
R2515 avss.n688 avss.n687 0.3083
R2516 avss.n687 avss.n686 0.3083
R2517 avss.n595 avss.n594 0.3083
R2518 avss.n594 avss.n593 0.3083
R2519 avss.n495 avss.n494 0.3083
R2520 avss.n494 avss.n493 0.3083
R2521 avss.n395 avss.n394 0.3083
R2522 avss.n394 avss.n393 0.3083
R2523 avss.n858 avss.n2 0.3002
R2524 avss.n1 avss.n0 0.252687
R2525 avss.n846 avss.n845 0.2165
R2526 avss.n771 avss.n770 0.2165
R2527 avss.n689 avss.n688 0.2165
R2528 avss.n596 avss.n595 0.2165
R2529 avss.n496 avss.n495 0.2165
R2530 avss.n396 avss.n395 0.2165
R2531 avss.n768 avss.n35 0.1748
R2532 avss.n593 avss.n592 0.1748
R2533 avss.n493 avss.n492 0.1748
R2534 avss.n393 avss.n392 0.1748
R2535 avss.n686 avss.n109 0.17465
R2536 avss.n849 avss.n848 0.1598
R2537 avss.n850 avss.n849 0.152487
R2538 avss.n845 avss.n844 0.148459
R2539 avss.n772 avss.n771 0.148459
R2540 avss.n690 avss.n689 0.148459
R2541 avss.n597 avss.n596 0.148459
R2542 avss.n497 avss.n496 0.148459
R2543 avss.n397 avss.n396 0.148459
R2544 avss.n136 avss.n109 0.13865
R2545 avss.n78 avss.n35 0.1385
R2546 avss.n592 avss.n591 0.1385
R2547 avss.n492 avss.n491 0.1385
R2548 avss.n392 avss.n391 0.1385
R2549 avss.n316 avss.n306 0.122607
R2550 avss.n417 avss.n264 0.122607
R2551 avss.n517 avss.n221 0.122607
R2552 avss.n617 avss.n178 0.122607
R2553 avss.n710 avss.n129 0.122607
R2554 avss.n67 avss.n59 0.122607
R2555 avss.n332 avss.n331 0.10457
R2556 avss.n432 avss.n431 0.10457
R2557 avss.n532 avss.n531 0.10457
R2558 avss.n632 avss.n631 0.10457
R2559 avss.n724 avss.n723 0.10457
R2560 avss.n796 avss.n795 0.10457
R2561 avss.n843 avss.n14 0.073981
R2562 avss.n773 avss.n89 0.073981
R2563 avss.n691 avss.n146 0.073981
R2564 avss.n598 avss.n189 0.073981
R2565 avss.n498 avss.n232 0.073981
R2566 avss.n398 avss.n275 0.073981
R2567 avss.n340 avss.n287 0.0679983
R2568 avss.n440 avss.n245 0.0679983
R2569 avss.n540 avss.n202 0.0679983
R2570 avss.n640 avss.n159 0.0679983
R2571 avss.n732 avss.n112 0.0679983
R2572 avss.n804 avss.n38 0.0679983
R2573 avss.n401 avss.n400 0.0635
R2574 avss.n501 avss.n500 0.0635
R2575 avss.n601 avss.n600 0.0635
R2576 avss.n694 avss.n693 0.0635
R2577 avss.n776 avss.n775 0.0635
R2578 avss.n841 avss.n840 0.0635
R2579 avss.n306 avss.n293 0.0622481
R2580 avss.n264 avss.n252 0.0622481
R2581 avss.n221 avss.n209 0.0622481
R2582 avss.n178 avss.n166 0.0622481
R2583 avss.n129 avss.n118 0.0622481
R2584 avss.n59 avss.n44 0.0622481
R2585 avss.n352 avss.n288 0.0568904
R2586 avss.n452 avss.n246 0.0568904
R2587 avss.n552 avss.n203 0.0568904
R2588 avss.n652 avss.n160 0.0568904
R2589 avss.n744 avss.n113 0.0568904
R2590 avss.n816 avss.n39 0.0568904
R2591 avss.n332 avss.n288 0.054837
R2592 avss.n432 avss.n246 0.054837
R2593 avss.n532 avss.n203 0.054837
R2594 avss.n632 avss.n160 0.054837
R2595 avss.n724 avss.n113 0.054837
R2596 avss.n796 avss.n39 0.054837
R2597 avss.n331 avss.n294 0.0466843
R2598 avss.n431 avss.n253 0.0466843
R2599 avss.n531 avss.n210 0.0466843
R2600 avss.n631 avss.n167 0.0466843
R2601 avss.n723 avss.n119 0.0466843
R2602 avss.n795 avss.n45 0.0466843
R2603 avss.n332 avss.n293 0.0415307
R2604 avss.n432 avss.n252 0.0415307
R2605 avss.n532 avss.n209 0.0415307
R2606 avss.n632 avss.n166 0.0415307
R2607 avss.n724 avss.n118 0.0415307
R2608 avss.n796 avss.n44 0.0415307
R2609 avss.n317 avss.n294 0.0405109
R2610 avss.n314 avss.n307 0.0405109
R2611 avss.n330 avss.n295 0.0405109
R2612 avss.n418 avss.n253 0.0405109
R2613 avss.n415 avss.n265 0.0405109
R2614 avss.n430 avss.n254 0.0405109
R2615 avss.n518 avss.n210 0.0405109
R2616 avss.n515 avss.n222 0.0405109
R2617 avss.n530 avss.n211 0.0405109
R2618 avss.n618 avss.n167 0.0405109
R2619 avss.n615 avss.n179 0.0405109
R2620 avss.n630 avss.n168 0.0405109
R2621 avss.n711 avss.n119 0.0405109
R2622 avss.n708 avss.n130 0.0405109
R2623 avss.n722 avss.n120 0.0405109
R2624 avss.n66 avss.n45 0.0405109
R2625 avss.n69 avss.n58 0.0405109
R2626 avss.n794 avss.n46 0.0405109
R2627 avss.n844 avss.n843 0.0389018
R2628 avss.n773 avss.n772 0.0389018
R2629 avss.n691 avss.n690 0.0389018
R2630 avss.n598 avss.n597 0.0389018
R2631 avss.n498 avss.n497 0.0389018
R2632 avss.n398 avss.n397 0.0389018
R2633 avss.n353 avss.n287 0.035635
R2634 avss.n453 avss.n245 0.035635
R2635 avss.n553 avss.n202 0.035635
R2636 avss.n653 avss.n159 0.035635
R2637 avss.n745 avss.n112 0.035635
R2638 avss.n817 avss.n38 0.035635
R2639 avss.n341 avss.n332 0.0349747
R2640 avss.n441 avss.n432 0.0349747
R2641 avss.n541 avss.n532 0.0349747
R2642 avss.n641 avss.n632 0.0349747
R2643 avss.n733 avss.n724 0.0349747
R2644 avss.n805 avss.n796 0.0349747
R2645 avss.n316 avss.n315 0.0322085
R2646 avss.n315 avss.n293 0.0322085
R2647 avss.n417 avss.n416 0.0322085
R2648 avss.n416 avss.n252 0.0322085
R2649 avss.n517 avss.n516 0.0322085
R2650 avss.n516 avss.n209 0.0322085
R2651 avss.n617 avss.n616 0.0322085
R2652 avss.n616 avss.n166 0.0322085
R2653 avss.n710 avss.n709 0.0322085
R2654 avss.n709 avss.n118 0.0322085
R2655 avss.n68 avss.n67 0.0322085
R2656 avss.n68 avss.n44 0.0322085
R2657 avss.n25 avss.n14 0.0258591
R2658 avss.n26 avss.n14 0.0258591
R2659 avss.n99 avss.n89 0.0258591
R2660 avss.n100 avss.n89 0.0258591
R2661 avss.n661 avss.n146 0.0258591
R2662 avss.n664 avss.n146 0.0258591
R2663 avss.n561 avss.n189 0.0258591
R2664 avss.n564 avss.n189 0.0258591
R2665 avss.n461 avss.n232 0.0258591
R2666 avss.n464 avss.n232 0.0258591
R2667 avss.n361 avss.n275 0.0258591
R2668 avss.n364 avss.n275 0.0258591
R2669 avss.n843 avss.n842 0.023066
R2670 avss.n774 avss.n773 0.023066
R2671 avss.n692 avss.n691 0.023066
R2672 avss.n599 avss.n598 0.023066
R2673 avss.n499 avss.n498 0.023066
R2674 avss.n399 avss.n398 0.023066
R2675 avss.n317 avss.n316 0.0214837
R2676 avss.n315 avss.n295 0.0214837
R2677 avss.n418 avss.n417 0.0214837
R2678 avss.n416 avss.n254 0.0214837
R2679 avss.n518 avss.n517 0.0214837
R2680 avss.n516 avss.n211 0.0214837
R2681 avss.n618 avss.n617 0.0214837
R2682 avss.n616 avss.n168 0.0214837
R2683 avss.n711 avss.n710 0.0214837
R2684 avss.n709 avss.n120 0.0214837
R2685 avss.n67 avss.n66 0.0214837
R2686 avss.n68 avss.n46 0.0214837
R2687 avss.n819 avss.n818 0.0196349
R2688 avss.n747 avss.n746 0.0196349
R2689 avss.n654 avss.n158 0.0196349
R2690 avss.n554 avss.n201 0.0196349
R2691 avss.n454 avss.n244 0.0196349
R2692 avss.n842 avss.n15 0.0163358
R2693 avss.n774 avss.n88 0.0163358
R2694 avss.n692 avss.n145 0.0163358
R2695 avss.n599 avss.n188 0.0163358
R2696 avss.n499 avss.n231 0.0163358
R2697 avss.n399 avss.n274 0.0163358
R2698 avss.n37 avss.n15 0.0139604
R2699 avss.n111 avss.n88 0.0139604
R2700 avss.n655 avss.n145 0.0139604
R2701 avss.n555 avss.n188 0.0139604
R2702 avss.n455 avss.n231 0.0139604
R2703 avss.n355 avss.n274 0.0139604
R2704 avss.n818 avss.n37 0.0130367
R2705 avss.n746 avss.n111 0.0130367
R2706 avss.n655 avss.n654 0.0130367
R2707 avss.n555 avss.n554 0.0130367
R2708 avss.n455 avss.n454 0.0130367
R2709 avss.n355 avss.n354 0.0130367
R2710 avss.n315 avss.n314 0.0121902
R2711 avss.n416 avss.n415 0.0121902
R2712 avss.n516 avss.n515 0.0121902
R2713 avss.n616 avss.n615 0.0121902
R2714 avss.n709 avss.n708 0.0121902
R2715 avss.n69 avss.n68 0.0121902
R2716 avss.n849 avss 0.0118245
R2717 avss.n307 avss.n306 0.00915761
R2718 avss.n265 avss.n264 0.00915761
R2719 avss.n222 avss.n221 0.00915761
R2720 avss.n179 avss.n178 0.00915761
R2721 avss.n130 avss.n129 0.00915761
R2722 avss.n59 avss.n58 0.00915761
R2723 avss.n331 avss.n330 0.00720109
R2724 avss.n431 avss.n430 0.00720109
R2725 avss.n531 avss.n530 0.00720109
R2726 avss.n631 avss.n630 0.00720109
R2727 avss.n723 avss.n722 0.00720109
R2728 avss.n795 avss.n794 0.00720109
R2729 avss.n353 avss.n352 0.00511663
R2730 avss.n453 avss.n452 0.00511663
R2731 avss.n553 avss.n552 0.00511663
R2732 avss.n653 avss.n652 0.00511663
R2733 avss.n745 avss.n744 0.00511663
R2734 avss.n817 avss.n816 0.00511663
R2735 avss.n341 avss.n340 0.000544599
R2736 avss.n441 avss.n440 0.000544599
R2737 avss.n541 avss.n540 0.000544599
R2738 avss.n641 avss.n640 0.000544599
R2739 avss.n733 avss.n732 0.000544599
R2740 avss.n805 avss.n804 0.000544599
R2741 a_48650_3501.n0 a_48650_3501.t4 34.1797
R2742 a_48650_3501.n0 a_48650_3501.t5 19.5798
R2743 a_48650_3501.t0 a_48650_3501.n3 18.7717
R2744 a_48650_3501.n3 a_48650_3501.t2 9.2885
R2745 a_48650_3501.n2 a_48650_3501.n0 4.93379
R2746 a_48650_3501.n1 a_48650_3501.t1 4.23346
R2747 a_48650_3501.n1 a_48650_3501.t3 3.85546
R2748 a_48650_3501.n3 a_48650_3501.n2 0.4055
R2749 a_48650_3501.n2 a_48650_3501.n1 0.352625
R2750 a_6520_1558.n2 a_6520_1558.t5 40.8177
R2751 a_6520_1558.n3 a_6520_1558.t4 40.6313
R2752 a_6520_1558.n3 a_6520_1558.t6 27.3166
R2753 a_6520_1558.n2 a_6520_1558.t7 27.1302
R2754 a_6520_1558.n4 a_6520_1558.n3 19.2576
R2755 a_6520_1558.t0 a_6520_1558.n5 10.0473
R2756 a_6520_1558.n1 a_6520_1558.t1 6.51042
R2757 a_6520_1558.n1 a_6520_1558.n0 6.04952
R2758 a_6520_1558.n4 a_6520_1558.n2 5.91752
R2759 a_6520_1558.n5 a_6520_1558.n4 4.89565
R2760 a_6520_1558.n5 a_6520_1558.n1 0.732092
R2761 a_6520_1558.n0 a_6520_1558.t3 0.7285
R2762 a_6520_1558.n0 a_6520_1558.t2 0.7285
R2763 a_6600_2510.n0 a_6600_2510.t4 41.0041
R2764 a_6600_2510.n1 a_6600_2510.t5 40.8177
R2765 a_6600_2510.n1 a_6600_2510.t7 27.1302
R2766 a_6600_2510.n0 a_6600_2510.t6 26.9438
R2767 a_6600_2510.n2 a_6600_2510.n1 22.5284
R2768 a_6600_2510.n3 a_6600_2510.n2 19.5781
R2769 a_6600_2510.n3 a_6600_2510.t1 10.0473
R2770 a_6600_2510.n4 a_6600_2510.t3 6.51042
R2771 a_6600_2510.n5 a_6600_2510.n4 6.04952
R2772 a_6600_2510.n2 a_6600_2510.n0 5.7305
R2773 a_6600_2510.n4 a_6600_2510.n3 0.732092
R2774 a_6600_2510.t0 a_6600_2510.n5 0.7285
R2775 a_6600_2510.n5 a_6600_2510.t2 0.7285
R2776 a_6520_3763.n1 a_6520_3763.t9 41.0041
R2777 a_6520_3763.n0 a_6520_3763.t5 40.8177
R2778 a_6520_3763.n2 a_6520_3763.t4 40.6313
R2779 a_6520_3763.n2 a_6520_3763.t7 27.3166
R2780 a_6520_3763.n0 a_6520_3763.t8 27.1302
R2781 a_6520_3763.n1 a_6520_3763.t6 26.9438
R2782 a_6520_3763.n3 a_6520_3763.n1 15.6312
R2783 a_6520_3763.n3 a_6520_3763.n2 15.046
R2784 a_6520_3763.n5 a_6520_3763.t3 10.0473
R2785 a_6520_3763.n6 a_6520_3763.t1 6.51042
R2786 a_6520_3763.n7 a_6520_3763.n6 6.04952
R2787 a_6520_3763.n4 a_6520_3763.n0 5.64619
R2788 a_6520_3763.n5 a_6520_3763.n4 5.17851
R2789 a_6520_3763.n4 a_6520_3763.n3 4.5005
R2790 a_6520_3763.n6 a_6520_3763.n5 0.732092
R2791 a_6520_3763.t0 a_6520_3763.n7 0.7285
R2792 a_6520_3763.n7 a_6520_3763.t2 0.7285
R2793 dffrs_1.Q.n3 dffrs_1.Q.t7 40.6313
R2794 dffrs_1.Q.n1 dffrs_1.Q.t4 34.1066
R2795 dffrs_1.Q.n3 dffrs_1.Q.t5 27.3166
R2796 dffrs_1.Q.n0 dffrs_1.Q.t6 19.673
R2797 dffrs_1.Q.n0 dffrs_1.Q.t8 19.4007
R2798 dffrs_1.Q.n7 dffrs_1.Q.n3 14.6967
R2799 dffrs_1.Q.n6 dffrs_1.Q.t3 10.0473
R2800 dffrs_1.Q.n7 dffrs_1.Q.n6 9.39565
R2801 dffrs_1.Q.n2 dffrs_1.Q.n1 6.70486
R2802 dffrs_1.Q.n5 dffrs_1.Q.t2 6.51042
R2803 dffrs_1.Q.n5 dffrs_1.Q.n4 6.04952
R2804 dffrs_1.Q dffrs_1.Q.n2 5.81354
R2805 dffrs_1.Q.n6 dffrs_1.Q.n5 0.732092
R2806 dffrs_1.Q.n4 dffrs_1.Q.t1 0.7285
R2807 dffrs_1.Q.n4 dffrs_1.Q.t0 0.7285
R2808 dffrs_1.Q dffrs_1.Q.n7 0.458082
R2809 dffrs_1.Q.n1 dffrs_1.Q.n0 0.252687
R2810 dffrs_1.Q.n2 2inmux_3.Bit 0.0519286
R2811 a_20234_3501.n0 a_20234_3501.t5 34.1797
R2812 a_20234_3501.n0 a_20234_3501.t4 19.5798
R2813 a_20234_3501.n3 a_20234_3501.t1 18.7717
R2814 a_20234_3501.t0 a_20234_3501.n3 9.2885
R2815 a_20234_3501.n2 a_20234_3501.n0 4.93379
R2816 a_20234_3501.n1 a_20234_3501.t2 4.23346
R2817 a_20234_3501.n1 a_20234_3501.t3 3.85546
R2818 a_20234_3501.n3 a_20234_3501.n2 0.4055
R2819 a_20234_3501.n2 a_20234_3501.n1 0.352625
R2820 2inmux_2.Bit.n3 2inmux_2.Bit.t6 40.6313
R2821 2inmux_2.Bit.n1 2inmux_2.Bit.t5 34.1066
R2822 2inmux_2.Bit.n3 2inmux_2.Bit.t8 27.3166
R2823 2inmux_2.Bit.n0 2inmux_2.Bit.t7 19.673
R2824 2inmux_2.Bit.n0 2inmux_2.Bit.t4 19.4007
R2825 2inmux_2.Bit.n7 2inmux_2.Bit.n3 14.6967
R2826 2inmux_2.Bit.n6 2inmux_2.Bit.t2 10.0473
R2827 2inmux_2.Bit.n7 2inmux_2.Bit.n6 9.39565
R2828 2inmux_2.Bit.n2 2inmux_2.Bit.n1 6.70486
R2829 2inmux_2.Bit.n5 2inmux_2.Bit.t1 6.51042
R2830 2inmux_2.Bit.n5 2inmux_2.Bit.n4 6.04952
R2831 dffrs_0.Q 2inmux_2.Bit.n2 5.81514
R2832 2inmux_2.Bit.n6 2inmux_2.Bit.n5 0.732092
R2833 2inmux_2.Bit.n4 2inmux_2.Bit.t3 0.7285
R2834 2inmux_2.Bit.n4 2inmux_2.Bit.t0 0.7285
R2835 dffrs_0.Q 2inmux_2.Bit.n7 0.458082
R2836 2inmux_2.Bit.n1 2inmux_2.Bit.n0 0.252687
R2837 2inmux_2.Bit.n2 2inmux_2.Bit 0.0519286
R2838 a_1290_3500.n0 a_1290_3500.t4 34.1797
R2839 a_1290_3500.n0 a_1290_3500.t5 19.5798
R2840 a_1290_3500.n3 a_1290_3500.t3 18.7717
R2841 a_1290_3500.t0 a_1290_3500.n3 9.2885
R2842 a_1290_3500.n2 a_1290_3500.n0 4.93379
R2843 a_1290_3500.n1 a_1290_3500.t1 4.23346
R2844 a_1290_3500.n1 a_1290_3500.t2 3.85546
R2845 a_1290_3500.n3 a_1290_3500.n2 0.4055
R2846 a_1290_3500.n2 a_1290_3500.n1 0.352625
R2847 clk.n3 clk.t18 41.0041
R2848 clk.n7 clk.t12 41.0041
R2849 clk.n11 clk.t1 41.0041
R2850 clk.n15 clk.t15 41.0041
R2851 clk.n19 clk.t3 41.0041
R2852 clk.n0 clk.t17 41.0041
R2853 clk.n4 clk.t2 40.8177
R2854 clk.n8 clk.t22 40.8177
R2855 clk.n12 clk.t11 40.8177
R2856 clk.n16 clk.t8 40.8177
R2857 clk.n20 clk.t20 40.8177
R2858 clk.n1 clk.t10 40.8177
R2859 clk.n4 clk.t13 27.1302
R2860 clk.n8 clk.t9 27.1302
R2861 clk.n12 clk.t23 27.1302
R2862 clk.n16 clk.t19 27.1302
R2863 clk.n20 clk.t5 27.1302
R2864 clk.n1 clk.t21 27.1302
R2865 clk.n3 clk.t7 26.9438
R2866 clk.n7 clk.t0 26.9438
R2867 clk.n11 clk.t14 26.9438
R2868 clk.n15 clk.t4 26.9438
R2869 clk.n19 clk.t16 26.9438
R2870 clk.n0 clk.t6 26.9438
R2871 dffrs_5.clk clk.n22 23.2034
R2872 clk.n10 clk.n6 13.9468
R2873 clk.n14 clk.n10 13.9463
R2874 clk.n22 clk.n18 13.9457
R2875 clk.n18 clk.n14 13.9457
R2876 clk.n6 dffrs_0.clk 9.25764
R2877 clk.n10 dffrs_1.clk 9.25764
R2878 clk.n14 dffrs_2.clk 9.25764
R2879 clk.n18 dffrs_3.clk 9.25764
R2880 clk.n22 dffrs_4.clk 9.25764
R2881 clk.n5 clk.n4 7.65746
R2882 clk.n9 clk.n8 7.65746
R2883 clk.n13 clk.n12 7.65746
R2884 clk.n17 clk.n16 7.65746
R2885 clk.n21 clk.n20 7.65746
R2886 clk.n2 clk.n1 7.65746
R2887 clk.n5 clk.n3 7.12229
R2888 clk.n9 clk.n7 7.12229
R2889 clk.n13 clk.n11 7.12229
R2890 clk.n17 clk.n15 7.12229
R2891 clk.n21 clk.n19 7.12229
R2892 clk.n2 clk.n0 7.12229
R2893 clk.n6 clk 3.54742
R2894 dffrs_0.clk clk.n5 0.611214
R2895 dffrs_1.clk clk.n9 0.611214
R2896 dffrs_2.clk clk.n13 0.611214
R2897 dffrs_3.clk clk.n17 0.611214
R2898 dffrs_4.clk clk.n21 0.611214
R2899 dffrs_5.clk clk.n2 0.611214
R2900 a_15992_3763.n1 a_15992_3763.t7 41.0041
R2901 a_15992_3763.n0 a_15992_3763.t5 40.8177
R2902 a_15992_3763.n2 a_15992_3763.t6 40.6313
R2903 a_15992_3763.n2 a_15992_3763.t9 27.3166
R2904 a_15992_3763.n0 a_15992_3763.t8 27.1302
R2905 a_15992_3763.n1 a_15992_3763.t4 26.9438
R2906 a_15992_3763.n3 a_15992_3763.n1 15.6312
R2907 a_15992_3763.n3 a_15992_3763.n2 15.046
R2908 a_15992_3763.n5 a_15992_3763.t3 10.0473
R2909 a_15992_3763.n6 a_15992_3763.t2 6.51042
R2910 a_15992_3763.n7 a_15992_3763.n6 6.04952
R2911 a_15992_3763.n4 a_15992_3763.n0 5.64619
R2912 a_15992_3763.n5 a_15992_3763.n4 5.17851
R2913 a_15992_3763.n4 a_15992_3763.n3 4.5005
R2914 a_15992_3763.n6 a_15992_3763.n5 0.732092
R2915 a_15992_3763.t0 a_15992_3763.n7 0.7285
R2916 a_15992_3763.n7 a_15992_3763.t1 0.7285
R2917 2inmux_1.Bit.n3 2inmux_1.Bit.t8 40.6313
R2918 2inmux_1.Bit.n1 2inmux_1.Bit.t7 34.1066
R2919 2inmux_1.Bit.n3 2inmux_1.Bit.t5 27.3166
R2920 2inmux_1.Bit.n0 2inmux_1.Bit.t4 19.673
R2921 2inmux_1.Bit.n0 2inmux_1.Bit.t6 19.4007
R2922 2inmux_1.Bit.n7 2inmux_1.Bit.n3 14.6967
R2923 2inmux_1.Bit.n6 2inmux_1.Bit.t1 10.0473
R2924 2inmux_1.Bit.n7 2inmux_1.Bit.n6 9.39565
R2925 2inmux_1.Bit.n2 2inmux_1.Bit.n1 6.70486
R2926 2inmux_1.Bit.n5 2inmux_1.Bit.t0 6.51042
R2927 2inmux_1.Bit.n5 2inmux_1.Bit.n4 6.04952
R2928 dffrs_4.Q 2inmux_1.Bit.n2 5.81514
R2929 2inmux_1.Bit.n6 2inmux_1.Bit.n5 0.732092
R2930 2inmux_1.Bit.n4 2inmux_1.Bit.t3 0.7285
R2931 2inmux_1.Bit.n4 2inmux_1.Bit.t2 0.7285
R2932 dffrs_4.Q 2inmux_1.Bit.n7 0.458082
R2933 2inmux_1.Bit.n1 2inmux_1.Bit.n0 0.252687
R2934 2inmux_1.Bit.n2 2inmux_1.Bit 0.0519286
R2935 a_15992_5968.n0 a_15992_5968.t5 40.6313
R2936 a_15992_5968.n0 a_15992_5968.t4 27.3166
R2937 a_15992_5968.n1 a_15992_5968.n0 24.1527
R2938 a_15992_5968.n1 a_15992_5968.t1 10.0473
R2939 a_15992_5968.t0 a_15992_5968.n3 6.51042
R2940 a_15992_5968.n3 a_15992_5968.n2 6.04952
R2941 a_15992_5968.n3 a_15992_5968.n1 0.732092
R2942 a_15992_5968.n2 a_15992_5968.t3 0.7285
R2943 a_15992_5968.n2 a_15992_5968.t2 0.7285
R2944 load.n4 load.t17 34.2529
R2945 load.n10 load.t23 34.2529
R2946 load.n16 load.t28 34.2529
R2947 load.n22 load.t13 34.2529
R2948 load.n28 load.t0 34.2529
R2949 load.n1 load.t9 34.2529
R2950 load.n6 load.t20 34.1797
R2951 load.n12 load.t19 34.1797
R2952 load.n18 load.t14 34.1797
R2953 load.n24 load.t1 34.1797
R2954 load.n30 load.t26 34.1797
R2955 load.n2 load.t3 34.1797
R2956 load.n3 load.t2 19.673
R2957 load.n9 load.t5 19.673
R2958 load.n15 load.t4 19.673
R2959 load.n21 load.t18 19.673
R2960 load.n27 load.t7 19.673
R2961 load.n0 load.t25 19.673
R2962 load.n6 load.t12 19.5798
R2963 load.n12 load.t11 19.5798
R2964 load.n18 load.t6 19.5798
R2965 load.n24 load.t22 19.5798
R2966 load.n30 load.t16 19.5798
R2967 load.n2 load.t24 19.5798
R2968 load.n3 load.t15 19.4007
R2969 load.n9 load.t21 19.4007
R2970 load.n15 load.t27 19.4007
R2971 load.n21 load.t10 19.4007
R2972 load.n27 load.t29 19.4007
R2973 load.n0 load.t8 19.4007
R2974 load.n33 load.n32 15.5531
R2975 load.n8 load.n7 8.46371
R2976 load.n20 load.n19 8.37371
R2977 load.n14 load.n13 8.32871
R2978 load.n26 load.n25 8.32871
R2979 load.n32 load.n31 8.32871
R2980 load.n5 load.n4 7.87164
R2981 load.n11 load.n10 7.87164
R2982 load.n17 load.n16 7.87164
R2983 load.n23 load.n22 7.87164
R2984 load.n29 load.n28 7.87164
R2985 load.n34 load.n1 7.87164
R2986 load.n14 load.n8 7.26762
R2987 load.n32 load.n26 7.22491
R2988 load.n26 load.n20 7.22491
R2989 load.n20 load.n14 7.22491
R2990 load.n7 load.n6 5.00771
R2991 load.n19 load.n18 5.00771
R2992 load.n13 load.n12 4.96432
R2993 load.n25 load.n24 4.96432
R2994 load.n31 load.n30 4.96432
R2995 load.n33 load.n2 4.96432
R2996 load.n13 load.n11 2.11068
R2997 load.n25 load.n23 2.11068
R2998 load.n31 load.n29 2.11068
R2999 load.n34 load.n33 2.11068
R3000 load.n7 load.n5 2.06729
R3001 load.n19 load.n17 2.06729
R3002 load.n5 2inmux_0.Load 0.2255
R3003 load.n11 2inmux_2.Load 0.2255
R3004 load.n17 2inmux_3.Load 0.2255
R3005 load.n23 2inmux_4.Load 0.2255
R3006 load.n29 2inmux_5.Load 0.2255
R3007 2inmux_1.Load load.n34 0.2255
R3008 load.n8 load 0.211008
R3009 load.n4 load.n3 0.106438
R3010 load.n10 load.n9 0.106438
R3011 load.n16 load.n15 0.106438
R3012 load.n22 load.n21 0.106438
R3013 load.n28 load.n27 0.106438
R3014 load.n1 load.n0 0.106438
R3015 a_39178_3501.n0 a_39178_3501.t5 34.1797
R3016 a_39178_3501.n0 a_39178_3501.t4 19.5798
R3017 a_39178_3501.n1 a_39178_3501.t2 18.7717
R3018 a_39178_3501.n1 a_39178_3501.t1 9.2885
R3019 a_39178_3501.n2 a_39178_3501.n0 4.93379
R3020 a_39178_3501.n3 a_39178_3501.t3 4.23346
R3021 a_39178_3501.t0 a_39178_3501.n3 3.85546
R3022 a_39178_3501.n2 a_39178_3501.n1 0.4055
R3023 a_39178_3501.n3 a_39178_3501.n2 0.352625
R3024 dffrs_2.Q.n3 dffrs_2.Q.t8 40.6313
R3025 dffrs_2.Q.n1 dffrs_2.Q.t7 34.1066
R3026 dffrs_2.Q.n3 dffrs_2.Q.t5 27.3166
R3027 dffrs_2.Q.n0 dffrs_2.Q.t4 19.673
R3028 dffrs_2.Q.n0 dffrs_2.Q.t6 19.4007
R3029 dffrs_2.Q.n7 dffrs_2.Q.n3 14.6967
R3030 dffrs_2.Q.n6 dffrs_2.Q.t1 10.0473
R3031 dffrs_2.Q.n7 dffrs_2.Q.n6 9.39565
R3032 dffrs_2.Q.n2 dffrs_2.Q.n1 6.70486
R3033 dffrs_2.Q.n5 dffrs_2.Q.t0 6.51042
R3034 dffrs_2.Q.n5 dffrs_2.Q.n4 6.04952
R3035 dffrs_2.Q dffrs_2.Q.n2 5.81514
R3036 dffrs_2.Q.n6 dffrs_2.Q.n5 0.732092
R3037 dffrs_2.Q.n4 dffrs_2.Q.t3 0.7285
R3038 dffrs_2.Q.n4 dffrs_2.Q.t2 0.7285
R3039 dffrs_2.Q dffrs_2.Q.n7 0.458082
R3040 dffrs_2.Q.n1 dffrs_2.Q.n0 0.252687
R3041 dffrs_2.Q.n2 2inmux_4.Bit 0.0519286
R3042 a_48650_1161.n0 a_48650_1161.t5 34.1797
R3043 a_48650_1161.n0 a_48650_1161.t4 19.5798
R3044 a_48650_1161.n1 a_48650_1161.t1 18.7717
R3045 a_48650_1161.n1 a_48650_1161.t3 9.2885
R3046 a_48650_1161.n2 a_48650_1161.n0 4.93379
R3047 a_48650_1161.t0 a_48650_1161.n3 4.23346
R3048 a_48650_1161.n3 a_48650_1161.t2 3.85546
R3049 a_48650_1161.n2 a_48650_1161.n1 0.4055
R3050 a_48650_1161.n3 a_48650_1161.n2 0.352625
R3051 a_50878_1605.n0 a_50878_1605.t5 34.1797
R3052 a_50878_1605.n0 a_50878_1605.t4 19.5798
R3053 a_50878_1605.n1 a_50878_1605.t3 10.3401
R3054 a_50878_1605.n1 a_50878_1605.t2 9.2885
R3055 a_50878_1605.n2 a_50878_1605.n0 4.93379
R3056 a_50878_1605.t1 a_50878_1605.n3 4.09202
R3057 a_50878_1605.n3 a_50878_1605.t0 3.95079
R3058 a_50878_1605.n2 a_50878_1605.n1 0.599711
R3059 a_50878_1605.n3 a_50878_1605.n2 0.296375
R3060 2inmux_1.OUT.n0 2inmux_1.OUT.t2 41.0041
R3061 2inmux_1.OUT.n0 2inmux_1.OUT.t3 26.9438
R3062 2inmux_1.OUT.n1 2inmux_1.OUT.t1 9.6935
R3063 dffrs_5.d 2inmux_1.OUT.n0 6.55979
R3064 2inmux_1.OUT dffrs_5.d 4.883
R3065 2inmux_1.OUT.n1 2inmux_1.OUT.t0 4.35383
R3066 2inmux_1.OUT 2inmux_1.OUT.n1 0.350857
R3067 a_22462_1605.n0 a_22462_1605.t5 34.1797
R3068 a_22462_1605.n0 a_22462_1605.t4 19.5798
R3069 a_22462_1605.n1 a_22462_1605.t3 10.3401
R3070 a_22462_1605.n1 a_22462_1605.t2 9.2885
R3071 a_22462_1605.n2 a_22462_1605.n0 4.93379
R3072 a_22462_1605.n3 a_22462_1605.t0 4.09202
R3073 a_22462_1605.t1 a_22462_1605.n3 3.95079
R3074 a_22462_1605.n2 a_22462_1605.n1 0.599711
R3075 a_22462_1605.n3 a_22462_1605.n2 0.296375
R3076 a_34936_1559.n0 a_34936_1559.t5 40.8177
R3077 a_34936_1559.n1 a_34936_1559.t6 40.6313
R3078 a_34936_1559.n1 a_34936_1559.t4 27.3166
R3079 a_34936_1559.n0 a_34936_1559.t7 27.1302
R3080 a_34936_1559.n2 a_34936_1559.n1 19.2576
R3081 a_34936_1559.n3 a_34936_1559.t2 10.0473
R3082 a_34936_1559.n4 a_34936_1559.t3 6.51042
R3083 a_34936_1559.n5 a_34936_1559.n4 6.04952
R3084 a_34936_1559.n2 a_34936_1559.n0 5.91752
R3085 a_34936_1559.n3 a_34936_1559.n2 4.89565
R3086 a_34936_1559.n4 a_34936_1559.n3 0.732092
R3087 a_34936_1559.n5 a_34936_1559.t1 0.7285
R3088 a_34936_1559.t0 a_34936_1559.n5 0.7285
R3089 a_34936_3764.n1 a_34936_3764.t8 41.0041
R3090 a_34936_3764.n0 a_34936_3764.t6 40.8177
R3091 a_34936_3764.n2 a_34936_3764.t7 40.6313
R3092 a_34936_3764.n2 a_34936_3764.t4 27.3166
R3093 a_34936_3764.n0 a_34936_3764.t9 27.1302
R3094 a_34936_3764.n1 a_34936_3764.t5 26.9438
R3095 a_34936_3764.n3 a_34936_3764.n1 15.6312
R3096 a_34936_3764.n3 a_34936_3764.n2 15.046
R3097 a_34936_3764.n5 a_34936_3764.t2 10.0473
R3098 a_34936_3764.n6 a_34936_3764.t3 6.51042
R3099 a_34936_3764.n7 a_34936_3764.n6 6.04952
R3100 a_34936_3764.n4 a_34936_3764.n0 5.64619
R3101 a_34936_3764.n5 a_34936_3764.n4 5.17851
R3102 a_34936_3764.n4 a_34936_3764.n3 4.5005
R3103 a_34936_3764.n6 a_34936_3764.n5 0.732092
R3104 a_34936_3764.t0 a_34936_3764.n7 0.7285
R3105 a_34936_3764.n7 a_34936_3764.t1 0.7285
R3106 a_3518_1604.n0 a_3518_1604.t5 34.1797
R3107 a_3518_1604.n0 a_3518_1604.t4 19.5798
R3108 a_3518_1604.n1 a_3518_1604.t3 10.3401
R3109 a_3518_1604.n1 a_3518_1604.t2 9.2885
R3110 a_3518_1604.n2 a_3518_1604.n0 4.93379
R3111 a_3518_1604.t1 a_3518_1604.n3 4.09202
R3112 a_3518_1604.n3 a_3518_1604.t0 3.95079
R3113 a_3518_1604.n2 a_3518_1604.n1 0.599711
R3114 a_3518_1604.n3 a_3518_1604.n2 0.296375
R3115 2inmux_0.OUT.n0 2inmux_0.OUT.t2 41.0041
R3116 2inmux_0.OUT.n0 2inmux_0.OUT.t3 26.9438
R3117 2inmux_0.OUT.n1 2inmux_0.OUT.t1 9.6935
R3118 dffrs_0.d 2inmux_0.OUT.n0 6.55979
R3119 2inmux_0.OUT dffrs_0.d 4.883
R3120 2inmux_0.OUT.n1 2inmux_0.OUT.t0 4.35383
R3121 2inmux_0.OUT 2inmux_0.OUT.n1 0.350857
R3122 a_44408_3764.n1 a_44408_3764.t6 41.0041
R3123 a_44408_3764.n0 a_44408_3764.t5 40.8177
R3124 a_44408_3764.n2 a_44408_3764.t4 40.6313
R3125 a_44408_3764.n2 a_44408_3764.t7 27.3166
R3126 a_44408_3764.n0 a_44408_3764.t9 27.1302
R3127 a_44408_3764.n1 a_44408_3764.t8 26.9438
R3128 a_44408_3764.n3 a_44408_3764.n1 15.6312
R3129 a_44408_3764.n3 a_44408_3764.n2 15.046
R3130 a_44408_3764.n5 a_44408_3764.t2 10.0473
R3131 a_44408_3764.n6 a_44408_3764.t3 6.51042
R3132 a_44408_3764.n7 a_44408_3764.n6 6.04952
R3133 a_44408_3764.n4 a_44408_3764.n0 5.64619
R3134 a_44408_3764.n5 a_44408_3764.n4 5.17851
R3135 a_44408_3764.n4 a_44408_3764.n3 4.5005
R3136 a_44408_3764.n6 a_44408_3764.n5 0.732092
R3137 a_44408_3764.t0 a_44408_3764.n7 0.7285
R3138 a_44408_3764.n7 a_44408_3764.t1 0.7285
R3139 a_20234_1161.n0 a_20234_1161.t4 34.1797
R3140 a_20234_1161.n0 a_20234_1161.t5 19.5798
R3141 a_20234_1161.n1 a_20234_1161.t3 18.7717
R3142 a_20234_1161.n1 a_20234_1161.t2 9.2885
R3143 a_20234_1161.n2 a_20234_1161.n0 4.93379
R3144 a_20234_1161.t0 a_20234_1161.n3 4.23346
R3145 a_20234_1161.n3 a_20234_1161.t1 3.85546
R3146 a_20234_1161.n2 a_20234_1161.n1 0.4055
R3147 a_20234_1161.n3 a_20234_1161.n2 0.352625
R3148 a_29706_1161.n0 a_29706_1161.t4 34.1797
R3149 a_29706_1161.n0 a_29706_1161.t5 19.5798
R3150 a_29706_1161.n1 a_29706_1161.t2 18.7717
R3151 a_29706_1161.n1 a_29706_1161.t1 9.2885
R3152 a_29706_1161.n2 a_29706_1161.n0 4.93379
R3153 a_29706_1161.t0 a_29706_1161.n3 4.23346
R3154 a_29706_1161.n3 a_29706_1161.t3 3.85546
R3155 a_29706_1161.n2 a_29706_1161.n1 0.4055
R3156 a_29706_1161.n3 a_29706_1161.n2 0.352625
R3157 a_25464_3764.n1 a_25464_3764.t5 41.0041
R3158 a_25464_3764.n0 a_25464_3764.t4 40.8177
R3159 a_25464_3764.n2 a_25464_3764.t6 40.6313
R3160 a_25464_3764.n2 a_25464_3764.t9 27.3166
R3161 a_25464_3764.n0 a_25464_3764.t8 27.1302
R3162 a_25464_3764.n1 a_25464_3764.t7 26.9438
R3163 a_25464_3764.n3 a_25464_3764.n1 15.6312
R3164 a_25464_3764.n3 a_25464_3764.n2 15.046
R3165 a_25464_3764.n5 a_25464_3764.t2 10.0473
R3166 a_25464_3764.n6 a_25464_3764.t3 6.51042
R3167 a_25464_3764.n7 a_25464_3764.n6 6.04952
R3168 a_25464_3764.n4 a_25464_3764.n0 5.64619
R3169 a_25464_3764.n5 a_25464_3764.n4 5.17851
R3170 a_25464_3764.n4 a_25464_3764.n3 4.5005
R3171 a_25464_3764.n6 a_25464_3764.n5 0.732092
R3172 a_25464_3764.t0 a_25464_3764.n7 0.7285
R3173 a_25464_3764.n7 a_25464_3764.t1 0.7285
R3174 B6.n1 B6.t1 34.2529
R3175 B6.n0 B6.t0 19.673
R3176 B6.n0 B6.t2 19.4007
R3177 B6.n2 B6.n1 8.05164
R3178 B6.n2 B6 1.87121
R3179 B6.n1 B6.n0 0.106438
R3180 2inmux_0.In B6.n2 0.0455
R3181 a_1290_1160.n0 a_1290_1160.t5 34.1797
R3182 a_1290_1160.n0 a_1290_1160.t4 19.5798
R3183 a_1290_1160.n1 a_1290_1160.t3 18.7717
R3184 a_1290_1160.n1 a_1290_1160.t2 9.2885
R3185 a_1290_1160.n2 a_1290_1160.n0 4.93379
R3186 a_1290_1160.t0 a_1290_1160.n3 4.23346
R3187 a_1290_1160.n3 a_1290_1160.t1 3.85546
R3188 a_1290_1160.n2 a_1290_1160.n1 0.4055
R3189 a_1290_1160.n3 a_1290_1160.n2 0.352625
R3190 a_10762_3500.n0 a_10762_3500.t5 34.1797
R3191 a_10762_3500.n0 a_10762_3500.t4 19.5798
R3192 a_10762_3500.t1 a_10762_3500.n3 18.7717
R3193 a_10762_3500.n3 a_10762_3500.t0 9.2885
R3194 a_10762_3500.n2 a_10762_3500.n0 4.93379
R3195 a_10762_3500.n1 a_10762_3500.t3 4.23346
R3196 a_10762_3500.n1 a_10762_3500.t2 3.85546
R3197 a_10762_3500.n3 a_10762_3500.n2 0.4055
R3198 a_10762_3500.n2 a_10762_3500.n1 0.352625
R3199 a_35016_2511.n0 a_35016_2511.t5 41.0041
R3200 a_35016_2511.n1 a_35016_2511.t6 40.8177
R3201 a_35016_2511.n1 a_35016_2511.t4 27.1302
R3202 a_35016_2511.n0 a_35016_2511.t7 26.9438
R3203 a_35016_2511.n2 a_35016_2511.n1 22.5284
R3204 a_35016_2511.n3 a_35016_2511.n2 19.5781
R3205 a_35016_2511.n3 a_35016_2511.t3 10.0473
R3206 a_35016_2511.n4 a_35016_2511.t2 6.51042
R3207 a_35016_2511.n5 a_35016_2511.n4 6.04952
R3208 a_35016_2511.n2 a_35016_2511.n0 5.7305
R3209 a_35016_2511.n4 a_35016_2511.n3 0.732092
R3210 a_35016_2511.n5 a_35016_2511.t1 0.7285
R3211 a_35016_2511.t0 a_35016_2511.n5 0.7285
R3212 a_41406_1605.n0 a_41406_1605.t5 34.1797
R3213 a_41406_1605.n0 a_41406_1605.t4 19.5798
R3214 a_41406_1605.t0 a_41406_1605.n3 10.3401
R3215 a_41406_1605.n3 a_41406_1605.t1 9.2885
R3216 a_41406_1605.n2 a_41406_1605.n0 4.93379
R3217 a_41406_1605.n1 a_41406_1605.t2 4.09202
R3218 a_41406_1605.n1 a_41406_1605.t3 3.95079
R3219 a_41406_1605.n3 a_41406_1605.n2 0.599711
R3220 a_41406_1605.n2 a_41406_1605.n1 0.296375
R3221 a_44488_2511.n0 a_44488_2511.t7 41.0041
R3222 a_44488_2511.n1 a_44488_2511.t4 40.8177
R3223 a_44488_2511.n1 a_44488_2511.t6 27.1302
R3224 a_44488_2511.n0 a_44488_2511.t5 26.9438
R3225 a_44488_2511.n2 a_44488_2511.n1 22.5284
R3226 a_44488_2511.n3 a_44488_2511.n2 19.5781
R3227 a_44488_2511.n3 a_44488_2511.t1 10.0473
R3228 a_44488_2511.n4 a_44488_2511.t2 6.51042
R3229 a_44488_2511.n5 a_44488_2511.n4 6.04952
R3230 a_44488_2511.n2 a_44488_2511.n0 5.7305
R3231 a_44488_2511.n4 a_44488_2511.n3 0.732092
R3232 a_44488_2511.t0 a_44488_2511.n5 0.7285
R3233 a_44488_2511.n5 a_44488_2511.t3 0.7285
R3234 a_44408_5969.n0 a_44408_5969.t4 40.6313
R3235 a_44408_5969.n0 a_44408_5969.t5 27.3166
R3236 a_44408_5969.n1 a_44408_5969.n0 24.1527
R3237 a_44408_5969.n1 a_44408_5969.t2 10.0473
R3238 a_44408_5969.n2 a_44408_5969.t3 6.51042
R3239 a_44408_5969.n3 a_44408_5969.n2 6.04952
R3240 a_44408_5969.n2 a_44408_5969.n1 0.732092
R3241 a_44408_5969.n3 a_44408_5969.t1 0.7285
R3242 a_44408_5969.t0 a_44408_5969.n3 0.7285
R3243 a_25464_1559.n2 a_25464_1559.t4 40.8177
R3244 a_25464_1559.n3 a_25464_1559.t5 40.6313
R3245 a_25464_1559.n3 a_25464_1559.t7 27.3166
R3246 a_25464_1559.n2 a_25464_1559.t6 27.1302
R3247 a_25464_1559.n4 a_25464_1559.n3 19.2576
R3248 a_25464_1559.t0 a_25464_1559.n5 10.0473
R3249 a_25464_1559.n1 a_25464_1559.t1 6.51042
R3250 a_25464_1559.n1 a_25464_1559.n0 6.04952
R3251 a_25464_1559.n4 a_25464_1559.n2 5.91752
R3252 a_25464_1559.n5 a_25464_1559.n4 4.89565
R3253 a_25464_1559.n5 a_25464_1559.n1 0.732092
R3254 a_25464_1559.n0 a_25464_1559.t3 0.7285
R3255 a_25464_1559.n0 a_25464_1559.t2 0.7285
R3256 a_29706_3501.n0 a_29706_3501.t5 34.1797
R3257 a_29706_3501.n0 a_29706_3501.t4 19.5798
R3258 a_29706_3501.n3 a_29706_3501.t0 18.7717
R3259 a_29706_3501.t1 a_29706_3501.n3 9.2885
R3260 a_29706_3501.n2 a_29706_3501.n0 4.93379
R3261 a_29706_3501.n1 a_29706_3501.t3 4.23346
R3262 a_29706_3501.n1 a_29706_3501.t2 3.85546
R3263 a_29706_3501.n3 a_29706_3501.n2 0.4055
R3264 a_29706_3501.n2 a_29706_3501.n1 0.352625
R3265 dffrs_3.Q.n3 dffrs_3.Q.t6 40.6313
R3266 dffrs_3.Q.n1 dffrs_3.Q.t5 34.1066
R3267 dffrs_3.Q.n3 dffrs_3.Q.t7 27.3166
R3268 dffrs_3.Q.n0 dffrs_3.Q.t8 19.673
R3269 dffrs_3.Q.n0 dffrs_3.Q.t4 19.4007
R3270 dffrs_3.Q.n7 dffrs_3.Q.n3 14.6967
R3271 dffrs_3.Q.n6 dffrs_3.Q.t3 10.0473
R3272 dffrs_3.Q.n7 dffrs_3.Q.n6 9.39565
R3273 dffrs_3.Q.n2 dffrs_3.Q.n1 6.70486
R3274 dffrs_3.Q.n5 dffrs_3.Q.t2 6.51042
R3275 dffrs_3.Q.n5 dffrs_3.Q.n4 6.04952
R3276 dffrs_3.Q dffrs_3.Q.n2 5.81514
R3277 dffrs_3.Q.n6 dffrs_3.Q.n5 0.732092
R3278 dffrs_3.Q.n4 dffrs_3.Q.t0 0.7285
R3279 dffrs_3.Q.n4 dffrs_3.Q.t1 0.7285
R3280 dffrs_3.Q dffrs_3.Q.n7 0.458082
R3281 dffrs_3.Q.n1 dffrs_3.Q.n0 0.252687
R3282 dffrs_3.Q.n2 2inmux_5.Bit 0.0519286
R3283 2inmux_3.OUT.n0 2inmux_3.OUT.t3 41.0041
R3284 2inmux_3.OUT.n0 2inmux_3.OUT.t2 26.9438
R3285 2inmux_3.OUT.n1 2inmux_3.OUT.t1 9.6935
R3286 dffrs_2.d 2inmux_3.OUT.n0 6.55979
R3287 2inmux_3.OUT dffrs_2.d 4.883
R3288 2inmux_3.OUT.n1 2inmux_3.OUT.t0 4.35383
R3289 2inmux_3.OUT 2inmux_3.OUT.n1 0.350857
R3290 a_12990_1604.n0 a_12990_1604.t5 34.1797
R3291 a_12990_1604.n0 a_12990_1604.t4 19.5798
R3292 a_12990_1604.n1 a_12990_1604.t3 10.3401
R3293 a_12990_1604.n1 a_12990_1604.t2 9.2885
R3294 a_12990_1604.n2 a_12990_1604.n0 4.93379
R3295 a_12990_1604.n3 a_12990_1604.t0 4.09202
R3296 a_12990_1604.t1 a_12990_1604.n3 3.95079
R3297 a_12990_1604.n2 a_12990_1604.n1 0.599711
R3298 a_12990_1604.n3 a_12990_1604.n2 0.296375
R3299 a_25464_5969.n0 a_25464_5969.t5 40.6313
R3300 a_25464_5969.n0 a_25464_5969.t4 27.3166
R3301 a_25464_5969.n1 a_25464_5969.n0 24.1527
R3302 a_25464_5969.n1 a_25464_5969.t2 10.0473
R3303 a_25464_5969.n2 a_25464_5969.t3 6.51042
R3304 a_25464_5969.n3 a_25464_5969.n2 6.04952
R3305 a_25464_5969.n2 a_25464_5969.n1 0.732092
R3306 a_25464_5969.n3 a_25464_5969.t1 0.7285
R3307 a_25464_5969.t0 a_25464_5969.n3 0.7285
R3308 a_44408_1559.n0 a_44408_1559.t5 40.8177
R3309 a_44408_1559.n1 a_44408_1559.t4 40.6313
R3310 a_44408_1559.n1 a_44408_1559.t6 27.3166
R3311 a_44408_1559.n0 a_44408_1559.t7 27.1302
R3312 a_44408_1559.n2 a_44408_1559.n1 19.2576
R3313 a_44408_1559.n3 a_44408_1559.t2 10.0473
R3314 a_44408_1559.n4 a_44408_1559.t1 6.51042
R3315 a_44408_1559.n5 a_44408_1559.n4 6.04952
R3316 a_44408_1559.n2 a_44408_1559.n0 5.91752
R3317 a_44408_1559.n3 a_44408_1559.n2 4.89565
R3318 a_44408_1559.n4 a_44408_1559.n3 0.732092
R3319 a_44408_1559.t0 a_44408_1559.n5 0.7285
R3320 a_44408_1559.n5 a_44408_1559.t3 0.7285
R3321 a_53880_1559.n2 a_53880_1559.t6 40.8177
R3322 a_53880_1559.n3 a_53880_1559.t7 40.6313
R3323 a_53880_1559.n3 a_53880_1559.t5 27.3166
R3324 a_53880_1559.n2 a_53880_1559.t4 27.1302
R3325 a_53880_1559.n4 a_53880_1559.n3 19.2576
R3326 a_53880_1559.t0 a_53880_1559.n5 10.0473
R3327 a_53880_1559.n1 a_53880_1559.t2 6.51042
R3328 a_53880_1559.n1 a_53880_1559.n0 6.04952
R3329 a_53880_1559.n4 a_53880_1559.n2 5.91752
R3330 a_53880_1559.n5 a_53880_1559.n4 4.89565
R3331 a_53880_1559.n5 a_53880_1559.n1 0.732092
R3332 a_53880_1559.n0 a_53880_1559.t3 0.7285
R3333 a_53880_1559.n0 a_53880_1559.t1 0.7285
R3334 a_53960_2511.n0 a_53960_2511.t5 41.0041
R3335 a_53960_2511.n1 a_53960_2511.t6 40.8177
R3336 a_53960_2511.n1 a_53960_2511.t4 27.1302
R3337 a_53960_2511.n0 a_53960_2511.t7 26.9438
R3338 a_53960_2511.n2 a_53960_2511.n1 22.5284
R3339 a_53960_2511.n3 a_53960_2511.n2 19.5781
R3340 a_53960_2511.n3 a_53960_2511.t1 10.0473
R3341 a_53960_2511.n4 a_53960_2511.t2 6.51042
R3342 a_53960_2511.n5 a_53960_2511.n4 6.04952
R3343 a_53960_2511.n2 a_53960_2511.n0 5.7305
R3344 a_53960_2511.n4 a_53960_2511.n3 0.732092
R3345 a_53960_2511.n5 a_53960_2511.t3 0.7285
R3346 a_53960_2511.t0 a_53960_2511.n5 0.7285
R3347 a_53880_3764.n1 a_53880_3764.t8 41.0041
R3348 a_53880_3764.n0 a_53880_3764.t7 40.8177
R3349 a_53880_3764.n2 a_53880_3764.t9 40.6313
R3350 a_53880_3764.n2 a_53880_3764.t6 27.3166
R3351 a_53880_3764.n0 a_53880_3764.t4 27.1302
R3352 a_53880_3764.n1 a_53880_3764.t5 26.9438
R3353 a_53880_3764.n3 a_53880_3764.n1 15.6312
R3354 a_53880_3764.n3 a_53880_3764.n2 15.046
R3355 a_53880_3764.n5 a_53880_3764.t2 10.0473
R3356 a_53880_3764.n6 a_53880_3764.t3 6.51042
R3357 a_53880_3764.n7 a_53880_3764.n6 6.04952
R3358 a_53880_3764.n4 a_53880_3764.n0 5.64619
R3359 a_53880_3764.n5 a_53880_3764.n4 5.17851
R3360 a_53880_3764.n4 a_53880_3764.n3 4.5005
R3361 a_53880_3764.n6 a_53880_3764.n5 0.732092
R3362 a_53880_3764.t0 a_53880_3764.n7 0.7285
R3363 a_53880_3764.n7 a_53880_3764.t1 0.7285
R3364 2inmux_2.OUT.n0 2inmux_2.OUT.t2 41.0041
R3365 2inmux_2.OUT.n0 2inmux_2.OUT.t3 26.9438
R3366 2inmux_2.OUT.n1 2inmux_2.OUT.t1 9.6935
R3367 dffrs_1.d 2inmux_2.OUT.n0 6.55979
R3368 2inmux_2.OUT dffrs_1.d 4.883
R3369 2inmux_2.OUT.n1 2inmux_2.OUT.t0 4.35383
R3370 2inmux_2.OUT 2inmux_2.OUT.n1 0.350857
R3371 a_16072_2510.n0 a_16072_2510.t4 41.0041
R3372 a_16072_2510.n1 a_16072_2510.t5 40.8177
R3373 a_16072_2510.n1 a_16072_2510.t7 27.1302
R3374 a_16072_2510.n0 a_16072_2510.t6 26.9438
R3375 a_16072_2510.n2 a_16072_2510.n1 22.5284
R3376 a_16072_2510.n3 a_16072_2510.n2 19.5781
R3377 a_16072_2510.n3 a_16072_2510.t1 10.0473
R3378 a_16072_2510.n4 a_16072_2510.t2 6.51042
R3379 a_16072_2510.n5 a_16072_2510.n4 6.04952
R3380 a_16072_2510.n2 a_16072_2510.n0 5.7305
R3381 a_16072_2510.n4 a_16072_2510.n3 0.732092
R3382 a_16072_2510.t0 a_16072_2510.n5 0.7285
R3383 a_16072_2510.n5 a_16072_2510.t3 0.7285
R3384 a_34936_5969.n0 a_34936_5969.t5 40.6313
R3385 a_34936_5969.n0 a_34936_5969.t4 27.3166
R3386 a_34936_5969.n1 a_34936_5969.n0 24.1527
R3387 a_34936_5969.n1 a_34936_5969.t2 10.0473
R3388 a_34936_5969.n2 a_34936_5969.t1 6.51042
R3389 a_34936_5969.n3 a_34936_5969.n2 6.04952
R3390 a_34936_5969.n2 a_34936_5969.n1 0.732092
R3391 a_34936_5969.t0 a_34936_5969.n3 0.7285
R3392 a_34936_5969.n3 a_34936_5969.t3 0.7285
R3393 a_15992_1558.n0 a_15992_1558.t4 40.8177
R3394 a_15992_1558.n1 a_15992_1558.t5 40.6313
R3395 a_15992_1558.n1 a_15992_1558.t7 27.3166
R3396 a_15992_1558.n0 a_15992_1558.t6 27.1302
R3397 a_15992_1558.n2 a_15992_1558.n1 19.2576
R3398 a_15992_1558.n3 a_15992_1558.t2 10.0473
R3399 a_15992_1558.n4 a_15992_1558.t1 6.51042
R3400 a_15992_1558.n5 a_15992_1558.n4 6.04952
R3401 a_15992_1558.n2 a_15992_1558.n0 5.91752
R3402 a_15992_1558.n3 a_15992_1558.n2 4.89565
R3403 a_15992_1558.n4 a_15992_1558.n3 0.732092
R3404 a_15992_1558.n5 a_15992_1558.t3 0.7285
R3405 a_15992_1558.t0 a_15992_1558.n5 0.7285
R3406 a_53880_5969.n2 a_53880_5969.t4 40.6313
R3407 a_53880_5969.n2 a_53880_5969.t5 27.3166
R3408 a_53880_5969.n3 a_53880_5969.n2 24.1527
R3409 a_53880_5969.t0 a_53880_5969.n3 10.0473
R3410 a_53880_5969.n1 a_53880_5969.t1 6.51042
R3411 a_53880_5969.n1 a_53880_5969.n0 6.04952
R3412 a_53880_5969.n3 a_53880_5969.n1 0.732092
R3413 a_53880_5969.n0 a_53880_5969.t2 0.7285
R3414 a_53880_5969.n0 a_53880_5969.t3 0.7285
R3415 a_31934_1605.n0 a_31934_1605.t5 34.1797
R3416 a_31934_1605.n0 a_31934_1605.t4 19.5798
R3417 a_31934_1605.n1 a_31934_1605.t3 10.3401
R3418 a_31934_1605.n1 a_31934_1605.t2 9.2885
R3419 a_31934_1605.n2 a_31934_1605.n0 4.93379
R3420 a_31934_1605.n3 a_31934_1605.t0 4.09202
R3421 a_31934_1605.t1 a_31934_1605.n3 3.95079
R3422 a_31934_1605.n2 a_31934_1605.n1 0.599711
R3423 a_31934_1605.n3 a_31934_1605.n2 0.296375
R3424 2inmux_4.OUT.n0 2inmux_4.OUT.t2 41.0041
R3425 2inmux_4.OUT.n0 2inmux_4.OUT.t3 26.9438
R3426 2inmux_4.OUT.n1 2inmux_4.OUT.t1 9.6935
R3427 dffrs_3.d 2inmux_4.OUT.n0 6.55979
R3428 2inmux_4.OUT dffrs_3.d 4.883
R3429 2inmux_4.OUT.n1 2inmux_4.OUT.t0 4.35383
R3430 2inmux_4.OUT 2inmux_4.OUT.n1 0.350857
R3431 a_25544_2511.n0 a_25544_2511.t6 41.0041
R3432 a_25544_2511.n1 a_25544_2511.t7 40.8177
R3433 a_25544_2511.n1 a_25544_2511.t5 27.1302
R3434 a_25544_2511.n0 a_25544_2511.t4 26.9438
R3435 a_25544_2511.n2 a_25544_2511.n1 22.5284
R3436 a_25544_2511.n3 a_25544_2511.n2 19.5781
R3437 a_25544_2511.n3 a_25544_2511.t2 10.0473
R3438 a_25544_2511.n4 a_25544_2511.t1 6.51042
R3439 a_25544_2511.n5 a_25544_2511.n4 6.04952
R3440 a_25544_2511.n2 a_25544_2511.n0 5.7305
R3441 a_25544_2511.n4 a_25544_2511.n3 0.732092
R3442 a_25544_2511.n5 a_25544_2511.t3 0.7285
R3443 a_25544_2511.t0 a_25544_2511.n5 0.7285
R3444 B5.n1 B5.t0 34.2529
R3445 B5.n0 B5.t1 19.673
R3446 B5.n0 B5.t2 19.4007
R3447 B5.n2 B5.n1 8.05164
R3448 B5.n2 B5 1.87121
R3449 B5.n1 B5.n0 0.106438
R3450 2inmux_2.In B5.n2 0.0455
R3451 a_10762_1160.n0 a_10762_1160.t5 34.1797
R3452 a_10762_1160.n0 a_10762_1160.t4 19.5798
R3453 a_10762_1160.n1 a_10762_1160.t2 18.7717
R3454 a_10762_1160.n1 a_10762_1160.t1 9.2885
R3455 a_10762_1160.n2 a_10762_1160.n0 4.93379
R3456 a_10762_1160.t0 a_10762_1160.n3 4.23346
R3457 a_10762_1160.n3 a_10762_1160.t3 3.85546
R3458 a_10762_1160.n2 a_10762_1160.n1 0.4055
R3459 a_10762_1160.n3 a_10762_1160.n2 0.352625
R3460 a_6520_5968.n0 a_6520_5968.t4 40.6313
R3461 a_6520_5968.n0 a_6520_5968.t5 27.3166
R3462 a_6520_5968.n1 a_6520_5968.n0 24.1527
R3463 a_6520_5968.n1 a_6520_5968.t3 10.0473
R3464 a_6520_5968.n2 a_6520_5968.t2 6.51042
R3465 a_6520_5968.n3 a_6520_5968.n2 6.04952
R3466 a_6520_5968.n2 a_6520_5968.n1 0.732092
R3467 a_6520_5968.n3 a_6520_5968.t1 0.7285
R3468 a_6520_5968.t0 a_6520_5968.n3 0.7285
R3469 serial_out.n0 serial_out.t4 40.6313
R3470 serial_out.n0 serial_out.t5 27.3166
R3471 serial_out.n4 serial_out.n0 14.6967
R3472 serial_out.n3 serial_out.t3 10.0473
R3473 serial_out.n4 serial_out.n3 9.39565
R3474 serial_out.n2 serial_out.t2 6.51042
R3475 serial_out.n2 serial_out.n1 6.04952
R3476 dffrs_5.Q serial_out 5.90514
R3477 serial_out.n3 serial_out.n2 0.732092
R3478 serial_out.n1 serial_out.t0 0.7285
R3479 serial_out.n1 serial_out.t1 0.7285
R3480 dffrs_5.Q serial_out.n4 0.458082
R3481 B2.n1 B2.t2 34.2529
R3482 B2.n0 B2.t0 19.673
R3483 B2.n0 B2.t1 19.4007
R3484 B2.n2 B2.n1 8.05164
R3485 B2.n2 B2 1.87121
R3486 B2.n1 B2.n0 0.106438
R3487 2inmux_5.In B2.n2 0.0455
R3488 a_39178_1161.n0 a_39178_1161.t5 34.1797
R3489 a_39178_1161.n0 a_39178_1161.t4 19.5798
R3490 a_39178_1161.n1 a_39178_1161.t2 18.7717
R3491 a_39178_1161.n1 a_39178_1161.t1 9.2885
R3492 a_39178_1161.n2 a_39178_1161.n0 4.93379
R3493 a_39178_1161.n3 a_39178_1161.t3 4.23346
R3494 a_39178_1161.t0 a_39178_1161.n3 3.85546
R3495 a_39178_1161.n2 a_39178_1161.n1 0.4055
R3496 a_39178_1161.n3 a_39178_1161.n2 0.352625
R3497 2inmux_5.OUT.n0 2inmux_5.OUT.t3 41.0041
R3498 2inmux_5.OUT.n0 2inmux_5.OUT.t2 26.9438
R3499 2inmux_5.OUT.n1 2inmux_5.OUT.t1 9.6935
R3500 dffrs_4.d 2inmux_5.OUT.n0 6.55979
R3501 2inmux_5.OUT dffrs_4.d 4.883
R3502 2inmux_5.OUT.n1 2inmux_5.OUT.t0 4.35383
R3503 2inmux_5.OUT 2inmux_5.OUT.n1 0.350857
R3504 B4.n1 B4.t1 34.2529
R3505 B4.n0 B4.t0 19.673
R3506 B4.n0 B4.t2 19.4007
R3507 B4.n2 B4.n1 8.05164
R3508 B4.n2 B4 1.87282
R3509 B4.n1 B4.n0 0.106438
R3510 2inmux_3.In B4.n2 0.0455
R3511 B1.n1 B1.t1 34.2529
R3512 B1.n0 B1.t0 19.673
R3513 B1.n0 B1.t2 19.4007
R3514 B1.n2 B1.n1 8.05164
R3515 B1.n2 B1 1.87121
R3516 B1.n1 B1.n0 0.106438
R3517 2inmux_1.In B1.n2 0.0455
R3518 B3.n1 B3.t1 34.2529
R3519 B3.n0 B3.t0 19.673
R3520 B3.n0 B3.t2 19.4007
R3521 B3.n2 B3.n1 8.05164
R3522 B3.n2 B3 1.87121
R3523 B3.n1 B3.n0 0.106438
R3524 2inmux_4.In B3.n2 0.0455
C0 2inmux_5.OUT.t3 0 0.27468f **FLOATING
C1 2inmux_5.OUT.t2 0 0.14601f **FLOATING
C2 2inmux_5.OUT.n0 0 0.52483f **FLOATING
C3 dffrs_4.d 0 0.51316f **FLOATING
C4 2inmux_5.OUT.t0 0 0.3775f **FLOATING
C5 2inmux_5.OUT.t1 0 0.1155f **FLOATING
C6 2inmux_5.OUT.n1 0 0.62644f **FLOATING
C7 2inmux_5.OUT 0 0.12188f **FLOATING
C8 a_39178_1161.t5 0 0.15843f **FLOATING
C9 a_39178_1161.t4 0 0.07081f **FLOATING
C10 a_39178_1161.n0 0 0.20989f **FLOATING
C11 a_39178_1161.t2 0 0.08492f **FLOATING
C12 a_39178_1161.t1 0 0.04534f **FLOATING
C13 a_39178_1161.n1 0 0.14994f **FLOATING
C14 a_39178_1161.n2 0 0.12745f **FLOATING
C15 a_39178_1161.t3 0 0.18548f **FLOATING
C16 a_39178_1161.n3 0 0.92376f **FLOATING
C17 a_39178_1161.t0 0 0.144f **FLOATING
C18 serial_out 0 0.25909f **FLOATING
C19 serial_out.t4 0 0.098f **FLOATING
C20 serial_out.t5 0 0.05344f **FLOATING
C21 serial_out.n0 0 0.38053f **FLOATING
C22 serial_out.t0 0 0.03269f **FLOATING
C23 serial_out.t1 0 0.03269f **FLOATING
C24 serial_out.n1 0 0.11684f **FLOATING
C25 serial_out.t2 0 0.14452f **FLOATING
C26 serial_out.n2 0 0.20435f **FLOATING
C27 serial_out.t3 0 0.05218f **FLOATING
C28 serial_out.n3 0 0.1756f **FLOATING
C29 serial_out.n4 0 0.36768f **FLOATING
C30 dffrs_5.Q 0 0.2824f **FLOATING
C31 a_6520_5968.t1 0 0.05581f **FLOATING
C32 a_6520_5968.t3 0 0.0891f **FLOATING
C33 a_6520_5968.t4 0 0.16734f **FLOATING
C34 a_6520_5968.t5 0 0.09125f **FLOATING
C35 a_6520_5968.n0 0 0.88217f **FLOATING
C36 a_6520_5968.n1 0 0.66334f **FLOATING
C37 a_6520_5968.t2 0 0.24676f **FLOATING
C38 a_6520_5968.n2 0 0.34892f **FLOATING
C39 a_6520_5968.n3 0 0.1995f **FLOATING
C40 a_6520_5968.t0 0 0.05581f **FLOATING
C41 a_10762_1160.t5 0 0.15843f **FLOATING
C42 a_10762_1160.t4 0 0.07081f **FLOATING
C43 a_10762_1160.n0 0 0.20989f **FLOATING
C44 a_10762_1160.t2 0 0.08492f **FLOATING
C45 a_10762_1160.t1 0 0.04534f **FLOATING
C46 a_10762_1160.n1 0 0.14994f **FLOATING
C47 a_10762_1160.n2 0 0.12745f **FLOATING
C48 a_10762_1160.t3 0 0.144f **FLOATING
C49 a_10762_1160.n3 0 0.92376f **FLOATING
C50 a_10762_1160.t0 0 0.18548f **FLOATING
C51 a_25544_2511.t3 0 0.04533f **FLOATING
C52 a_25544_2511.t2 0 0.07236f **FLOATING
C53 a_25544_2511.t6 0 0.13696f **FLOATING
C54 a_25544_2511.t4 0 0.07281f **FLOATING
C55 a_25544_2511.n0 0 0.23752f **FLOATING
C56 a_25544_2511.t7 0 0.13638f **FLOATING
C57 a_25544_2511.t5 0 0.07339f **FLOATING
C58 a_25544_2511.n1 0 0.71031f **FLOATING
C59 a_25544_2511.n2 0 1.37628f **FLOATING
C60 a_25544_2511.n3 0 0.44756f **FLOATING
C61 a_25544_2511.t1 0 0.2004f **FLOATING
C62 a_25544_2511.n4 0 0.28337f **FLOATING
C63 a_25544_2511.n5 0 0.16202f **FLOATING
C64 a_25544_2511.t0 0 0.04533f **FLOATING
C65 2inmux_4.OUT.t2 0 0.27468f **FLOATING
C66 2inmux_4.OUT.t3 0 0.14601f **FLOATING
C67 2inmux_4.OUT.n0 0 0.52483f **FLOATING
C68 dffrs_3.d 0 0.51316f **FLOATING
C69 2inmux_4.OUT.t0 0 0.3775f **FLOATING
C70 2inmux_4.OUT.t1 0 0.1155f **FLOATING
C71 2inmux_4.OUT.n1 0 0.62644f **FLOATING
C72 2inmux_4.OUT 0 0.12188f **FLOATING
C73 a_31934_1605.t5 0 0.1705f **FLOATING
C74 a_31934_1605.t4 0 0.0762f **FLOATING
C75 a_31934_1605.n0 0 0.22588f **FLOATING
C76 a_31934_1605.t3 0 0.06122f **FLOATING
C77 a_31934_1605.t2 0 0.0488f **FLOATING
C78 a_31934_1605.n1 0 0.29156f **FLOATING
C79 a_31934_1605.n2 0 0.15481f **FLOATING
C80 a_31934_1605.t0 0 0.21992f **FLOATING
C81 a_31934_1605.n3 0 0.54012f **FLOATING
C82 a_31934_1605.t1 0 0.21101f **FLOATING
C83 a_53880_5969.t2 0 0.05581f **FLOATING
C84 a_53880_5969.t3 0 0.05581f **FLOATING
C85 a_53880_5969.n0 0 0.1995f **FLOATING
C86 a_53880_5969.t1 0 0.24676f **FLOATING
C87 a_53880_5969.n1 0 0.34892f **FLOATING
C88 a_53880_5969.t4 0 0.16734f **FLOATING
C89 a_53880_5969.t5 0 0.09125f **FLOATING
C90 a_53880_5969.n2 0 0.88217f **FLOATING
C91 a_53880_5969.n3 0 0.66334f **FLOATING
C92 a_53880_5969.t0 0 0.0891f **FLOATING
C93 a_15992_1558.t3 0 0.06293f **FLOATING
C94 a_15992_1558.t2 0 0.10047f **FLOATING
C95 a_15992_1558.t4 0 0.18936f **FLOATING
C96 a_15992_1558.t6 0 0.10189f **FLOATING
C97 a_15992_1558.n0 0 0.33658f **FLOATING
C98 a_15992_1558.t5 0 0.18869f **FLOATING
C99 a_15992_1558.t7 0 0.1029f **FLOATING
C100 a_15992_1558.n1 0 0.87879f **FLOATING
C101 a_15992_1558.n2 0 0.78698f **FLOATING
C102 a_15992_1558.n3 0 0.29183f **FLOATING
C103 a_15992_1558.t1 0 0.27825f **FLOATING
C104 a_15992_1558.n4 0 0.39345f **FLOATING
C105 a_15992_1558.n5 0 0.22496f **FLOATING
C106 a_15992_1558.t0 0 0.06293f **FLOATING
C107 a_34936_5969.t3 0 0.05581f **FLOATING
C108 a_34936_5969.t2 0 0.0891f **FLOATING
C109 a_34936_5969.t5 0 0.16734f **FLOATING
C110 a_34936_5969.t4 0 0.09125f **FLOATING
C111 a_34936_5969.n0 0 0.88217f **FLOATING
C112 a_34936_5969.n1 0 0.66334f **FLOATING
C113 a_34936_5969.t1 0 0.24676f **FLOATING
C114 a_34936_5969.n2 0 0.34892f **FLOATING
C115 a_34936_5969.n3 0 0.1995f **FLOATING
C116 a_34936_5969.t0 0 0.05581f **FLOATING
C117 a_16072_2510.t3 0 0.04533f **FLOATING
C118 a_16072_2510.t1 0 0.07236f **FLOATING
C119 a_16072_2510.t4 0 0.13696f **FLOATING
C120 a_16072_2510.t6 0 0.07281f **FLOATING
C121 a_16072_2510.n0 0 0.23752f **FLOATING
C122 a_16072_2510.t5 0 0.13638f **FLOATING
C123 a_16072_2510.t7 0 0.07339f **FLOATING
C124 a_16072_2510.n1 0 0.71031f **FLOATING
C125 a_16072_2510.n2 0 1.37628f **FLOATING
C126 a_16072_2510.n3 0 0.44756f **FLOATING
C127 a_16072_2510.t2 0 0.2004f **FLOATING
C128 a_16072_2510.n4 0 0.28337f **FLOATING
C129 a_16072_2510.n5 0 0.16202f **FLOATING
C130 a_16072_2510.t0 0 0.04533f **FLOATING
C131 2inmux_2.OUT.t2 0 0.27468f **FLOATING
C132 2inmux_2.OUT.t3 0 0.14601f **FLOATING
C133 2inmux_2.OUT.n0 0 0.52483f **FLOATING
C134 dffrs_1.d 0 0.51316f **FLOATING
C135 2inmux_2.OUT.t0 0 0.3775f **FLOATING
C136 2inmux_2.OUT.t1 0 0.1155f **FLOATING
C137 2inmux_2.OUT.n1 0 0.62644f **FLOATING
C138 2inmux_2.OUT 0 0.12188f **FLOATING
C139 a_53880_3764.t1 0 0.04005f **FLOATING
C140 a_53880_3764.t2 0 0.06394f **FLOATING
C141 a_53880_3764.t7 0 0.12051f **FLOATING
C142 a_53880_3764.t4 0 0.06484f **FLOATING
C143 a_53880_3764.n0 0 0.20809f **FLOATING
C144 a_53880_3764.t8 0 0.12102f **FLOATING
C145 a_53880_3764.t5 0 0.06433f **FLOATING
C146 a_53880_3764.n1 0 0.50381f **FLOATING
C147 a_53880_3764.t9 0 0.12008f **FLOATING
C148 a_53880_3764.t6 0 0.06549f **FLOATING
C149 a_53880_3764.n2 0 0.48367f **FLOATING
C150 a_53880_3764.n3 0 0.84489f **FLOATING
C151 a_53880_3764.n4 0 0.19941f **FLOATING
C152 a_53880_3764.n5 0 0.18919f **FLOATING
C153 a_53880_3764.t3 0 0.17708f **FLOATING
C154 a_53880_3764.n6 0 0.25039f **FLOATING
C155 a_53880_3764.n7 0 0.14316f **FLOATING
C156 a_53880_3764.t0 0 0.04005f **FLOATING
C157 a_53960_2511.t3 0 0.04533f **FLOATING
C158 a_53960_2511.t1 0 0.07236f **FLOATING
C159 a_53960_2511.t5 0 0.13696f **FLOATING
C160 a_53960_2511.t7 0 0.07281f **FLOATING
C161 a_53960_2511.n0 0 0.23752f **FLOATING
C162 a_53960_2511.t6 0 0.13638f **FLOATING
C163 a_53960_2511.t4 0 0.07339f **FLOATING
C164 a_53960_2511.n1 0 0.71031f **FLOATING
C165 a_53960_2511.n2 0 1.37628f **FLOATING
C166 a_53960_2511.n3 0 0.44756f **FLOATING
C167 a_53960_2511.t2 0 0.2004f **FLOATING
C168 a_53960_2511.n4 0 0.28337f **FLOATING
C169 a_53960_2511.n5 0 0.16202f **FLOATING
C170 a_53960_2511.t0 0 0.04533f **FLOATING
C171 a_53880_1559.t3 0 0.06293f **FLOATING
C172 a_53880_1559.t1 0 0.06293f **FLOATING
C173 a_53880_1559.n0 0 0.22496f **FLOATING
C174 a_53880_1559.t2 0 0.27825f **FLOATING
C175 a_53880_1559.n1 0 0.39345f **FLOATING
C176 a_53880_1559.t6 0 0.18936f **FLOATING
C177 a_53880_1559.t4 0 0.10189f **FLOATING
C178 a_53880_1559.n2 0 0.33658f **FLOATING
C179 a_53880_1559.t7 0 0.18869f **FLOATING
C180 a_53880_1559.t5 0 0.1029f **FLOATING
C181 a_53880_1559.n3 0 0.87879f **FLOATING
C182 a_53880_1559.n4 0 0.78698f **FLOATING
C183 a_53880_1559.n5 0 0.29183f **FLOATING
C184 a_53880_1559.t0 0 0.10047f **FLOATING
C185 a_44408_1559.t3 0 0.06293f **FLOATING
C186 a_44408_1559.t2 0 0.10047f **FLOATING
C187 a_44408_1559.t5 0 0.18936f **FLOATING
C188 a_44408_1559.t7 0 0.10189f **FLOATING
C189 a_44408_1559.n0 0 0.33658f **FLOATING
C190 a_44408_1559.t4 0 0.18869f **FLOATING
C191 a_44408_1559.t6 0 0.1029f **FLOATING
C192 a_44408_1559.n1 0 0.87879f **FLOATING
C193 a_44408_1559.n2 0 0.78698f **FLOATING
C194 a_44408_1559.n3 0 0.29183f **FLOATING
C195 a_44408_1559.t1 0 0.27825f **FLOATING
C196 a_44408_1559.n4 0 0.39345f **FLOATING
C197 a_44408_1559.n5 0 0.22496f **FLOATING
C198 a_44408_1559.t0 0 0.06293f **FLOATING
C199 a_25464_5969.t1 0 0.05581f **FLOATING
C200 a_25464_5969.t2 0 0.0891f **FLOATING
C201 a_25464_5969.t5 0 0.16734f **FLOATING
C202 a_25464_5969.t4 0 0.09125f **FLOATING
C203 a_25464_5969.n0 0 0.88217f **FLOATING
C204 a_25464_5969.n1 0 0.66334f **FLOATING
C205 a_25464_5969.t3 0 0.24676f **FLOATING
C206 a_25464_5969.n2 0 0.34892f **FLOATING
C207 a_25464_5969.n3 0 0.1995f **FLOATING
C208 a_25464_5969.t0 0 0.05581f **FLOATING
C209 a_12990_1604.t5 0 0.1705f **FLOATING
C210 a_12990_1604.t4 0 0.0762f **FLOATING
C211 a_12990_1604.n0 0 0.22588f **FLOATING
C212 a_12990_1604.t3 0 0.06122f **FLOATING
C213 a_12990_1604.t2 0 0.0488f **FLOATING
C214 a_12990_1604.n1 0 0.29156f **FLOATING
C215 a_12990_1604.n2 0 0.15481f **FLOATING
C216 a_12990_1604.t0 0 0.21992f **FLOATING
C217 a_12990_1604.n3 0 0.54012f **FLOATING
C218 a_12990_1604.t1 0 0.21101f **FLOATING
C219 2inmux_3.OUT.t3 0 0.27468f **FLOATING
C220 2inmux_3.OUT.t2 0 0.14601f **FLOATING
C221 2inmux_3.OUT.n0 0 0.52483f **FLOATING
C222 dffrs_2.d 0 0.51316f **FLOATING
C223 2inmux_3.OUT.t0 0 0.3775f **FLOATING
C224 2inmux_3.OUT.t1 0 0.1155f **FLOATING
C225 2inmux_3.OUT.n1 0 0.62644f **FLOATING
C226 2inmux_3.OUT 0 0.12188f **FLOATING
C227 dffrs_3.Q.t5 0 0.14856f **FLOATING
C228 dffrs_3.Q.t8 0 0.06654f **FLOATING
C229 dffrs_3.Q.t4 0 0.06601f **FLOATING
C230 dffrs_3.Q.n0 0 0.10908f **FLOATING
C231 dffrs_3.Q.n1 0 0.1562f **FLOATING
C232 2inmux_5.Bit 0 0.00243f **FLOATING
C233 dffrs_3.Q.n2 0 0.46007f **FLOATING
C234 dffrs_3.Q.t6 0 0.1058f **FLOATING
C235 dffrs_3.Q.t7 0 0.0577f **FLOATING
C236 dffrs_3.Q.n3 0 0.41081f **FLOATING
C237 dffrs_3.Q.t0 0 0.03529f **FLOATING
C238 dffrs_3.Q.t1 0 0.03529f **FLOATING
C239 dffrs_3.Q.n4 0 0.12614f **FLOATING
C240 dffrs_3.Q.t2 0 0.15602f **FLOATING
C241 dffrs_3.Q.n5 0 0.22061f **FLOATING
C242 dffrs_3.Q.t3 0 0.05633f **FLOATING
C243 dffrs_3.Q.n6 0 0.18958f **FLOATING
C244 dffrs_3.Q.n7 0 0.39693f **FLOATING
C245 dffrs_3.Q 0 0.30061f **FLOATING
C246 a_29706_3501.t5 0 0.16597f **FLOATING
C247 a_29706_3501.t4 0 0.07418f **FLOATING
C248 a_29706_3501.n0 0 0.21988f **FLOATING
C249 a_29706_3501.t2 0 0.15085f **FLOATING
C250 a_29706_3501.t3 0 0.19431f **FLOATING
C251 a_29706_3501.n1 0 0.96775f **FLOATING
C252 a_29706_3501.n2 0 0.13352f **FLOATING
C253 a_29706_3501.t0 0 0.08896f **FLOATING
C254 a_29706_3501.n3 0 0.15708f **FLOATING
C255 a_29706_3501.t1 0 0.0475f **FLOATING
C256 a_25464_1559.t3 0 0.06293f **FLOATING
C257 a_25464_1559.t2 0 0.06293f **FLOATING
C258 a_25464_1559.n0 0 0.22496f **FLOATING
C259 a_25464_1559.t1 0 0.27825f **FLOATING
C260 a_25464_1559.n1 0 0.39345f **FLOATING
C261 a_25464_1559.t4 0 0.18936f **FLOATING
C262 a_25464_1559.t6 0 0.10189f **FLOATING
C263 a_25464_1559.n2 0 0.33658f **FLOATING
C264 a_25464_1559.t5 0 0.18869f **FLOATING
C265 a_25464_1559.t7 0 0.1029f **FLOATING
C266 a_25464_1559.n3 0 0.87879f **FLOATING
C267 a_25464_1559.n4 0 0.78698f **FLOATING
C268 a_25464_1559.n5 0 0.29183f **FLOATING
C269 a_25464_1559.t0 0 0.10047f **FLOATING
C270 a_44408_5969.t1 0 0.05581f **FLOATING
C271 a_44408_5969.t2 0 0.0891f **FLOATING
C272 a_44408_5969.t4 0 0.16734f **FLOATING
C273 a_44408_5969.t5 0 0.09125f **FLOATING
C274 a_44408_5969.n0 0 0.88217f **FLOATING
C275 a_44408_5969.n1 0 0.66334f **FLOATING
C276 a_44408_5969.t3 0 0.24676f **FLOATING
C277 a_44408_5969.n2 0 0.34892f **FLOATING
C278 a_44408_5969.n3 0 0.1995f **FLOATING
C279 a_44408_5969.t0 0 0.05581f **FLOATING
C280 a_44488_2511.t3 0 0.04533f **FLOATING
C281 a_44488_2511.t1 0 0.07236f **FLOATING
C282 a_44488_2511.t7 0 0.13696f **FLOATING
C283 a_44488_2511.t5 0 0.07281f **FLOATING
C284 a_44488_2511.n0 0 0.23752f **FLOATING
C285 a_44488_2511.t4 0 0.13638f **FLOATING
C286 a_44488_2511.t6 0 0.07339f **FLOATING
C287 a_44488_2511.n1 0 0.71031f **FLOATING
C288 a_44488_2511.n2 0 1.37628f **FLOATING
C289 a_44488_2511.n3 0 0.44756f **FLOATING
C290 a_44488_2511.t2 0 0.2004f **FLOATING
C291 a_44488_2511.n4 0 0.28337f **FLOATING
C292 a_44488_2511.n5 0 0.16202f **FLOATING
C293 a_44488_2511.t0 0 0.04533f **FLOATING
C294 a_41406_1605.t5 0 0.1705f **FLOATING
C295 a_41406_1605.t4 0 0.0762f **FLOATING
C296 a_41406_1605.n0 0 0.22588f **FLOATING
C297 a_41406_1605.t3 0 0.21101f **FLOATING
C298 a_41406_1605.t2 0 0.21992f **FLOATING
C299 a_41406_1605.n1 0 0.54012f **FLOATING
C300 a_41406_1605.n2 0 0.15481f **FLOATING
C301 a_41406_1605.t1 0 0.0488f **FLOATING
C302 a_41406_1605.n3 0 0.29156f **FLOATING
C303 a_41406_1605.t0 0 0.06122f **FLOATING
C304 a_35016_2511.t1 0 0.04533f **FLOATING
C305 a_35016_2511.t3 0 0.07236f **FLOATING
C306 a_35016_2511.t5 0 0.13696f **FLOATING
C307 a_35016_2511.t7 0 0.07281f **FLOATING
C308 a_35016_2511.n0 0 0.23752f **FLOATING
C309 a_35016_2511.t6 0 0.13638f **FLOATING
C310 a_35016_2511.t4 0 0.07339f **FLOATING
C311 a_35016_2511.n1 0 0.71031f **FLOATING
C312 a_35016_2511.n2 0 1.37628f **FLOATING
C313 a_35016_2511.n3 0 0.44756f **FLOATING
C314 a_35016_2511.t2 0 0.2004f **FLOATING
C315 a_35016_2511.n4 0 0.28337f **FLOATING
C316 a_35016_2511.n5 0 0.16202f **FLOATING
C317 a_35016_2511.t0 0 0.04533f **FLOATING
C318 a_10762_3500.t5 0 0.16597f **FLOATING
C319 a_10762_3500.t4 0 0.07418f **FLOATING
C320 a_10762_3500.n0 0 0.21988f **FLOATING
C321 a_10762_3500.t2 0 0.15085f **FLOATING
C322 a_10762_3500.t3 0 0.19431f **FLOATING
C323 a_10762_3500.n1 0 0.96775f **FLOATING
C324 a_10762_3500.n2 0 0.13352f **FLOATING
C325 a_10762_3500.t0 0 0.0475f **FLOATING
C326 a_10762_3500.n3 0 0.15708f **FLOATING
C327 a_10762_3500.t1 0 0.08896f **FLOATING
C328 a_1290_1160.t5 0 0.15843f **FLOATING
C329 a_1290_1160.t4 0 0.07081f **FLOATING
C330 a_1290_1160.n0 0 0.20989f **FLOATING
C331 a_1290_1160.t3 0 0.08492f **FLOATING
C332 a_1290_1160.t2 0 0.04534f **FLOATING
C333 a_1290_1160.n1 0 0.14994f **FLOATING
C334 a_1290_1160.n2 0 0.12745f **FLOATING
C335 a_1290_1160.t1 0 0.144f **FLOATING
C336 a_1290_1160.n3 0 0.92376f **FLOATING
C337 a_1290_1160.t0 0 0.18548f **FLOATING
C338 a_25464_3764.t1 0 0.04005f **FLOATING
C339 a_25464_3764.t2 0 0.06394f **FLOATING
C340 a_25464_3764.t4 0 0.12051f **FLOATING
C341 a_25464_3764.t8 0 0.06484f **FLOATING
C342 a_25464_3764.n0 0 0.20809f **FLOATING
C343 a_25464_3764.t5 0 0.12102f **FLOATING
C344 a_25464_3764.t7 0 0.06433f **FLOATING
C345 a_25464_3764.n1 0 0.50381f **FLOATING
C346 a_25464_3764.t6 0 0.12008f **FLOATING
C347 a_25464_3764.t9 0 0.06549f **FLOATING
C348 a_25464_3764.n2 0 0.48367f **FLOATING
C349 a_25464_3764.n3 0 0.84489f **FLOATING
C350 a_25464_3764.n4 0 0.19941f **FLOATING
C351 a_25464_3764.n5 0 0.18919f **FLOATING
C352 a_25464_3764.t3 0 0.17708f **FLOATING
C353 a_25464_3764.n6 0 0.25039f **FLOATING
C354 a_25464_3764.n7 0 0.14316f **FLOATING
C355 a_25464_3764.t0 0 0.04005f **FLOATING
C356 a_29706_1161.t4 0 0.15843f **FLOATING
C357 a_29706_1161.t5 0 0.07081f **FLOATING
C358 a_29706_1161.n0 0 0.20989f **FLOATING
C359 a_29706_1161.t2 0 0.08492f **FLOATING
C360 a_29706_1161.t1 0 0.04534f **FLOATING
C361 a_29706_1161.n1 0 0.14994f **FLOATING
C362 a_29706_1161.n2 0 0.12745f **FLOATING
C363 a_29706_1161.t3 0 0.144f **FLOATING
C364 a_29706_1161.n3 0 0.92376f **FLOATING
C365 a_29706_1161.t0 0 0.18548f **FLOATING
C366 a_20234_1161.t4 0 0.15843f **FLOATING
C367 a_20234_1161.t5 0 0.07081f **FLOATING
C368 a_20234_1161.n0 0 0.20989f **FLOATING
C369 a_20234_1161.t3 0 0.08492f **FLOATING
C370 a_20234_1161.t2 0 0.04534f **FLOATING
C371 a_20234_1161.n1 0 0.14994f **FLOATING
C372 a_20234_1161.n2 0 0.12745f **FLOATING
C373 a_20234_1161.t1 0 0.144f **FLOATING
C374 a_20234_1161.n3 0 0.92376f **FLOATING
C375 a_20234_1161.t0 0 0.18548f **FLOATING
C376 a_44408_3764.t1 0 0.04005f **FLOATING
C377 a_44408_3764.t2 0 0.06394f **FLOATING
C378 a_44408_3764.t5 0 0.12051f **FLOATING
C379 a_44408_3764.t9 0 0.06484f **FLOATING
C380 a_44408_3764.n0 0 0.20809f **FLOATING
C381 a_44408_3764.t6 0 0.12102f **FLOATING
C382 a_44408_3764.t8 0 0.06433f **FLOATING
C383 a_44408_3764.n1 0 0.50381f **FLOATING
C384 a_44408_3764.t4 0 0.12008f **FLOATING
C385 a_44408_3764.t7 0 0.06549f **FLOATING
C386 a_44408_3764.n2 0 0.48367f **FLOATING
C387 a_44408_3764.n3 0 0.84489f **FLOATING
C388 a_44408_3764.n4 0 0.19941f **FLOATING
C389 a_44408_3764.n5 0 0.18919f **FLOATING
C390 a_44408_3764.t3 0 0.17708f **FLOATING
C391 a_44408_3764.n6 0 0.25039f **FLOATING
C392 a_44408_3764.n7 0 0.14316f **FLOATING
C393 a_44408_3764.t0 0 0.04005f **FLOATING
C394 2inmux_0.OUT.t2 0 0.27468f **FLOATING
C395 2inmux_0.OUT.t3 0 0.14601f **FLOATING
C396 2inmux_0.OUT.n0 0 0.52483f **FLOATING
C397 dffrs_0.d 0 0.51316f **FLOATING
C398 2inmux_0.OUT.t0 0 0.3775f **FLOATING
C399 2inmux_0.OUT.t1 0 0.1155f **FLOATING
C400 2inmux_0.OUT.n1 0 0.62644f **FLOATING
C401 2inmux_0.OUT 0 0.12188f **FLOATING
C402 a_3518_1604.t5 0 0.1705f **FLOATING
C403 a_3518_1604.t4 0 0.0762f **FLOATING
C404 a_3518_1604.n0 0 0.22588f **FLOATING
C405 a_3518_1604.t3 0 0.06122f **FLOATING
C406 a_3518_1604.t2 0 0.0488f **FLOATING
C407 a_3518_1604.n1 0 0.29156f **FLOATING
C408 a_3518_1604.n2 0 0.15481f **FLOATING
C409 a_3518_1604.t0 0 0.21101f **FLOATING
C410 a_3518_1604.n3 0 0.54012f **FLOATING
C411 a_3518_1604.t1 0 0.21992f **FLOATING
C412 a_34936_3764.t1 0 0.04005f **FLOATING
C413 a_34936_3764.t2 0 0.06394f **FLOATING
C414 a_34936_3764.t6 0 0.12051f **FLOATING
C415 a_34936_3764.t9 0 0.06484f **FLOATING
C416 a_34936_3764.n0 0 0.20809f **FLOATING
C417 a_34936_3764.t8 0 0.12102f **FLOATING
C418 a_34936_3764.t5 0 0.06433f **FLOATING
C419 a_34936_3764.n1 0 0.50381f **FLOATING
C420 a_34936_3764.t7 0 0.12008f **FLOATING
C421 a_34936_3764.t4 0 0.06549f **FLOATING
C422 a_34936_3764.n2 0 0.48367f **FLOATING
C423 a_34936_3764.n3 0 0.84489f **FLOATING
C424 a_34936_3764.n4 0 0.19941f **FLOATING
C425 a_34936_3764.n5 0 0.18919f **FLOATING
C426 a_34936_3764.t3 0 0.17708f **FLOATING
C427 a_34936_3764.n6 0 0.25039f **FLOATING
C428 a_34936_3764.n7 0 0.14316f **FLOATING
C429 a_34936_3764.t0 0 0.04005f **FLOATING
C430 a_34936_1559.t1 0 0.06293f **FLOATING
C431 a_34936_1559.t2 0 0.10047f **FLOATING
C432 a_34936_1559.t5 0 0.18936f **FLOATING
C433 a_34936_1559.t7 0 0.10189f **FLOATING
C434 a_34936_1559.n0 0 0.33658f **FLOATING
C435 a_34936_1559.t6 0 0.18869f **FLOATING
C436 a_34936_1559.t4 0 0.1029f **FLOATING
C437 a_34936_1559.n1 0 0.87879f **FLOATING
C438 a_34936_1559.n2 0 0.78698f **FLOATING
C439 a_34936_1559.n3 0 0.29183f **FLOATING
C440 a_34936_1559.t3 0 0.27825f **FLOATING
C441 a_34936_1559.n4 0 0.39345f **FLOATING
C442 a_34936_1559.n5 0 0.22496f **FLOATING
C443 a_34936_1559.t0 0 0.06293f **FLOATING
C444 a_22462_1605.t5 0 0.1705f **FLOATING
C445 a_22462_1605.t4 0 0.0762f **FLOATING
C446 a_22462_1605.n0 0 0.22588f **FLOATING
C447 a_22462_1605.t3 0 0.06122f **FLOATING
C448 a_22462_1605.t2 0 0.0488f **FLOATING
C449 a_22462_1605.n1 0 0.29156f **FLOATING
C450 a_22462_1605.n2 0 0.15481f **FLOATING
C451 a_22462_1605.t0 0 0.21992f **FLOATING
C452 a_22462_1605.n3 0 0.54012f **FLOATING
C453 a_22462_1605.t1 0 0.21101f **FLOATING
C454 2inmux_1.OUT.t2 0 0.27468f **FLOATING
C455 2inmux_1.OUT.t3 0 0.14601f **FLOATING
C456 2inmux_1.OUT.n0 0 0.52483f **FLOATING
C457 dffrs_5.d 0 0.51316f **FLOATING
C458 2inmux_1.OUT.t0 0 0.3775f **FLOATING
C459 2inmux_1.OUT.t1 0 0.1155f **FLOATING
C460 2inmux_1.OUT.n1 0 0.62644f **FLOATING
C461 2inmux_1.OUT 0 0.12188f **FLOATING
C462 a_50878_1605.t5 0 0.1705f **FLOATING
C463 a_50878_1605.t4 0 0.0762f **FLOATING
C464 a_50878_1605.n0 0 0.22588f **FLOATING
C465 a_50878_1605.t3 0 0.06122f **FLOATING
C466 a_50878_1605.t2 0 0.0488f **FLOATING
C467 a_50878_1605.n1 0 0.29156f **FLOATING
C468 a_50878_1605.n2 0 0.15481f **FLOATING
C469 a_50878_1605.t0 0 0.21101f **FLOATING
C470 a_50878_1605.n3 0 0.54012f **FLOATING
C471 a_50878_1605.t1 0 0.21992f **FLOATING
C472 a_48650_1161.t5 0 0.15843f **FLOATING
C473 a_48650_1161.t4 0 0.07081f **FLOATING
C474 a_48650_1161.n0 0 0.20989f **FLOATING
C475 a_48650_1161.t1 0 0.08492f **FLOATING
C476 a_48650_1161.t3 0 0.04534f **FLOATING
C477 a_48650_1161.n1 0 0.14994f **FLOATING
C478 a_48650_1161.n2 0 0.12745f **FLOATING
C479 a_48650_1161.t2 0 0.144f **FLOATING
C480 a_48650_1161.n3 0 0.92376f **FLOATING
C481 a_48650_1161.t0 0 0.18548f **FLOATING
C482 dffrs_2.Q.t7 0 0.14856f **FLOATING
C483 dffrs_2.Q.t4 0 0.06654f **FLOATING
C484 dffrs_2.Q.t6 0 0.06601f **FLOATING
C485 dffrs_2.Q.n0 0 0.10908f **FLOATING
C486 dffrs_2.Q.n1 0 0.1562f **FLOATING
C487 2inmux_4.Bit 0 0.00243f **FLOATING
C488 dffrs_2.Q.n2 0 0.46007f **FLOATING
C489 dffrs_2.Q.t8 0 0.1058f **FLOATING
C490 dffrs_2.Q.t5 0 0.0577f **FLOATING
C491 dffrs_2.Q.n3 0 0.41081f **FLOATING
C492 dffrs_2.Q.t3 0 0.03529f **FLOATING
C493 dffrs_2.Q.t2 0 0.03529f **FLOATING
C494 dffrs_2.Q.n4 0 0.12614f **FLOATING
C495 dffrs_2.Q.t0 0 0.15602f **FLOATING
C496 dffrs_2.Q.n5 0 0.22061f **FLOATING
C497 dffrs_2.Q.t1 0 0.05633f **FLOATING
C498 dffrs_2.Q.n6 0 0.18958f **FLOATING
C499 dffrs_2.Q.n7 0 0.39693f **FLOATING
C500 dffrs_2.Q 0 0.30061f **FLOATING
C501 a_39178_3501.t5 0 0.16597f **FLOATING
C502 a_39178_3501.t4 0 0.07418f **FLOATING
C503 a_39178_3501.n0 0 0.21988f **FLOATING
C504 a_39178_3501.t2 0 0.08896f **FLOATING
C505 a_39178_3501.t1 0 0.0475f **FLOATING
C506 a_39178_3501.n1 0 0.15708f **FLOATING
C507 a_39178_3501.n2 0 0.13352f **FLOATING
C508 a_39178_3501.t3 0 0.19431f **FLOATING
C509 a_39178_3501.n3 0 0.96775f **FLOATING
C510 a_39178_3501.t0 0 0.15085f **FLOATING
C511 load.t9 0 0.04173f **FLOATING
C512 load.t25 0 0.01863f **FLOATING
C513 load.t8 0 0.01849f **FLOATING
C514 load.n0 0 0.02486f **FLOATING
C515 load.n1 0 0.06282f **FLOATING
C516 load.t3 0 0.04166f **FLOATING
C517 load.t24 0 0.01862f **FLOATING
C518 load.n2 0 0.05528f **FLOATING
C519 load 0 0.01238f **FLOATING
C520 load.t17 0 0.04173f **FLOATING
C521 load.t2 0 0.01863f **FLOATING
C522 load.t15 0 0.01849f **FLOATING
C523 load.n3 0 0.02486f **FLOATING
C524 load.n4 0 0.06282f **FLOATING
C525 2inmux_0.Load 0 0.00298f **FLOATING
C526 load.n5 0 0.10183f **FLOATING
C527 load.t20 0 0.04166f **FLOATING
C528 load.t12 0 0.01862f **FLOATING
C529 load.n6 0 0.0554f **FLOATING
C530 load.n7 0 0.12541f **FLOATING
C531 load.n8 0 0.46572f **FLOATING
C532 load.t23 0 0.04173f **FLOATING
C533 load.t5 0 0.01863f **FLOATING
C534 load.t21 0 0.01849f **FLOATING
C535 load.n9 0 0.02486f **FLOATING
C536 load.n10 0 0.06282f **FLOATING
C537 2inmux_2.Load 0 0.00298f **FLOATING
C538 load.n11 0 0.1024f **FLOATING
C539 load.t19 0 0.04166f **FLOATING
C540 load.t11 0 0.01862f **FLOATING
C541 load.n12 0 0.05528f **FLOATING
C542 load.n13 0 0.1239f **FLOATING
C543 load.n14 0 0.87684f **FLOATING
C544 load.t28 0 0.04173f **FLOATING
C545 load.t4 0 0.01863f **FLOATING
C546 load.t27 0 0.01849f **FLOATING
C547 load.n15 0 0.02486f **FLOATING
C548 load.n16 0 0.06282f **FLOATING
C549 2inmux_3.Load 0 0.00298f **FLOATING
C550 load.n17 0 0.10183f **FLOATING
C551 load.t14 0 0.04166f **FLOATING
C552 load.t6 0 0.01862f **FLOATING
C553 load.n18 0 0.0554f **FLOATING
C554 load.n19 0 0.12391f **FLOATING
C555 load.n20 0 0.87477f **FLOATING
C556 load.t13 0 0.04173f **FLOATING
C557 load.t18 0 0.01863f **FLOATING
C558 load.t10 0 0.01849f **FLOATING
C559 load.n21 0 0.02486f **FLOATING
C560 load.n22 0 0.06282f **FLOATING
C561 2inmux_4.Load 0 0.00298f **FLOATING
C562 load.n23 0 0.1024f **FLOATING
C563 load.t1 0 0.04166f **FLOATING
C564 load.t22 0 0.01862f **FLOATING
C565 load.n24 0 0.05528f **FLOATING
C566 load.n25 0 0.1239f **FLOATING
C567 load.n26 0 0.87433f **FLOATING
C568 load.t0 0 0.04173f **FLOATING
C569 load.t7 0 0.01863f **FLOATING
C570 load.t29 0 0.01849f **FLOATING
C571 load.n27 0 0.02486f **FLOATING
C572 load.n28 0 0.06282f **FLOATING
C573 2inmux_5.Load 0 0.00298f **FLOATING
C574 load.n29 0 0.1024f **FLOATING
C575 load.t26 0 0.04166f **FLOATING
C576 load.t16 0 0.01862f **FLOATING
C577 load.n30 0 0.05528f **FLOATING
C578 load.n31 0 0.1239f **FLOATING
C579 load.n32 0 1.11686f **FLOATING
C580 load.n33 0 0.33428f **FLOATING
C581 load.n34 0 0.1024f **FLOATING
C582 2inmux_1.Load 0 0.00298f **FLOATING
C583 a_15992_5968.t1 0 0.0891f **FLOATING
C584 a_15992_5968.t5 0 0.16734f **FLOATING
C585 a_15992_5968.t4 0 0.09125f **FLOATING
C586 a_15992_5968.n0 0 0.88217f **FLOATING
C587 a_15992_5968.n1 0 0.66334f **FLOATING
C588 a_15992_5968.t3 0 0.05581f **FLOATING
C589 a_15992_5968.t2 0 0.05581f **FLOATING
C590 a_15992_5968.n2 0 0.1995f **FLOATING
C591 a_15992_5968.n3 0 0.34892f **FLOATING
C592 a_15992_5968.t0 0 0.24676f **FLOATING
C593 2inmux_1.Bit.t7 0 0.14856f **FLOATING
C594 2inmux_1.Bit.t4 0 0.06654f **FLOATING
C595 2inmux_1.Bit.t6 0 0.06601f **FLOATING
C596 2inmux_1.Bit.n0 0 0.10908f **FLOATING
C597 2inmux_1.Bit.n1 0 0.1562f **FLOATING
C598 2inmux_1.Bit 0 0.00243f **FLOATING
C599 2inmux_1.Bit.n2 0 0.46007f **FLOATING
C600 2inmux_1.Bit.t8 0 0.1058f **FLOATING
C601 2inmux_1.Bit.t5 0 0.0577f **FLOATING
C602 2inmux_1.Bit.n3 0 0.41081f **FLOATING
C603 2inmux_1.Bit.t3 0 0.03529f **FLOATING
C604 2inmux_1.Bit.t2 0 0.03529f **FLOATING
C605 2inmux_1.Bit.n4 0 0.12614f **FLOATING
C606 2inmux_1.Bit.t0 0 0.15602f **FLOATING
C607 2inmux_1.Bit.n5 0 0.22061f **FLOATING
C608 2inmux_1.Bit.t1 0 0.05633f **FLOATING
C609 2inmux_1.Bit.n6 0 0.18958f **FLOATING
C610 2inmux_1.Bit.n7 0 0.39693f **FLOATING
C611 dffrs_4.Q 0 0.30061f **FLOATING
C612 a_15992_3763.t1 0 0.04005f **FLOATING
C613 a_15992_3763.t3 0 0.06394f **FLOATING
C614 a_15992_3763.t5 0 0.12051f **FLOATING
C615 a_15992_3763.t8 0 0.06484f **FLOATING
C616 a_15992_3763.n0 0 0.20809f **FLOATING
C617 a_15992_3763.t7 0 0.12102f **FLOATING
C618 a_15992_3763.t4 0 0.06433f **FLOATING
C619 a_15992_3763.n1 0 0.50381f **FLOATING
C620 a_15992_3763.t6 0 0.12008f **FLOATING
C621 a_15992_3763.t9 0 0.06549f **FLOATING
C622 a_15992_3763.n2 0 0.48367f **FLOATING
C623 a_15992_3763.n3 0 0.84489f **FLOATING
C624 a_15992_3763.n4 0 0.19941f **FLOATING
C625 a_15992_3763.n5 0 0.18919f **FLOATING
C626 a_15992_3763.t2 0 0.17708f **FLOATING
C627 a_15992_3763.n6 0 0.25039f **FLOATING
C628 a_15992_3763.n7 0 0.14316f **FLOATING
C629 a_15992_3763.t0 0 0.04005f **FLOATING
C630 clk.t17 0 0.07668f **FLOATING
C631 clk.t6 0 0.04076f **FLOATING
C632 clk.n0 0 0.15813f **FLOATING
C633 clk.t10 0 0.07635f **FLOATING
C634 clk.t21 0 0.04108f **FLOATING
C635 clk.n1 0 0.1701f **FLOATING
C636 clk.n2 0 0.35106f **FLOATING
C637 clk 0 0.14314f **FLOATING
C638 clk.t18 0 0.07668f **FLOATING
C639 clk.t7 0 0.04076f **FLOATING
C640 clk.n3 0 0.15813f **FLOATING
C641 clk.t2 0 0.07635f **FLOATING
C642 clk.t13 0 0.04108f **FLOATING
C643 clk.n4 0 0.1701f **FLOATING
C644 clk.n5 0 0.35106f **FLOATING
C645 dffrs_0.clk 0 0.05372f **FLOATING
C646 clk.n6 0 0.71832f **FLOATING
C647 clk.t12 0 0.07668f **FLOATING
C648 clk.t0 0 0.04076f **FLOATING
C649 clk.n7 0 0.15813f **FLOATING
C650 clk.t22 0 0.07635f **FLOATING
C651 clk.t9 0 0.04108f **FLOATING
C652 clk.n8 0 0.1701f **FLOATING
C653 clk.n9 0 0.35106f **FLOATING
C654 dffrs_1.clk 0 0.05372f **FLOATING
C655 clk.n10 0 1.13795f **FLOATING
C656 clk.t1 0 0.07668f **FLOATING
C657 clk.t14 0 0.04076f **FLOATING
C658 clk.n11 0 0.15813f **FLOATING
C659 clk.t11 0 0.07635f **FLOATING
C660 clk.t23 0 0.04108f **FLOATING
C661 clk.n12 0 0.1701f **FLOATING
C662 clk.n13 0 0.35106f **FLOATING
C663 dffrs_2.clk 0 0.05372f **FLOATING
C664 clk.n14 0 1.13815f **FLOATING
C665 clk.t15 0 0.07668f **FLOATING
C666 clk.t4 0 0.04076f **FLOATING
C667 clk.n15 0 0.15813f **FLOATING
C668 clk.t8 0 0.07635f **FLOATING
C669 clk.t19 0 0.04108f **FLOATING
C670 clk.n16 0 0.1701f **FLOATING
C671 clk.n17 0 0.35106f **FLOATING
C672 dffrs_3.clk 0 0.05372f **FLOATING
C673 clk.n18 0 1.13813f **FLOATING
C674 clk.t3 0 0.07668f **FLOATING
C675 clk.t16 0 0.04076f **FLOATING
C676 clk.n19 0 0.15813f **FLOATING
C677 clk.t20 0 0.07635f **FLOATING
C678 clk.t5 0 0.04108f **FLOATING
C679 clk.n20 0 0.1701f **FLOATING
C680 clk.n21 0 0.35106f **FLOATING
C681 dffrs_4.clk 0 0.05372f **FLOATING
C682 clk.n22 0 1.36908f **FLOATING
C683 dffrs_5.clk 0 0.40161f **FLOATING
C684 a_1290_3500.t4 0 0.15843f **FLOATING
C685 a_1290_3500.t5 0 0.07081f **FLOATING
C686 a_1290_3500.n0 0 0.20989f **FLOATING
C687 a_1290_3500.t2 0 0.144f **FLOATING
C688 a_1290_3500.t1 0 0.18548f **FLOATING
C689 a_1290_3500.n1 0 0.92376f **FLOATING
C690 a_1290_3500.n2 0 0.12745f **FLOATING
C691 a_1290_3500.t3 0 0.08492f **FLOATING
C692 a_1290_3500.n3 0 0.14994f **FLOATING
C693 a_1290_3500.t0 0 0.04534f **FLOATING
C694 2inmux_2.Bit.t5 0 0.14856f **FLOATING
C695 2inmux_2.Bit.t7 0 0.06654f **FLOATING
C696 2inmux_2.Bit.t4 0 0.06601f **FLOATING
C697 2inmux_2.Bit.n0 0 0.10908f **FLOATING
C698 2inmux_2.Bit.n1 0 0.1562f **FLOATING
C699 2inmux_2.Bit 0 0.00243f **FLOATING
C700 2inmux_2.Bit.n2 0 0.46007f **FLOATING
C701 2inmux_2.Bit.t6 0 0.1058f **FLOATING
C702 2inmux_2.Bit.t8 0 0.0577f **FLOATING
C703 2inmux_2.Bit.n3 0 0.41081f **FLOATING
C704 2inmux_2.Bit.t3 0 0.03529f **FLOATING
C705 2inmux_2.Bit.t0 0 0.03529f **FLOATING
C706 2inmux_2.Bit.n4 0 0.12614f **FLOATING
C707 2inmux_2.Bit.t1 0 0.15602f **FLOATING
C708 2inmux_2.Bit.n5 0 0.22061f **FLOATING
C709 2inmux_2.Bit.t2 0 0.05633f **FLOATING
C710 2inmux_2.Bit.n6 0 0.18958f **FLOATING
C711 2inmux_2.Bit.n7 0 0.39693f **FLOATING
C712 dffrs_0.Q 0 0.30061f **FLOATING
C713 a_20234_3501.t5 0 0.16597f **FLOATING
C714 a_20234_3501.t4 0 0.07418f **FLOATING
C715 a_20234_3501.n0 0 0.21988f **FLOATING
C716 a_20234_3501.t3 0 0.15085f **FLOATING
C717 a_20234_3501.t2 0 0.19431f **FLOATING
C718 a_20234_3501.n1 0 0.96775f **FLOATING
C719 a_20234_3501.n2 0 0.13352f **FLOATING
C720 a_20234_3501.t1 0 0.08896f **FLOATING
C721 a_20234_3501.n3 0 0.15708f **FLOATING
C722 a_20234_3501.t0 0 0.0475f **FLOATING
C723 dffrs_1.Q.t4 0 0.14858f **FLOATING
C724 dffrs_1.Q.t6 0 0.06654f **FLOATING
C725 dffrs_1.Q.t8 0 0.06602f **FLOATING
C726 dffrs_1.Q.n0 0 0.10909f **FLOATING
C727 dffrs_1.Q.n1 0 0.15622f **FLOATING
C728 2inmux_3.Bit 0 0.00243f **FLOATING
C729 dffrs_1.Q.n2 0 0.45988f **FLOATING
C730 dffrs_1.Q.t7 0 0.10581f **FLOATING
C731 dffrs_1.Q.t5 0 0.0577f **FLOATING
C732 dffrs_1.Q.n3 0 0.41085f **FLOATING
C733 dffrs_1.Q.t1 0 0.03529f **FLOATING
C734 dffrs_1.Q.t0 0 0.03529f **FLOATING
C735 dffrs_1.Q.n4 0 0.12615f **FLOATING
C736 dffrs_1.Q.t2 0 0.15603f **FLOATING
C737 dffrs_1.Q.n5 0 0.22063f **FLOATING
C738 dffrs_1.Q.t3 0 0.05634f **FLOATING
C739 dffrs_1.Q.n6 0 0.18959f **FLOATING
C740 dffrs_1.Q.n7 0 0.39697f **FLOATING
C741 dffrs_1.Q 0 0.30057f **FLOATING
C742 a_6520_3763.t2 0 0.04005f **FLOATING
C743 a_6520_3763.t3 0 0.06394f **FLOATING
C744 a_6520_3763.t5 0 0.12051f **FLOATING
C745 a_6520_3763.t8 0 0.06484f **FLOATING
C746 a_6520_3763.n0 0 0.20809f **FLOATING
C747 a_6520_3763.t9 0 0.12102f **FLOATING
C748 a_6520_3763.t6 0 0.06433f **FLOATING
C749 a_6520_3763.n1 0 0.50381f **FLOATING
C750 a_6520_3763.t4 0 0.12008f **FLOATING
C751 a_6520_3763.t7 0 0.06549f **FLOATING
C752 a_6520_3763.n2 0 0.48367f **FLOATING
C753 a_6520_3763.n3 0 0.84489f **FLOATING
C754 a_6520_3763.n4 0 0.19941f **FLOATING
C755 a_6520_3763.n5 0 0.18919f **FLOATING
C756 a_6520_3763.t1 0 0.17708f **FLOATING
C757 a_6520_3763.n6 0 0.25039f **FLOATING
C758 a_6520_3763.n7 0 0.14316f **FLOATING
C759 a_6520_3763.t0 0 0.04005f **FLOATING
C760 a_6600_2510.t2 0 0.04533f **FLOATING
C761 a_6600_2510.t1 0 0.07236f **FLOATING
C762 a_6600_2510.t4 0 0.13696f **FLOATING
C763 a_6600_2510.t6 0 0.07281f **FLOATING
C764 a_6600_2510.n0 0 0.23752f **FLOATING
C765 a_6600_2510.t5 0 0.13638f **FLOATING
C766 a_6600_2510.t7 0 0.07339f **FLOATING
C767 a_6600_2510.n1 0 0.71031f **FLOATING
C768 a_6600_2510.n2 0 1.37628f **FLOATING
C769 a_6600_2510.n3 0 0.44756f **FLOATING
C770 a_6600_2510.t3 0 0.2004f **FLOATING
C771 a_6600_2510.n4 0 0.28337f **FLOATING
C772 a_6600_2510.n5 0 0.16202f **FLOATING
C773 a_6600_2510.t0 0 0.04533f **FLOATING
C774 a_6520_1558.t3 0 0.06293f **FLOATING
C775 a_6520_1558.t2 0 0.06293f **FLOATING
C776 a_6520_1558.n0 0 0.22496f **FLOATING
C777 a_6520_1558.t1 0 0.27825f **FLOATING
C778 a_6520_1558.n1 0 0.39345f **FLOATING
C779 a_6520_1558.t5 0 0.18936f **FLOATING
C780 a_6520_1558.t7 0 0.10189f **FLOATING
C781 a_6520_1558.n2 0 0.33658f **FLOATING
C782 a_6520_1558.t4 0 0.18869f **FLOATING
C783 a_6520_1558.t6 0 0.1029f **FLOATING
C784 a_6520_1558.n3 0 0.87879f **FLOATING
C785 a_6520_1558.n4 0 0.78698f **FLOATING
C786 a_6520_1558.n5 0 0.29183f **FLOATING
C787 a_6520_1558.t0 0 0.10047f **FLOATING
C788 a_48650_3501.t4 0 0.16597f **FLOATING
C789 a_48650_3501.t5 0 0.07418f **FLOATING
C790 a_48650_3501.n0 0 0.21988f **FLOATING
C791 a_48650_3501.t3 0 0.15085f **FLOATING
C792 a_48650_3501.t1 0 0.19431f **FLOATING
C793 a_48650_3501.n1 0 0.96775f **FLOATING
C794 a_48650_3501.n2 0 0.13352f **FLOATING
C795 a_48650_3501.t2 0 0.0475f **FLOATING
C796 a_48650_3501.n3 0 0.15708f **FLOATING
C797 a_48650_3501.t0 0 0.08896f **FLOATING
C798 avdd.t86 0 0.01935f **FLOATING
C799 avdd.t407 0 0.01055f **FLOATING
C800 avdd.n0 0 0.09149f **FLOATING
C801 avdd.t92 0 0.01935f **FLOATING
C802 avdd.t404 0 0.01055f **FLOATING
C803 avdd.n1 0 0.03208f **FLOATING
C804 avdd.n2 0 0.13216f **FLOATING
C805 avdd.t29 0 0.00645f **FLOATING
C806 avdd.t15 0 0.00645f **FLOATING
C807 avdd.n3 0 0.02312f **FLOATING
C808 avdd.n4 0 0.14951f **FLOATING
C809 avdd.t28 0 0.09482f **FLOATING
C810 avdd.t14 0 0.08403f **FLOATING
C811 avdd.t93 0 0.09482f **FLOATING
C812 avdd.n5 0 0.13889f **FLOATING
C813 avdd.t94 0 0.01613f **FLOATING
C814 avdd.n6 0 0.03079f **FLOATING
C815 avdd.n7 0 0.06566f **FLOATING
C816 avdd.t301 0 0.00645f **FLOATING
C817 avdd.t309 0 0.00645f **FLOATING
C818 avdd.n8 0 0.02312f **FLOATING
C819 avdd.n9 0 0.14951f **FLOATING
C820 avdd.t300 0 0.09482f **FLOATING
C821 avdd.t308 0 0.08403f **FLOATING
C822 avdd.t87 0 0.09482f **FLOATING
C823 avdd.n10 0 0.13889f **FLOATING
C824 avdd.t88 0 0.01613f **FLOATING
C825 avdd.n11 0 0.03079f **FLOATING
C826 avdd.n12 0 0.06443f **FLOATING
C827 avdd.t217 0 0.01909f **FLOATING
C828 avdd.n13 0 0.08303f **FLOATING
C829 avdd.t137 0 0.01909f **FLOATING
C830 avdd.t136 0 0.14751f **FLOATING
C831 avdd.n14 0 0.32056f **FLOATING
C832 avdd.t339 0 0.01861f **FLOATING
C833 avdd.n15 0 0.0584f **FLOATING
C834 avdd.t35 0 0.01861f **FLOATING
C835 avdd.n16 0 0.0584f **FLOATING
C836 avdd.t37 0 0.01861f **FLOATING
C837 avdd.n17 0 0.0584f **FLOATING
C838 avdd.t229 0 0.01861f **FLOATING
C839 avdd.n18 0 0.0584f **FLOATING
C840 avdd.n19 0 0.03619f **FLOATING
C841 avdd.n20 0 0.03619f **FLOATING
C842 avdd.t36 0 0.1124f **FLOATING
C843 avdd.n21 0 0.03973f **FLOATING
C844 avdd.t34 0 0.11271f **FLOATING
C845 avdd.n22 0 0.13168f **FLOATING
C846 avdd.n23 0 0.03973f **FLOATING
C847 avdd.n24 0 0.0148f **FLOATING
C848 avdd.n25 0 0.12152f **FLOATING
C849 avdd.t8 0 0.1124f **FLOATING
C850 avdd.t9 0 0.1124f **FLOATING
C851 avdd.n26 0 0.0148f **FLOATING
C852 avdd.n27 0 0.12152f **FLOATING
C853 avdd.t228 0 0.12182f **FLOATING
C854 avdd.n28 0 0.13388f **FLOATING
C855 avdd.t351 0 0.01909f **FLOATING
C856 avdd.n29 0 0.08303f **FLOATING
C857 avdd.t337 0 0.01909f **FLOATING
C858 avdd.t336 0 0.14751f **FLOATING
C859 avdd.n30 0 0.32056f **FLOATING
C860 avdd.t369 0 0.01861f **FLOATING
C861 avdd.n31 0 0.0584f **FLOATING
C862 avdd.t145 0 0.01861f **FLOATING
C863 avdd.n32 0 0.0584f **FLOATING
C864 avdd.t143 0 0.01861f **FLOATING
C865 avdd.n33 0 0.0584f **FLOATING
C866 avdd.t223 0 0.01861f **FLOATING
C867 avdd.n34 0 0.0584f **FLOATING
C868 avdd.n35 0 0.03619f **FLOATING
C869 avdd.n36 0 0.03619f **FLOATING
C870 avdd.t142 0 0.1124f **FLOATING
C871 avdd.n37 0 0.03973f **FLOATING
C872 avdd.t144 0 0.11271f **FLOATING
C873 avdd.n38 0 0.13168f **FLOATING
C874 avdd.n39 0 0.03973f **FLOATING
C875 avdd.n40 0 0.0148f **FLOATING
C876 avdd.n41 0 0.12152f **FLOATING
C877 avdd.t24 0 0.1124f **FLOATING
C878 avdd.t25 0 0.1124f **FLOATING
C879 avdd.n42 0 0.0148f **FLOATING
C880 avdd.n43 0 0.12152f **FLOATING
C881 avdd.t222 0 0.12182f **FLOATING
C882 avdd.n44 0 0.13388f **FLOATING
C883 avdd.t293 0 0.01909f **FLOATING
C884 avdd.n45 0 0.08303f **FLOATING
C885 avdd.t151 0 0.01909f **FLOATING
C886 avdd.t150 0 0.14751f **FLOATING
C887 avdd.n46 0 0.32056f **FLOATING
C888 avdd.t305 0 0.01861f **FLOATING
C889 avdd.n47 0 0.0584f **FLOATING
C890 avdd.t297 0 0.01861f **FLOATING
C891 avdd.n48 0 0.0584f **FLOATING
C892 avdd.t299 0 0.01861f **FLOATING
C893 avdd.n49 0 0.0584f **FLOATING
C894 avdd.t373 0 0.01861f **FLOATING
C895 avdd.n50 0 0.0584f **FLOATING
C896 avdd.n51 0 0.03619f **FLOATING
C897 avdd.n52 0 0.03619f **FLOATING
C898 avdd.t298 0 0.1124f **FLOATING
C899 avdd.n53 0 0.03973f **FLOATING
C900 avdd.t296 0 0.11271f **FLOATING
C901 avdd.n54 0 0.13168f **FLOATING
C902 avdd.n55 0 0.03973f **FLOATING
C903 avdd.n56 0 0.0148f **FLOATING
C904 avdd.n57 0 0.12152f **FLOATING
C905 avdd.t128 0 0.1124f **FLOATING
C906 avdd.t129 0 0.1124f **FLOATING
C907 avdd.n58 0 0.0148f **FLOATING
C908 avdd.n59 0 0.12152f **FLOATING
C909 avdd.t372 0 0.12182f **FLOATING
C910 avdd.n60 0 0.13388f **FLOATING
C911 avdd.t271 0 0.01909f **FLOATING
C912 avdd.n61 0 0.08303f **FLOATING
C913 avdd.t235 0 0.01909f **FLOATING
C914 avdd.t234 0 0.14751f **FLOATING
C915 avdd.n62 0 0.32056f **FLOATING
C916 avdd.t237 0 0.01861f **FLOATING
C917 avdd.n63 0 0.0584f **FLOATING
C918 avdd.t227 0 0.01861f **FLOATING
C919 avdd.n64 0 0.0584f **FLOATING
C920 avdd.t225 0 0.01861f **FLOATING
C921 avdd.n65 0 0.0584f **FLOATING
C922 avdd.t169 0 0.01861f **FLOATING
C923 avdd.n66 0 0.0584f **FLOATING
C924 avdd.n67 0 0.03619f **FLOATING
C925 avdd.n68 0 0.03619f **FLOATING
C926 avdd.t224 0 0.1124f **FLOATING
C927 avdd.n69 0 0.03973f **FLOATING
C928 avdd.t226 0 0.11271f **FLOATING
C929 avdd.n70 0 0.13168f **FLOATING
C930 avdd.n71 0 0.03973f **FLOATING
C931 avdd.n72 0 0.0148f **FLOATING
C932 avdd.n73 0 0.12152f **FLOATING
C933 avdd.t310 0 0.1124f **FLOATING
C934 avdd.t311 0 0.1124f **FLOATING
C935 avdd.n74 0 0.0148f **FLOATING
C936 avdd.n75 0 0.12152f **FLOATING
C937 avdd.t168 0 0.12182f **FLOATING
C938 avdd.n76 0 0.13388f **FLOATING
C939 avdd.t353 0 0.01909f **FLOATING
C940 avdd.n77 0 0.08303f **FLOATING
C941 avdd.t321 0 0.01909f **FLOATING
C942 avdd.t320 0 0.14751f **FLOATING
C943 avdd.n78 0 0.32056f **FLOATING
C944 avdd.t5 0 0.01861f **FLOATING
C945 avdd.n79 0 0.0584f **FLOATING
C946 avdd.t211 0 0.01861f **FLOATING
C947 avdd.n80 0 0.0584f **FLOATING
C948 avdd.t209 0 0.01861f **FLOATING
C949 avdd.n81 0 0.0584f **FLOATING
C950 avdd.t213 0 0.01861f **FLOATING
C951 avdd.n82 0 0.0584f **FLOATING
C952 avdd.n83 0 0.03619f **FLOATING
C953 avdd.n84 0 0.03619f **FLOATING
C954 avdd.t208 0 0.1124f **FLOATING
C955 avdd.n85 0 0.03973f **FLOATING
C956 avdd.t210 0 0.11271f **FLOATING
C957 avdd.n86 0 0.13168f **FLOATING
C958 avdd.n87 0 0.03973f **FLOATING
C959 avdd.n88 0 0.0148f **FLOATING
C960 avdd.n89 0 0.12152f **FLOATING
C961 avdd.t21 0 0.1124f **FLOATING
C962 avdd.t20 0 0.1124f **FLOATING
C963 avdd.n90 0 0.0148f **FLOATING
C964 avdd.n91 0 0.12152f **FLOATING
C965 avdd.t212 0 0.12182f **FLOATING
C966 avdd.n92 0 0.13388f **FLOATING
C967 avdd.t98 0 0.01935f **FLOATING
C968 avdd.t403 0 0.01055f **FLOATING
C969 avdd.n93 0 0.09149f **FLOATING
C970 avdd.t104 0 0.01935f **FLOATING
C971 avdd.t399 0 0.01055f **FLOATING
C972 avdd.n94 0 0.03208f **FLOATING
C973 avdd.n95 0 0.13216f **FLOATING
C974 dffrs_5.setb 0 0.00111f **FLOATING
C975 avdd.n96 0 0.01325f **FLOATING
C976 avdd.t193 0 0.00645f **FLOATING
C977 avdd.t189 0 0.00645f **FLOATING
C978 avdd.n97 0 0.02312f **FLOATING
C979 avdd.n98 0 0.14951f **FLOATING
C980 avdd.t192 0 0.09482f **FLOATING
C981 avdd.t188 0 0.08403f **FLOATING
C982 avdd.t105 0 0.09482f **FLOATING
C983 avdd.n99 0 0.13889f **FLOATING
C984 avdd.t106 0 0.01613f **FLOATING
C985 avdd.n100 0 0.03079f **FLOATING
C986 avdd.n101 0 0.06566f **FLOATING
C987 avdd.n102 0 2.80882f **FLOATING
C988 avdd.t139 0 0.00645f **FLOATING
C989 avdd.t191 0 0.00645f **FLOATING
C990 avdd.n103 0 0.02312f **FLOATING
C991 avdd.n104 0 0.14951f **FLOATING
C992 avdd.t138 0 0.09482f **FLOATING
C993 avdd.t190 0 0.08403f **FLOATING
C994 avdd.t99 0 0.09482f **FLOATING
C995 avdd.n105 0 0.13889f **FLOATING
C996 avdd.t100 0 0.01613f **FLOATING
C997 avdd.n106 0 0.03079f **FLOATING
C998 avdd.n107 0 0.06443f **FLOATING
C999 avdd.t131 0 0.00645f **FLOATING
C1000 avdd.t73 0 0.00645f **FLOATING
C1001 avdd.n108 0 0.02312f **FLOATING
C1002 avdd.n109 0 0.14951f **FLOATING
C1003 avdd.t130 0 0.09482f **FLOATING
C1004 avdd.t72 0 0.08403f **FLOATING
C1005 avdd.t202 0 0.09482f **FLOATING
C1006 avdd.n110 0 0.13889f **FLOATING
C1007 avdd.t203 0 0.01613f **FLOATING
C1008 avdd.n111 0 0.03079f **FLOATING
C1009 avdd.n112 0 0.06443f **FLOATING
C1010 avdd.n113 0 2.85645f **FLOATING
C1011 avdd.t58 0 0.00645f **FLOATING
C1012 avdd.t173 0 0.00645f **FLOATING
C1013 avdd.n114 0 0.02312f **FLOATING
C1014 avdd.n115 0 0.14951f **FLOATING
C1015 avdd.t57 0 0.09482f **FLOATING
C1016 avdd.t172 0 0.08403f **FLOATING
C1017 avdd.t166 0 0.09482f **FLOATING
C1018 avdd.n116 0 0.13889f **FLOATING
C1019 avdd.t167 0 0.01613f **FLOATING
C1020 avdd.n117 0 0.03079f **FLOATING
C1021 avdd.n118 0 0.06443f **FLOATING
C1022 avdd.n119 0 1.80909f **FLOATING
C1023 avdd.t197 0 0.00645f **FLOATING
C1024 avdd.t273 0 0.00645f **FLOATING
C1025 avdd.n120 0 0.02312f **FLOATING
C1026 avdd.n121 0 0.14951f **FLOATING
C1027 avdd.t196 0 0.09482f **FLOATING
C1028 avdd.t272 0 0.08403f **FLOATING
C1029 avdd.t194 0 0.09482f **FLOATING
C1030 avdd.n122 0 0.13889f **FLOATING
C1031 avdd.t195 0 0.01613f **FLOATING
C1032 avdd.n123 0 0.03079f **FLOATING
C1033 avdd.n124 0 0.06443f **FLOATING
C1034 avdd.n125 0 1.28162f **FLOATING
C1035 avdd.t56 0 0.0195f **FLOATING
C1036 avdd.t387 0 0.01037f **FLOATING
C1037 avdd.n126 0 0.08453f **FLOATING
C1038 avdd.t71 0 0.01942f **FLOATING
C1039 avdd.t381 0 0.01045f **FLOATING
C1040 avdd.n127 0 0.07805f **FLOATING
C1041 avdd.t95 0 0.01942f **FLOATING
C1042 avdd.t402 0 0.01045f **FLOATING
C1043 avdd.n128 0 0.04661f **FLOATING
C1044 avdd.n129 0 0.14749f **FLOATING
C1045 avdd.n130 0 0.11028f **FLOATING
C1046 dffrs_5.resetb 0 0.01446f **FLOATING
C1047 avdd.t149 0 0.00645f **FLOATING
C1048 avdd.t97 0 0.00645f **FLOATING
C1049 avdd.n131 0 0.02312f **FLOATING
C1050 avdd.n132 0 0.14951f **FLOATING
C1051 avdd.t148 0 0.09482f **FLOATING
C1052 avdd.t96 0 0.08403f **FLOATING
C1053 avdd.t170 0 0.09482f **FLOATING
C1054 avdd.n133 0 0.13889f **FLOATING
C1055 avdd.t171 0 0.01613f **FLOATING
C1056 avdd.n134 0 0.03079f **FLOATING
C1057 avdd.n135 0 0.06443f **FLOATING
C1058 avdd.n136 0 3.87524f **FLOATING
C1059 avdd.n137 0 2.36436f **FLOATING
C1060 avdd.n138 0 0.54101f **FLOATING
C1061 avdd.n139 0 0.22311f **FLOATING
C1062 avdd.n140 0 0.13505f **FLOATING
C1063 avdd.t279 0 0.01861f **FLOATING
C1064 avdd.n141 0 0.0584f **FLOATING
C1065 avdd.t295 0 0.01909f **FLOATING
C1066 avdd.n142 0 0.04054f **FLOATING
C1067 avdd.n143 0 0.04054f **FLOATING
C1068 avdd.t278 0 0.12182f **FLOATING
C1069 avdd.n144 0 0.0148f **FLOATING
C1070 avdd.n145 0 0.12152f **FLOATING
C1071 avdd.t294 0 0.12182f **FLOATING
C1072 avdd.n146 0 0.12417f **FLOATING
C1073 avdd.n147 0 0.08303f **FLOATING
C1074 avdd.t11 0 0.01909f **FLOATING
C1075 avdd.t10 0 0.14751f **FLOATING
C1076 avdd.n148 0 0.32056f **FLOATING
C1077 avdd.n149 0 0.11564f **FLOATING
C1078 avdd.n150 0 0.04514f **FLOATING
C1079 avdd.n151 0 0.40282f **FLOATING
C1080 avdd.n152 0 1.36009f **FLOATING
C1081 avdd.n153 0 0.32215f **FLOATING
C1082 avdd.n154 0 0.29609f **FLOATING
C1083 avdd.n155 0 0.04054f **FLOATING
C1084 avdd.n156 0 0.04054f **FLOATING
C1085 avdd.n157 0 0.12417f **FLOATING
C1086 avdd.t352 0 0.12182f **FLOATING
C1087 avdd.n158 0 0.0148f **FLOATING
C1088 avdd.n159 0 0.12152f **FLOATING
C1089 avdd.t4 0 0.12182f **FLOATING
C1090 avdd.n160 0 0.13228f **FLOATING
C1091 avdd.n161 0 0.05291f **FLOATING
C1092 avdd.n162 0 0.06202f **FLOATING
C1093 avdd.n163 0 0.22294f **FLOATING
C1094 avdd.t346 0 0.12368f **FLOATING
C1095 avdd.t347 0 0.04896f **FLOATING
C1096 avdd.n164 0 0.28487f **FLOATING
C1097 avdd.n165 0 0.71105f **FLOATING
C1098 avdd.t41 0 0.01935f **FLOATING
C1099 avdd.t386 0 0.01055f **FLOATING
C1100 avdd.n166 0 0.09149f **FLOATING
C1101 avdd.t80 0 0.01935f **FLOATING
C1102 avdd.t378 0 0.01055f **FLOATING
C1103 avdd.n167 0 0.03208f **FLOATING
C1104 avdd.n168 0 0.13216f **FLOATING
C1105 dffrs_4.setb 0 0.00111f **FLOATING
C1106 avdd.n169 0 0.01325f **FLOATING
C1107 avdd.t263 0 0.00645f **FLOATING
C1108 avdd.t187 0 0.00645f **FLOATING
C1109 avdd.n170 0 0.02312f **FLOATING
C1110 avdd.n171 0 0.14951f **FLOATING
C1111 avdd.t262 0 0.09482f **FLOATING
C1112 avdd.t186 0 0.08403f **FLOATING
C1113 avdd.t81 0 0.09482f **FLOATING
C1114 avdd.n172 0 0.13889f **FLOATING
C1115 avdd.t82 0 0.01613f **FLOATING
C1116 avdd.n173 0 0.03079f **FLOATING
C1117 avdd.n174 0 0.06566f **FLOATING
C1118 avdd.n175 0 2.80882f **FLOATING
C1119 avdd.t31 0 0.00645f **FLOATING
C1120 avdd.t261 0 0.00645f **FLOATING
C1121 avdd.n176 0 0.02312f **FLOATING
C1122 avdd.n177 0 0.14951f **FLOATING
C1123 avdd.t30 0 0.09482f **FLOATING
C1124 avdd.t260 0 0.08403f **FLOATING
C1125 avdd.t42 0 0.09482f **FLOATING
C1126 avdd.n178 0 0.13889f **FLOATING
C1127 avdd.t43 0 0.01613f **FLOATING
C1128 avdd.n179 0 0.03079f **FLOATING
C1129 avdd.n180 0 0.06443f **FLOATING
C1130 avdd.t359 0 0.00645f **FLOATING
C1131 avdd.t127 0 0.00645f **FLOATING
C1132 avdd.n181 0 0.02312f **FLOATING
C1133 avdd.n182 0 0.14951f **FLOATING
C1134 avdd.t358 0 0.09482f **FLOATING
C1135 avdd.t126 0 0.08403f **FLOATING
C1136 avdd.t158 0 0.09482f **FLOATING
C1137 avdd.n183 0 0.13889f **FLOATING
C1138 avdd.t159 0 0.01613f **FLOATING
C1139 avdd.n184 0 0.03079f **FLOATING
C1140 avdd.n185 0 0.06443f **FLOATING
C1141 avdd.n186 0 2.85645f **FLOATING
C1142 avdd.t79 0 0.00645f **FLOATING
C1143 avdd.t287 0 0.00645f **FLOATING
C1144 avdd.n187 0 0.02312f **FLOATING
C1145 avdd.n188 0 0.14951f **FLOATING
C1146 avdd.t78 0 0.09482f **FLOATING
C1147 avdd.t286 0 0.08403f **FLOATING
C1148 avdd.t322 0 0.09482f **FLOATING
C1149 avdd.n189 0 0.13889f **FLOATING
C1150 avdd.t323 0 0.01613f **FLOATING
C1151 avdd.n190 0 0.03079f **FLOATING
C1152 avdd.n191 0 0.06443f **FLOATING
C1153 avdd.n192 0 1.80909f **FLOATING
C1154 avdd.t361 0 0.00645f **FLOATING
C1155 avdd.t135 0 0.00645f **FLOATING
C1156 avdd.n193 0 0.02312f **FLOATING
C1157 avdd.n194 0 0.14951f **FLOATING
C1158 avdd.t360 0 0.09482f **FLOATING
C1159 avdd.t134 0 0.08403f **FLOATING
C1160 avdd.t258 0 0.09482f **FLOATING
C1161 avdd.n195 0 0.13889f **FLOATING
C1162 avdd.t259 0 0.01613f **FLOATING
C1163 avdd.n196 0 0.03079f **FLOATING
C1164 avdd.n197 0 0.06443f **FLOATING
C1165 avdd.n198 0 1.28162f **FLOATING
C1166 avdd.t77 0 0.0195f **FLOATING
C1167 avdd.t379 0 0.01037f **FLOATING
C1168 avdd.n199 0 0.08453f **FLOATING
C1169 avdd.t125 0 0.01942f **FLOATING
C1170 avdd.t394 0 0.01045f **FLOATING
C1171 avdd.n200 0 0.07805f **FLOATING
C1172 avdd.t59 0 0.01942f **FLOATING
C1173 avdd.t384 0 0.01045f **FLOATING
C1174 avdd.n201 0 0.04661f **FLOATING
C1175 avdd.n202 0 0.14749f **FLOATING
C1176 avdd.n203 0 0.11028f **FLOATING
C1177 dffrs_4.resetb 0 0.01446f **FLOATING
C1178 avdd.t199 0 0.00645f **FLOATING
C1179 avdd.t61 0 0.00645f **FLOATING
C1180 avdd.n204 0 0.02312f **FLOATING
C1181 avdd.n205 0 0.14951f **FLOATING
C1182 avdd.t198 0 0.09482f **FLOATING
C1183 avdd.t60 0 0.08403f **FLOATING
C1184 avdd.t284 0 0.09482f **FLOATING
C1185 avdd.n206 0 0.13889f **FLOATING
C1186 avdd.t285 0 0.01613f **FLOATING
C1187 avdd.n207 0 0.03079f **FLOATING
C1188 avdd.n208 0 0.06443f **FLOATING
C1189 avdd.n209 0 3.87524f **FLOATING
C1190 avdd.n210 0 2.89876f **FLOATING
C1191 avdd.n211 0 0.54101f **FLOATING
C1192 avdd.n212 0 0.22311f **FLOATING
C1193 avdd.n213 0 0.13505f **FLOATING
C1194 avdd.t163 0 0.01861f **FLOATING
C1195 avdd.n214 0 0.0584f **FLOATING
C1196 avdd.t165 0 0.01909f **FLOATING
C1197 avdd.n215 0 0.04054f **FLOATING
C1198 avdd.n216 0 0.04054f **FLOATING
C1199 avdd.t162 0 0.12182f **FLOATING
C1200 avdd.n217 0 0.0148f **FLOATING
C1201 avdd.n218 0 0.12152f **FLOATING
C1202 avdd.t164 0 0.12182f **FLOATING
C1203 avdd.n219 0 0.12417f **FLOATING
C1204 avdd.n220 0 0.08303f **FLOATING
C1205 avdd.t155 0 0.01909f **FLOATING
C1206 avdd.t154 0 0.14751f **FLOATING
C1207 avdd.n221 0 0.32056f **FLOATING
C1208 avdd.n222 0 0.11564f **FLOATING
C1209 avdd.n223 0 0.04514f **FLOATING
C1210 avdd.n224 0 0.40282f **FLOATING
C1211 avdd.n225 0 1.36009f **FLOATING
C1212 avdd.n226 0 0.32215f **FLOATING
C1213 avdd.n227 0 0.29609f **FLOATING
C1214 avdd.n228 0 0.04054f **FLOATING
C1215 avdd.n229 0 0.04054f **FLOATING
C1216 avdd.n230 0 0.12417f **FLOATING
C1217 avdd.t270 0 0.12182f **FLOATING
C1218 avdd.n231 0 0.0148f **FLOATING
C1219 avdd.n232 0 0.12152f **FLOATING
C1220 avdd.t236 0 0.12182f **FLOATING
C1221 avdd.n233 0 0.13228f **FLOATING
C1222 avdd.n234 0 0.05291f **FLOATING
C1223 avdd.n235 0 0.06202f **FLOATING
C1224 avdd.n236 0 0.22294f **FLOATING
C1225 avdd.t174 0 0.12368f **FLOATING
C1226 avdd.t175 0 0.04896f **FLOATING
C1227 avdd.n237 0 0.28487f **FLOATING
C1228 avdd.n238 0 0.71105f **FLOATING
C1229 avdd.t110 0 0.01935f **FLOATING
C1230 avdd.t400 0 0.01055f **FLOATING
C1231 avdd.n239 0 0.09149f **FLOATING
C1232 avdd.t44 0 0.01935f **FLOATING
C1233 avdd.t391 0 0.01055f **FLOATING
C1234 avdd.n240 0 0.03208f **FLOATING
C1235 avdd.n241 0 0.13216f **FLOATING
C1236 dffrs_3.setb 0 0.00111f **FLOATING
C1237 avdd.n242 0 0.01325f **FLOATING
C1238 avdd.t291 0 0.00645f **FLOATING
C1239 avdd.t341 0 0.00645f **FLOATING
C1240 avdd.n243 0 0.02312f **FLOATING
C1241 avdd.n244 0 0.14951f **FLOATING
C1242 avdd.t290 0 0.09482f **FLOATING
C1243 avdd.t340 0 0.08403f **FLOATING
C1244 avdd.t45 0 0.09482f **FLOATING
C1245 avdd.n245 0 0.13889f **FLOATING
C1246 avdd.t46 0 0.01613f **FLOATING
C1247 avdd.n246 0 0.03079f **FLOATING
C1248 avdd.n247 0 0.06566f **FLOATING
C1249 avdd.n248 0 2.80882f **FLOATING
C1250 avdd.t315 0 0.00645f **FLOATING
C1251 avdd.t181 0 0.00645f **FLOATING
C1252 avdd.n249 0 0.02312f **FLOATING
C1253 avdd.n250 0 0.14951f **FLOATING
C1254 avdd.t314 0 0.09482f **FLOATING
C1255 avdd.t180 0 0.08403f **FLOATING
C1256 avdd.t111 0 0.09482f **FLOATING
C1257 avdd.n251 0 0.13889f **FLOATING
C1258 avdd.t112 0 0.01613f **FLOATING
C1259 avdd.n252 0 0.03079f **FLOATING
C1260 avdd.n253 0 0.06443f **FLOATING
C1261 avdd.t19 0 0.00645f **FLOATING
C1262 avdd.t76 0 0.00645f **FLOATING
C1263 avdd.n254 0 0.02312f **FLOATING
C1264 avdd.n255 0 0.14951f **FLOATING
C1265 avdd.t18 0 0.09482f **FLOATING
C1266 avdd.t75 0 0.08403f **FLOATING
C1267 avdd.t250 0 0.09482f **FLOATING
C1268 avdd.n256 0 0.13889f **FLOATING
C1269 avdd.t251 0 0.01613f **FLOATING
C1270 avdd.n257 0 0.03079f **FLOATING
C1271 avdd.n258 0 0.06443f **FLOATING
C1272 avdd.n259 0 2.85645f **FLOATING
C1273 avdd.t40 0 0.00645f **FLOATING
C1274 avdd.t375 0 0.00645f **FLOATING
C1275 avdd.n260 0 0.02312f **FLOATING
C1276 avdd.n261 0 0.14951f **FLOATING
C1277 avdd.t39 0 0.09482f **FLOATING
C1278 avdd.t374 0 0.08403f **FLOATING
C1279 avdd.t256 0 0.09482f **FLOATING
C1280 avdd.n262 0 0.13889f **FLOATING
C1281 avdd.t257 0 0.01613f **FLOATING
C1282 avdd.n263 0 0.03079f **FLOATING
C1283 avdd.n264 0 0.06443f **FLOATING
C1284 avdd.n265 0 1.80909f **FLOATING
C1285 avdd.t343 0 0.00645f **FLOATING
C1286 avdd.t269 0 0.00645f **FLOATING
C1287 avdd.n266 0 0.02312f **FLOATING
C1288 avdd.n267 0 0.14951f **FLOATING
C1289 avdd.t342 0 0.09482f **FLOATING
C1290 avdd.t268 0 0.08403f **FLOATING
C1291 avdd.t288 0 0.09482f **FLOATING
C1292 avdd.n268 0 0.13889f **FLOATING
C1293 avdd.t289 0 0.01613f **FLOATING
C1294 avdd.n269 0 0.03079f **FLOATING
C1295 avdd.n270 0 0.06443f **FLOATING
C1296 avdd.n271 0 1.28162f **FLOATING
C1297 avdd.t38 0 0.0195f **FLOATING
C1298 avdd.t392 0 0.01037f **FLOATING
C1299 avdd.n272 0 0.08453f **FLOATING
C1300 avdd.t74 0 0.01942f **FLOATING
C1301 avdd.t380 0 0.01045f **FLOATING
C1302 avdd.n273 0 0.07805f **FLOATING
C1303 avdd.t107 0 0.01942f **FLOATING
C1304 avdd.t398 0 0.01045f **FLOATING
C1305 avdd.n274 0 0.04661f **FLOATING
C1306 avdd.n275 0 0.14749f **FLOATING
C1307 avdd.n276 0 0.11028f **FLOATING
C1308 dffrs_3.resetb 0 0.01446f **FLOATING
C1309 avdd.t205 0 0.00645f **FLOATING
C1310 avdd.t109 0 0.00645f **FLOATING
C1311 avdd.n277 0 0.02312f **FLOATING
C1312 avdd.n278 0 0.14951f **FLOATING
C1313 avdd.t204 0 0.09482f **FLOATING
C1314 avdd.t108 0 0.08403f **FLOATING
C1315 avdd.t376 0 0.09482f **FLOATING
C1316 avdd.n279 0 0.13889f **FLOATING
C1317 avdd.t377 0 0.01613f **FLOATING
C1318 avdd.n280 0 0.03079f **FLOATING
C1319 avdd.n281 0 0.06443f **FLOATING
C1320 avdd.n282 0 3.87524f **FLOATING
C1321 avdd.n283 0 2.89876f **FLOATING
C1322 avdd.n284 0 0.54101f **FLOATING
C1323 avdd.n285 0 0.22311f **FLOATING
C1324 avdd.n286 0 0.13505f **FLOATING
C1325 avdd.t313 0 0.01861f **FLOATING
C1326 avdd.n287 0 0.0584f **FLOATING
C1327 avdd.t333 0 0.01909f **FLOATING
C1328 avdd.n288 0 0.04054f **FLOATING
C1329 avdd.n289 0 0.04054f **FLOATING
C1330 avdd.t312 0 0.12182f **FLOATING
C1331 avdd.n290 0 0.0148f **FLOATING
C1332 avdd.n291 0 0.12152f **FLOATING
C1333 avdd.t332 0 0.12182f **FLOATING
C1334 avdd.n292 0 0.12417f **FLOATING
C1335 avdd.n293 0 0.08303f **FLOATING
C1336 avdd.t27 0 0.01909f **FLOATING
C1337 avdd.t26 0 0.14751f **FLOATING
C1338 avdd.n294 0 0.32056f **FLOATING
C1339 avdd.n295 0 0.11564f **FLOATING
C1340 avdd.n296 0 0.04514f **FLOATING
C1341 avdd.n297 0 0.40282f **FLOATING
C1342 avdd.n298 0 1.36009f **FLOATING
C1343 avdd.n299 0 0.32215f **FLOATING
C1344 avdd.n300 0 0.29609f **FLOATING
C1345 avdd.n301 0 0.04054f **FLOATING
C1346 avdd.n302 0 0.04054f **FLOATING
C1347 avdd.n303 0 0.12417f **FLOATING
C1348 avdd.t292 0 0.12182f **FLOATING
C1349 avdd.n304 0 0.0148f **FLOATING
C1350 avdd.n305 0 0.12152f **FLOATING
C1351 avdd.t304 0 0.12182f **FLOATING
C1352 avdd.n306 0 0.13228f **FLOATING
C1353 avdd.n307 0 0.05291f **FLOATING
C1354 avdd.n308 0 0.06202f **FLOATING
C1355 avdd.n309 0 0.22294f **FLOATING
C1356 avdd.t344 0 0.12368f **FLOATING
C1357 avdd.t345 0 0.04896f **FLOATING
C1358 avdd.n310 0 0.28487f **FLOATING
C1359 avdd.n311 0 0.71105f **FLOATING
C1360 avdd.t68 0 0.01935f **FLOATING
C1361 avdd.t383 0 0.01055f **FLOATING
C1362 avdd.n312 0 0.09149f **FLOATING
C1363 avdd.t65 0 0.01935f **FLOATING
C1364 avdd.t382 0 0.01055f **FLOATING
C1365 avdd.n313 0 0.03208f **FLOATING
C1366 avdd.n314 0 0.13216f **FLOATING
C1367 dffrs_2.setb 0 0.00111f **FLOATING
C1368 avdd.n315 0 0.01325f **FLOATING
C1369 avdd.t241 0 0.00645f **FLOATING
C1370 avdd.t177 0 0.00645f **FLOATING
C1371 avdd.n316 0 0.02312f **FLOATING
C1372 avdd.n317 0 0.14951f **FLOATING
C1373 avdd.t240 0 0.09482f **FLOATING
C1374 avdd.t176 0 0.08403f **FLOATING
C1375 avdd.t66 0 0.09482f **FLOATING
C1376 avdd.n318 0 0.13889f **FLOATING
C1377 avdd.t67 0 0.01613f **FLOATING
C1378 avdd.n319 0 0.03079f **FLOATING
C1379 avdd.n320 0 0.06566f **FLOATING
C1380 avdd.n321 0 2.80882f **FLOATING
C1381 avdd.t1 0 0.00645f **FLOATING
C1382 avdd.t239 0 0.00645f **FLOATING
C1383 avdd.n322 0 0.02312f **FLOATING
C1384 avdd.n323 0 0.14951f **FLOATING
C1385 avdd.t0 0 0.09482f **FLOATING
C1386 avdd.t238 0 0.08403f **FLOATING
C1387 avdd.t69 0 0.09482f **FLOATING
C1388 avdd.n324 0 0.13889f **FLOATING
C1389 avdd.t70 0 0.01613f **FLOATING
C1390 avdd.n325 0 0.03079f **FLOATING
C1391 avdd.n326 0 0.06443f **FLOATING
C1392 avdd.t355 0 0.00645f **FLOATING
C1393 avdd.t64 0 0.00645f **FLOATING
C1394 avdd.n327 0 0.02312f **FLOATING
C1395 avdd.n328 0 0.14951f **FLOATING
C1396 avdd.t354 0 0.09482f **FLOATING
C1397 avdd.t63 0 0.08403f **FLOATING
C1398 avdd.t206 0 0.09482f **FLOATING
C1399 avdd.n329 0 0.13889f **FLOATING
C1400 avdd.t207 0 0.01613f **FLOATING
C1401 avdd.n330 0 0.03079f **FLOATING
C1402 avdd.n331 0 0.06443f **FLOATING
C1403 avdd.n332 0 2.85645f **FLOATING
C1404 avdd.t115 0 0.00645f **FLOATING
C1405 avdd.t219 0 0.00645f **FLOATING
C1406 avdd.n333 0 0.02312f **FLOATING
C1407 avdd.n334 0 0.14951f **FLOATING
C1408 avdd.t114 0 0.09482f **FLOATING
C1409 avdd.t218 0 0.08403f **FLOATING
C1410 avdd.t152 0 0.09482f **FLOATING
C1411 avdd.n335 0 0.13889f **FLOATING
C1412 avdd.t153 0 0.01613f **FLOATING
C1413 avdd.n336 0 0.03079f **FLOATING
C1414 avdd.n337 0 0.06443f **FLOATING
C1415 avdd.n338 0 1.80909f **FLOATING
C1416 avdd.t179 0 0.00645f **FLOATING
C1417 avdd.t275 0 0.00645f **FLOATING
C1418 avdd.n339 0 0.02312f **FLOATING
C1419 avdd.n340 0 0.14951f **FLOATING
C1420 avdd.t178 0 0.09482f **FLOATING
C1421 avdd.t274 0 0.08403f **FLOATING
C1422 avdd.t242 0 0.09482f **FLOATING
C1423 avdd.n341 0 0.13889f **FLOATING
C1424 avdd.t243 0 0.01613f **FLOATING
C1425 avdd.n342 0 0.03079f **FLOATING
C1426 avdd.n343 0 0.06443f **FLOATING
C1427 avdd.n344 0 1.28162f **FLOATING
C1428 avdd.t113 0 0.0195f **FLOATING
C1429 avdd.t397 0 0.01037f **FLOATING
C1430 avdd.n345 0 0.08453f **FLOATING
C1431 avdd.t62 0 0.01942f **FLOATING
C1432 avdd.t385 0 0.01045f **FLOATING
C1433 avdd.n346 0 0.07805f **FLOATING
C1434 avdd.t83 0 0.01942f **FLOATING
C1435 avdd.t405 0 0.01045f **FLOATING
C1436 avdd.n347 0 0.04661f **FLOATING
C1437 avdd.n348 0 0.14749f **FLOATING
C1438 avdd.n349 0 0.11028f **FLOATING
C1439 dffrs_2.resetb 0 0.01446f **FLOATING
C1440 avdd.t249 0 0.00645f **FLOATING
C1441 avdd.t85 0 0.00645f **FLOATING
C1442 avdd.n350 0 0.02312f **FLOATING
C1443 avdd.n351 0 0.14951f **FLOATING
C1444 avdd.t248 0 0.09482f **FLOATING
C1445 avdd.t84 0 0.08403f **FLOATING
C1446 avdd.t220 0 0.09482f **FLOATING
C1447 avdd.n352 0 0.13889f **FLOATING
C1448 avdd.t221 0 0.01613f **FLOATING
C1449 avdd.n353 0 0.03079f **FLOATING
C1450 avdd.n354 0 0.06443f **FLOATING
C1451 avdd.n355 0 3.87524f **FLOATING
C1452 avdd.n356 0 2.89876f **FLOATING
C1453 avdd.n357 0 0.54101f **FLOATING
C1454 avdd.n358 0 0.22311f **FLOATING
C1455 avdd.n359 0 0.13505f **FLOATING
C1456 avdd.t245 0 0.01861f **FLOATING
C1457 avdd.n360 0 0.0584f **FLOATING
C1458 avdd.t7 0 0.01909f **FLOATING
C1459 avdd.n361 0 0.04054f **FLOATING
C1460 avdd.n362 0 0.04054f **FLOATING
C1461 avdd.t244 0 0.12182f **FLOATING
C1462 avdd.n363 0 0.0148f **FLOATING
C1463 avdd.n364 0 0.12152f **FLOATING
C1464 avdd.t6 0 0.12182f **FLOATING
C1465 avdd.n365 0 0.12417f **FLOATING
C1466 avdd.n366 0 0.08303f **FLOATING
C1467 avdd.t3 0 0.01909f **FLOATING
C1468 avdd.t2 0 0.14751f **FLOATING
C1469 avdd.n367 0 0.32056f **FLOATING
C1470 avdd.n368 0 0.11564f **FLOATING
C1471 avdd.n369 0 0.04514f **FLOATING
C1472 avdd.n370 0 0.40282f **FLOATING
C1473 avdd.n371 0 1.36009f **FLOATING
C1474 avdd.n372 0 0.32215f **FLOATING
C1475 avdd.n373 0 0.29609f **FLOATING
C1476 avdd.n374 0 0.04054f **FLOATING
C1477 avdd.n375 0 0.04054f **FLOATING
C1478 avdd.n376 0 0.12417f **FLOATING
C1479 avdd.t350 0 0.12182f **FLOATING
C1480 avdd.n377 0 0.0148f **FLOATING
C1481 avdd.n378 0 0.12152f **FLOATING
C1482 avdd.t368 0 0.12182f **FLOATING
C1483 avdd.n379 0 0.13228f **FLOATING
C1484 avdd.n380 0 0.05291f **FLOATING
C1485 avdd.n381 0 0.06202f **FLOATING
C1486 avdd.n382 0 0.22294f **FLOATING
C1487 avdd.t214 0 0.12368f **FLOATING
C1488 avdd.t215 0 0.04896f **FLOATING
C1489 avdd.n383 0 0.28487f **FLOATING
C1490 avdd.n384 0 0.71105f **FLOATING
C1491 avdd.t50 0 0.01935f **FLOATING
C1492 avdd.t390 0 0.01055f **FLOATING
C1493 avdd.n385 0 0.09149f **FLOATING
C1494 avdd.t53 0 0.01935f **FLOATING
C1495 avdd.t388 0 0.01055f **FLOATING
C1496 avdd.n386 0 0.03208f **FLOATING
C1497 avdd.n387 0 0.13216f **FLOATING
C1498 dffrs_1.setb 0 0.00111f **FLOATING
C1499 avdd.n388 0 0.01325f **FLOATING
C1500 avdd.t283 0 0.00645f **FLOATING
C1501 avdd.t233 0 0.00645f **FLOATING
C1502 avdd.n389 0 0.02312f **FLOATING
C1503 avdd.n390 0 0.14951f **FLOATING
C1504 avdd.t282 0 0.09482f **FLOATING
C1505 avdd.t232 0 0.08403f **FLOATING
C1506 avdd.t54 0 0.09482f **FLOATING
C1507 avdd.n391 0 0.13889f **FLOATING
C1508 avdd.t55 0 0.01613f **FLOATING
C1509 avdd.n392 0 0.03079f **FLOATING
C1510 avdd.n393 0 0.06566f **FLOATING
C1511 avdd.n394 0 2.80882f **FLOATING
C1512 avdd.t363 0 0.00645f **FLOATING
C1513 avdd.t303 0 0.00645f **FLOATING
C1514 avdd.n395 0 0.02312f **FLOATING
C1515 avdd.n396 0 0.14951f **FLOATING
C1516 avdd.t362 0 0.09482f **FLOATING
C1517 avdd.t302 0 0.08403f **FLOATING
C1518 avdd.t51 0 0.09482f **FLOATING
C1519 avdd.n397 0 0.13889f **FLOATING
C1520 avdd.t52 0 0.01613f **FLOATING
C1521 avdd.n398 0 0.03079f **FLOATING
C1522 avdd.n399 0 0.06443f **FLOATING
C1523 avdd.t277 0 0.00645f **FLOATING
C1524 avdd.t118 0 0.00645f **FLOATING
C1525 avdd.n400 0 0.02312f **FLOATING
C1526 avdd.n401 0 0.14951f **FLOATING
C1527 avdd.t276 0 0.09482f **FLOATING
C1528 avdd.t117 0 0.08403f **FLOATING
C1529 avdd.t264 0 0.09482f **FLOATING
C1530 avdd.n402 0 0.13889f **FLOATING
C1531 avdd.t265 0 0.01613f **FLOATING
C1532 avdd.n403 0 0.03079f **FLOATING
C1533 avdd.n404 0 0.06443f **FLOATING
C1534 avdd.n405 0 2.85645f **FLOATING
C1535 avdd.t103 0 0.00645f **FLOATING
C1536 avdd.t253 0 0.00645f **FLOATING
C1537 avdd.n406 0 0.02312f **FLOATING
C1538 avdd.n407 0 0.14951f **FLOATING
C1539 avdd.t102 0 0.09482f **FLOATING
C1540 avdd.t252 0 0.08403f **FLOATING
C1541 avdd.t334 0 0.09482f **FLOATING
C1542 avdd.n408 0 0.13889f **FLOATING
C1543 avdd.t335 0 0.01613f **FLOATING
C1544 avdd.n409 0 0.03079f **FLOATING
C1545 avdd.n410 0 0.06443f **FLOATING
C1546 avdd.n411 0 1.80909f **FLOATING
C1547 avdd.t231 0 0.00645f **FLOATING
C1548 avdd.t331 0 0.00645f **FLOATING
C1549 avdd.n412 0 0.02312f **FLOATING
C1550 avdd.n413 0 0.14951f **FLOATING
C1551 avdd.t230 0 0.09482f **FLOATING
C1552 avdd.t330 0 0.08403f **FLOATING
C1553 avdd.t280 0 0.09482f **FLOATING
C1554 avdd.n414 0 0.13889f **FLOATING
C1555 avdd.t281 0 0.01613f **FLOATING
C1556 avdd.n415 0 0.03079f **FLOATING
C1557 avdd.n416 0 0.06443f **FLOATING
C1558 avdd.n417 0 1.2808f **FLOATING
C1559 avdd.n418 0 1.81212f **FLOATING
C1560 avdd.t101 0 0.0195f **FLOATING
C1561 avdd.t401 0 0.01037f **FLOATING
C1562 avdd.n419 0 0.08453f **FLOATING
C1563 avdd.t116 0 0.01942f **FLOATING
C1564 avdd.t396 0 0.01045f **FLOATING
C1565 avdd.n420 0 0.07805f **FLOATING
C1566 avdd.t47 0 0.01942f **FLOATING
C1567 avdd.t389 0 0.01045f **FLOATING
C1568 avdd.n421 0 0.04661f **FLOATING
C1569 avdd.n422 0 0.14749f **FLOATING
C1570 avdd.n423 0 0.11028f **FLOATING
C1571 dffrs_1.resetb 0 0.01446f **FLOATING
C1572 avdd.t371 0 0.00645f **FLOATING
C1573 avdd.t49 0 0.00645f **FLOATING
C1574 avdd.n424 0 0.02312f **FLOATING
C1575 avdd.n425 0 0.14951f **FLOATING
C1576 avdd.t370 0 0.09482f **FLOATING
C1577 avdd.t48 0 0.08403f **FLOATING
C1578 avdd.t254 0 0.09482f **FLOATING
C1579 avdd.n426 0 0.13889f **FLOATING
C1580 avdd.t255 0 0.01613f **FLOATING
C1581 avdd.n427 0 0.03079f **FLOATING
C1582 avdd.n428 0 0.06443f **FLOATING
C1583 avdd.n429 0 3.87524f **FLOATING
C1584 avdd.n430 0 1.08746f **FLOATING
C1585 avdd.n431 0 0.54101f **FLOATING
C1586 avdd.n432 0 0.22311f **FLOATING
C1587 avdd.n433 0 0.13505f **FLOATING
C1588 avdd.t157 0 0.01861f **FLOATING
C1589 avdd.n434 0 0.0584f **FLOATING
C1590 avdd.t185 0 0.01909f **FLOATING
C1591 avdd.n435 0 0.04054f **FLOATING
C1592 avdd.n436 0 0.04054f **FLOATING
C1593 avdd.t156 0 0.12182f **FLOATING
C1594 avdd.n437 0 0.0148f **FLOATING
C1595 avdd.n438 0 0.12152f **FLOATING
C1596 avdd.t184 0 0.12182f **FLOATING
C1597 avdd.n439 0 0.12417f **FLOATING
C1598 avdd.n440 0 0.08303f **FLOATING
C1599 avdd.t33 0 0.01909f **FLOATING
C1600 avdd.t32 0 0.14751f **FLOATING
C1601 avdd.n441 0 0.32056f **FLOATING
C1602 avdd.n442 0 0.11564f **FLOATING
C1603 avdd.n443 0 0.04514f **FLOATING
C1604 avdd.n444 0 0.40282f **FLOATING
C1605 avdd.n445 0 1.36009f **FLOATING
C1606 avdd.n446 0 0.32215f **FLOATING
C1607 avdd.n447 0 0.29609f **FLOATING
C1608 avdd.n448 0 0.04054f **FLOATING
C1609 avdd.n449 0 0.04054f **FLOATING
C1610 avdd.n450 0 0.12417f **FLOATING
C1611 avdd.t216 0 0.12182f **FLOATING
C1612 avdd.n451 0 0.0148f **FLOATING
C1613 avdd.n452 0 0.12152f **FLOATING
C1614 avdd.t338 0 0.12182f **FLOATING
C1615 avdd.n453 0 0.13228f **FLOATING
C1616 avdd.n454 0 0.05291f **FLOATING
C1617 avdd.n455 0 0.06202f **FLOATING
C1618 avdd.n456 0 0.22294f **FLOATING
C1619 avdd.t328 0 0.12368f **FLOATING
C1620 avdd.t329 0 0.04896f **FLOATING
C1621 avdd.n457 0 0.28487f **FLOATING
C1622 avdd.n458 0 0.71105f **FLOATING
C1623 avdd.t119 0 0.0195f **FLOATING
C1624 avdd.t395 0 0.01037f **FLOATING
C1625 avdd.n459 0 0.08453f **FLOATING
C1626 avdd.t89 0 0.01942f **FLOATING
C1627 avdd.t406 0 0.01045f **FLOATING
C1628 avdd.n460 0 0.07805f **FLOATING
C1629 avdd.t122 0 0.01942f **FLOATING
C1630 avdd.t393 0 0.01045f **FLOATING
C1631 avdd.n461 0 0.04661f **FLOATING
C1632 avdd.n462 0 0.14749f **FLOATING
C1633 avdd.n463 0 0.11028f **FLOATING
C1634 dffrs_0.resetb 0 0.01446f **FLOATING
C1635 avdd.t201 0 0.00645f **FLOATING
C1636 avdd.t124 0 0.00645f **FLOATING
C1637 avdd.n464 0 0.02312f **FLOATING
C1638 avdd.n465 0 0.14951f **FLOATING
C1639 avdd.t200 0 0.09482f **FLOATING
C1640 avdd.t123 0 0.08403f **FLOATING
C1641 avdd.t316 0 0.09482f **FLOATING
C1642 avdd.n466 0 0.13889f **FLOATING
C1643 avdd.t317 0 0.01613f **FLOATING
C1644 avdd.n467 0 0.03079f **FLOATING
C1645 avdd.n468 0 0.06443f **FLOATING
C1646 avdd.n469 0 3.87524f **FLOATING
C1647 avdd.n470 0 0.13388f **FLOATING
C1648 avdd.t183 0 0.01861f **FLOATING
C1649 avdd.n471 0 0.0584f **FLOATING
C1650 avdd.t367 0 0.01861f **FLOATING
C1651 avdd.n472 0 0.0584f **FLOATING
C1652 avdd.t365 0 0.01861f **FLOATING
C1653 avdd.n473 0 0.03973f **FLOATING
C1654 avdd.n474 0 0.03973f **FLOATING
C1655 avdd.t182 0 0.12182f **FLOATING
C1656 avdd.n475 0 0.03619f **FLOATING
C1657 avdd.n476 0 0.03619f **FLOATING
C1658 avdd.n477 0 0.0148f **FLOATING
C1659 avdd.n478 0 0.12152f **FLOATING
C1660 avdd.t16 0 0.1124f **FLOATING
C1661 avdd.t17 0 0.1124f **FLOATING
C1662 avdd.n479 0 0.0148f **FLOATING
C1663 avdd.n480 0 0.12152f **FLOATING
C1664 avdd.t366 0 0.1124f **FLOATING
C1665 avdd.t364 0 0.11271f **FLOATING
C1666 avdd.n481 0 0.13168f **FLOATING
C1667 avdd.n482 0 0.0584f **FLOATING
C1668 avdd.n483 0 0.06202f **FLOATING
C1669 avdd.n484 0 0.04054f **FLOATING
C1670 avdd.n485 0 0.04054f **FLOATING
C1671 avdd.t327 0 0.01909f **FLOATING
C1672 avdd.t325 0 0.01909f **FLOATING
C1673 avdd.t324 0 0.14751f **FLOATING
C1674 avdd.n486 0 0.32056f **FLOATING
C1675 avdd 0 0.01754f **FLOATING
C1676 avdd.t348 0 0.12368f **FLOATING
C1677 avdd.t349 0 0.04896f **FLOATING
C1678 avdd.n487 0 0.34759f **FLOATING
C1679 avdd.n488 0 0.50217f **FLOATING
C1680 avdd.n489 0 0.19964f **FLOATING
C1681 avdd.n490 0 0.08303f **FLOATING
C1682 avdd.n491 0 0.12417f **FLOATING
C1683 avdd.t326 0 0.12182f **FLOATING
C1684 avdd.t141 0 0.01861f **FLOATING
C1685 avdd.n492 0 0.0584f **FLOATING
C1686 avdd.n493 0 0.0148f **FLOATING
C1687 avdd.n494 0 0.12152f **FLOATING
C1688 avdd.t140 0 0.12182f **FLOATING
C1689 avdd.n495 0 0.13228f **FLOATING
C1690 avdd.n496 0 0.05291f **FLOATING
C1691 avdd.n497 0 0.29609f **FLOATING
C1692 avdd.n498 0 0.32215f **FLOATING
C1693 avdd.n499 0 0.13505f **FLOATING
C1694 avdd.t267 0 0.01861f **FLOATING
C1695 avdd.n500 0 0.0584f **FLOATING
C1696 avdd.t247 0 0.01909f **FLOATING
C1697 avdd.n501 0 0.04054f **FLOATING
C1698 avdd.n502 0 0.04054f **FLOATING
C1699 avdd.t266 0 0.12182f **FLOATING
C1700 avdd.n503 0 0.0148f **FLOATING
C1701 avdd.n504 0 0.12152f **FLOATING
C1702 avdd.t246 0 0.12182f **FLOATING
C1703 avdd.n505 0 0.12417f **FLOATING
C1704 avdd.n506 0 0.08303f **FLOATING
C1705 avdd.t23 0 0.01909f **FLOATING
C1706 avdd.t22 0 0.14751f **FLOATING
C1707 avdd.n507 0 0.32056f **FLOATING
C1708 avdd.n508 0 0.11564f **FLOATING
C1709 avdd.n509 0 0.04514f **FLOATING
C1710 avdd.n510 0 0.40282f **FLOATING
C1711 avdd.n511 0 1.36009f **FLOATING
C1712 avdd.n512 0 0.22311f **FLOATING
C1713 avdd.n513 0 0.54101f **FLOATING
C1714 avdd.n514 0 2.89876f **FLOATING
C1715 avdd.t13 0 0.00645f **FLOATING
C1716 avdd.t357 0 0.00645f **FLOATING
C1717 avdd.n515 0 0.02312f **FLOATING
C1718 avdd.n516 0 0.14951f **FLOATING
C1719 avdd.t12 0 0.09482f **FLOATING
C1720 avdd.t356 0 0.08403f **FLOATING
C1721 avdd.t306 0 0.09482f **FLOATING
C1722 avdd.n517 0 0.13889f **FLOATING
C1723 avdd.t307 0 0.01613f **FLOATING
C1724 avdd.n518 0 0.03079f **FLOATING
C1725 avdd.n519 0 0.06443f **FLOATING
C1726 avdd.n520 0 1.28162f **FLOATING
C1727 avdd.t121 0 0.00645f **FLOATING
C1728 avdd.t319 0 0.00645f **FLOATING
C1729 avdd.n521 0 0.02312f **FLOATING
C1730 avdd.n522 0 0.14951f **FLOATING
C1731 avdd.t120 0 0.09482f **FLOATING
C1732 avdd.t318 0 0.08403f **FLOATING
C1733 avdd.t146 0 0.09482f **FLOATING
C1734 avdd.n523 0 0.13889f **FLOATING
C1735 avdd.t147 0 0.01613f **FLOATING
C1736 avdd.n524 0 0.03079f **FLOATING
C1737 avdd.n525 0 0.06443f **FLOATING
C1738 avdd.n526 0 1.80909f **FLOATING
C1739 avdd.t133 0 0.00645f **FLOATING
C1740 avdd.t91 0 0.00645f **FLOATING
C1741 avdd.n527 0 0.02312f **FLOATING
C1742 avdd.n528 0 0.14951f **FLOATING
C1743 avdd.t132 0 0.09482f **FLOATING
C1744 avdd.t90 0 0.08403f **FLOATING
C1745 avdd.t160 0 0.09482f **FLOATING
C1746 avdd.n529 0 0.13889f **FLOATING
C1747 avdd.t161 0 0.01613f **FLOATING
C1748 avdd.n530 0 0.03079f **FLOATING
C1749 avdd.n531 0 0.06443f **FLOATING
C1750 avdd.n532 0 2.85645f **FLOATING
C1751 avdd.n533 0 2.80882f **FLOATING
C1752 avdd.n534 0 0.01325f **FLOATING
C1753 dffrs_0.setb 0 0.00111f **FLOATING
