magic
tech gf180mcuD
magscale 1 10
timestamp 1757675420
<< nwell >>
rect 5150 -850 5730 322
<< pwell >>
rect 5150 -1650 5730 -878
<< nmos >>
rect 5400 -1488 5480 -1088
<< pmos >>
rect 5400 -640 5480 160
<< ndiff >>
rect 5312 -1101 5400 -1088
rect 5312 -1475 5325 -1101
rect 5371 -1475 5400 -1101
rect 5312 -1488 5400 -1475
rect 5480 -1101 5568 -1088
rect 5480 -1475 5509 -1101
rect 5555 -1475 5568 -1101
rect 5480 -1488 5568 -1475
<< pdiff >>
rect 5312 147 5400 160
rect 5312 -627 5325 147
rect 5371 -627 5400 147
rect 5312 -640 5400 -627
rect 5480 147 5568 160
rect 5480 -627 5509 147
rect 5555 -627 5568 147
rect 5480 -640 5568 -627
<< ndiffc >>
rect 5325 -1475 5371 -1101
rect 5509 -1475 5555 -1101
<< pdiffc >>
rect 5325 -627 5371 147
rect 5509 -627 5555 147
<< psubdiff >>
rect 5174 -974 5706 -902
rect 5174 -1554 5246 -974
rect 5634 -1554 5706 -974
rect 5174 -1567 5706 -1554
rect 5174 -1613 5290 -1567
rect 5590 -1613 5706 -1567
rect 5174 -1626 5706 -1613
<< nsubdiff >>
rect 5174 285 5706 298
rect 5174 239 5290 285
rect 5590 239 5706 285
rect 5174 226 5706 239
rect 5174 -754 5246 226
rect 5634 -754 5706 226
rect 5174 -826 5706 -754
<< psubdiffcont >>
rect 5290 -1613 5590 -1567
<< nsubdiffcont >>
rect 5290 239 5590 285
<< polysilicon >>
rect 5400 160 5480 204
rect 5400 -673 5480 -640
rect 5400 -719 5413 -673
rect 5467 -719 5480 -673
rect 5400 -732 5480 -719
rect 5400 -1009 5480 -996
rect 5400 -1055 5413 -1009
rect 5467 -1055 5480 -1009
rect 5400 -1088 5480 -1055
rect 5400 -1532 5480 -1488
<< polycontact >>
rect 5413 -719 5467 -673
rect 5413 -1055 5467 -1009
<< metal1 >>
rect 5279 284 5290 285
rect 5208 239 5290 284
rect 5590 284 5601 285
rect 5590 239 5658 284
rect 5208 232 5658 239
rect 5216 224 5658 232
rect 5316 147 5376 224
rect 5316 0 5325 147
rect 5371 0 5376 147
rect 5509 156 5555 158
rect 5509 147 5592 156
rect 5325 -638 5371 -627
rect 5555 -627 5592 147
rect 5509 -638 5592 -627
rect 5402 -700 5413 -673
rect 5400 -719 5413 -700
rect 5467 -700 5478 -673
rect 5467 -719 5480 -700
rect 5400 -1009 5480 -719
rect 5400 -1020 5413 -1009
rect 5402 -1055 5413 -1020
rect 5467 -1020 5480 -1009
rect 5528 -756 5592 -638
rect 5467 -1055 5478 -1020
rect 5528 -1090 5596 -756
rect 5325 -1101 5371 -1090
rect 5324 -1475 5325 -1392
rect 5509 -1101 5596 -1090
rect 5371 -1475 5372 -1392
rect 5324 -1560 5372 -1475
rect 5555 -1472 5596 -1101
rect 5509 -1486 5555 -1475
rect 5280 -1564 5610 -1560
rect 5208 -1567 5658 -1564
rect 5208 -1613 5290 -1567
rect 5590 -1613 5658 -1567
rect 5208 -1624 5658 -1613
<< labels >>
rlabel metal1 5208 252 5208 252 7 avdd
port 0 w
rlabel metal1 5212 -1604 5212 -1604 7 avss
port 1 w
rlabel metal1 5412 -876 5412 -876 7 in
port 2 w
rlabel metal1 5564 -872 5564 -872 7 out
port 3 w
<< end >>
