magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< nwell >>
rect -702 -11254 702 11254
<< pmos >>
rect -452 9044 -52 11044
rect 52 9044 452 11044
rect -452 6812 -52 8812
rect 52 6812 452 8812
rect -452 4580 -52 6580
rect 52 4580 452 6580
rect -452 2348 -52 4348
rect 52 2348 452 4348
rect -452 116 -52 2116
rect 52 116 452 2116
rect -452 -2116 -52 -116
rect 52 -2116 452 -116
rect -452 -4348 -52 -2348
rect 52 -4348 452 -2348
rect -452 -6580 -52 -4580
rect 52 -6580 452 -4580
rect -452 -8812 -52 -6812
rect 52 -8812 452 -6812
rect -452 -11044 -52 -9044
rect 52 -11044 452 -9044
<< pdiff >>
rect -540 11031 -452 11044
rect -540 9057 -527 11031
rect -481 9057 -452 11031
rect -540 9044 -452 9057
rect -52 11031 52 11044
rect -52 9057 -23 11031
rect 23 9057 52 11031
rect -52 9044 52 9057
rect 452 11031 540 11044
rect 452 9057 481 11031
rect 527 9057 540 11031
rect 452 9044 540 9057
rect -540 8799 -452 8812
rect -540 6825 -527 8799
rect -481 6825 -452 8799
rect -540 6812 -452 6825
rect -52 8799 52 8812
rect -52 6825 -23 8799
rect 23 6825 52 8799
rect -52 6812 52 6825
rect 452 8799 540 8812
rect 452 6825 481 8799
rect 527 6825 540 8799
rect 452 6812 540 6825
rect -540 6567 -452 6580
rect -540 4593 -527 6567
rect -481 4593 -452 6567
rect -540 4580 -452 4593
rect -52 6567 52 6580
rect -52 4593 -23 6567
rect 23 4593 52 6567
rect -52 4580 52 4593
rect 452 6567 540 6580
rect 452 4593 481 6567
rect 527 4593 540 6567
rect 452 4580 540 4593
rect -540 4335 -452 4348
rect -540 2361 -527 4335
rect -481 2361 -452 4335
rect -540 2348 -452 2361
rect -52 4335 52 4348
rect -52 2361 -23 4335
rect 23 2361 52 4335
rect -52 2348 52 2361
rect 452 4335 540 4348
rect 452 2361 481 4335
rect 527 2361 540 4335
rect 452 2348 540 2361
rect -540 2103 -452 2116
rect -540 129 -527 2103
rect -481 129 -452 2103
rect -540 116 -452 129
rect -52 2103 52 2116
rect -52 129 -23 2103
rect 23 129 52 2103
rect -52 116 52 129
rect 452 2103 540 2116
rect 452 129 481 2103
rect 527 129 540 2103
rect 452 116 540 129
rect -540 -129 -452 -116
rect -540 -2103 -527 -129
rect -481 -2103 -452 -129
rect -540 -2116 -452 -2103
rect -52 -129 52 -116
rect -52 -2103 -23 -129
rect 23 -2103 52 -129
rect -52 -2116 52 -2103
rect 452 -129 540 -116
rect 452 -2103 481 -129
rect 527 -2103 540 -129
rect 452 -2116 540 -2103
rect -540 -2361 -452 -2348
rect -540 -4335 -527 -2361
rect -481 -4335 -452 -2361
rect -540 -4348 -452 -4335
rect -52 -2361 52 -2348
rect -52 -4335 -23 -2361
rect 23 -4335 52 -2361
rect -52 -4348 52 -4335
rect 452 -2361 540 -2348
rect 452 -4335 481 -2361
rect 527 -4335 540 -2361
rect 452 -4348 540 -4335
rect -540 -4593 -452 -4580
rect -540 -6567 -527 -4593
rect -481 -6567 -452 -4593
rect -540 -6580 -452 -6567
rect -52 -4593 52 -4580
rect -52 -6567 -23 -4593
rect 23 -6567 52 -4593
rect -52 -6580 52 -6567
rect 452 -4593 540 -4580
rect 452 -6567 481 -4593
rect 527 -6567 540 -4593
rect 452 -6580 540 -6567
rect -540 -6825 -452 -6812
rect -540 -8799 -527 -6825
rect -481 -8799 -452 -6825
rect -540 -8812 -452 -8799
rect -52 -6825 52 -6812
rect -52 -8799 -23 -6825
rect 23 -8799 52 -6825
rect -52 -8812 52 -8799
rect 452 -6825 540 -6812
rect 452 -8799 481 -6825
rect 527 -8799 540 -6825
rect 452 -8812 540 -8799
rect -540 -9057 -452 -9044
rect -540 -11031 -527 -9057
rect -481 -11031 -452 -9057
rect -540 -11044 -452 -11031
rect -52 -9057 52 -9044
rect -52 -11031 -23 -9057
rect 23 -11031 52 -9057
rect -52 -11044 52 -11031
rect 452 -9057 540 -9044
rect 452 -11031 481 -9057
rect 527 -11031 540 -9057
rect 452 -11044 540 -11031
<< pdiffc >>
rect -527 9057 -481 11031
rect -23 9057 23 11031
rect 481 9057 527 11031
rect -527 6825 -481 8799
rect -23 6825 23 8799
rect 481 6825 527 8799
rect -527 4593 -481 6567
rect -23 4593 23 6567
rect 481 4593 527 6567
rect -527 2361 -481 4335
rect -23 2361 23 4335
rect 481 2361 527 4335
rect -527 129 -481 2103
rect -23 129 23 2103
rect 481 129 527 2103
rect -527 -2103 -481 -129
rect -23 -2103 23 -129
rect 481 -2103 527 -129
rect -527 -4335 -481 -2361
rect -23 -4335 23 -2361
rect 481 -4335 527 -2361
rect -527 -6567 -481 -4593
rect -23 -6567 23 -4593
rect 481 -6567 527 -4593
rect -527 -8799 -481 -6825
rect -23 -8799 23 -6825
rect 481 -8799 527 -6825
rect -527 -11031 -481 -9057
rect -23 -11031 23 -9057
rect 481 -11031 527 -9057
<< nsubdiff >>
rect -678 11158 678 11230
rect -678 11114 -606 11158
rect -678 -11114 -665 11114
rect -619 -11114 -606 11114
rect 606 11114 678 11158
rect -678 -11158 -606 -11114
rect 606 -11114 619 11114
rect 665 -11114 678 11114
rect 606 -11158 678 -11114
rect -678 -11230 678 -11158
<< nsubdiffcont >>
rect -665 -11114 -619 11114
rect 619 -11114 665 11114
<< polysilicon >>
rect -452 11123 -52 11136
rect -452 11077 -439 11123
rect -65 11077 -52 11123
rect -452 11044 -52 11077
rect 52 11123 452 11136
rect 52 11077 65 11123
rect 439 11077 452 11123
rect 52 11044 452 11077
rect -452 9011 -52 9044
rect -452 8965 -439 9011
rect -65 8965 -52 9011
rect -452 8952 -52 8965
rect 52 9011 452 9044
rect 52 8965 65 9011
rect 439 8965 452 9011
rect 52 8952 452 8965
rect -452 8891 -52 8904
rect -452 8845 -439 8891
rect -65 8845 -52 8891
rect -452 8812 -52 8845
rect 52 8891 452 8904
rect 52 8845 65 8891
rect 439 8845 452 8891
rect 52 8812 452 8845
rect -452 6779 -52 6812
rect -452 6733 -439 6779
rect -65 6733 -52 6779
rect -452 6720 -52 6733
rect 52 6779 452 6812
rect 52 6733 65 6779
rect 439 6733 452 6779
rect 52 6720 452 6733
rect -452 6659 -52 6672
rect -452 6613 -439 6659
rect -65 6613 -52 6659
rect -452 6580 -52 6613
rect 52 6659 452 6672
rect 52 6613 65 6659
rect 439 6613 452 6659
rect 52 6580 452 6613
rect -452 4547 -52 4580
rect -452 4501 -439 4547
rect -65 4501 -52 4547
rect -452 4488 -52 4501
rect 52 4547 452 4580
rect 52 4501 65 4547
rect 439 4501 452 4547
rect 52 4488 452 4501
rect -452 4427 -52 4440
rect -452 4381 -439 4427
rect -65 4381 -52 4427
rect -452 4348 -52 4381
rect 52 4427 452 4440
rect 52 4381 65 4427
rect 439 4381 452 4427
rect 52 4348 452 4381
rect -452 2315 -52 2348
rect -452 2269 -439 2315
rect -65 2269 -52 2315
rect -452 2256 -52 2269
rect 52 2315 452 2348
rect 52 2269 65 2315
rect 439 2269 452 2315
rect 52 2256 452 2269
rect -452 2195 -52 2208
rect -452 2149 -439 2195
rect -65 2149 -52 2195
rect -452 2116 -52 2149
rect 52 2195 452 2208
rect 52 2149 65 2195
rect 439 2149 452 2195
rect 52 2116 452 2149
rect -452 83 -52 116
rect -452 37 -439 83
rect -65 37 -52 83
rect -452 24 -52 37
rect 52 83 452 116
rect 52 37 65 83
rect 439 37 452 83
rect 52 24 452 37
rect -452 -37 -52 -24
rect -452 -83 -439 -37
rect -65 -83 -52 -37
rect -452 -116 -52 -83
rect 52 -37 452 -24
rect 52 -83 65 -37
rect 439 -83 452 -37
rect 52 -116 452 -83
rect -452 -2149 -52 -2116
rect -452 -2195 -439 -2149
rect -65 -2195 -52 -2149
rect -452 -2208 -52 -2195
rect 52 -2149 452 -2116
rect 52 -2195 65 -2149
rect 439 -2195 452 -2149
rect 52 -2208 452 -2195
rect -452 -2269 -52 -2256
rect -452 -2315 -439 -2269
rect -65 -2315 -52 -2269
rect -452 -2348 -52 -2315
rect 52 -2269 452 -2256
rect 52 -2315 65 -2269
rect 439 -2315 452 -2269
rect 52 -2348 452 -2315
rect -452 -4381 -52 -4348
rect -452 -4427 -439 -4381
rect -65 -4427 -52 -4381
rect -452 -4440 -52 -4427
rect 52 -4381 452 -4348
rect 52 -4427 65 -4381
rect 439 -4427 452 -4381
rect 52 -4440 452 -4427
rect -452 -4501 -52 -4488
rect -452 -4547 -439 -4501
rect -65 -4547 -52 -4501
rect -452 -4580 -52 -4547
rect 52 -4501 452 -4488
rect 52 -4547 65 -4501
rect 439 -4547 452 -4501
rect 52 -4580 452 -4547
rect -452 -6613 -52 -6580
rect -452 -6659 -439 -6613
rect -65 -6659 -52 -6613
rect -452 -6672 -52 -6659
rect 52 -6613 452 -6580
rect 52 -6659 65 -6613
rect 439 -6659 452 -6613
rect 52 -6672 452 -6659
rect -452 -6733 -52 -6720
rect -452 -6779 -439 -6733
rect -65 -6779 -52 -6733
rect -452 -6812 -52 -6779
rect 52 -6733 452 -6720
rect 52 -6779 65 -6733
rect 439 -6779 452 -6733
rect 52 -6812 452 -6779
rect -452 -8845 -52 -8812
rect -452 -8891 -439 -8845
rect -65 -8891 -52 -8845
rect -452 -8904 -52 -8891
rect 52 -8845 452 -8812
rect 52 -8891 65 -8845
rect 439 -8891 452 -8845
rect 52 -8904 452 -8891
rect -452 -8965 -52 -8952
rect -452 -9011 -439 -8965
rect -65 -9011 -52 -8965
rect -452 -9044 -52 -9011
rect 52 -8965 452 -8952
rect 52 -9011 65 -8965
rect 439 -9011 452 -8965
rect 52 -9044 452 -9011
rect -452 -11077 -52 -11044
rect -452 -11123 -439 -11077
rect -65 -11123 -52 -11077
rect -452 -11136 -52 -11123
rect 52 -11077 452 -11044
rect 52 -11123 65 -11077
rect 439 -11123 452 -11077
rect 52 -11136 452 -11123
<< polycontact >>
rect -439 11077 -65 11123
rect 65 11077 439 11123
rect -439 8965 -65 9011
rect 65 8965 439 9011
rect -439 8845 -65 8891
rect 65 8845 439 8891
rect -439 6733 -65 6779
rect 65 6733 439 6779
rect -439 6613 -65 6659
rect 65 6613 439 6659
rect -439 4501 -65 4547
rect 65 4501 439 4547
rect -439 4381 -65 4427
rect 65 4381 439 4427
rect -439 2269 -65 2315
rect 65 2269 439 2315
rect -439 2149 -65 2195
rect 65 2149 439 2195
rect -439 37 -65 83
rect 65 37 439 83
rect -439 -83 -65 -37
rect 65 -83 439 -37
rect -439 -2195 -65 -2149
rect 65 -2195 439 -2149
rect -439 -2315 -65 -2269
rect 65 -2315 439 -2269
rect -439 -4427 -65 -4381
rect 65 -4427 439 -4381
rect -439 -4547 -65 -4501
rect 65 -4547 439 -4501
rect -439 -6659 -65 -6613
rect 65 -6659 439 -6613
rect -439 -6779 -65 -6733
rect 65 -6779 439 -6733
rect -439 -8891 -65 -8845
rect 65 -8891 439 -8845
rect -439 -9011 -65 -8965
rect 65 -9011 439 -8965
rect -439 -11123 -65 -11077
rect 65 -11123 439 -11077
<< metal1 >>
rect -665 11171 665 11217
rect -665 11114 -619 11171
rect -450 11077 -439 11123
rect -65 11077 -54 11123
rect 54 11077 65 11123
rect 439 11077 450 11123
rect 619 11114 665 11171
rect -527 11031 -481 11042
rect -527 9046 -481 9057
rect -23 11031 23 11042
rect -23 9046 23 9057
rect 481 11031 527 11042
rect 481 9046 527 9057
rect -450 8965 -439 9011
rect -65 8965 -54 9011
rect 54 8965 65 9011
rect 439 8965 450 9011
rect -450 8845 -439 8891
rect -65 8845 -54 8891
rect 54 8845 65 8891
rect 439 8845 450 8891
rect -527 8799 -481 8810
rect -527 6814 -481 6825
rect -23 8799 23 8810
rect -23 6814 23 6825
rect 481 8799 527 8810
rect 481 6814 527 6825
rect -450 6733 -439 6779
rect -65 6733 -54 6779
rect 54 6733 65 6779
rect 439 6733 450 6779
rect -450 6613 -439 6659
rect -65 6613 -54 6659
rect 54 6613 65 6659
rect 439 6613 450 6659
rect -527 6567 -481 6578
rect -527 4582 -481 4593
rect -23 6567 23 6578
rect -23 4582 23 4593
rect 481 6567 527 6578
rect 481 4582 527 4593
rect -450 4501 -439 4547
rect -65 4501 -54 4547
rect 54 4501 65 4547
rect 439 4501 450 4547
rect -450 4381 -439 4427
rect -65 4381 -54 4427
rect 54 4381 65 4427
rect 439 4381 450 4427
rect -527 4335 -481 4346
rect -527 2350 -481 2361
rect -23 4335 23 4346
rect -23 2350 23 2361
rect 481 4335 527 4346
rect 481 2350 527 2361
rect -450 2269 -439 2315
rect -65 2269 -54 2315
rect 54 2269 65 2315
rect 439 2269 450 2315
rect -450 2149 -439 2195
rect -65 2149 -54 2195
rect 54 2149 65 2195
rect 439 2149 450 2195
rect -527 2103 -481 2114
rect -527 118 -481 129
rect -23 2103 23 2114
rect -23 118 23 129
rect 481 2103 527 2114
rect 481 118 527 129
rect -450 37 -439 83
rect -65 37 -54 83
rect 54 37 65 83
rect 439 37 450 83
rect -450 -83 -439 -37
rect -65 -83 -54 -37
rect 54 -83 65 -37
rect 439 -83 450 -37
rect -527 -129 -481 -118
rect -527 -2114 -481 -2103
rect -23 -129 23 -118
rect -23 -2114 23 -2103
rect 481 -129 527 -118
rect 481 -2114 527 -2103
rect -450 -2195 -439 -2149
rect -65 -2195 -54 -2149
rect 54 -2195 65 -2149
rect 439 -2195 450 -2149
rect -450 -2315 -439 -2269
rect -65 -2315 -54 -2269
rect 54 -2315 65 -2269
rect 439 -2315 450 -2269
rect -527 -2361 -481 -2350
rect -527 -4346 -481 -4335
rect -23 -2361 23 -2350
rect -23 -4346 23 -4335
rect 481 -2361 527 -2350
rect 481 -4346 527 -4335
rect -450 -4427 -439 -4381
rect -65 -4427 -54 -4381
rect 54 -4427 65 -4381
rect 439 -4427 450 -4381
rect -450 -4547 -439 -4501
rect -65 -4547 -54 -4501
rect 54 -4547 65 -4501
rect 439 -4547 450 -4501
rect -527 -4593 -481 -4582
rect -527 -6578 -481 -6567
rect -23 -4593 23 -4582
rect -23 -6578 23 -6567
rect 481 -4593 527 -4582
rect 481 -6578 527 -6567
rect -450 -6659 -439 -6613
rect -65 -6659 -54 -6613
rect 54 -6659 65 -6613
rect 439 -6659 450 -6613
rect -450 -6779 -439 -6733
rect -65 -6779 -54 -6733
rect 54 -6779 65 -6733
rect 439 -6779 450 -6733
rect -527 -6825 -481 -6814
rect -527 -8810 -481 -8799
rect -23 -6825 23 -6814
rect -23 -8810 23 -8799
rect 481 -6825 527 -6814
rect 481 -8810 527 -8799
rect -450 -8891 -439 -8845
rect -65 -8891 -54 -8845
rect 54 -8891 65 -8845
rect 439 -8891 450 -8845
rect -450 -9011 -439 -8965
rect -65 -9011 -54 -8965
rect 54 -9011 65 -8965
rect 439 -9011 450 -8965
rect -527 -9057 -481 -9046
rect -527 -11042 -481 -11031
rect -23 -9057 23 -9046
rect -23 -11042 23 -11031
rect 481 -9057 527 -9046
rect 481 -11042 527 -11031
rect -665 -11171 -619 -11114
rect -450 -11123 -439 -11077
rect -65 -11123 -54 -11077
rect 54 -11123 65 -11077
rect 439 -11123 450 -11077
rect 619 -11171 665 -11114
rect -665 -11217 665 -11171
<< properties >>
string FIXED_BBOX -642 -11194 642 11194
string gencell pfet_03v3
string library gf180mcu
string parameters w 10.0 l 2.0 m 10 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
