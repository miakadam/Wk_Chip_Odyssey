magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 221 -23 267
rect 134 221 145 267
rect -118 129 -107 175
rect 50 129 61 175
rect 218 129 229 175
rect -34 37 -23 83
rect 134 37 145 83
<< nwell >>
rect -206 -22 376 366
<< pmos >>
rect -28 130 28 174
rect 140 130 196 174
<< pdiff >>
rect -120 175 -48 188
rect -120 129 -107 175
rect -61 174 -48 175
rect 48 175 120 188
rect 48 174 61 175
rect -61 130 -28 174
rect 28 130 61 174
rect -61 129 -48 130
rect -120 116 -48 129
rect 48 129 61 130
rect 107 174 120 175
rect 216 175 288 188
rect 216 174 229 175
rect 107 130 140 174
rect 196 130 229 174
rect 107 129 120 130
rect 48 116 120 129
rect 216 129 229 130
rect 275 129 288 175
rect 216 116 288 129
<< pdiffc >>
rect -107 129 -61 175
rect 61 129 107 175
rect 229 129 275 175
<< polysilicon >>
rect -36 267 36 280
rect -36 221 -23 267
rect 23 221 36 267
rect -36 208 36 221
rect 132 267 204 280
rect 132 221 145 267
rect 191 221 204 267
rect 132 208 204 221
rect -28 174 28 208
rect -28 96 28 130
rect 140 174 196 208
rect 140 96 196 130
rect -36 83 36 96
rect -36 37 -23 83
rect 23 37 36 83
rect -36 24 36 37
rect 132 83 204 96
rect 132 37 145 83
rect 191 37 204 83
rect 132 24 204 37
<< polycontact >>
rect -23 221 23 267
rect 145 221 191 267
rect -23 37 23 83
rect 145 37 191 83
<< metal1 >>
rect -34 221 -23 267
rect 23 221 34 267
rect 134 221 145 267
rect 191 221 202 267
rect -118 129 -107 175
rect -61 129 -50 175
rect 50 129 61 175
rect 107 129 118 175
rect 218 129 229 175
rect 275 129 286 175
rect -34 37 -23 83
rect 23 37 34 83
rect 134 37 145 83
rect 191 37 202 83
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.220 l 0.280 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
