** sch_path: /foss/designs/FinalBlocksLayout/nor2/nor2.sch
.subckt nor2 VDD VSS OUT A B
*.PININFO VDD:B VSS:B B:B A:B OUT:B
XM1 OUT A VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=1
XM2 OUT B VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=1
XM3 OUT B net1 VDD pfet_03v3 L=0.5u W=3u nf=1 m=2
XM4 net1 A VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=2
.ends
