magic
tech gf180mcuD
magscale 1 10
timestamp 1757546838
<< error_s >>
rect 5394 -447 5528 -418
rect 5592 -447 5686 -418
rect 5394 -464 5403 -447
rect 5440 -654 5449 -464
rect 5633 -576 5640 -541
rect 5440 -664 5526 -654
rect 5679 -664 5686 -576
rect 5495 -864 5526 -664
rect 5368 -1020 5440 -1018
rect 5368 -1064 5403 -1020
rect 5440 -1064 5449 -1020
rect 5414 -1264 5449 -1064
rect 5440 -1401 5449 -1264
rect 5679 -1332 5686 -818
rect 5482 -1374 5570 -1332
rect 5650 -1374 5738 -1332
rect 5368 -1432 5440 -1418
rect 5510 -1432 5710 -1388
rect 5368 -1440 5778 -1432
rect 5368 -1447 5544 -1440
rect 5368 -1464 5403 -1447
rect 5416 -1460 5544 -1447
rect 5550 -1460 5778 -1440
rect 5440 -1464 5449 -1460
rect 5414 -1501 5449 -1464
rect 5570 -1466 5650 -1460
rect 5524 -1508 5644 -1488
rect 5377 -1518 5414 -1514
rect 5484 -1518 5684 -1508
rect 5377 -1547 5768 -1518
rect 5400 -1560 5768 -1547
rect 5414 -1664 5423 -1624
rect 5653 -1664 5686 -1624
rect 5318 -1764 5326 -1732
rect 4788 -1847 5080 -1818
rect 4788 -1864 4797 -1847
rect 4834 -2064 4843 -1864
rect 5027 -1976 5034 -1941
rect 5073 -2064 5080 -1976
rect 4788 -2264 4797 -2218
rect 4834 -2455 4843 -2264
rect 5073 -2372 5080 -2218
rect 4834 -2464 5034 -2455
rect 5318 -2560 5874 -1764
rect 5320 -2584 5874 -2560
<< metal1 >>
rect 5208 232 5658 284
rect 5216 224 5658 232
rect 5316 0 5376 224
rect 5400 -1020 5480 -700
rect 5528 -756 5592 156
rect 5528 -1252 5596 -756
rect 5324 -1560 5372 -1392
rect 5532 -1472 5596 -1252
rect 5280 -1564 5610 -1560
rect 5208 -1624 5658 -1564
use nfet_03v3_Q7US5R  XM3
timestamp 1757546837
transform 1 0 5440 0 1 -1264
box -120 -1320 460 200
use pfet_03v3_YXHA8C  XM4
timestamp 1757546838
transform 1 0 5440 0 1 -264
box -120 -1320 460 200
use nfet_03v3_Q7US5R  XXM3
timestamp 1757546837
transform 1 0 4834 0 1 -1264
box -120 -1320 460 200
use pfet_03v3_YXHA8C  XXM4
timestamp 1757546838
transform 1 0 5414 0 1 -1264
box -120 -1320 460 200
<< labels >>
rlabel metal1 5208 252 5208 252 7 avdd
port 0 w
rlabel metal1 5212 -1604 5212 -1604 7 avss
port 1 w
rlabel metal1 5412 -876 5412 -876 7 in
port 2 w
rlabel metal1 5564 -872 5564 -872 7 out
port 3 w
<< end >>
