** sch_path: /foss/designs/comparator/final_magic/buffer/gf180mcu_osu_sc_gp9t3v3__buf_2.sch
.subckt gf180mcu_osu_sc_gp9t3v3__buf_2 VDD A Y VSS
*.PININFO A:I Y:O VDD:I VSS:I
XM1 net1 A VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 net1 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM3 Y net1 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=2
XM4 Y net1 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=2
.ends
