* NGSPICE file created from comp_SAR_final.ext - technology: (null)

.subckt comp_SAR_final Vdd Vss Clk Vin1 Vin2 Comp_out Reset SAR_in Clk_piso Load Piso_out
X0 Vdd.t89 adc_PISO_0.B4.t4 SARlogic_0.dffrs_7.nand3_8.C.t2 Vdd.t88 pfet_03v3
**devattr s=26000,604 d=26000,604
X1 a_5803_9634 SARlogic_0.dffrs_4.d.t4 Vss.t16 Vss.t15 nfet_03v3
**devattr s=17600,576 d=10400,304
X2 adc_PISO_0.dffrs_4.Qb Vdd.t600 Vdd.t602 Vdd.t601 pfet_03v3
**devattr s=26000,604 d=44000,1176
X3 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t4 Vdd.t866 Vdd.t865 pfet_03v3
**devattr s=26000,604 d=44000,1176
X4 a_37687_30440 inv2_0.out.t2 a_37499_31160.t1 Vss.t231 nfet_03v3
**devattr s=17600,576 d=10400,304
X5 a_n7937_n2793 a_n8017_n2885 a_n9429_n2007.t10 Vss.t201 nfet_03v3
**devattr s=8320,264 d=14080,496
X6 a_28027_28820.t2 adc_PISO_0.B2.t4 Vdd.t772 Vdd.t771 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X7 Vss.t173 a_8377_29020 a_9271_28100 Vss.t172 nfet_03v3
**devattr s=10400,304 d=17600,576
X8 Vdd.t393 Reset.t0 SARlogic_0.dffrs_14.nand3_6.C.t3 Vdd.t392 pfet_03v3
**devattr s=26000,604 d=26000,604
X9 a_n7809_21417 SARlogic_0.dffrs_14.nand3_1.C Vss.t324 Vss.t323 nfet_03v3
**devattr s=17600,576 d=10400,304
X10 SARlogic_0.dffrs_2.nand3_1.C.t0 SARlogic_0.dffrs_2.nand3_6.C.t4 a_459_14043 Vss.t316 nfet_03v3
**devattr s=10400,304 d=17600,576
X11 adc_PISO_0.B4.t3 SARlogic_0.dffrs_1.Qb.t4 Vdd.t271 Vdd.t270 pfet_03v3
**devattr s=44000,1176 d=26000,604
X12 SARlogic_0.dffrs_4.nand3_8.C.t0 SARlogic_0.dffrs_4.nand3_8.Z.t4 a_8543_9633 Vss.t514 nfet_03v3
**devattr s=10400,304 d=17600,576
X13 Vdd.t145 SARlogic_0.dffrs_1.nand3_8.C.t4 SARlogic_0.dffrs_1.Qb.t0 Vdd.t144 pfet_03v3
**devattr s=26000,604 d=26000,604
X14 adc_PISO_0.dffrs_0.Qb Vdd.t597 Vdd.t599 Vdd.t598 pfet_03v3
**devattr s=26000,604 d=44000,1176
X15 a_12401_7428 SARlogic_0.dffrs_5.nand3_8.C.t4 Vss.t46 Vss.t45 nfet_03v3
**devattr s=17600,576 d=10400,304
X16 SARlogic_0.dffrs_3.nand3_8.C.t1 SARlogic_0.dffrs_3.nand3_8.Z.t4 Vdd.t63 Vdd.t62 pfet_03v3
**devattr s=26000,604 d=44000,1176
X17 Vdd.t596 Vdd.t594 a_33257_31423.t2 Vdd.t595 pfet_03v3
**devattr s=26000,604 d=26000,604
X18 SARlogic_0.dffrs_5.nand3_8.C.t2 SARlogic_0.dffrs_5.nand3_6.C.t4 Vdd.t255 Vdd.t254 pfet_03v3
**devattr s=44000,1176 d=26000,604
X19 a_14071_9634 SARlogic_0.dffrs_5.nand3_8.C.t5 a_13887_9634 Vss.t47 nfet_03v3
**devattr s=10400,304 d=10400,304
X20 SARlogic_0.dffrs_1.Qb.t2 Reset.t1 Vdd.t862 Vdd.t861 pfet_03v3
**devattr s=26000,604 d=44000,1176
X21 a_18113_19210 SARlogic_0.dffrs_12.nand3_8.C.t4 a_17929_19210 Vss.t643 nfet_03v3
**devattr s=10400,304 d=10400,304
X22 Vdd.t686 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t7 Vdd.t685 pfet_03v3
**devattr s=10400,304 d=10400,304
X23 a_10029_9634 SARlogic_0.dffrs_4.nand3_8.C.t4 a_9845_9634 Vss.t479 nfet_03v3
**devattr s=10400,304 d=10400,304
X24 SARlogic_0.dffrs_1.nand3_6.C.t1 Clk.t0 a_n3583_11838 Vss.t509 nfet_03v3
**devattr s=10400,304 d=17600,576
X25 a_n4367_29309 Vdd.t943 a_n4551_29309 Vss.t458 nfet_03v3
**devattr s=10400,304 d=10400,304
X26 SARlogic_0.dffrs_9.Qb adc_PISO_0.B3.t4 Vdd.t924 Vdd.t923 pfet_03v3
**devattr s=44000,1176 d=26000,604
X27 a_4841_33627.t0 a_4841_31422.t4 Vdd.t307 Vdd.t306 pfet_03v3
**devattr s=26000,604 d=44000,1176
X28 Vdd.t918 adc_PISO_0.2inmux_1.Bit.t4 a_37499_31160.t3 Vdd.t917 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X29 SARlogic_0.dffrs_5.nand3_6.C.t0 SARlogic_0.dffrs_5.nand3_1.C.t4 Vdd.t189 Vdd.t188 pfet_03v3
**devattr s=44000,1176 d=26000,604
X30 SARlogic_0.dffrs_4.d.t2 Vdd.t591 Vdd.t593 Vdd.t592 pfet_03v3
**devattr s=44000,1176 d=26000,604
X31 SARlogic_0.dffrs_3.nand3_6.C.t2 Clk.t1 Vdd.t702 Vdd.t701 pfet_03v3
**devattr s=26000,604 d=44000,1176
X32 Vdd.t864 Reset.t2 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t863 pfet_03v3
**devattr s=26000,604 d=26000,604
X33 Vdd.t886 a_33337_30170.t4 a_33257_33628.t0 Vdd.t885 pfet_03v3
**devattr s=26000,604 d=26000,604
X34 SARlogic_0.dffrs_13.Qb.t0 SARlogic_0.dffrs_0.d.t4 Vdd.t179 Vdd.t178 pfet_03v3
**devattr s=44000,1176 d=26000,604
X35 Vdd.t301 a_n10831_4320 Comp_out.t7 Vdd.t300 pfet_03v3
**devattr s=18700,450 d=18700,450
X36 a_10639_28100 a_9083_28820.t4 Vdd.t896 Vdd.t895 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X37 a_5987_21414 SARlogic_0.dffrs_9.nand3_6.C.t4 a_5803_21414 Vss.t644 nfet_03v3
**devattr s=10400,304 d=10400,304
X38 a_275_7428 SARlogic_0.dffrs_2.nand3_8.C.t4 Vss.t175 Vss.t174 nfet_03v3
**devattr s=17600,576 d=10400,304
X39 adc_PISO_0.2inmux_5.OUT.t0 a_30255_29264.t4 Vss.t184 Vss.t183 nfet_03v3
**devattr s=17600,576 d=17600,576
X40 SARlogic_0.dffrs_10.nand3_6.C.t2 adc_PISO_0.B1.t4 Vdd.t796 Vdd.t795 pfet_03v3
**devattr s=26000,604 d=44000,1176
X41 adc_PISO_0.B2.t1 SARlogic_0.dffrs_3.Qb.t4 Vdd.t211 Vdd.t210 pfet_03v3
**devattr s=44000,1176 d=26000,604
X42 a_12585_21414 Reset.t3 a_12401_21414 Vss.t616 nfet_03v3
**devattr s=10400,304 d=10400,304
X43 SARlogic_0.dffrs_3.Qb.t2 Reset.t4 a_5987_9634 Vss.t609 nfet_03v3
**devattr s=10400,304 d=17600,576
X44 SARlogic_0.dffrs_12.nand3_6.C.t0 SARlogic_0.dffrs_12.nand3_1.C Vdd.t47 Vdd.t46 pfet_03v3
**devattr s=44000,1176 d=26000,604
X45 SARlogic_0.dffrs_1.Qb.t3 Reset.t5 a_n2097_9634 Vss.t610 nfet_03v3
**devattr s=10400,304 d=17600,576
X46 a_n11637_11838 Vdd.t944 a_n11821_11838 Vss.t457 nfet_03v3
**devattr s=10400,304 d=10400,304
X47 a_n4551_35924 Vdd.t945 Vss.t456 Vss.t455 nfet_03v3
**devattr s=17600,576 d=10400,304
X48 SARlogic_0.dffrs_4.nand3_8.Z.t2 SARlogic_0.dffrs_4.nand3_8.C.t5 Vdd.t638 Vdd.t637 pfet_03v3
**devattr s=44000,1176 d=26000,604
X49 a_1761_19210 adc_PISO_0.B4.t5 Vss.t74 Vss.t73 nfet_03v3
**devattr s=17600,576 d=10400,304
X50 a_14393_33720 a_14313_33628.t4 Vss.t243 Vss.t242 nfet_03v3
**devattr s=17600,576 d=10400,304
X51 a_9271_28100 adc_PISO_0.B4.t6 a_9083_28820.t1 Vss.t72 nfet_03v3
**devattr s=17600,576 d=10400,304
X52 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t4 Vdd.t371 Vdd.t370 pfet_03v3
**devattr s=26000,604 d=44000,1176
X53 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_5.Qb.t4 Vdd.t103 Vdd.t102 pfet_03v3
**devattr s=44000,1176 d=26000,604
X54 a_12585_23619 SARlogic_0.dffrs_11.nand3_8.Z a_12401_23619 Vss.t152 nfet_03v3
**devattr s=10400,304 d=10400,304
X55 adc_PISO_0.dffrs_1.Qb adc_PISO_0.dffrs_1.Q.t4 Vdd.t107 Vdd.t106 pfet_03v3
**devattr s=44000,1176 d=26000,604
X56 Vdd.t774 SARlogic_0.dffrs_14.nand3_6.C.t4 adc_PISO_0.B6.t0 Vdd.t773 pfet_03v3
**devattr s=26000,604 d=26000,604
X57 a_275_14043 Vdd.t946 Vss.t454 Vss.t453 nfet_03v3
**devattr s=17600,576 d=10400,304
X58 a_33257_29218.t0 a_33337_30170.t5 a_33521_31515 Vss.t624 nfet_03v3
**devattr s=10400,304 d=17600,576
X59 SARlogic_0.dffrs_0.Qb.t3 Reset.t6 a_n6139_9634 Vss.t611 nfet_03v3
**devattr s=10400,304 d=17600,576
X60 a_14393_35925 Vdd.t947 Vss.t452 Vss.t451 nfet_03v3
**devattr s=17600,576 d=10400,304
X61 SARlogic_0.dffrs_3.nand3_8.C.t3 SARlogic_0.dffrs_3.nand3_6.C.t4 Vdd.t694 Vdd.t693 pfet_03v3
**devattr s=44000,1176 d=26000,604
X62 a_9083_31160.t2 inv2_0.out.t3 a_9271_30440 Vss.t232 nfet_03v3
**devattr s=10400,304 d=17600,576
X63 a_23865_30170.t0 a_23785_29218.t4 Vdd.t99 Vdd.t98 pfet_03v3
**devattr s=44000,1176 d=26000,604
X64 a_18743_28100 a_17849_29020 Vss.t67 Vss.t66 nfet_03v3
**devattr s=17600,576 d=10400,304
X65 a_9845_19210 adc_PISO_0.B2.t5 Vss.t531 Vss.t530 nfet_03v3
**devattr s=17600,576 d=10400,304
X66 SARlogic_0.dffrs_3.nand3_6.C.t0 SARlogic_0.dffrs_3.nand3_1.C.t4 Vdd.t41 Vdd.t40 pfet_03v3
**devattr s=44000,1176 d=26000,604
X67 a_42729_31423.t1 a_42729_33628.t4 Vdd.t830 Vdd.t829 pfet_03v3
**devattr s=44000,1176 d=26000,604
X68 a_29583_30440 a_28027_31160.t4 Vdd.t91 Vdd.t90 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X69 SARlogic_0.dffrs_13.Qb.t2 Vdd.t588 Vdd.t590 Vdd.t589 pfet_03v3
**devattr s=26000,604 d=44000,1176
X70 a_23785_29218.t2 a_23785_31423.t4 Vdd.t932 Vdd.t931 pfet_03v3
**devattr s=44000,1176 d=26000,604
X71 Vdd.t157 a_20111_30440 a_20971_29984 Vdd.t156 pfet_03v3
**devattr s=31200,704 d=52800,1376
X72 a_n9429_n2007.t1 Vin1.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t12 Vss.t159 nfet_03v3
**devattr s=15600,404 d=15600,404
X73 a_28027_31160.t2 inv2_0.out.t4 a_28215_30440 Vss.t233 nfet_03v3
**devattr s=10400,304 d=17600,576
X74 SARlogic_0.dffrs_10.nand3_6.C.t0 SARlogic_0.dffrs_10.nand3_1.C Vdd.t291 Vdd.t290 pfet_03v3
**devattr s=44000,1176 d=26000,604
X75 a_42729_33628.t2 Vdd.t585 Vdd.t587 Vdd.t586 pfet_03v3
**devattr s=44000,1176 d=26000,604
X76 a_n4631_33627.t1 a_n4631_31422.t4 a_n4367_35924 Vss.t278 nfet_03v3
**devattr s=10400,304 d=17600,576
X77 a_12401_17004 SARlogic_0.dffrs_11.nand3_8.C.t4 Vss.t538 Vss.t537 nfet_03v3
**devattr s=17600,576 d=10400,304
X78 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t0 a_4501_17004 Vss.t247 nfet_03v3
**devattr s=10400,304 d=17600,576
X79 a_n8305_30439 a_n9861_31159.t4 Vdd.t225 Vdd.t224 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X80 a_n6139_19213 SARlogic_0.dffrs_14.nand3_8.C.t4 a_n6323_19213 Vss.t542 nfet_03v3
**devattr s=10400,304 d=10400,304
X81 a_n201_28099 a_n1095_29019 Vss.t9 Vss.t8 nfet_03v3
**devattr s=17600,576 d=10400,304
X82 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_3.Qb.t5 Vdd.t213 Vdd.t212 pfet_03v3
**devattr s=44000,1176 d=26000,604
X83 adc_PISO_0.B2.t3 SARlogic_0.dffrs_10.Qb Vdd.t435 Vdd.t434 pfet_03v3
**devattr s=26000,604 d=44000,1176
X84 Vdd.t584 Vdd.t582 SARlogic_0.dffrs_13.nand3_8.Z.t3 Vdd.t583 pfet_03v3
**devattr s=26000,604 d=26000,604
X85 SARlogic_0.dffrs_5.Qb.t3 Reset.t7 Vdd.t858 Vdd.t857 pfet_03v3
**devattr s=26000,604 d=44000,1176
X86 a_1167_30439 a_n389_31159.t4 Vdd.t381 Vdd.t380 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X87 SARlogic_0.dffrs_9.nand3_8.C.t2 SARlogic_0.dffrs_9.nand3_8.Z a_4501_19209 Vss.t462 nfet_03v3
**devattr s=10400,304 d=17600,576
X88 SARlogic_0.dffrs_0.nand3_8.C.t0 SARlogic_0.dffrs_0.nand3_6.C.t4 Vdd.t419 Vdd.t418 pfet_03v3
**devattr s=44000,1176 d=26000,604
X89 a_12401_19209 SARlogic_0.dffrs_11.nand3_6.C.t4 Vss.t308 Vss.t307 nfet_03v3
**devattr s=17600,576 d=10400,304
X90 a_33337_31515 a_33257_31423.t4 Vss.t146 Vss.t145 nfet_03v3
**devattr s=17600,576 d=10400,304
X91 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_13.Qb.t4 Vdd.t369 Vdd.t368 pfet_03v3
**devattr s=44000,1176 d=26000,604
X92 SARlogic_0.dffrs_3.nand3_8.C.t0 SARlogic_0.dffrs_3.nand3_8.Z.t5 a_4501_9633 Vss.t48 nfet_03v3
**devattr s=10400,304 d=17600,576
X93 a_10639_30440 a_9083_31160.t4 Vss.t78 Vss.t77 nfet_03v3
**devattr s=17600,576 d=17600,576
X94 Vdd.t59 SARlogic_0.dffrs_5.nand3_8.C.t6 SARlogic_0.dffrs_5.Qb.t1 Vdd.t58 pfet_03v3
**devattr s=26000,604 d=26000,604
X95 Vss.t117 a_29583_30440 a_30255_29264.t3 Vss.t116 nfet_03v3
**devattr s=17600,576 d=17600,576
X96 Vss.t654 adc_PISO_0.2inmux_1.Bit.t5 a_37687_30440 Vss.t653 nfet_03v3
**devattr s=10400,304 d=17600,576
X97 SARlogic_0.dffrs_8.nand3_6.C.t2 adc_PISO_0.B3.t5 Vdd.t926 Vdd.t925 pfet_03v3
**devattr s=26000,604 d=44000,1176
X98 Vdd.t17 a_n1095_29019 a_n389_28819.t0 Vdd.t16 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X99 Vss.t266 a_1167_30439 a_1839_29263.t3 Vss.t265 nfet_03v3
**devattr s=17600,576 d=17600,576
X100 a_5987_9634 SARlogic_0.dffrs_3.nand3_8.C.t4 a_5803_9634 Vss.t142 nfet_03v3
**devattr s=10400,304 d=10400,304
X101 SARlogic_0.dffrs_0.nand3_6.C.t0 SARlogic_0.dffrs_0.nand3_1.C.t4 Vdd.t319 Vdd.t318 pfet_03v3
**devattr s=44000,1176 d=26000,604
X102 SARlogic_0.dffrs_5.nand3_1.C.t3 Vdd.t579 Vdd.t581 Vdd.t580 pfet_03v3
**devattr s=44000,1176 d=26000,604
X103 SARlogic_0.dffrs_3.nand3_1.C.t2 SARlogic_0.dffrs_3.nand3_6.C.t5 Vdd.t832 Vdd.t831 pfet_03v3
**devattr s=26000,604 d=44000,1176
X104 a_20971_29984 a_20111_28100 a_20783_29264.t2 Vdd.t289 pfet_03v3
**devattr s=52800,1376 d=31200,704
X105 a_n3065_31515 adc_PISO_0.2inmux_2.Bit.t4 Vss.t18 Vss.t17 nfet_03v3
**devattr s=17600,576 d=10400,304
X106 SARlogic_0.dffrs_12.Q.t2 SARlogic_0.dffrs_12.Qb Vdd.t159 Vdd.t158 pfet_03v3
**devattr s=26000,604 d=44000,1176
X107 SARlogic_0.dffrs_12.nand3_8.Z Vss.t677 Vdd.t762 Vdd.t761 pfet_03v3
**devattr s=26000,604 d=44000,1176
X108 a_4921_30169.t1 adc_PISO_0.2inmux_2.OUT.t2 a_5105_29309 Vss.t97 nfet_03v3
**devattr s=10400,304 d=17600,576
X109 Vdd.t802 a_27321_29020 a_28027_28820.t3 Vdd.t801 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X110 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t4 Vdd.t219 Vdd.t218 pfet_03v3
**devattr s=26000,604 d=44000,1176
X111 a_n2881_31515 a_n4631_29217.t4 a_n3065_31515 Vss.t623 nfet_03v3
**devattr s=10400,304 d=10400,304
X112 a_12585_7428 Reset.t8 a_12401_7428 Vss.t612 nfet_03v3
**devattr s=10400,304 d=10400,304
X113 SARlogic_0.dffrs_10.Qb Reset.t9 a_10029_19210 Vss.t613 nfet_03v3
**devattr s=10400,304 d=17600,576
X114 a_17849_29020 inv2_0.out.t5 Vdd.t131 Vdd.t130 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X115 SARlogic_0.dffrs_3.nand3_8.Z.t0 SARlogic_0.dffrs_3.nand3_8.C.t5 Vdd.t161 Vdd.t160 pfet_03v3
**devattr s=44000,1176 d=26000,604
X116 a_4317_17004 SARlogic_0.dffrs_9.nand3_8.C.t4 Vss.t190 Vss.t189 nfet_03v3
**devattr s=17600,576 d=10400,304
X117 Vdd.t860 Reset.t10 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t859 pfet_03v3
**devattr s=26000,604 d=26000,604
X118 SARlogic_0.dffrs_7.nand3_8.C.t3 SARlogic_0.dffrs_7.nand3_6.C.t4 Vdd.t149 Vdd.t148 pfet_03v3
**devattr s=44000,1176 d=26000,604
X119 adc_PISO_0.B4.t0 SARlogic_0.dffrs_8.Qb Vdd.t77 Vdd.t76 pfet_03v3
**devattr s=26000,604 d=44000,1176
X120 Vdd.t315 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t6 Vdd.t314 pfet_03v3
**devattr s=10400,304 d=10400,304
X121 a_14393_30170.t0 adc_PISO_0.2inmux_3.OUT.t2 Vdd.t451 Vdd.t450 pfet_03v3
**devattr s=26000,604 d=44000,1176
X122 Vdd.t221 SARlogic_0.dffrs_8.nand3_6.C.t5 adc_PISO_0.B4.t2 Vdd.t220 pfet_03v3
**devattr s=26000,604 d=26000,604
X123 a_4317_19209 SARlogic_0.dffrs_9.nand3_6.C.t5 Vss.t634 Vss.t633 nfet_03v3
**devattr s=17600,576 d=10400,304
X124 a_459_7428 Reset.t11 a_275_7428 Vss.t614 nfet_03v3
**devattr s=10400,304 d=10400,304
X125 a_n9429_n2007.t0 Vin2.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t153 nfet_03v3
**devattr s=15600,404 d=15600,404
X126 Vdd.t704 Clk.t2 SARlogic_0.dffrs_5.nand3_8.C.t3 Vdd.t703 pfet_03v3
**devattr s=26000,604 d=26000,604
X127 a_33257_31423.t3 Clk_piso.t0 Vdd.t642 Vdd.t641 pfet_03v3
**devattr s=26000,604 d=44000,1176
X128 adc_PISO_0.2inmux_1.Bit.t1 Vdd.t576 Vdd.t578 Vdd.t577 pfet_03v3
**devattr s=44000,1176 d=26000,604
X129 SARlogic_0.dffrs_8.nand3_6.C.t0 SARlogic_0.dffrs_8.nand3_1.C Vdd.t51 Vdd.t50 pfet_03v3
**devattr s=44000,1176 d=26000,604
X130 SARlogic_0.dffrs_12.Qb Reset.t12 a_18113_19210 Vss.t615 nfet_03v3
**devattr s=10400,304 d=17600,576
X131 a_14313_29218.t2 a_14393_30170.t4 Vdd.t936 Vdd.t935 pfet_03v3
**devattr s=26000,604 d=44000,1176
X132 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t0 a_n7971_249 a_n8059_341 Vss.t227 nfet_03v3
**devattr s=35200,976 d=20800,504
X133 SARlogic_0.dffrs_3.nand3_1.C.t3 Vdd.t573 Vdd.t575 Vdd.t574 pfet_03v3
**devattr s=44000,1176 d=26000,604
X134 Vdd.t209 SARlogic_0.dffrs_9.nand3_8.C.t5 SARlogic_0.dffrs_9.Qb Vdd.t208 pfet_03v3
**devattr s=26000,604 d=26000,604
X135 SARlogic_0.dffrs_5.nand3_6.C.t2 Clk.t3 a_12585_11838 Vss.t510 nfet_03v3
**devattr s=10400,304 d=17600,576
X136 Vdd.t804 Reset.t13 SARlogic_0.dffrs_5.nand3_6.C.t3 Vdd.t803 pfet_03v3
**devattr s=26000,604 d=26000,604
X137 Vdd.t834 SARlogic_0.dffrs_3.nand3_6.C.t6 SARlogic_0.dffrs_4.d.t3 Vdd.t833 pfet_03v3
**devattr s=26000,604 d=26000,604
X138 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_8.C.t5 Vdd.t884 Vdd.t883 pfet_03v3
**devattr s=44000,1176 d=26000,604
X139 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t1 Vdd.t275 Vdd.t274 pfet_03v3
**devattr s=26000,604 d=44000,1176
X140 a_33257_33628.t1 a_33257_31423.t5 Vdd.t237 Vdd.t236 pfet_03v3
**devattr s=26000,604 d=44000,1176
X141 a_6591_31515 a_4841_29217.t4 a_6407_31515 Vss.t486 nfet_03v3
**devattr s=10400,304 d=10400,304
X142 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_1.Qb.t5 Vdd.t273 Vdd.t272 pfet_03v3
**devattr s=44000,1176 d=26000,604
X143 SARlogic_0.dffrs_14.nand3_6.C.t0 adc_PISO_0.B5.t4 a_n7625_21417 Vss.t298 nfet_03v3
**devattr s=10400,304 d=17600,576
X144 a_n6323_21417 SARlogic_0.dffrs_13.Qb.t5 Vss.t306 Vss.t305 nfet_03v3
**devattr s=17600,576 d=10400,304
X145 a_13887_21414 SARlogic_0.dffrs_4.Qb.t4 Vss.t193 Vss.t192 nfet_03v3
**devattr s=17600,576 d=10400,304
X146 Vdd.t199 SARlogic_0.dffrs_10.nand3_6.C.t5 adc_PISO_0.B2.t0 Vdd.t198 pfet_03v3
**devattr s=26000,604 d=26000,604
X147 Vdd.t806 Reset.t14 SARlogic_0.dffrs_12.nand3_6.C.t3 Vdd.t805 pfet_03v3
**devattr s=26000,604 d=26000,604
X148 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t1 a_n9429_n2007.t7 Vss.t160 nfet_03v3
**devattr s=15600,404 d=15600,404
X149 a_n3583_9633 Clk.t4 a_n3767_9633 Vss.t511 nfet_03v3
**devattr s=10400,304 d=10400,304
X150 a_n6139_9634 SARlogic_0.dffrs_0.nand3_8.C.t4 a_n6323_9634 Vss.t217 nfet_03v3
**devattr s=10400,304 d=10400,304
X151 SARlogic_0.dffrs_8.Qb Reset.t15 a_1945_19210 Vss.t560 nfet_03v3
**devattr s=10400,304 d=17600,576
X152 a_44295_33720 Vdd.t948 Vss.t450 Vss.t449 nfet_03v3
**devattr s=17600,576 d=10400,304
X153 a_n7445_29983 a_n8305_30439 Vdd.t55 Vdd.t54 pfet_03v3
**devattr s=52800,1376 d=31200,704
X154 a_23785_29218.t3 a_23865_30170.t4 a_24049_31515 Vss.t668 nfet_03v3
**devattr s=10400,304 d=17600,576
X155 a_1945_19210 SARlogic_0.dffrs_8.nand3_8.C.t4 a_1761_19210 Vss.t275 nfet_03v3
**devattr s=10400,304 d=10400,304
X156 a_5105_35924 a_4921_30169.t4 a_4921_35924 Vss.t572 nfet_03v3
**devattr s=10400,304 d=10400,304
X157 a_n201_30439 adc_PISO_0.2inmux_2.Bit.t5 Vss.t20 Vss.t19 nfet_03v3
**devattr s=17600,576 d=10400,304
X158 Vdd.t23 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_1.C Vdd.t22 pfet_03v3
**devattr s=26000,604 d=26000,604
X159 SARlogic_0.dffrs_7.nand3_8.C.t0 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t73 Vdd.t72 pfet_03v3
**devattr s=26000,604 d=44000,1176
X160 a_4501_11838 Reset.t16 a_4317_11838 Vss.t561 nfet_03v3
**devattr s=10400,304 d=10400,304
X161 a_42993_33720 Vdd.t949 a_42809_33720 Vss.t448 nfet_03v3
**devattr s=10400,304 d=10400,304
X162 a_4921_35924 Vdd.t950 Vss.t447 Vss.t446 nfet_03v3
**devattr s=17600,576 d=10400,304
X163 adc_PISO_0.dffrs_4.Qb adc_PISO_0.2inmux_1.Bit.t6 Vdd.t920 Vdd.t919 pfet_03v3
**devattr s=44000,1176 d=26000,604
X164 a_459_14043 SARlogic_0.dffrs_2.nand3_8.Z.t4 a_275_14043 Vss.t375 nfet_03v3
**devattr s=10400,304 d=10400,304
X165 a_28215_30440 adc_PISO_0.dffrs_3.Q.t4 Vss.t475 Vss.t474 nfet_03v3
**devattr s=17600,576 d=10400,304
X166 a_39727_29264.t2 a_39055_28100 a_39915_29984 Vdd.t261 pfet_03v3
**devattr s=31200,704 d=52800,1376
X167 a_8543_21414 Reset.t17 a_8359_21414 Vss.t562 nfet_03v3
**devattr s=10400,304 d=10400,304
X168 a_n7809_9633 SARlogic_0.dffrs_0.nand3_6.C.t5 Vss.t349 Vss.t348 nfet_03v3
**devattr s=17600,576 d=10400,304
X169 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq a_n9933_n2099 a_n10021_n2007 Vss.t228 nfet_03v3
**devattr s=26400,776 d=15600,404
X170 SARlogic_0.dffrs_0.nand3_1.C.t2 Vdd.t570 Vdd.t572 Vdd.t571 pfet_03v3
**devattr s=44000,1176 d=26000,604
X171 a_n7809_17007 SARlogic_0.dffrs_14.nand3_8.C.t5 Vss.t544 Vss.t543 nfet_03v3
**devattr s=17600,576 d=10400,304
X172 a_42993_35925 a_42809_30170.t4 a_42809_35925 Vss.t585 nfet_03v3
**devattr s=10400,304 d=10400,304
X173 a_33257_31423.t0 a_33257_33628.t4 Vdd.t217 Vdd.t216 pfet_03v3
**devattr s=44000,1176 d=26000,604
X174 a_28215_28100 adc_PISO_0.B2.t6 a_28027_28820.t1 Vss.t532 nfet_03v3
**devattr s=17600,576 d=10400,304
X175 Vdd.t569 Vdd.t567 a_23865_30170.t3 Vdd.t568 pfet_03v3
**devattr s=26000,604 d=26000,604
X176 a_8543_23619 SARlogic_0.dffrs_10.nand3_8.Z a_8359_23619 Vss.t221 nfet_03v3
**devattr s=10400,304 d=10400,304
X177 a_10029_19210 SARlogic_0.dffrs_10.nand3_8.C.t4 a_9845_19210 Vss.t600 nfet_03v3
**devattr s=10400,304 d=10400,304
X178 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_8.C.t5 Vdd.t850 Vdd.t849 pfet_03v3
**devattr s=44000,1176 d=26000,604
X179 a_33257_33628.t3 Vdd.t564 Vdd.t566 Vdd.t565 pfet_03v3
**devattr s=44000,1176 d=26000,604
X180 Vdd.t644 Clk_piso.t1 a_23785_29218.t1 Vdd.t643 pfet_03v3
**devattr s=26000,604 d=26000,604
X181 adc_PISO_0.B6.t3 SARlogic_0.dffrs_14.Qb a_n6139_21417 Vss.t248 nfet_03v3
**devattr s=10400,304 d=17600,576
X182 a_44295_31516 Piso_out.t4 Vss.t369 Vss.t368 nfet_03v3
**devattr s=17600,576 d=10400,304
X183 a_n4367_35924 a_n4551_30169.t4 a_n4551_35924 Vss.t330 nfet_03v3
**devattr s=10400,304 d=10400,304
X184 a_n4551_30169.t0 a_n4631_29217.t5 Vdd.t874 Vdd.t873 pfet_03v3
**devattr s=44000,1176 d=26000,604
X185 a_12585_17004 Reset.t18 a_12401_17004 Vss.t563 nfet_03v3
**devattr s=10400,304 d=10400,304
X186 a_8377_29020 inv2_0.out.t6 Vss.t110 Vss.t109 nfet_03v3
**devattr s=17600,576 d=17600,576
X187 SARlogic_0.dffrs_0.nand3_8.Z.t1 SARlogic_0.dffrs_0.d.t5 Vdd.t181 Vdd.t180 pfet_03v3
**devattr s=26000,604 d=44000,1176
X188 a_14393_29310 a_14313_29218.t4 Vss.t568 Vss.t567 nfet_03v3
**devattr s=17600,576 d=10400,304
X189 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t2 Vdd.t277 Vdd.t276 pfet_03v3
**devattr s=26000,604 d=44000,1176
X190 a_12585_19209 SARlogic_0.dffrs_12.Q.t4 a_12401_19209 Vss.t336 nfet_03v3
**devattr s=10400,304 d=10400,304
X191 a_39727_29264.t0 a_39055_28100 Vss.t230 Vss.t229 nfet_03v3
**devattr s=17600,576 d=17600,576
X192 a_11499_29984 a_10639_28100 a_11311_29264.t1 Vdd.t153 pfet_03v3
**devattr s=52800,1376 d=31200,704
X193 a_n6555_341 a_n6755_249 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t96 nfet_03v3
**devattr s=20800,504 d=35200,976
X194 Vdd.t3 SARlogic_0.dffrs_5.nand3_8.Z.t4 SARlogic_0.dffrs_5.nand3_1.C.t0 Vdd.t2 pfet_03v3
**devattr s=26000,604 d=26000,604
X195 a_n10151_9634 SARlogic_0.dffrs_13.nand3_8.C.t4 a_n10335_9634 Vss.t295 nfet_03v3
**devattr s=10400,304 d=10400,304
X196 adc_PISO_0.B3.t1 SARlogic_0.dffrs_9.Qb Vdd.t129 Vdd.t128 pfet_03v3
**devattr s=26000,604 d=44000,1176
X197 adc_PISO_0.2inmux_1.Bit.t3 adc_PISO_0.dffrs_4.Qb a_35007_33720 Vss.t670 nfet_03v3
**devattr s=10400,304 d=17600,576
X198 adc_PISO_0.2inmux_0.OUT.t1 a_n7633_29263.t4 Vdd.t403 Vdd.t402 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X199 adc_PISO_0.B5.t0 SARlogic_0.dffrs_0.Qb.t4 Vdd.t43 Vdd.t42 pfet_03v3
**devattr s=44000,1176 d=26000,604
X200 SARlogic_0.dffrs_0.nand3_8.C.t3 SARlogic_0.dffrs_0.nand3_8.Z.t4 Vdd.t892 Vdd.t891 pfet_03v3
**devattr s=26000,604 d=44000,1176
X201 a_36793_29020 inv2_0.out.t7 Vdd.t133 Vdd.t132 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X202 Vdd.t714 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t6 Vdd.t713 pfet_03v3
**devattr s=10400,304 d=10400,304
X203 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t5 Vdd.t776 Vdd.t775 pfet_03v3
**devattr s=26000,604 d=44000,1176
X204 SARlogic_0.dffrs_5.nand3_8.Z.t1 SARlogic_0.dffrs_4.Q.t4 Vdd.t439 Vdd.t438 pfet_03v3
**devattr s=26000,604 d=44000,1176
X205 a_n9429_n2007.t8 Vin2.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t161 nfet_03v3
**devattr s=15600,404 d=15600,404
X206 SARlogic_0.dffrs_0.nand3_6.C.t1 Clk.t5 Vdd.t726 Vdd.t725 pfet_03v3
**devattr s=26000,604 d=44000,1176
X207 a_n4551_30169.t3 adc_PISO_0.2inmux_0.OUT.t2 Vdd.t614 Vdd.t613 pfet_03v3
**devattr s=26000,604 d=44000,1176
X208 SARlogic_0.dffrs_0.Q.t3 Vdd.t561 Vdd.t563 Vdd.t562 pfet_03v3
**devattr s=44000,1176 d=26000,604
X209 adc_PISO_0.dffrs_3.Q.t3 Vdd.t558 Vdd.t560 Vdd.t559 pfet_03v3
**devattr s=44000,1176 d=26000,604
X210 a_18555_28820.t3 adc_PISO_0.B3.t6 Vdd.t928 Vdd.t927 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X211 a_18113_21414 SARlogic_0.dffrs_12.nand3_6.C.t5 a_17929_21414 Vss.t617 nfet_03v3
**devattr s=10400,304 d=10400,304
X212 a_23785_31423.t0 Clk_piso.t2 Vdd.t405 Vdd.t404 pfet_03v3
**devattr s=26000,604 d=44000,1176
X213 SARlogic_0.dffrs_13.nand3_8.Z.t0 Vss.t133 a_n11637_7428 Vss.t134 nfet_03v3
**devattr s=10400,304 d=17600,576
X214 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t67 Vdd.t66 pfet_03v3
**devattr s=17600,576 d=17600,576
X215 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_8.C.t5 Vdd.t323 Vdd.t322 pfet_03v3
**devattr s=44000,1176 d=26000,604
X216 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x3.out Vss.t149 Vss.t148 nfet_03v3
**devattr s=17600,576 d=17600,576
X217 SARlogic_0.dffrs_12.nand3_6.C.t1 Vss.t131 a_16627_21414 Vss.t132 nfet_03v3
**devattr s=10400,304 d=17600,576
X218 a_n3767_9633 SARlogic_0.dffrs_1.nand3_6.C.t4 Vss.t595 Vss.t594 nfet_03v3
**devattr s=17600,576 d=10400,304
X219 Vdd.t239 a_33257_31423.t6 adc_PISO_0.2inmux_1.Bit.t0 Vdd.t238 pfet_03v3
**devattr s=26000,604 d=26000,604
X220 SARlogic_0.dffrs_9.Qb Reset.t19 a_5987_19210 Vss.t564 nfet_03v3
**devattr s=10400,304 d=17600,576
X221 a_23785_33628.t2 a_23785_31423.t5 Vdd.t191 Vdd.t190 pfet_03v3
**devattr s=26000,604 d=44000,1176
X222 Vdd.t808 Reset.t20 SARlogic_0.dffrs_8.nand3_6.C.t1 Vdd.t807 pfet_03v3
**devattr s=26000,604 d=26000,604
X223 SARlogic_0.dffrs_14.Qb adc_PISO_0.B6.t4 Vdd.t930 Vdd.t929 pfet_03v3
**devattr s=44000,1176 d=26000,604
X224 a_n2281_19210 adc_PISO_0.B5.t5 Vss.t300 Vss.t299 nfet_03v3
**devattr s=17600,576 d=10400,304
X225 a_n3583_14043 SARlogic_0.dffrs_1.nand3_8.Z.t4 a_n3767_14043 Vss.t329 nfet_03v3
**devattr s=10400,304 d=10400,304
X226 a_n7633_29263.t2 a_n8305_28099 a_n7445_29983 Vdd.t123 pfet_03v3
**devattr s=31200,704 d=52800,1376
X227 SARlogic_0.dffrs_2.nand3_8.Z.t1 SARlogic_0.dffrs_2.d.t4 Vdd.t455 Vdd.t454 pfet_03v3
**devattr s=26000,604 d=44000,1176
X228 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t6 a_16627_23619 Vss.t618 nfet_03v3
**devattr s=10400,304 d=17600,576
X229 SARlogic_0.dffrs_11.Qb adc_PISO_0.B1.t5 Vdd.t798 Vdd.t797 pfet_03v3
**devattr s=44000,1176 d=26000,604
X230 adc_PISO_0.dffrs_4.Qb Vdd.t951 a_35007_31516 Vss.t445 nfet_03v3
**devattr s=10400,304 d=17600,576
X231 SARlogic_0.dffrs_5.Q.t3 Vdd.t555 Vdd.t557 Vdd.t556 pfet_03v3
**devattr s=44000,1176 d=26000,604
X232 Vdd.t810 Reset.t21 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t809 pfet_03v3
**devattr s=26000,604 d=26000,604
X233 a_n389_31159.t3 inv2_0.out.t8 Vdd.t135 Vdd.t134 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X234 a_n7625_21417 Reset.t22 a_n7809_21417 Vss.t494 nfet_03v3
**devattr s=10400,304 d=10400,304
X235 Vdd.t7 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_1.C Vdd.t6 pfet_03v3
**devattr s=26000,604 d=26000,604
X236 adc_PISO_0.dffrs_0.Qb Vdd.t952 a_n2881_31515 Vss.t444 nfet_03v3
**devattr s=10400,304 d=17600,576
X237 a_1761_21414 SARlogic_0.dffrs_1.Qb.t6 Vss.t35 Vss.t34 nfet_03v3
**devattr s=17600,576 d=10400,304
X238 a_n10567_29019 inv2_0.out.t9 Vss.t112 Vss.t111 nfet_03v3
**devattr s=17600,576 d=17600,576
X239 a_n201_28099 adc_PISO_0.B5.t6 a_n389_28819.t1 Vss.t154 nfet_03v3
**devattr s=17600,576 d=10400,304
X240 SARlogic_0.dffrs_12.Q.t0 SARlogic_0.dffrs_5.Qb.t5 Vdd.t37 Vdd.t36 pfet_03v3
**devattr s=44000,1176 d=26000,604
X241 a_n11821_14043 Reset.t23 Vss.t496 Vss.t495 nfet_03v3
**devattr s=17600,576 d=10400,304
X242 a_33521_33720 Vdd.t953 a_33337_33720 Vss.t443 nfet_03v3
**devattr s=10400,304 d=10400,304
X243 Vdd.t728 Clk.t6 SARlogic_0.dffrs_4.nand3_8.C.t3 Vdd.t727 pfet_03v3
**devattr s=26000,604 d=26000,604
X244 SARlogic_0.dffrs_1.nand3_8.Z.t1 SARlogic_0.dffrs_0.Q.t4 Vdd.t465 Vdd.t464 pfet_03v3
**devattr s=26000,604 d=44000,1176
X245 SARlogic_0.dffrs_0.Q.t0 SARlogic_0.dffrs_0.Qb.t5 Vdd.t45 Vdd.t44 pfet_03v3
**devattr s=26000,604 d=44000,1176
X246 adc_PISO_0.dffrs_3.Qb adc_PISO_0.dffrs_3.Q.t5 Vdd.t656 Vdd.t655 pfet_03v3
**devattr s=44000,1176 d=26000,604
X247 a_30255_29264.t1 a_29583_28100 a_30443_29984 Vdd.t11 pfet_03v3
**devattr s=31200,704 d=52800,1376
X248 a_5803_11838 Vdd.t954 Vss.t442 Vss.t441 nfet_03v3
**devattr s=17600,576 d=10400,304
X249 a_4841_33627.t1 a_4841_31422.t5 a_5105_35924 Vss.t267 nfet_03v3
**devattr s=10400,304 d=17600,576
X250 a_1839_29263.t1 a_1167_28099 a_2027_29983 Vdd.t109 pfet_03v3
**devattr s=31200,704 d=52800,1376
X251 a_12401_11838 SARlogic_0.dffrs_5.nand3_1.C.t5 Vss.t304 Vss.t303 nfet_03v3
**devattr s=17600,576 d=10400,304
X252 SARlogic_0.dffrs_3.nand3_6.C.t1 Clk.t7 a_4501_11838 Vss.t522 nfet_03v3
**devattr s=10400,304 d=17600,576
X253 Vdd.t668 Reset.t24 SARlogic_0.dffrs_4.nand3_6.C.t2 Vdd.t667 pfet_03v3
**devattr s=26000,604 d=26000,604
X254 a_33521_35925 a_33337_30170.t6 a_33337_35925 Vss.t626 nfet_03v3
**devattr s=10400,304 d=10400,304
X255 a_42809_30170.t1 adc_PISO_0.2inmux_1.OUT.t2 Vdd.t427 Vdd.t426 pfet_03v3
**devattr s=26000,604 d=44000,1176
X256 inv2_0.out.t0 Load.t0 Vss.t351 Vss.t350 nfet_03v3
**devattr s=17600,576 d=17600,576
X257 Vdd.t554 Vdd.t552 a_14393_30170.t2 Vdd.t553 pfet_03v3
**devattr s=26000,604 d=26000,604
X258 Comp_out.t3 a_n10831_4320 Vss.t264 Vss.t263 nfet_03v3
**devattr s=17000,540 d=9350,280
X259 Vdd.t263 a_33257_29218.t4 adc_PISO_0.dffrs_4.Qb Vdd.t262 pfet_03v3
**devattr s=26000,604 d=26000,604
X260 SARlogic_0.dffrs_11.nand3_8.C.t1 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t173 Vdd.t172 pfet_03v3
**devattr s=26000,604 d=44000,1176
X261 SARlogic_0.dffrs_10.nand3_6.C.t1 adc_PISO_0.B1.t6 a_8543_21414 Vss.t553 nfet_03v3
**devattr s=10400,304 d=17600,576
X262 a_9845_21414 SARlogic_0.dffrs_3.Qb.t6 Vss.t196 Vss.t195 nfet_03v3
**devattr s=17600,576 d=10400,304
X263 a_16443_21414 SARlogic_0.dffrs_12.nand3_1.C Vss.t33 Vss.t32 nfet_03v3
**devattr s=17600,576 d=10400,304
X264 a_42729_29218.t2 a_42809_30170.t5 Vdd.t836 Vdd.t835 pfet_03v3
**devattr s=26000,604 d=44000,1176
X265 a_8359_7428 SARlogic_0.dffrs_4.nand3_8.C.t6 Vss.t481 Vss.t480 nfet_03v3
**devattr s=17600,576 d=10400,304
X266 Vdd.t407 Clk_piso.t3 a_14313_29218.t0 Vdd.t406 pfet_03v3
**devattr s=26000,604 d=26000,604
X267 SARlogic_0.dffrs_14.Qb Reset.t25 Vdd.t670 Vdd.t669 pfet_03v3
**devattr s=26000,604 d=44000,1176
X268 inv2_0.out.t1 Load.t1 inv2_0.vdd inv2_0.vdd pfet_03v3
**devattr s=52800,1376 d=52800,1376
X269 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t6 a_8543_23619 Vss.t177 nfet_03v3
**devattr s=10400,304 d=17600,576
X270 a_16443_23619 SARlogic_0.dffrs_5.Qb.t6 Vss.t26 Vss.t25 nfet_03v3
**devattr s=17600,576 d=10400,304
X271 a_17929_19210 SARlogic_0.dffrs_12.Q.t5 Vss.t547 Vss.t546 nfet_03v3
**devattr s=17600,576 d=10400,304
X272 a_n9429_n2007.t9 Vin2.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t159 nfet_03v3
**devattr s=15600,404 d=15600,404
X273 a_6407_31515 adc_PISO_0.dffrs_1.Q.t5 Vss.t628 Vss.t627 nfet_03v3
**devattr s=17600,576 d=10400,304
X274 a_18555_31160.t2 inv2_0.out.t10 a_18743_30440 Vss.t113 nfet_03v3
**devattr s=10400,304 d=17600,576
X275 Vdd.t680 adc_PISO_0.B2.t7 SARlogic_0.dffrs_9.nand3_8.C.t1 Vdd.t679 pfet_03v3
**devattr s=26000,604 d=26000,604
X276 Vdd.t672 Reset.t26 SARlogic_0.dffrs_0.nand3_8.Z.t3 Vdd.t671 pfet_03v3
**devattr s=26000,604 d=26000,604
X277 a_n6139_21417 SARlogic_0.dffrs_14.nand3_6.C.t6 a_n6323_21417 Vss.t533 nfet_03v3
**devattr s=10400,304 d=10400,304
X278 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t11 Vss.t516 Vss.t515 nfet_03v3
**devattr s=35200,976 d=35200,976
X279 SARlogic_0.dffrs_13.nand3_1.C.t0 SARlogic_0.dffrs_13.nand3_6.C.t4 a_n11637_14043 Vss.t469 nfet_03v3
**devattr s=10400,304 d=17600,576
X280 SARlogic_0.dffrs_0.nand3_1.C.t0 SARlogic_0.dffrs_0.nand3_6.C.t6 Vdd.t421 Vdd.t420 pfet_03v3
**devattr s=26000,604 d=44000,1176
X281 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t3 a_n7625_17007 Vss.t313 nfet_03v3
**devattr s=10400,304 d=17600,576
X282 adc_PISO_0.2inmux_5.OUT.t1 a_30255_29264.t5 Vdd.t205 Vdd.t204 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X283 a_n10335_9634 SARlogic_0.dffrs_0.d.t6 Vss.t641 Vss.t640 nfet_03v3
**devattr s=17600,576 d=10400,304
X284 a_42809_33720 a_42729_33628.t5 Vss.t578 Vss.t577 nfet_03v3
**devattr s=17600,576 d=10400,304
X285 Vdd.t551 Vdd.t549 a_4921_30169.t3 Vdd.t550 pfet_03v3
**devattr s=26000,604 d=26000,604
X286 a_4317_11838 SARlogic_0.dffrs_3.nand3_1.C.t5 Vss.t31 Vss.t30 nfet_03v3
**devattr s=17600,576 d=10400,304
X287 a_23865_31515 a_23785_31423.t6 Vss.t168 Vss.t167 nfet_03v3
**devattr s=17600,576 d=10400,304
X288 a_4921_30169.t2 a_4841_29217.t5 Vdd.t441 Vdd.t440 pfet_03v3
**devattr s=44000,1176 d=26000,604
X289 a_42993_29310 Vdd.t955 a_42809_29310 Vss.t440 nfet_03v3
**devattr s=10400,304 d=10400,304
X290 Vss.t138 a_20111_30440 a_20783_29264.t0 Vss.t137 nfet_03v3
**devattr s=17600,576 d=17600,576
X291 a_8359_21414 SARlogic_0.dffrs_10.nand3_1.C Vss.t254 Vss.t253 nfet_03v3
**devattr s=17600,576 d=10400,304
X292 a_42809_35925 Vdd.t956 Vss.t439 Vss.t438 nfet_03v3
**devattr s=17600,576 d=10400,304
X293 a_n9673_28099 a_n10567_29019 Vss.t93 Vss.t92 nfet_03v3
**devattr s=17600,576 d=10400,304
X294 a_8543_17004 Reset.t27 a_8359_17004 Vss.t497 nfet_03v3
**devattr s=10400,304 d=10400,304
X295 adc_PISO_0.B2.t2 SARlogic_0.dffrs_10.Qb a_10029_21414 Vss.t358 nfet_03v3
**devattr s=10400,304 d=17600,576
X296 a_8359_23619 SARlogic_0.dffrs_3.Qb.t7 Vss.t198 Vss.t197 nfet_03v3
**devattr s=17600,576 d=10400,304
X297 a_n11637_7428 Vdd.t957 a_n11821_7428 Vss.t437 nfet_03v3
**devattr s=10400,304 d=10400,304
X298 Vdd.t79 a_17849_29020 a_18555_28820.t0 Vdd.t78 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X299 Vdd.t674 Reset.t28 SARlogic_0.dffrs_7.nand3_6.C.t3 Vdd.t673 pfet_03v3
**devattr s=26000,604 d=26000,604
X300 Vdd.t730 Clk.t8 SARlogic_0.dffrs_0.nand3_8.C.t2 Vdd.t729 pfet_03v3
**devattr s=26000,604 d=26000,604
X301 a_n201_30439 inv2_0.out.t11 a_n389_31159.t2 Vss.t114 nfet_03v3
**devattr s=17600,576 d=10400,304
X302 a_20111_28100 a_18555_28820.t4 Vss.t360 Vss.t359 nfet_03v3
**devattr s=17600,576 d=17600,576
X303 a_8543_19209 adc_PISO_0.B1.t7 a_8359_19209 Vss.t554 nfet_03v3
**devattr s=10400,304 d=10400,304
X304 Vdd.t111 a_n10567_29019 a_n9861_28819.t0 Vdd.t110 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X305 Vdd.t784 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_1.C Vdd.t783 pfet_03v3
**devattr s=26000,604 d=26000,604
X306 a_n7809_23622 SARlogic_0.dffrs_13.Qb.t6 Vss.t164 Vss.t163 nfet_03v3
**devattr s=17600,576 d=10400,304
X307 Vss.t630 adc_PISO_0.dffrs_1.Q.t6 a_9271_30440 Vss.t629 nfet_03v3
**devattr s=10400,304 d=17600,576
X308 a_37499_28820.t2 adc_PISO_0.B1.t8 a_37687_28100 Vss.t555 nfet_03v3
**devattr s=10400,304 d=17600,576
X309 Vdd.t71 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_1.C Vdd.t70 pfet_03v3
**devattr s=26000,604 d=26000,604
X310 SARlogic_0.dffrs_8.nand3_6.C.t3 adc_PISO_0.B3.t7 a_459_21414 Vss.t662 nfet_03v3
**devattr s=10400,304 d=17600,576
X311 Vdd.t95 SARlogic_0.dffrs_12.nand3_8.C.t6 SARlogic_0.dffrs_12.Qb Vdd.t94 pfet_03v3
**devattr s=26000,604 d=26000,604
X312 Vdd.t548 Vdd.t546 a_n4551_30169.t2 Vdd.t547 pfet_03v3
**devattr s=26000,604 d=26000,604
X313 a_12401_9633 SARlogic_0.dffrs_5.nand3_6.C.t5 Vss.t223 Vss.t222 nfet_03v3
**devattr s=17600,576 d=10400,304
X314 a_n7809_11838 SARlogic_0.dffrs_0.nand3_1.C.t5 Vss.t273 Vss.t272 nfet_03v3
**devattr s=17600,576 d=10400,304
X315 Vdd.t676 Reset.t29 SARlogic_0.dffrs_0.nand3_6.C.t3 Vdd.t675 pfet_03v3
**devattr s=26000,604 d=26000,604
X316 Vdd.t712 SARlogic_0.dffrs_4.nand3_8.Z.t5 SARlogic_0.dffrs_4.nand3_1.C.t0 Vdd.t711 pfet_03v3
**devattr s=26000,604 d=26000,604
X317 a_1761_9634 SARlogic_0.dffrs_2.Q.t4 Vss.t334 Vss.t333 nfet_03v3
**devattr s=17600,576 d=10400,304
X318 Vdd.t193 a_23785_31423.t7 adc_PISO_0.dffrs_3.Q.t0 Vdd.t192 pfet_03v3
**devattr s=26000,604 d=26000,604
X319 SARlogic_0.dffrs_12.Q.t1 SARlogic_0.dffrs_12.Qb a_18113_21414 Vss.t139 nfet_03v3
**devattr s=10400,304 d=17600,576
X320 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t6 a_459_23619 Vss.t202 nfet_03v3
**devattr s=10400,304 d=17600,576
X321 Vdd.t678 Reset.t30 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t677 pfet_03v3
**devattr s=26000,604 d=26000,604
X322 Vdd.t732 Clk.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vdd.t731 pfet_03v3
**devattr s=14080,496 d=14080,496
X323 a_275_9633 SARlogic_0.dffrs_2.nand3_6.C.t5 Vss.t318 Vss.t317 nfet_03v3
**devattr s=17600,576 d=10400,304
X324 adc_PISO_0.dffrs_1.Q.t0 adc_PISO_0.dffrs_1.Qb Vdd.t15 Vdd.t14 pfet_03v3
**devattr s=26000,604 d=44000,1176
X325 a_4317_7428 SARlogic_0.dffrs_3.nand3_8.C.t6 Vss.t144 Vss.t143 nfet_03v3
**devattr s=17600,576 d=10400,304
X326 a_n3767_14043 Vdd.t958 Vss.t436 Vss.t435 nfet_03v3
**devattr s=17600,576 d=10400,304
X327 SARlogic_0.dffrs_8.Qb adc_PISO_0.B4.t7 Vdd.t87 Vdd.t86 pfet_03v3
**devattr s=44000,1176 d=26000,604
X328 a_30443_29984 a_29583_30440 Vdd.t143 Vdd.t142 pfet_03v3
**devattr s=52800,1376 d=31200,704
X329 SARlogic_0.dffrs_2.Q.t1 Vdd.t543 Vdd.t545 Vdd.t544 pfet_03v3
**devattr s=44000,1176 d=26000,604
X330 adc_PISO_0.B4.t1 SARlogic_0.dffrs_8.Qb a_1945_21414 Vss.t63 nfet_03v3
**devattr s=10400,304 d=17600,576
X331 a_2027_29983 a_1167_30439 Vdd.t305 Vdd.t304 pfet_03v3
**devattr s=52800,1376 d=31200,704
X332 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t11 Vin1.t1 a_n9429_n2007.t2 Vss.t160 nfet_03v3
**devattr s=15600,404 d=15600,404
X333 a_9271_30440 inv2_0.out.t12 a_9083_31160.t1 Vss.t98 nfet_03v3
**devattr s=17600,576 d=10400,304
X334 a_39055_28100 a_37499_28820.t4 Vss.t460 Vss.t459 nfet_03v3
**devattr s=17600,576 d=17600,576
X335 Vdd.t151 SARlogic_0.dffrs_7.nand3_6.C.t5 adc_PISO_0.B5.t1 Vdd.t150 pfet_03v3
**devattr s=26000,604 d=26000,604
X336 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t3 Vss.t517 nfet_03v3
**devattr s=20800,504 d=20800,504
X337 a_n7633_29263.t3 a_n8305_28099 Vss.t105 Vss.t104 nfet_03v3
**devattr s=17600,576 d=17600,576
X338 a_1945_21414 SARlogic_0.dffrs_8.nand3_6.C.t7 a_1761_21414 Vss.t203 nfet_03v3
**devattr s=10400,304 d=10400,304
X339 SARlogic_0.dffrs_3.Qb.t0 SARlogic_0.dffrs_4.d.t5 Vdd.t878 Vdd.t877 pfet_03v3
**devattr s=44000,1176 d=26000,604
X340 a_33257_31423.t1 Clk_piso.t4 a_33521_33720 Vss.t339 nfet_03v3
**devattr s=10400,304 d=17600,576
X341 a_34823_33720 Vdd.t959 Vss.t434 Vss.t433 nfet_03v3
**devattr s=17600,576 d=10400,304
X342 adc_PISO_0.B5.t2 SARlogic_0.dffrs_7.Qb Vdd.t888 Vdd.t887 pfet_03v3
**devattr s=26000,604 d=44000,1176
X343 SARlogic_0.dffrs_4.nand3_8.C.t1 SARlogic_0.dffrs_4.nand3_8.Z.t6 Vdd.t401 Vdd.t400 pfet_03v3
**devattr s=26000,604 d=44000,1176
X344 a_14313_29218.t1 a_14393_30170.t5 a_14577_31515 Vss.t669 nfet_03v3
**devattr s=10400,304 d=17600,576
X345 a_275_21414 SARlogic_0.dffrs_8.nand3_1.C Vss.t40 Vss.t39 nfet_03v3
**devattr s=17600,576 d=10400,304
X346 a_9083_31160.t3 inv2_0.out.t13 Vdd.t117 Vdd.t116 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X347 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t10 Vdd.t229 Vdd.t228 pfet_03v3
**devattr s=10400,304 d=10400,304
X348 Vdd.t207 SARlogic_0.dffrs_0.nand3_6.C.t7 SARlogic_0.dffrs_0.Q.t2 Vdd.t206 pfet_03v3
**devattr s=26000,604 d=26000,604
X349 Vdd.t101 a_23785_29218.t5 adc_PISO_0.dffrs_3.Qb Vdd.t100 pfet_03v3
**devattr s=26000,604 d=26000,604
X350 SARlogic_0.dffrs_10.Qb adc_PISO_0.B2.t8 Vdd.t682 Vdd.t681 pfet_03v3
**devattr s=44000,1176 d=26000,604
X351 a_5987_11838 SARlogic_0.dffrs_3.nand3_6.C.t7 a_5803_11838 Vss.t579 nfet_03v3
**devattr s=10400,304 d=10400,304
X352 a_n1095_29019 inv2_0.out.t14 Vss.t100 Vss.t99 nfet_03v3
**devattr s=17600,576 d=17600,576
X353 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vss.t95 Vss.t94 nfet_03v3
**devattr s=9350,280 d=17000,540
X354 a_12585_11838 Reset.t31 a_12401_11838 Vss.t524 nfet_03v3
**devattr s=10400,304 d=10400,304
X355 SARlogic_0.dffrs_4.Q.t0 Vdd.t540 Vdd.t542 Vdd.t541 pfet_03v3
**devattr s=44000,1176 d=26000,604
X356 SARlogic_0.dffrs_4.nand3_6.C.t1 Clk.t10 Vdd.t734 Vdd.t733 pfet_03v3
**devattr s=26000,604 d=44000,1176
X357 a_33257_33628.t2 a_33257_31423.t7 a_33521_35925 Vss.t211 nfet_03v3
**devattr s=10400,304 d=17600,576
X358 a_18743_30440 adc_PISO_0.dffrs_2.Q.t4 Vss.t246 Vss.t245 nfet_03v3
**devattr s=17600,576 d=10400,304
X359 a_275_23619 SARlogic_0.dffrs_1.Qb.t7 Vss.t37 Vss.t36 nfet_03v3
**devattr s=17600,576 d=10400,304
X360 a_n6389_n1044 a_n6589_n1136 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t385 nfet_03v3
**devattr s=15600,404 d=26400,776
X361 a_23785_31423.t3 a_23785_33628.t4 Vdd.t654 Vdd.t653 pfet_03v3
**devattr s=44000,1176 d=26000,604
X362 a_28027_31160.t3 inv2_0.out.t15 Vdd.t119 Vdd.t118 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X363 a_10029_21414 SARlogic_0.dffrs_10.nand3_6.C.t7 a_9845_21414 Vss.t178 nfet_03v3
**devattr s=10400,304 d=10400,304
X364 a_16627_21414 Reset.t32 a_16443_21414 Vss.t525 nfet_03v3
**devattr s=10400,304 d=10400,304
X365 a_n9673_30439 Vss.t128 Vss.t130 Vss.t129 nfet_03v3
**devattr s=17600,576 d=10400,304
X366 Vdd.t786 SARlogic_0.dffrs_14.nand3_8.C.t6 SARlogic_0.dffrs_14.Qb Vdd.t785 pfet_03v3
**devattr s=26000,604 d=26000,604
X367 a_n2097_19210 SARlogic_0.dffrs_7.nand3_8.C.t4 a_n2281_19210 Vss.t647 nfet_03v3
**devattr s=10400,304 d=10400,304
X368 SARlogic_0.dffrs_1.nand3_1.C.t1 SARlogic_0.dffrs_1.nand3_6.C.t5 a_n3583_14043 Vss.t596 nfet_03v3
**devattr s=10400,304 d=17600,576
X369 SARlogic_0.dffrs_12.nand3_8.Z Vss.t126 a_16627_17004 Vss.t127 nfet_03v3
**devattr s=10400,304 d=17600,576
X370 a_23785_33628.t3 Vdd.t537 Vdd.t539 Vdd.t538 pfet_03v3
**devattr s=44000,1176 d=26000,604
X371 a_1839_29263.t2 a_1167_28099 Vss.t89 Vss.t88 nfet_03v3
**devattr s=17600,576 d=17600,576
X372 adc_PISO_0.2inmux_4.OUT.t0 a_20783_29264.t4 Vss.t216 Vss.t215 nfet_03v3
**devattr s=17600,576 d=17600,576
X373 a_16627_23619 SARlogic_0.dffrs_12.nand3_8.Z a_16443_23619 Vss.t13 nfet_03v3
**devattr s=10400,304 d=10400,304
X374 SARlogic_0.dffrs_7.Qb Reset.t33 a_n2097_19210 Vss.t526 nfet_03v3
**devattr s=10400,304 d=17600,576
X375 SARlogic_0.dffrs_9.nand3_8.C.t3 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t608 Vdd.t607 pfet_03v3
**devattr s=26000,604 d=44000,1176
X376 SARlogic_0.dffrs_11.nand3_8.C.t2 SARlogic_0.dffrs_11.nand3_6.C.t5 Vdd.t373 Vdd.t372 pfet_03v3
**devattr s=44000,1176 d=26000,604
X377 Vdd.t738 Reset.t34 SARlogic_0.dffrs_4.nand3_8.Z.t3 Vdd.t737 pfet_03v3
**devattr s=26000,604 d=26000,604
X378 a_34823_31516 adc_PISO_0.2inmux_1.Bit.t7 Vss.t656 Vss.t655 nfet_03v3
**devattr s=17600,576 d=10400,304
X379 a_9271_28100 a_8377_29020 Vss.t171 Vss.t170 nfet_03v3
**devattr s=17600,576 d=10400,304
X380 SARlogic_0.dffrs_12.nand3_8.C.t0 SARlogic_0.dffrs_12.nand3_8.Z a_16627_19209 Vss.t12 nfet_03v3
**devattr s=10400,304 d=17600,576
X381 Vdd.t894 SARlogic_0.dffrs_0.nand3_8.Z.t5 SARlogic_0.dffrs_0.nand3_1.C.t3 Vdd.t893 pfet_03v3
**devattr s=26000,604 d=26000,604
X382 a_10639_30440 a_9083_31160.t5 Vdd.t93 Vdd.t92 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X383 a_27321_29020 inv2_0.out.t16 Vss.t102 Vss.t101 nfet_03v3
**devattr s=17600,576 d=17600,576
X384 SARlogic_0.dffrs_4.nand3_8.C.t2 SARlogic_0.dffrs_4.nand3_6.C.t4 Vdd.t423 Vdd.t422 pfet_03v3
**devattr s=44000,1176 d=26000,604
X385 a_n11637_14043 SARlogic_0.dffrs_13.nand3_8.Z.t4 a_n11821_14043 Vss.t281 nfet_03v3
**devattr s=10400,304 d=10400,304
X386 a_n7625_17007 Reset.t35 a_n7809_17007 Vss.t527 nfet_03v3
**devattr s=10400,304 d=10400,304
X387 a_33337_33720 a_33257_33628.t5 Vss.t200 Vss.t199 nfet_03v3
**devattr s=17600,576 d=10400,304
X388 a_n9861_28819.t3 adc_PISO_0.B6.t5 a_n9673_28099 Vss.t573 nfet_03v3
**devattr s=10400,304 d=17600,576
X389 a_33521_29310 Vdd.t960 a_33337_29310 Vss.t432 nfet_03v3
**devattr s=10400,304 d=10400,304
X390 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t8 Clk.t11 Vdd.t736 Vdd.t735 pfet_03v3
**devattr s=14080,496 d=14080,496
X391 a_4921_30169.t0 adc_PISO_0.2inmux_2.OUT.t3 Vdd.t9 Vdd.t8 pfet_03v3
**devattr s=26000,604 d=44000,1176
X392 SARlogic_0.dffrs_4.nand3_6.C.t3 SARlogic_0.dffrs_4.nand3_1.C.t4 Vdd.t872 Vdd.t871 pfet_03v3
**devattr s=44000,1176 d=26000,604
X393 a_33337_35925 Vdd.t961 Vss.t431 Vss.t430 nfet_03v3
**devattr s=17600,576 d=10400,304
X394 a_24049_31515 Clk_piso.t5 a_23865_31515 Vss.t476 nfet_03v3
**devattr s=10400,304 d=10400,304
X395 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t14 Clk.t12 Vdd.t696 Vdd.t695 pfet_03v3
**devattr s=14080,496 d=14080,496
X396 a_n9861_28819.t1 adc_PISO_0.B6.t6 Vdd.t828 Vdd.t827 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X397 a_37687_28100 a_36793_29020 Vss.t58 Vss.t57 nfet_03v3
**devattr s=17600,576 d=10400,304
X398 SARlogic_0.dffrs_10.Qb Reset.t36 Vdd.t740 Vdd.t739 pfet_03v3
**devattr s=26000,604 d=44000,1176
X399 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t2 Vss.t206 nfet_03v3
**devattr s=20800,504 d=20800,504
X400 a_12585_9633 Clk.t13 a_12401_9633 Vss.t505 nfet_03v3
**devattr s=10400,304 d=10400,304
X401 SARlogic_0.dffrs_4.Q.t3 SARlogic_0.dffrs_4.Qb.t5 Vdd.t910 Vdd.t909 pfet_03v3
**devattr s=26000,604 d=44000,1176
X402 Vdd.t742 Reset.t37 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t741 pfet_03v3
**devattr s=26000,604 d=26000,604
X403 SARlogic_0.dffrs_2.nand3_8.C.t1 SARlogic_0.dffrs_2.nand3_8.Z.t5 Vdd.t453 Vdd.t452 pfet_03v3
**devattr s=26000,604 d=44000,1176
X404 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t4 a_8543_17004 Vss.t314 nfet_03v3
**devattr s=10400,304 d=17600,576
X405 a_16443_17004 SARlogic_0.dffrs_12.nand3_8.C.t7 Vss.t80 Vss.t79 nfet_03v3
**devattr s=17600,576 d=10400,304
X406 a_1945_9634 SARlogic_0.dffrs_2.nand3_8.C.t5 a_1761_9634 Vss.t176 nfet_03v3
**devattr s=10400,304 d=10400,304
X407 adc_PISO_0.B1.t1 SARlogic_0.dffrs_11.Qb Vdd.t169 Vdd.t168 pfet_03v3
**devattr s=26000,604 d=44000,1176
X408 a_13887_9634 SARlogic_0.dffrs_5.Q.t4 Vss.t11 Vss.t10 nfet_03v3
**devattr s=17600,576 d=10400,304
X409 SARlogic_0.dffrs_7.nand3_6.C.t2 SARlogic_0.dffrs_7.nand3_1.C Vdd.t125 Vdd.t124 pfet_03v3
**devattr s=44000,1176 d=26000,604
X410 SARlogic_0.dffrs_0.nand3_8.Z.t0 SARlogic_0.dffrs_0.d.t7 a_n7625_7428 Vss.t642 nfet_03v3
**devattr s=10400,304 d=17600,576
X411 SARlogic_0.dffrs_9.nand3_8.C.t0 SARlogic_0.dffrs_9.nand3_6.C.t6 Vdd.t900 Vdd.t899 pfet_03v3
**devattr s=44000,1176 d=26000,604
X412 SARlogic_0.dffrs_2.nand3_6.C.t0 Clk.t14 Vdd.t698 Vdd.t697 pfet_03v3
**devattr s=26000,604 d=44000,1176
X413 a_16443_19209 SARlogic_0.dffrs_12.nand3_6.C.t7 Vss.t620 Vss.t619 nfet_03v3
**devattr s=17600,576 d=10400,304
X414 SARlogic_0.dffrs_10.nand3_8.C.t1 SARlogic_0.dffrs_10.nand3_8.Z a_8543_19209 Vss.t220 nfet_03v3
**devattr s=10400,304 d=17600,576
X415 Vdd.t375 SARlogic_0.dffrs_11.nand3_6.C.t6 adc_PISO_0.B1.t3 Vdd.t374 pfet_03v3
**devattr s=26000,604 d=26000,604
X416 a_n9429_n2007.t3 Vin1.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t10 Vss.t161 nfet_03v3
**devattr s=15600,404 d=15600,404
X417 SARlogic_0.dffrs_12.Qb Reset.t38 Vdd.t744 Vdd.t743 pfet_03v3
**devattr s=26000,604 d=44000,1176
X418 a_459_9633 Clk.t15 a_275_9633 Vss.t506 nfet_03v3
**devattr s=10400,304 d=10400,304
X419 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_0.Qb.t6 Vdd.t265 Vdd.t264 pfet_03v3
**devattr s=44000,1176 d=26000,604
X420 SARlogic_0.dffrs_13.nand3_8.Z.t2 SARlogic_0.dffrs_13.nand3_8.C.t5 Vdd.t365 Vdd.t364 pfet_03v3
**devattr s=44000,1176 d=26000,604
X421 SARlogic_0.dffrs_4.nand3_1.C.t3 SARlogic_0.dffrs_4.nand3_6.C.t5 Vdd.t425 Vdd.t424 pfet_03v3
**devattr s=26000,604 d=44000,1176
X422 a_14313_31423.t1 Clk_piso.t6 Vdd.t636 Vdd.t635 pfet_03v3
**devattr s=26000,604 d=44000,1176
X423 Vss.t208 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t12 comparator_no_offsetcal_0.x5.out Vss.t207 nfet_03v3
**devattr s=35200,976 d=35200,976
X424 adc_PISO_0.dffrs_3.Q.t2 adc_PISO_0.dffrs_3.Qb Vdd.t269 Vdd.t268 pfet_03v3
**devattr s=26000,604 d=44000,1176
X425 adc_PISO_0.B3.t0 SARlogic_0.dffrs_9.Qb a_5987_21414 Vss.t108 nfet_03v3
**devattr s=10400,304 d=17600,576
X426 a_8377_29020 inv2_0.out.t17 Vdd.t121 Vdd.t120 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X427 a_n2281_21414 SARlogic_0.dffrs_0.Qb.t7 Vss.t238 Vss.t237 nfet_03v3
**devattr s=17600,576 d=10400,304
X428 Comp_out.t2 a_n10831_4320 Vss.t262 Vss.t261 nfet_03v3
**devattr s=9350,280 d=9350,280
X429 Comp_out.t6 a_n10831_4320 Vdd.t299 Vdd.t298 pfet_03v3
**devattr s=34000,880 d=18700,450
X430 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t7 a_n7625_23622 Vss.t534 nfet_03v3
**devattr s=10400,304 d=17600,576
X431 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t9 Vin1.t3 a_n9429_n2007.t4 Vss.t162 nfet_03v3
**devattr s=15600,404 d=15600,404
X432 a_14313_33628.t3 a_14313_31423.t4 Vdd.t852 Vdd.t851 pfet_03v3
**devattr s=26000,604 d=44000,1176
X433 a_42809_29310 a_42729_29218.t4 Vss.t341 Vss.t340 nfet_03v3
**devattr s=17600,576 d=10400,304
X434 SARlogic_0.dffrs_8.Qb Reset.t39 Vdd.t854 Vdd.t853 pfet_03v3
**devattr s=26000,604 d=44000,1176
X435 SARlogic_0.dffrs_5.nand3_8.Z.t2 SARlogic_0.dffrs_4.Q.t5 a_12585_7428 Vss.t361 nfet_03v3
**devattr s=10400,304 d=17600,576
X436 SARlogic_0.dffrs_5.Qb.t2 Reset.t40 a_14071_9634 Vss.t604 nfet_03v3
**devattr s=10400,304 d=17600,576
X437 SARlogic_0.dffrs_2.Q.t2 SARlogic_0.dffrs_2.Qb.t4 Vdd.t812 Vdd.t811 pfet_03v3
**devattr s=26000,604 d=44000,1176
X438 SARlogic_0.dffrs_11.Qb Reset.t41 a_14071_19210 Vss.t605 nfet_03v3
**devattr s=10400,304 d=17600,576
X439 a_39915_29984 a_39055_28100 a_39727_29264.t1 Vdd.t260 pfet_03v3
**devattr s=52800,1376 d=31200,704
X440 a_n6323_11838 Vdd.t962 Vss.t429 Vss.t428 nfet_03v3
**devattr s=17600,576 d=10400,304
X441 SARlogic_0.dffrs_0.nand3_6.C.t2 Clk.t16 a_n7625_11838 Vss.t507 nfet_03v3
**devattr s=10400,304 d=17600,576
X442 a_29583_28100 a_28027_28820.t4 Vss.t186 Vss.t185 nfet_03v3
**devattr s=17600,576 d=17600,576
X443 Vdd.t325 SARlogic_0.dffrs_8.nand3_8.C.t6 SARlogic_0.dffrs_8.Qb Vdd.t324 pfet_03v3
**devattr s=26000,604 d=26000,604
X444 SARlogic_0.dffrs_2.nand3_8.C.t0 SARlogic_0.dffrs_2.nand3_6.C.t6 Vdd.t385 Vdd.t384 pfet_03v3
**devattr s=44000,1176 d=26000,604
X445 a_8359_17004 SARlogic_0.dffrs_10.nand3_8.C.t6 Vss.t602 Vss.t601 nfet_03v3
**devattr s=17600,576 d=10400,304
X446 Vdd.t27 adc_PISO_0.2inmux_2.Bit.t6 a_n389_31159.t0 Vdd.t26 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X447 Vdd.t387 SARlogic_0.dffrs_2.nand3_6.C.t7 SARlogic_0.dffrs_2.Q.t0 Vdd.t386 pfet_03v3
**devattr s=26000,604 d=26000,604
X448 a_14071_19210 SARlogic_0.dffrs_11.nand3_8.C.t5 a_13887_19210 Vss.t539 nfet_03v3
**devattr s=10400,304 d=10400,304
X449 a_23785_31423.t1 Clk_piso.t7 a_24049_33720 Vss.t354 nfet_03v3
**devattr s=10400,304 d=17600,576
X450 a_25351_33720 Vdd.t963 Vss.t427 Vss.t426 nfet_03v3
**devattr s=17600,576 d=10400,304
X451 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t13 Vdd.t716 Vdd.t715 pfet_03v3
**devattr s=10400,304 d=10400,304
X452 SARlogic_0.dffrs_7.nand3_6.C.t0 adc_PISO_0.B4.t8 Vdd.t85 Vdd.t84 pfet_03v3
**devattr s=26000,604 d=44000,1176
X453 Vdd.t856 Reset.t42 SARlogic_0.dffrs_3.nand3_8.Z.t2 Vdd.t855 pfet_03v3
**devattr s=26000,604 d=26000,604
X454 SARlogic_0.dffrs_2.nand3_6.C.t3 SARlogic_0.dffrs_2.nand3_1.C.t4 Vdd.t914 Vdd.t913 pfet_03v3
**devattr s=44000,1176 d=26000,604
X455 a_8359_19209 SARlogic_0.dffrs_10.nand3_6.C.t8 Vss.t180 Vss.t179 nfet_03v3
**devattr s=17600,576 d=10400,304
X456 a_35007_33720 a_33257_31423.t8 a_34823_33720 Vss.t212 nfet_03v3
**devattr s=10400,304 d=10400,304
X457 Vdd.t658 adc_PISO_0.dffrs_3.Q.t6 a_28027_31160.t0 Vdd.t657 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X458 a_n2097_9634 SARlogic_0.dffrs_1.nand3_8.C.t5 a_n2281_9634 Vss.t118 nfet_03v3
**devattr s=10400,304 d=10400,304
X459 Vdd.t163 SARlogic_0.dffrs_3.nand3_8.C.t7 SARlogic_0.dffrs_3.Qb.t1 Vdd.t162 pfet_03v3
**devattr s=26000,604 d=26000,604
X460 a_23785_33628.t1 a_23785_31423.t8 a_24049_35925 Vss.t169 nfet_03v3
**devattr s=10400,304 d=17600,576
X461 a_n9861_31159.t2 inv2_0.out.t18 a_n9673_30439 Vss.t103 nfet_03v3
**devattr s=10400,304 d=17600,576
X462 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t6 Vdd.t57 Vdd.t56 pfet_03v3
**devattr s=26000,604 d=44000,1176
X463 a_459_21414 Reset.t43 a_275_21414 Vss.t606 nfet_03v3
**devattr s=10400,304 d=10400,304
X464 a_n7809_19212 SARlogic_0.dffrs_14.nand3_6.C.t8 Vss.t536 Vss.t535 nfet_03v3
**devattr s=17600,576 d=10400,304
X465 Vss.t559 a_27321_29020 a_28215_28100 Vss.t558 nfet_03v3
**devattr s=10400,304 d=17600,576
X466 SARlogic_0.dffrs_2.nand3_8.Z.t2 SARlogic_0.dffrs_2.d.t5 a_459_7428 Vss.t376 nfet_03v3
**devattr s=10400,304 d=17600,576
X467 SARlogic_0.dffrs_4.nand3_1.C.t1 Vdd.t534 Vdd.t536 Vdd.t535 pfet_03v3
**devattr s=44000,1176 d=26000,604
X468 adc_PISO_0.dffrs_3.Qb Vdd.t531 Vdd.t533 Vdd.t532 pfet_03v3
**devattr s=26000,604 d=44000,1176
X469 Vdd.t848 SARlogic_0.dffrs_10.nand3_8.C.t7 SARlogic_0.dffrs_10.Qb Vdd.t847 pfet_03v3
**devattr s=26000,604 d=26000,604
X470 a_13887_11838 Vdd.t964 Vss.t425 Vss.t424 nfet_03v3
**devattr s=17600,576 d=10400,304
X471 a_28215_30440 inv2_0.out.t19 a_28027_31160.t1 Vss.t528 nfet_03v3
**devattr s=17600,576 d=10400,304
X472 Vdd.t618 SARlogic_0.dffrs_4.nand3_6.C.t6 SARlogic_0.dffrs_4.Q.t1 Vdd.t617 pfet_03v3
**devattr s=26000,604 d=26000,604
X473 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t5 a_459_17004 Vss.t315 nfet_03v3
**devattr s=10400,304 d=17600,576
X474 SARlogic_0.dffrs_4.nand3_8.Z.t1 SARlogic_0.dffrs_4.d.t6 Vdd.t876 Vdd.t875 pfet_03v3
**devattr s=26000,604 d=44000,1176
X475 a_459_23619 SARlogic_0.dffrs_8.nand3_8.Z a_275_23619 Vss.t2 nfet_03v3
**devattr s=10400,304 d=10400,304
X476 Vdd.t530 Vdd.t528 a_23785_31423.t2 Vdd.t529 pfet_03v3
**devattr s=26000,604 d=26000,604
X477 a_17929_21414 SARlogic_0.dffrs_5.Qb.t7 Vss.t28 Vss.t27 nfet_03v3
**devattr s=17600,576 d=10400,304
X478 adc_PISO_0.2inmux_1.OUT.t0 a_39727_29264.t4 Vss.t672 Vss.t671 nfet_03v3
**devattr s=17600,576 d=17600,576
X479 SARlogic_0.dffrs_8.nand3_8.C.t0 SARlogic_0.dffrs_8.nand3_8.Z a_459_19209 Vss.t1 nfet_03v3
**devattr s=10400,304 d=17600,576
X480 SARlogic_0.dffrs_1.nand3_8.Z.t2 SARlogic_0.dffrs_0.Q.t5 a_n3583_7428 Vss.t342 nfet_03v3
**devattr s=10400,304 d=17600,576
X481 a_25351_31516 adc_PISO_0.dffrs_3.Q.t7 Vss.t488 Vss.t487 nfet_03v3
**devattr s=17600,576 d=10400,304
X482 SARlogic_0.dffrs_0.Q.t1 SARlogic_0.dffrs_0.Qb.t8 a_n6139_11838 Vss.t239 nfet_03v3
**devattr s=10400,304 d=17600,576
X483 a_n4631_29217.t0 a_n4631_31422.t5 Vdd.t329 Vdd.t328 pfet_03v3
**devattr s=44000,1176 d=26000,604
X484 a_n6323_9634 SARlogic_0.dffrs_0.Q.t6 Vss.t344 Vss.t343 nfet_03v3
**devattr s=17600,576 d=10400,304
X485 Vdd.t934 a_23865_30170.t5 a_23785_33628.t0 Vdd.t933 pfet_03v3
**devattr s=26000,604 d=26000,604
X486 a_8543_11838 Reset.t44 a_8359_11838 Vss.t607 nfet_03v3
**devattr s=10400,304 d=10400,304
X487 SARlogic_0.dffrs_5.nand3_1.C.t1 SARlogic_0.dffrs_5.nand3_6.C.t6 a_12585_14043 Vss.t224 nfet_03v3
**devattr s=10400,304 d=17600,576
X488 SARlogic_0.dffrs_2.nand3_1.C.t1 SARlogic_0.dffrs_2.nand3_6.C.t8 Vdd.t389 Vdd.t388 pfet_03v3
**devattr s=26000,604 d=44000,1176
X489 a_14393_30170.t3 a_14313_29218.t5 Vdd.t814 Vdd.t813 pfet_03v3
**devattr s=44000,1176 d=26000,604
X490 Vdd.t790 SARlogic_0.dffrs_12.Q.t6 SARlogic_0.dffrs_11.nand3_8.C.t3 Vdd.t789 pfet_03v3
**devattr s=26000,604 d=26000,604
X491 a_35007_31516 a_33257_29218.t5 a_34823_31516 Vss.t234 nfet_03v3
**devattr s=10400,304 d=10400,304
X492 a_n4631_31422.t1 a_n4631_33627.t4 Vdd.t415 Vdd.t414 pfet_03v3
**devattr s=44000,1176 d=26000,604
X493 a_42729_29218.t1 a_42809_30170.t6 a_42993_31515 Vss.t586 nfet_03v3
**devattr s=10400,304 d=17600,576
X494 a_14313_29218.t3 a_14313_31423.t5 Vdd.t880 Vdd.t879 pfet_03v3
**devattr s=44000,1176 d=26000,604
X495 a_14577_31515 Clk_piso.t8 a_14393_31515 Vss.t355 nfet_03v3
**devattr s=10400,304 d=10400,304
X496 a_n10567_29019 inv2_0.out.t20 Vdd.t752 Vdd.t751 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X497 a_33337_30170.t3 adc_PISO_0.2inmux_5.OUT.t2 a_33521_29310 Vss.t489 nfet_03v3
**devattr s=10400,304 d=17600,576
X498 a_4501_14043 SARlogic_0.dffrs_3.nand3_8.Z.t6 a_4317_14043 Vss.t49 nfet_03v3
**devattr s=10400,304 d=10400,304
X499 a_275_17004 SARlogic_0.dffrs_8.nand3_8.C.t7 Vss.t666 Vss.t665 nfet_03v3
**devattr s=17600,576 d=10400,304
X500 a_n7625_7428 Reset.t45 a_n7809_7428 Vss.t608 nfet_03v3
**devattr s=10400,304 d=10400,304
X501 a_275_19209 SARlogic_0.dffrs_8.nand3_6.C.t8 Vss.t214 Vss.t213 nfet_03v3
**devattr s=17600,576 d=10400,304
X502 Vdd.t231 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t2 Vdd.t230 pfet_03v3
**devattr s=10400,304 d=10400,304
X503 SARlogic_0.dffrs_4.Qb.t3 Reset.t46 a_10029_9634 Vss.t290 nfet_03v3
**devattr s=10400,304 d=17600,576
X504 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_8.C.t5 Vdd.t908 Vdd.t907 pfet_03v3
**devattr s=44000,1176 d=26000,604
X505 a_16627_17004 Reset.t47 a_16443_17004 Vss.t291 nfet_03v3
**devattr s=10400,304 d=10400,304
X506 a_n4631_29217.t2 a_n4551_30169.t5 Vdd.t624 Vdd.t623 pfet_03v3
**devattr s=26000,604 d=44000,1176
X507 Vdd.t53 a_n8305_30439 a_n7445_29983 Vdd.t52 pfet_03v3
**devattr s=31200,704 d=52800,1376
X508 SARlogic_0.dffrs_2.nand3_1.C.t2 Vdd.t525 Vdd.t527 Vdd.t526 pfet_03v3
**devattr s=44000,1176 d=26000,604
X509 SARlogic_0.dffrs_13.nand3_8.C.t0 SARlogic_0.dffrs_13.nand3_8.Z.t5 a_n11637_9633 Vss.t115 nfet_03v3
**devattr s=10400,304 d=17600,576
X510 a_16627_19209 Vss.t124 a_16443_19209 Vss.t125 nfet_03v3
**devattr s=10400,304 d=10400,304
X511 a_n4631_31422.t3 Clk_piso.t9 Vdd.t610 Vdd.t609 pfet_03v3
**devattr s=26000,604 d=44000,1176
X512 adc_PISO_0.2inmux_2.Bit.t3 Vdd.t522 Vdd.t524 Vdd.t523 pfet_03v3
**devattr s=44000,1176 d=26000,604
X513 adc_PISO_0.dffrs_2.Q.t0 adc_PISO_0.dffrs_2.Qb Vdd.t461 Vdd.t460 pfet_03v3
**devattr s=26000,604 d=44000,1176
X514 SARlogic_0.dffrs_9.Qb Reset.t48 Vdd.t359 Vdd.t358 pfet_03v3
**devattr s=26000,604 d=44000,1176
X515 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t482 nfet_03v3
**devattr s=20800,504 d=20800,504
X516 SARlogic_0.dffrs_7.Qb adc_PISO_0.B5.t7 Vdd.t175 Vdd.t174 pfet_03v3
**devattr s=44000,1176 d=26000,604
X517 SARlogic_0.dffrs_4.d.t1 SARlogic_0.dffrs_3.Qb.t8 Vdd.t215 Vdd.t214 pfet_03v3
**devattr s=26000,604 d=44000,1176
X518 Piso_out.t0 adc_PISO_0.dffrs_5.Qb Vdd.t321 Vdd.t320 pfet_03v3
**devattr s=26000,604 d=44000,1176
X519 SARlogic_0.dffrs_2.d.t3 Vdd.t519 Vdd.t521 Vdd.t520 pfet_03v3
**devattr s=44000,1176 d=26000,604
X520 Vdd.t331 a_n4631_31422.t6 adc_PISO_0.2inmux_2.Bit.t0 Vdd.t330 pfet_03v3
**devattr s=26000,604 d=26000,604
X521 Vdd.t882 a_14313_31423.t6 adc_PISO_0.dffrs_2.Q.t3 Vdd.t881 pfet_03v3
**devattr s=26000,604 d=26000,604
X522 a_33337_29310 a_33257_29218.t6 Vss.t236 Vss.t235 nfet_03v3
**devattr s=17600,576 d=10400,304
X523 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vdd.t115 Vdd.t114 pfet_03v3
**devattr s=18700,450 d=34000,880
X524 a_n3583_21414 Reset.t49 a_n3767_21414 Vss.t292 nfet_03v3
**devattr s=10400,304 d=10400,304
X525 SARlogic_0.dffrs_3.nand3_8.Z.t1 SARlogic_0.dffrs_2.Q.t5 Vdd.t399 Vdd.t398 pfet_03v3
**devattr s=26000,604 d=44000,1176
X526 SARlogic_0.dffrs_0.Qb.t1 SARlogic_0.dffrs_0.Q.t7 Vdd.t413 Vdd.t412 pfet_03v3
**devattr s=44000,1176 d=26000,604
X527 a_n7625_23622 SARlogic_0.dffrs_14.nand3_8.Z a_n7809_23622 Vss.t541 nfet_03v3
**devattr s=10400,304 d=10400,304
X528 a_n3583_23619 SARlogic_0.dffrs_7.nand3_8.Z a_n3767_23619 Vss.t62 nfet_03v3
**devattr s=10400,304 d=10400,304
X529 a_20971_29984 a_20111_30440 Vdd.t155 Vdd.t154 pfet_03v3
**devattr s=52800,1376 d=31200,704
X530 Vdd.t700 Clk.t17 SARlogic_0.dffrs_2.nand3_8.C.t3 Vdd.t699 pfet_03v3
**devattr s=26000,604 d=26000,604
X531 a_n7625_11838 Reset.t50 a_n7809_11838 Vss.t293 nfet_03v3
**devattr s=10400,304 d=10400,304
X532 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t6 Vdd.t383 Vdd.t382 pfet_03v3
**devattr s=26000,604 d=44000,1176
X533 a_25535_33720 a_23785_31423.t9 a_25351_33720 Vss.t366 nfet_03v3
**devattr s=10400,304 d=10400,304
X534 Vss.t513 a_39055_30440 a_39727_29264.t3 Vss.t512 nfet_03v3
**devattr s=17600,576 d=17600,576
X535 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t15 a_n9767_249 a_n9855_341 Vss.t545 nfet_03v3
**devattr s=35200,976 d=20800,504
X536 Vdd.t361 Reset.t51 SARlogic_0.dffrs_2.nand3_6.C.t2 Vdd.t360 pfet_03v3
**devattr s=26000,604 d=26000,604
X537 adc_PISO_0.dffrs_2.Qb Vdd.t516 Vdd.t518 Vdd.t517 pfet_03v3
**devattr s=26000,604 d=44000,1176
X538 adc_PISO_0.dffrs_5.Qb Vdd.t513 Vdd.t515 Vdd.t514 pfet_03v3
**devattr s=26000,604 d=44000,1176
X539 a_20111_28100 a_18555_28820.t5 Vdd.t437 Vdd.t436 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X540 SARlogic_0.dffrs_11.nand3_6.C.t3 SARlogic_0.dffrs_12.Q.t7 Vdd.t792 Vdd.t791 pfet_03v3
**devattr s=26000,604 d=44000,1176
X541 SARlogic_0.dffrs_5.Qb.t0 SARlogic_0.dffrs_5.Q.t5 Vdd.t19 Vdd.t18 pfet_03v3
**devattr s=44000,1176 d=26000,604
X542 Vdd.t309 a_4841_31422.t6 adc_PISO_0.dffrs_1.Q.t2 Vdd.t308 pfet_03v3
**devattr s=26000,604 d=26000,604
X543 adc_PISO_0.dffrs_1.Q.t1 adc_PISO_0.dffrs_1.Qb a_6591_33719 Vss.t5 nfet_03v3
**devattr s=10400,304 d=17600,576
X544 Vdd.t816 a_14313_29218.t6 adc_PISO_0.dffrs_2.Qb Vdd.t815 pfet_03v3
**devattr s=26000,604 d=26000,604
X545 a_37499_28820.t3 adc_PISO_0.B1.t9 Vdd.t800 Vdd.t799 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X546 a_42729_31423.t3 Clk_piso.t10 Vdd.t612 Vdd.t611 pfet_03v3
**devattr s=26000,604 d=44000,1176
X547 a_8359_9633 SARlogic_0.dffrs_4.nand3_6.C.t7 Vss.t467 Vss.t466 nfet_03v3
**devattr s=17600,576 d=10400,304
X548 Vdd.t512 Vdd.t510 a_14313_31423.t3 Vdd.t511 pfet_03v3
**devattr s=26000,604 d=26000,604
X549 SARlogic_0.dffrs_12.Qb SARlogic_0.dffrs_12.Q.t8 Vdd.t794 Vdd.t793 pfet_03v3
**devattr s=44000,1176 d=26000,604
X550 a_1761_11838 Vdd.t965 Vss.t423 Vss.t422 nfet_03v3
**devattr s=17600,576 d=10400,304
X551 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t7 Vdd.t203 Vdd.t202 pfet_03v3
**devattr s=26000,604 d=44000,1176
X552 a_n6389_n2007 a_n6589_n2099 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t13 Vss.t385 nfet_03v3
**devattr s=15600,404 d=26400,776
X553 a_18555_31160.t3 inv2_0.out.t21 Vdd.t754 Vdd.t753 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X554 adc_PISO_0.2inmux_2.OUT.t0 a_1839_29263.t4 Vss.t674 Vss.t673 nfet_03v3
**devattr s=17600,576 d=17600,576
X555 a_n2097_21414 SARlogic_0.dffrs_7.nand3_6.C.t7 a_n2281_21414 Vss.t43 nfet_03v3
**devattr s=10400,304 d=10400,304
X556 SARlogic_0.dffrs_0.Qb.t2 Reset.t52 Vdd.t363 Vdd.t362 pfet_03v3
**devattr s=26000,604 d=44000,1176
X557 a_42729_33628.t0 a_42729_31423.t4 Vdd.t281 Vdd.t280 pfet_03v3
**devattr s=26000,604 d=44000,1176
X558 Vdd.t349 Reset.t53 SARlogic_0.dffrs_9.nand3_6.C.t3 Vdd.t348 pfet_03v3
**devattr s=26000,604 d=26000,604
X559 Vdd.t105 a_14393_30170.t6 a_14313_33628.t0 Vdd.t104 pfet_03v3
**devattr s=26000,604 d=26000,604
X560 adc_PISO_0.B5.t3 SARlogic_0.dffrs_7.Qb a_n2097_21414 Vss.t625 nfet_03v3
**devattr s=10400,304 d=17600,576
X561 Vdd.t622 SARlogic_0.dffrs_13.nand3_6.C.t5 SARlogic_0.dffrs_0.d.t2 Vdd.t621 pfet_03v3
**devattr s=26000,604 d=26000,604
X562 SARlogic_0.dffrs_14.nand3_8.C.t3 SARlogic_0.dffrs_14.nand3_8.Z a_n7625_19212 Vss.t540 nfet_03v3
**devattr s=10400,304 d=17600,576
X563 a_n6139_11838 SARlogic_0.dffrs_0.nand3_6.C.t8 a_n6323_11838 Vss.t187 nfet_03v3
**devattr s=10400,304 d=10400,304
X564 a_n8351_341 a_n8551_249 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t7 Vss.t367 nfet_03v3
**devattr s=20800,504 d=35200,976
X565 adc_PISO_0.2inmux_3.OUT.t0 a_11311_29264.t4 Vss.t326 Vss.t325 nfet_03v3
**devattr s=17600,576 d=17600,576
X566 a_25535_31516 a_23785_29218.t6 a_25351_31516 Vss.t85 nfet_03v3
**devattr s=10400,304 d=10400,304
X567 Vdd.t606 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_1.C Vdd.t605 pfet_03v3
**devattr s=26000,604 d=26000,604
X568 SARlogic_0.dffrs_4.nand3_6.C.t0 Clk.t18 a_8543_11838 Vss.t508 nfet_03v3
**devattr s=10400,304 d=17600,576
X569 a_9845_11838 Vdd.t966 Vss.t421 Vss.t420 nfet_03v3
**devattr s=17600,576 d=10400,304
X570 a_18743_28100 adc_PISO_0.B3.t8 a_18555_28820.t2 Vss.t663 nfet_03v3
**devattr s=17600,576 d=10400,304
X571 Vdd.t351 Reset.t54 SARlogic_0.dffrs_1.nand3_8.Z.t3 Vdd.t350 pfet_03v3
**devattr s=26000,604 d=26000,604
X572 Vdd.t646 Clk_piso.t11 a_4841_29217.t0 Vdd.t645 pfet_03v3
**devattr s=26000,604 d=26000,604
X573 Vdd.t509 Vdd.t507 a_42809_30170.t3 Vdd.t508 pfet_03v3
**devattr s=26000,604 d=26000,604
X574 a_39055_28100 a_37499_28820.t5 Vdd.t604 Vdd.t603 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X575 a_23865_30170.t1 adc_PISO_0.2inmux_4.OUT.t2 a_24049_29310 Vss.t83 nfet_03v3
**devattr s=10400,304 d=17600,576
X576 Vdd.t303 a_1167_30439 a_2027_29983 Vdd.t302 pfet_03v3
**devattr s=31200,704 d=52800,1376
X577 a_23865_33720 a_23785_33628.t5 Vss.t485 Vss.t484 nfet_03v3
**devattr s=17600,576 d=10400,304
X578 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t15 Vdd.t650 Vdd.t649 pfet_03v3
**devattr s=10400,304 d=10400,304
X579 a_n7445_29983 a_n8305_28099 a_n7633_29263.t1 Vdd.t122 pfet_03v3
**devattr s=52800,1376 d=31200,704
X580 a_4841_29217.t1 a_4841_31422.t7 Vdd.t311 Vdd.t310 pfet_03v3
**devattr s=44000,1176 d=26000,604
X581 a_n9429_n2007.t14 Vin2.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t372 nfet_03v3
**devattr s=15600,404 d=15600,404
X582 Vdd.t506 Vdd.t504 a_4841_31422.t1 Vdd.t505 pfet_03v3
**devattr s=26000,604 d=26000,604
X583 Vdd.t648 Clk_piso.t12 a_42729_29218.t0 Vdd.t647 pfet_03v3
**devattr s=26000,604 d=26000,604
X584 a_459_17004 Reset.t55 a_275_17004 Vss.t288 nfet_03v3
**devattr s=10400,304 d=10400,304
X585 SARlogic_0.dffrs_3.nand3_1.C.t1 SARlogic_0.dffrs_3.nand3_6.C.t8 a_4501_14043 Vss.t580 nfet_03v3
**devattr s=10400,304 d=17600,576
X586 a_12401_14043 Vdd.t968 Vss.t417 Vss.t416 nfet_03v3
**devattr s=17600,576 d=10400,304
X587 Vdd.t820 a_10639_30440 a_11499_29984 Vdd.t819 pfet_03v3
**devattr s=31200,704 d=52800,1376
X588 a_23865_35925 Vdd.t967 Vss.t419 Vss.t418 nfet_03v3
**devattr s=17600,576 d=10400,304
X589 Comp_out.t5 a_n10831_4320 Vdd.t297 Vdd.t296 pfet_03v3
**devattr s=18700,450 d=18700,450
X590 a_8543_7428 Reset.t56 a_8359_7428 Vss.t289 nfet_03v3
**devattr s=10400,304 d=10400,304
X591 a_4841_31422.t3 a_4841_33627.t4 Vdd.t916 Vdd.t915 pfet_03v3
**devattr s=44000,1176 d=26000,604
X592 SARlogic_0.dffrs_0.nand3_8.Z.t2 SARlogic_0.dffrs_0.nand3_8.C.t5 Vdd.t247 Vdd.t246 pfet_03v3
**devattr s=44000,1176 d=26000,604
X593 Vdd.t391 adc_PISO_0.B1.t10 SARlogic_0.dffrs_10.nand3_8.C.t3 Vdd.t390 pfet_03v3
**devattr s=26000,604 d=26000,604
X594 a_n1095_29019 inv2_0.out.t22 Vdd.t756 Vdd.t755 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X595 a_n11637_9633 Clk.t19 a_n11821_9633 Vss.t520 nfet_03v3
**devattr s=10400,304 d=10400,304
X596 a_459_19209 adc_PISO_0.B3.t9 a_275_19209 Vss.t664 nfet_03v3
**devattr s=10400,304 d=10400,304
X597 a_20111_30440 a_18555_31160.t4 Vss.t389 Vss.t388 nfet_03v3
**devattr s=17600,576 d=17600,576
X598 a_37499_31160.t0 inv2_0.out.t23 a_37687_30440 Vss.t529 nfet_03v3
**devattr s=10400,304 d=17600,576
X599 a_30255_29264.t2 a_29583_28100 Vss.t4 Vss.t3 nfet_03v3
**devattr s=17600,576 d=17600,576
X600 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t5 a_n9429_n2007.t15 Vss.t373 nfet_03v3
**devattr s=15600,404 d=15600,404
X601 Vdd.t417 Clk_piso.t13 a_n4631_29217.t1 Vdd.t416 pfet_03v3
**devattr s=26000,604 d=26000,604
X602 Vdd.t634 SARlogic_0.dffrs_2.nand3_8.Z.t6 SARlogic_0.dffrs_2.nand3_1.C.t3 Vdd.t633 pfet_03v3
**devattr s=26000,604 d=26000,604
X603 a_8359_11838 SARlogic_0.dffrs_4.nand3_1.C.t5 Vss.t622 Vss.t621 nfet_03v3
**devattr s=17600,576 d=10400,304
X604 Vss.t584 a_n8385_n2885 a_n8473_n2793 Vss.t583 nfet_03v3
**devattr s=14080,496 d=8320,264
X605 Vdd.t718 Clk.t20 SARlogic_0.dffrs_1.nand3_8.C.t2 Vdd.t717 pfet_03v3
**devattr s=26000,604 d=26000,604
X606 adc_PISO_0.2inmux_4.OUT.t1 a_20783_29264.t5 Vdd.t245 Vdd.t244 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X607 a_2027_29983 a_1167_28099 a_1839_29263.t0 Vdd.t108 pfet_03v3
**devattr s=52800,1376 d=31200,704
X608 SARlogic_0.dffrs_4.Q.t2 SARlogic_0.dffrs_4.Qb.t6 a_10029_11838 Vss.t648 nfet_03v3
**devattr s=10400,304 d=17600,576
X609 Vdd.t503 Vdd.t501 a_n4631_31422.t2 Vdd.t502 pfet_03v3
**devattr s=26000,604 d=26000,604
X610 Vdd.t195 a_8377_29020 a_9083_28820.t3 Vdd.t194 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X611 Vdd.t353 Reset.t57 SARlogic_0.dffrs_1.nand3_6.C.t3 Vdd.t352 pfet_03v3
**devattr s=26000,604 d=26000,604
X612 a_27321_29020 inv2_0.out.t24 Vdd.t758 Vdd.t757 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X613 a_4317_9633 SARlogic_0.dffrs_3.nand3_6.C.t9 Vss.t582 Vss.t581 nfet_03v3
**devattr s=17600,576 d=10400,304
X614 a_4317_14043 Vdd.t969 Vss.t415 Vss.t414 nfet_03v3
**devattr s=17600,576 d=10400,304
X615 SARlogic_0.dffrs_13.nand3_8.C.t2 SARlogic_0.dffrs_13.nand3_6.C.t6 Vdd.t628 Vdd.t627 pfet_03v3
**devattr s=44000,1176 d=26000,604
X616 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t6 a_n9429_n2007.t16 Vss.t166 nfet_03v3
**devattr s=15600,404 d=15600,404
X617 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t7 a_n9429_n2007.t11 Vss.t162 nfet_03v3
**devattr s=15600,404 d=15600,404
X618 adc_PISO_0.B1.t0 SARlogic_0.dffrs_11.Qb a_14071_21414 Vss.t150 nfet_03v3
**devattr s=10400,304 d=17600,576
X619 a_n3767_21414 SARlogic_0.dffrs_7.nand3_1.C Vss.t107 Vss.t106 nfet_03v3
**devattr s=17600,576 d=10400,304
X620 Vss.t7 a_n1095_29019 a_n201_28099 Vss.t6 nfet_03v3
**devattr s=10400,304 d=17600,576
X621 Vss.t570 a_10639_30440 a_11311_29264.t3 Vss.t569 nfet_03v3
**devattr s=17600,576 d=17600,576
X622 SARlogic_0.dffrs_2.nand3_6.C.t1 Clk.t21 a_459_11838 Vss.t521 nfet_03v3
**devattr s=10400,304 d=17600,576
X623 a_14071_21414 SARlogic_0.dffrs_11.nand3_6.C.t8 a_13887_21414 Vss.t181 nfet_03v3
**devattr s=10400,304 d=10400,304
X624 SARlogic_0.dffrs_13.nand3_6.C.t1 SARlogic_0.dffrs_13.nand3_1.C.t4 Vdd.t616 Vdd.t615 pfet_03v3
**devattr s=44000,1176 d=26000,604
X625 a_n11821_7428 SARlogic_0.dffrs_13.nand3_8.C.t6 Vss.t297 Vss.t296 nfet_03v3
**devattr s=17600,576 d=10400,304
X626 a_n3767_23619 SARlogic_0.dffrs_0.Qb.t9 Vss.t241 Vss.t240 nfet_03v3
**devattr s=17600,576 d=10400,304
X627 a_39055_30440 a_37499_31160.t4 Vss.t650 Vss.t649 nfet_03v3
**devattr s=17600,576 d=17600,576
X628 Vdd.t69 a_36793_29020 a_37499_28820.t0 Vdd.t68 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X629 a_14313_31423.t0 Clk_piso.t14 a_14577_33720 Vss.t347 nfet_03v3
**devattr s=10400,304 d=17600,576
X630 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t7 Vdd.t377 Vdd.t376 pfet_03v3
**devattr s=26000,604 d=44000,1176
X631 a_n9429_n2007.t17 Vin1.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t8 Vss.t362 nfet_03v3
**devattr s=15600,404 d=15600,404
X632 adc_PISO_0.dffrs_3.Q.t1 adc_PISO_0.dffrs_3.Qb a_25535_33720 Vss.t244 nfet_03v3
**devattr s=10400,304 d=17600,576
X633 adc_PISO_0.dffrs_1.Qb Vdd.t498 Vdd.t500 Vdd.t499 pfet_03v3
**devattr s=26000,604 d=44000,1176
X634 Vdd.t31 adc_PISO_0.dffrs_2.Q.t5 a_18555_31160.t0 Vdd.t30 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X635 SARlogic_0.dffrs_2.Qb.t1 SARlogic_0.dffrs_2.Q.t6 Vdd.t822 Vdd.t821 pfet_03v3
**devattr s=44000,1176 d=26000,604
X636 a_14313_33628.t2 a_14313_31423.t7 a_14577_35925 Vss.t550 nfet_03v3
**devattr s=10400,304 d=17600,576
X637 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t16 Vdd.t652 Vdd.t651 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X638 SARlogic_0.dffrs_2.Q.t3 SARlogic_0.dffrs_2.Qb.t5 a_1945_11838 Vss.t565 nfet_03v3
**devattr s=10400,304 d=17600,576
X639 Vdd.t764 Vss.t678 a_n9861_31159.t0 Vdd.t763 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X640 a_n7809_14043 Vdd.t970 Vss.t413 Vss.t412 nfet_03v3
**devattr s=17600,576 d=10400,304
X641 Vdd.t906 SARlogic_0.dffrs_7.nand3_8.C.t6 SARlogic_0.dffrs_7.Qb Vdd.t905 pfet_03v3
**devattr s=26000,604 d=26000,604
X642 Vss.t65 a_17849_29020 a_18743_28100 Vss.t64 nfet_03v3
**devattr s=10400,304 d=17600,576
X643 Vdd.t283 a_42729_31423.t5 Piso_out.t3 Vdd.t282 pfet_03v3
**devattr s=26000,604 d=26000,604
X644 Vdd.t840 SARlogic_0.dffrs_1.nand3_6.C.t6 SARlogic_0.dffrs_2.d.t0 Vdd.t839 pfet_03v3
**devattr s=26000,604 d=26000,604
X645 Vdd.t355 Reset.t58 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t354 pfet_03v3
**devattr s=26000,604 d=26000,604
X646 a_1945_11838 SARlogic_0.dffrs_2.nand3_6.C.t9 a_1761_11838 Vss.t319 nfet_03v3
**devattr s=10400,304 d=10400,304
X647 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t7 Vin1.t5 a_n9429_n2007.t18 Vss.t363 nfet_03v3
**devattr s=15600,404 d=15600,404
X648 Vdd.t720 Clk.t22 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t8 Vdd.t719 pfet_03v3
**devattr s=14080,496 d=14080,496
X649 adc_PISO_0.dffrs_2.Q.t2 Vdd.t495 Vdd.t497 Vdd.t496 pfet_03v3
**devattr s=44000,1176 d=26000,604
X650 adc_PISO_0.2inmux_2.Bit.t2 adc_PISO_0.dffrs_0.Qb Vdd.t81 Vdd.t80 pfet_03v3
**devattr s=26000,604 d=44000,1176
X651 SARlogic_0.dffrs_13.nand3_8.C.t1 SARlogic_0.dffrs_13.nand3_8.Z.t6 Vdd.t137 Vdd.t136 pfet_03v3
**devattr s=26000,604 d=44000,1176
X652 SARlogic_0.dffrs_7.Qb Reset.t59 Vdd.t357 Vdd.t356 pfet_03v3
**devattr s=26000,604 d=44000,1176
X653 SARlogic_0.dffrs_2.d.t1 SARlogic_0.dffrs_1.Qb.t8 Vdd.t49 Vdd.t48 pfet_03v3
**devattr s=26000,604 d=44000,1176
X654 a_4501_7428 Reset.t60 a_4317_7428 Vss.t286 nfet_03v3
**devattr s=10400,304 d=10400,304
X655 SARlogic_0.dffrs_7.nand3_6.C.t1 adc_PISO_0.B4.t9 a_n3583_21414 Vss.t71 nfet_03v3
**devattr s=10400,304 d=17600,576
X656 a_275_11838 SARlogic_0.dffrs_2.nand3_1.C.t5 Vss.t120 Vss.t119 nfet_03v3
**devattr s=17600,576 d=10400,304
X657 Vdd.t249 SARlogic_0.dffrs_0.nand3_8.C.t6 SARlogic_0.dffrs_0.Qb.t0 Vdd.t248 pfet_03v3
**devattr s=26000,604 d=26000,604
X658 SARlogic_0.dffrs_1.nand3_8.Z.t0 SARlogic_0.dffrs_1.nand3_8.C.t6 Vdd.t147 Vdd.t146 pfet_03v3
**devattr s=44000,1176 d=26000,604
X659 SARlogic_0.dffrs_12.nand3_8.C.t1 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t21 Vdd.t20 pfet_03v3
**devattr s=26000,604 d=44000,1176
X660 SARlogic_0.dffrs_11.nand3_6.C.t0 SARlogic_0.dffrs_11.nand3_1.C Vdd.t313 Vdd.t312 pfet_03v3
**devattr s=44000,1176 d=26000,604
X661 adc_PISO_0.B3.t2 SARlogic_0.dffrs_2.Qb.t6 Vdd.t746 Vdd.t745 pfet_03v3
**devattr s=44000,1176 d=26000,604
X662 SARlogic_0.dffrs_9.nand3_6.C.t2 adc_PISO_0.B2.t9 Vdd.t684 Vdd.t683 pfet_03v3
**devattr s=26000,604 d=44000,1176
X663 a_n3583_17004 Reset.t61 a_n3767_17004 Vss.t287 nfet_03v3
**devattr s=10400,304 d=10400,304
X664 SARlogic_0.dffrs_13.nand3_6.C.t3 Clk.t23 Vdd.t722 Vdd.t721 pfet_03v3
**devattr s=26000,604 d=44000,1176
X665 SARlogic_0.dffrs_4.Qb.t1 SARlogic_0.dffrs_4.Q.t6 Vdd.t433 Vdd.t432 pfet_03v3
**devattr s=44000,1176 d=26000,604
X666 SARlogic_0.dffrs_0.d.t3 Reset.t62 Vdd.t339 Vdd.t338 pfet_03v3
**devattr s=44000,1176 d=26000,604
X667 a_n7625_19212 adc_PISO_0.B5.t8 a_n7809_19212 Vss.t155 nfet_03v3
**devattr s=10400,304 d=10400,304
X668 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t8 a_n3583_23619 Vss.t44 nfet_03v3
**devattr s=10400,304 d=17600,576
X669 a_37687_28100 adc_PISO_0.B1.t11 a_37499_28820.t1 Vss.t320 nfet_03v3
**devattr s=17600,576 d=10400,304
X670 a_9271_30440 adc_PISO_0.dffrs_1.Q.t7 Vss.t632 Vss.t631 nfet_03v3
**devattr s=17600,576 d=10400,304
X671 Vdd.t494 Vdd.t492 a_33337_30170.t2 Vdd.t493 pfet_03v3
**devattr s=26000,604 d=26000,604
X672 adc_PISO_0.dffrs_3.Qb Vdd.t971 a_25535_31516 Vss.t411 nfet_03v3
**devattr s=10400,304 d=17600,576
X673 a_10029_11838 SARlogic_0.dffrs_4.nand3_6.C.t8 a_9845_11838 Vss.t370 nfet_03v3
**devattr s=10400,304 d=10400,304
X674 Vdd.t25 a_n9629_1405 a_n9717_1497 Vdd.t24 pfet_03v3
**devattr s=17600,576 d=10400,304
X675 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_4.Qb.t7 Vdd.t912 Vdd.t911 pfet_03v3
**devattr s=44000,1176 d=26000,604
X676 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t7 Vdd.t902 Vdd.t901 pfet_03v3
**devattr s=26000,604 d=44000,1176
X677 a_n8305_28099 a_n9861_28819.t4 Vss.t328 Vss.t327 nfet_03v3
**devattr s=17600,576 d=17600,576
X678 a_n3583_19209 adc_PISO_0.B4.t10 a_n3767_19209 Vss.t70 nfet_03v3
**devattr s=10400,304 d=10400,304
X679 a_29583_28100 a_28027_28820.t5 Vdd.t750 Vdd.t749 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X680 SARlogic_0.dffrs_4.nand3_8.Z.t0 SARlogic_0.dffrs_4.d.t7 a_8543_7428 Vss.t14 nfet_03v3
**devattr s=10400,304 d=17600,576
X681 a_4841_29217.t2 a_4921_30169.t5 Vdd.t824 Vdd.t823 pfet_03v3
**devattr s=26000,604 d=44000,1176
X682 a_1167_28099 a_n389_28819.t4 Vss.t271 Vss.t270 nfet_03v3
**devattr s=17600,576 d=17600,576
X683 Vdd.t445 Clk_piso.t15 a_33257_29218.t3 Vdd.t444 pfet_03v3
**devattr s=26000,604 d=26000,604
X684 Vdd.t397 SARlogic_0.dffrs_1.nand3_8.Z.t5 SARlogic_0.dffrs_1.nand3_1.C.t0 Vdd.t396 pfet_03v3
**devattr s=26000,604 d=26000,604
X685 a_24049_33720 Vdd.t972 a_23865_33720 Vss.t410 nfet_03v3
**devattr s=10400,304 d=10400,304
X686 Vdd.t409 a_42729_29218.t5 adc_PISO_0.dffrs_5.Qb Vdd.t408 pfet_03v3
**devattr s=26000,604 d=26000,604
X687 a_n8305_28099 a_n9861_28819.t5 Vdd.t75 Vdd.t74 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X688 adc_PISO_0.dffrs_2.Qb adc_PISO_0.dffrs_2.Q.t6 Vdd.t33 Vdd.t32 pfet_03v3
**devattr s=44000,1176 d=26000,604
X689 adc_PISO_0.dffrs_1.Q.t3 Vdd.t489 Vdd.t491 Vdd.t490 pfet_03v3
**devattr s=44000,1176 d=26000,604
X690 a_20783_29264.t1 a_20111_28100 a_20971_29984 Vdd.t288 pfet_03v3
**devattr s=31200,704 d=52800,1376
X691 a_4841_31422.t0 Clk_piso.t16 Vdd.t447 Vdd.t446 pfet_03v3
**devattr s=26000,604 d=44000,1176
X692 a_5803_19210 adc_PISO_0.B3.t10 Vss.t660 Vss.t659 nfet_03v3
**devattr s=17600,576 d=10400,304
X693 a_37687_30440 adc_PISO_0.2inmux_1.Bit.t8 Vss.t658 Vss.t657 nfet_03v3
**devattr s=17600,576 d=10400,304
X694 a_n4551_31514 a_n4631_31422.t7 Vss.t280 Vss.t279 nfet_03v3
**devattr s=17600,576 d=10400,304
X695 a_12585_14043 SARlogic_0.dffrs_5.nand3_8.Z.t5 a_12401_14043 Vss.t0 nfet_03v3
**devattr s=10400,304 d=10400,304
X696 Vss.t676 adc_PISO_0.2inmux_2.Bit.t7 a_n201_30439 Vss.t675 nfet_03v3
**devattr s=10400,304 d=17600,576
X697 a_24049_35925 a_23865_30170.t6 a_23865_35925 Vss.t250 nfet_03v3
**devattr s=10400,304 d=10400,304
X698 a_1167_28099 a_n389_28819.t5 Vdd.t317 Vdd.t316 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X699 SARlogic_0.dffrs_13.nand3_1.C.t3 Reset.t63 Vdd.t341 Vdd.t340 pfet_03v3
**devattr s=44000,1176 d=26000,604
X700 SARlogic_0.dffrs_12.nand3_8.C.t3 SARlogic_0.dffrs_12.nand3_6.C.t8 Vdd.t868 Vdd.t867 pfet_03v3
**devattr s=44000,1176 d=26000,604
X701 SARlogic_0.dffrs_10.nand3_8.C.t2 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t253 Vdd.t252 pfet_03v3
**devattr s=26000,604 d=44000,1176
X702 SARlogic_0.dffrs_0.nand3_8.C.t1 SARlogic_0.dffrs_0.nand3_8.Z.t6 a_n7625_9633 Vss.t477 nfet_03v3
**devattr s=10400,304 d=17600,576
X703 SARlogic_0.dffrs_9.nand3_6.C.t0 SARlogic_0.dffrs_9.nand3_1.C Vdd.t367 Vdd.t366 pfet_03v3
**devattr s=44000,1176 d=26000,604
X704 a_n4551_33719 a_n4631_33627.t5 Vss.t346 Vss.t345 nfet_03v3
**devattr s=17600,576 d=10400,304
X705 SARlogic_0.dffrs_0.d.t0 SARlogic_0.dffrs_13.Qb.t7 Vdd.t185 Vdd.t184 pfet_03v3
**devattr s=26000,604 d=44000,1176
X706 a_14393_31515 a_14313_31423.t8 Vss.t552 Vss.t551 nfet_03v3
**devattr s=17600,576 d=10400,304
X707 adc_PISO_0.2inmux_1.OUT.t1 a_39727_29264.t5 Vdd.t940 Vdd.t939 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X708 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_2.Qb.t7 Vdd.t748 Vdd.t747 pfet_03v3
**devattr s=44000,1176 d=26000,604
X709 SARlogic_0.dffrs_4.Qb.t2 Reset.t64 Vdd.t343 Vdd.t342 pfet_03v3
**devattr s=26000,604 d=44000,1176
X710 SARlogic_0.dffrs_1.nand3_8.C.t3 SARlogic_0.dffrs_1.nand3_6.C.t7 Vdd.t842 Vdd.t841 pfet_03v3
**devattr s=44000,1176 d=26000,604
X711 a_9083_28820.t0 adc_PISO_0.B4.t11 a_9271_28100 Vss.t69 nfet_03v3
**devattr s=10400,304 d=17600,576
X712 a_42809_30170.t0 a_42729_29218.t6 Vdd.t411 Vdd.t410 pfet_03v3
**devattr s=44000,1176 d=26000,604
X713 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t1 Vss.t209 nfet_03v3
**devattr s=20800,504 d=20800,504
X714 SARlogic_0.dffrs_11.Qb Reset.t65 Vdd.t345 Vdd.t344 pfet_03v3
**devattr s=26000,604 d=44000,1176
X715 SARlogic_0.dffrs_5.Q.t0 SARlogic_0.dffrs_5.Qb.t8 Vdd.t39 Vdd.t38 pfet_03v3
**devattr s=26000,604 d=44000,1176
X716 SARlogic_0.dffrs_5.nand3_8.C.t0 SARlogic_0.dffrs_5.nand3_8.Z.t6 a_12585_9633 Vss.t24 nfet_03v3
**devattr s=10400,304 d=17600,576
X717 SARlogic_0.dffrs_1.nand3_6.C.t0 SARlogic_0.dffrs_1.nand3_1.C.t4 Vdd.t1 Vdd.t0 pfet_03v3
**devattr s=44000,1176 d=26000,604
X718 a_23865_29310 a_23785_29218.t7 Vss.t87 Vss.t86 nfet_03v3
**devattr s=17600,576 d=10400,304
X719 Vdd.t780 SARlogic_0.dffrs_11.nand3_8.C.t6 SARlogic_0.dffrs_11.Qb Vdd.t779 pfet_03v3
**devattr s=26000,604 d=26000,604
X720 Vdd.t710 a_39055_30440 a_39915_29984 Vdd.t709 pfet_03v3
**devattr s=31200,704 d=52800,1376
X721 a_42729_29218.t3 a_42729_31423.t6 Vdd.t285 Vdd.t284 pfet_03v3
**devattr s=44000,1176 d=26000,604
X722 Vdd.t257 SARlogic_0.dffrs_5.nand3_6.C.t7 SARlogic_0.dffrs_5.Q.t2 Vdd.t256 pfet_03v3
**devattr s=26000,604 d=26000,604
X723 a_28027_28820.t0 adc_PISO_0.B2.t10 a_28215_28100 Vss.t498 nfet_03v3
**devattr s=10400,304 d=17600,576
X724 a_n4631_29217.t3 a_n4551_30169.t6 a_n4367_31514 Vss.t470 nfet_03v3
**devattr s=10400,304 d=17600,576
X725 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t17 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t1 Vss.t483 nfet_03v3
**devattr s=20800,504 d=20800,504
X726 a_29583_30440 a_28027_31160.t5 Vss.t76 Vss.t75 nfet_03v3
**devattr s=17600,576 d=17600,576
X727 SARlogic_0.dffrs_13.nand3_1.C.t1 SARlogic_0.dffrs_13.nand3_6.C.t7 Vdd.t630 Vdd.t629 pfet_03v3
**devattr s=26000,604 d=44000,1176
X728 SARlogic_0.dffrs_10.nand3_8.C.t0 SARlogic_0.dffrs_10.nand3_6.C.t9 Vdd.t201 Vdd.t200 pfet_03v3
**devattr s=44000,1176 d=26000,604
X729 a_n4631_31422.t0 Clk_piso.t17 a_n4367_33719 Vss.t81 nfet_03v3
**devattr s=10400,304 d=17600,576
X730 SARlogic_0.dffrs_4.d.t0 SARlogic_0.dffrs_3.Qb.t9 a_5987_11838 Vss.t194 nfet_03v3
**devattr s=10400,304 d=17600,576
X731 adc_PISO_0.dffrs_2.Q.t1 adc_PISO_0.dffrs_2.Qb a_16063_33720 Vss.t384 nfet_03v3
**devattr s=10400,304 d=17600,576
X732 a_n3065_33719 Vdd.t973 Vss.t409 Vss.t408 nfet_03v3
**devattr s=17600,576 d=10400,304
X733 SARlogic_0.dffrs_14.nand3_8.C.t1 SARlogic_0.dffrs_14.nand3_6.C.t9 Vdd.t778 Vdd.t777 pfet_03v3
**devattr s=44000,1176 d=26000,604
X734 a_n9861_31159.t3 inv2_0.out.t25 Vdd.t760 Vdd.t759 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X735 Piso_out.t1 adc_PISO_0.dffrs_5.Qb a_44479_33720 Vss.t274 nfet_03v3
**devattr s=10400,304 d=17600,576
X736 a_n2281_11838 Vdd.t974 Vss.t407 Vss.t406 nfet_03v3
**devattr s=17600,576 d=10400,304
X737 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t15 Vdd.t233 Vdd.t232 pfet_03v3
**devattr s=10400,304 d=10400,304
X738 a_n8305_30439 a_n9861_31159.t5 Vss.t205 Vss.t204 nfet_03v3
**devattr s=17600,576 d=17600,576
X739 a_16063_33720 a_14313_31423.t9 a_15879_33720 Vss.t603 nfet_03v3
**devattr s=10400,304 d=10400,304
X740 a_n2881_33719 a_n4631_31422.t8 a_n3065_33719 Vss.t158 nfet_03v3
**devattr s=10400,304 d=10400,304
X741 SARlogic_0.dffrs_2.nand3_8.C.t2 SARlogic_0.dffrs_2.nand3_8.Z.t7 a_459_9633 Vss.t473 nfet_03v3
**devattr s=10400,304 d=17600,576
X742 SARlogic_0.dffrs_2.Qb.t3 Reset.t66 Vdd.t347 Vdd.t346 pfet_03v3
**devattr s=26000,604 d=44000,1176
X743 Vss.t260 a_n10831_4320 Comp_out.t1 Vss.t259 nfet_03v3
**devattr s=9350,280 d=9350,280
X744 a_10639_28100 a_9083_28820.t5 Vss.t60 Vss.t59 nfet_03v3
**devattr s=17600,576 d=17600,576
X745 SARlogic_0.dffrs_1.nand3_8.C.t0 SARlogic_0.dffrs_1.nand3_8.Z.t6 Vdd.t620 Vdd.t619 pfet_03v3
**devattr s=26000,604 d=44000,1176
X746 SARlogic_0.dffrs_3.nand3_8.Z.t3 SARlogic_0.dffrs_2.Q.t7 a_4501_7428 Vss.t571 nfet_03v3
**devattr s=10400,304 d=17600,576
X747 SARlogic_0.dffrs_14.nand3_6.C.t1 SARlogic_0.dffrs_14.nand3_1.C Vdd.t395 Vdd.t394 pfet_03v3
**devattr s=44000,1176 d=26000,604
X748 Vss.t226 adc_PISO_0.dffrs_3.Q.t8 a_28215_30440 Vss.t225 nfet_03v3
**devattr s=10400,304 d=17600,576
X749 Vss.t56 a_36793_29020 a_37687_28100 Vss.t55 nfet_03v3
**devattr s=10400,304 d=17600,576
X750 a_1167_30439 a_n389_31159.t5 Vss.t312 Vss.t311 nfet_03v3
**devattr s=17600,576 d=17600,576
X751 Vdd.t197 SARlogic_0.dffrs_2.nand3_8.C.t6 SARlogic_0.dffrs_2.Qb.t0 Vdd.t196 pfet_03v3
**devattr s=26000,604 d=26000,604
X752 SARlogic_0.dffrs_5.nand3_8.Z.t0 SARlogic_0.dffrs_5.nand3_8.C.t7 Vdd.t61 Vdd.t60 pfet_03v3
**devattr s=44000,1176 d=26000,604
X753 SARlogic_0.dffrs_8.nand3_8.C.t1 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t5 Vdd.t4 pfet_03v3
**devattr s=26000,604 d=44000,1176
X754 SARlogic_0.dffrs_1.nand3_6.C.t2 Clk.t24 Vdd.t724 Vdd.t723 pfet_03v3
**devattr s=26000,604 d=44000,1176
X755 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t8 Vdd.t379 Vdd.t378 pfet_03v3
**devattr s=26000,604 d=44000,1176
X756 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_8.C.t7 Vdd.t227 Vdd.t226 pfet_03v3
**devattr s=44000,1176 d=26000,604
X757 Vdd.t688 Clk.t25 SARlogic_0.dffrs_13.nand3_8.C.t3 Vdd.t687 pfet_03v3
**devattr s=26000,604 d=26000,604
X758 SARlogic_0.dffrs_1.nand3_8.C.t1 SARlogic_0.dffrs_1.nand3_8.Z.t7 a_n3583_9633 Vss.t468 nfet_03v3
**devattr s=10400,304 d=17600,576
X759 a_459_11838 Reset.t67 a_275_11838 Vss.t282 nfet_03v3
**devattr s=10400,304 d=10400,304
X760 SARlogic_0.dffrs_2.nand3_8.Z.t0 SARlogic_0.dffrs_2.nand3_8.C.t7 Vdd.t223 Vdd.t222 pfet_03v3
**devattr s=44000,1176 d=26000,604
X761 SARlogic_0.dffrs_11.nand3_6.C.t1 SARlogic_0.dffrs_12.Q.t9 a_12585_21414 Vss.t465 nfet_03v3
**devattr s=10400,304 d=17600,576
X762 Vdd.t333 Reset.t68 SARlogic_0.dffrs_11.nand3_6.C.t2 Vdd.t332 pfet_03v3
**devattr s=26000,604 d=26000,604
X763 Vdd.t904 SARlogic_0.dffrs_9.nand3_6.C.t8 adc_PISO_0.B3.t3 Vdd.t903 pfet_03v3
**devattr s=26000,604 d=26000,604
X764 adc_PISO_0.dffrs_2.Qb Vdd.t975 a_16063_31516 Vss.t405 nfet_03v3
**devattr s=10400,304 d=17600,576
X765 a_n3767_17004 SARlogic_0.dffrs_7.nand3_8.C.t7 Vss.t646 Vss.t645 nfet_03v3
**devattr s=17600,576 d=10400,304
X766 Vdd.t488 Vdd.t486 SARlogic_0.dffrs_13.nand3_6.C.t0 Vdd.t487 pfet_03v3
**devattr s=26000,604 d=26000,604
X767 Vdd.t640 SARlogic_0.dffrs_4.nand3_8.C.t7 SARlogic_0.dffrs_4.Qb.t0 Vdd.t639 pfet_03v3
**devattr s=26000,604 d=26000,604
X768 adc_PISO_0.dffrs_5.Qb Vdd.t976 a_44479_31516 Vss.t404 nfet_03v3
**devattr s=10400,304 d=17600,576
X769 a_16063_31516 a_14313_29218.t7 a_15879_31516 Vss.t667 nfet_03v3
**devattr s=10400,304 d=10400,304
X770 a_6591_33719 a_4841_31422.t8 a_6407_33719 Vss.t50 nfet_03v3
**devattr s=10400,304 d=10400,304
X771 a_n4631_33627.t2 Vdd.t483 Vdd.t485 Vdd.t484 pfet_03v3
**devattr s=44000,1176 d=26000,604
X772 SARlogic_0.dffrs_0.nand3_1.C.t1 SARlogic_0.dffrs_0.nand3_6.C.t9 a_n7625_14043 Vss.t188 nfet_03v3
**devattr s=10400,304 d=17600,576
X773 a_42729_31423.t0 Clk_piso.t18 a_42993_33720 Vss.t82 nfet_03v3
**devattr s=10400,304 d=17600,576
X774 a_33337_30170.t0 adc_PISO_0.2inmux_5.OUT.t3 Vdd.t13 Vdd.t12 pfet_03v3
**devattr s=26000,604 d=44000,1176
X775 a_n3767_19209 SARlogic_0.dffrs_7.nand3_6.C.t9 Vss.t549 Vss.t548 nfet_03v3
**devattr s=17600,576 d=10400,304
X776 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t9 a_12585_23619 Vss.t182 nfet_03v3
**devattr s=10400,304 d=17600,576
X777 Vdd.t171 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_1.C Vdd.t170 pfet_03v3
**devattr s=26000,604 d=26000,604
X778 a_14577_33720 Vdd.t977 a_14393_33720 Vss.t403 nfet_03v3
**devattr s=10400,304 d=10400,304
X779 a_14313_31423.t2 a_14313_33628.t5 Vdd.t267 Vdd.t266 pfet_03v3
**devattr s=44000,1176 d=26000,604
X780 a_n2281_9634 SARlogic_0.dffrs_2.d.t6 Vss.t378 Vss.t377 nfet_03v3
**devattr s=17600,576 d=10400,304
X781 a_n7625_9633 Clk.t26 a_n7809_9633 Vss.t501 nfet_03v3
**devattr s=10400,304 d=10400,304
X782 a_14393_30170.t1 adc_PISO_0.2inmux_3.OUT.t3 a_14577_29310 Vss.t374 nfet_03v3
**devattr s=10400,304 d=17600,576
X783 a_11311_29264.t0 a_10639_28100 a_11499_29984 Vdd.t152 pfet_03v3
**devattr s=31200,704 d=52800,1376
X784 a_42729_33628.t1 a_42729_31423.t7 a_42993_35925 Vss.t249 nfet_03v3
**devattr s=10400,304 d=17600,576
X785 a_4501_21414 Reset.t69 a_4317_21414 Vss.t283 nfet_03v3
**devattr s=10400,304 d=10400,304
X786 a_33257_29218.t1 a_33337_30170.t7 Vdd.t890 Vdd.t889 pfet_03v3
**devattr s=26000,604 d=44000,1176
X787 SARlogic_0.dffrs_1.nand3_1.C.t3 Vdd.t477 Vdd.t479 Vdd.t478 pfet_03v3
**devattr s=44000,1176 d=26000,604
X788 a_n9429_n2007.t19 Vin1.t6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t6 Vss.t372 nfet_03v3
**devattr s=15600,404 d=15600,404
X789 SARlogic_0.dffrs_8.nand3_8.C.t2 SARlogic_0.dffrs_8.nand3_6.C.t9 Vdd.t243 Vdd.t242 pfet_03v3
**devattr s=44000,1176 d=26000,604
X790 a_39915_29984 a_39055_30440 Vdd.t708 Vdd.t707 pfet_03v3
**devattr s=52800,1376 d=31200,704
X791 a_14577_35925 a_14393_30170.t7 a_14393_35925 Vss.t84 nfet_03v3
**devattr s=10400,304 d=10400,304
X792 a_14313_33628.t1 Vdd.t480 Vdd.t482 Vdd.t481 pfet_03v3
**devattr s=44000,1176 d=26000,604
X793 a_n10151_11838 SARlogic_0.dffrs_13.nand3_6.C.t8 a_n10335_11838 Vss.t471 nfet_03v3
**devattr s=10400,304 d=10400,304
X794 a_5987_19210 SARlogic_0.dffrs_9.nand3_8.C.t6 a_5803_19210 Vss.t191 nfet_03v3
**devattr s=10400,304 d=10400,304
X795 a_4501_23619 SARlogic_0.dffrs_9.nand3_8.Z a_4317_23619 Vss.t461 nfet_03v3
**devattr s=10400,304 d=10400,304
X796 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_8.C.t7 Vdd.t259 Vdd.t258 pfet_03v3
**devattr s=44000,1176 d=26000,604
X797 Vdd.t235 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t16 comparator_no_offsetcal_0.x5.out Vdd.t234 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X798 a_n3583_7428 Reset.t70 a_n3767_7428 Vss.t284 nfet_03v3
**devattr s=10400,304 d=10400,304
X799 Vdd.t766 Vss.t679 SARlogic_0.dffrs_12.nand3_8.C.t2 Vdd.t765 pfet_03v3
**devattr s=26000,604 d=26000,604
X800 a_5105_31514 Clk_piso.t19 a_4921_31514 Vss.t331 nfet_03v3
**devattr s=10400,304 d=10400,304
X801 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t9 a_n3583_17004 Vss.t309 nfet_03v3
**devattr s=10400,304 d=17600,576
X802 adc_PISO_0.2inmux_2.OUT.t1 a_1839_29263.t5 Vdd.t706 Vdd.t705 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X803 a_4921_31514 a_4841_31422.t9 Vss.t52 Vss.t51 nfet_03v3
**devattr s=17600,576 d=10400,304
X804 a_20783_29264.t3 a_20111_28100 Vss.t252 Vss.t251 nfet_03v3
**devattr s=17600,576 d=17600,576
X805 a_5105_33719 Vdd.t978 a_4921_33719 Vss.t402 nfet_03v3
**devattr s=10400,304 d=10400,304
X806 a_n4631_33627.t0 a_n4631_31422.t9 Vdd.t183 Vdd.t182 pfet_03v3
**devattr s=26000,604 d=44000,1176
X807 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t5 Vin1.t7 a_n9429_n2007.t20 Vss.t373 nfet_03v3
**devattr s=15600,404 d=15600,404
X808 SARlogic_0.dffrs_2.Qb.t2 Reset.t71 a_1945_9634 Vss.t285 nfet_03v3
**devattr s=10400,304 d=17600,576
X809 a_33337_30170.t1 a_33257_29218.t7 Vdd.t29 Vdd.t28 pfet_03v3
**devattr s=44000,1176 d=26000,604
X810 a_42993_31515 Clk_piso.t20 a_42809_31515 Vss.t332 nfet_03v3
**devattr s=10400,304 d=10400,304
X811 a_8543_14043 SARlogic_0.dffrs_4.nand3_8.Z.t7 a_8359_14043 Vss.t335 nfet_03v3
**devattr s=10400,304 d=10400,304
X812 SARlogic_0.dffrs_7.nand3_8.C.t1 SARlogic_0.dffrs_7.nand3_8.Z a_n3583_19209 Vss.t61 nfet_03v3
**devattr s=10400,304 d=17600,576
X813 a_28215_28100 a_27321_29020 Vss.t557 Vss.t556 nfet_03v3
**devattr s=17600,576 d=10400,304
X814 adc_PISO_0.2inmux_3.OUT.t1 a_11311_29264.t5 Vdd.t431 Vdd.t430 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X815 a_4921_33719 a_4841_33627.t5 Vss.t652 Vss.t651 nfet_03v3
**devattr s=17600,576 d=10400,304
X816 a_n7809_7428 SARlogic_0.dffrs_0.nand3_8.C.t7 Vss.t219 Vss.t218 nfet_03v3
**devattr s=17600,576 d=10400,304
X817 Vss.t258 a_n10831_4320 Comp_out.t0 Vss.t257 nfet_03v3
**devattr s=9350,280 d=9350,280
X818 SARlogic_0.dffrs_13.Qb.t1 Vdd.t979 a_n10151_9634 Vss.t401 nfet_03v3
**devattr s=10400,304 d=17600,576
X819 SARlogic_0.dffrs_1.nand3_1.C.t2 SARlogic_0.dffrs_1.nand3_6.C.t8 Vdd.t844 Vdd.t843 pfet_03v3
**devattr s=26000,604 d=44000,1176
X820 a_17849_29020 inv2_0.out.t26 Vss.t588 Vss.t587 nfet_03v3
**devattr s=17600,576 d=17600,576
X821 a_33257_29218.t2 a_33257_31423.t9 Vdd.t241 Vdd.t240 pfet_03v3
**devattr s=44000,1176 d=26000,604
X822 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t4 Vin1.t8 a_n9429_n2007.t5 Vss.t166 nfet_03v3
**devattr s=15600,404 d=15600,404
X823 a_24049_29310 Vdd.t980 a_23865_29310 Vss.t400 nfet_03v3
**devattr s=10400,304 d=10400,304
X824 a_n4367_31514 Clk_piso.t21 a_n4551_31514 Vss.t386 nfet_03v3
**devattr s=10400,304 d=10400,304
X825 adc_PISO_0.dffrs_0.Qb adc_PISO_0.2inmux_2.Bit.t8 Vdd.t942 Vdd.t941 pfet_03v3
**devattr s=44000,1176 d=26000,604
X826 SARlogic_0.dffrs_3.Qb.t3 Reset.t72 Vdd.t335 Vdd.t334 pfet_03v3
**devattr s=26000,604 d=44000,1176
X827 a_n9429_n2007.t21 Clk.t27 Vss.t503 Vss.t502 nfet_03v3
**devattr s=8320,264 d=8320,264
X828 SARlogic_0.dffrs_1.Qb.t1 SARlogic_0.dffrs_2.d.t7 Vdd.t429 Vdd.t428 pfet_03v3
**devattr s=44000,1176 d=26000,604
X829 a_n389_28819.t2 adc_PISO_0.B5.t9 a_n201_28099 Vss.t379 nfet_03v3
**devattr s=10400,304 d=17600,576
X830 Vdd.t139 SARlogic_0.dffrs_13.nand3_8.Z.t7 SARlogic_0.dffrs_13.nand3_1.C.t2 Vdd.t138 pfet_03v3
**devattr s=26000,604 d=26000,604
X831 Vdd.t293 a_n4631_29217.t6 adc_PISO_0.dffrs_0.Qb Vdd.t292 pfet_03v3
**devattr s=26000,604 d=26000,604
X832 Vdd.t337 Reset.t73 SARlogic_0.dffrs_5.nand3_8.Z.t3 Vdd.t336 pfet_03v3
**devattr s=26000,604 d=26000,604
X833 a_n4367_33719 Vdd.t981 a_n4551_33719 Vss.t399 nfet_03v3
**devattr s=10400,304 d=10400,304
X834 a_n3583_11838 Reset.t74 a_n3767_11838 Vss.t490 nfet_03v3
**devattr s=10400,304 d=10400,304
X835 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_8.C.t7 Vdd.t788 Vdd.t787 pfet_03v3
**devattr s=44000,1176 d=26000,604
X836 a_n4551_29309 a_n4631_29217.t7 Vss.t256 Vss.t255 nfet_03v3
**devattr s=17600,576 d=10400,304
X837 a_n9429_n2007.t12 Vin2.t8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t362 nfet_03v3
**devattr s=15600,404 d=15600,404
X838 a_n389_28819.t3 adc_PISO_0.B5.t10 Vdd.t457 Vdd.t456 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X839 a_30443_29984 a_29583_28100 a_30255_29264.t0 Vdd.t10 pfet_03v3
**devattr s=52800,1376 d=31200,704
X840 Vdd.t660 Reset.t75 SARlogic_0.dffrs_2.nand3_8.Z.t3 Vdd.t659 pfet_03v3
**devattr s=26000,604 d=26000,604
X841 a_n11821_11838 SARlogic_0.dffrs_13.nand3_1.C.t5 Vss.t464 Vss.t463 nfet_03v3
**devattr s=17600,576 d=10400,304
X842 SARlogic_0.dffrs_5.nand3_8.C.t1 SARlogic_0.dffrs_5.nand3_8.Z.t7 Vdd.t35 Vdd.t34 pfet_03v3
**devattr s=26000,604 d=44000,1176
X843 Vss.t42 a_n8305_30439 a_n7633_29263.t0 Vss.t41 nfet_03v3
**devattr s=17600,576 d=17600,576
X844 SARlogic_0.dffrs_14.nand3_8.C.t2 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t782 Vdd.t781 pfet_03v3
**devattr s=26000,604 d=44000,1176
X845 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t9 a_n9429_n2007.t13 Vss.t363 nfet_03v3
**devattr s=15600,404 d=15600,404
X846 Vdd.t662 Reset.t76 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t661 pfet_03v3
**devattr s=26000,604 d=26000,604
X847 SARlogic_0.dffrs_5.nand3_6.C.t1 Clk.t28 Vdd.t690 Vdd.t689 pfet_03v3
**devattr s=26000,604 d=44000,1176
X848 SARlogic_0.dffrs_14.nand3_6.C.t2 adc_PISO_0.B5.t11 Vdd.t459 Vdd.t458 pfet_03v3
**devattr s=26000,604 d=44000,1176
X849 adc_PISO_0.B6.t1 SARlogic_0.dffrs_13.Qb.t8 Vdd.t187 Vdd.t186 pfet_03v3
**devattr s=44000,1176 d=26000,604
X850 Vdd.t113 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t112 pfet_03v3
**devattr s=17600,576 d=17600,576
X851 a_n9673_28099 adc_PISO_0.B6.t7 a_n9861_28819.t2 Vss.t574 nfet_03v3
**devattr s=17600,576 d=10400,304
X852 adc_PISO_0.dffrs_1.Qb Vdd.t982 a_6591_31515 Vss.t398 nfet_03v3
**devattr s=10400,304 d=17600,576
X853 Vdd.t443 a_4841_29217.t6 adc_PISO_0.dffrs_1.Qb Vdd.t442 pfet_03v3
**devattr s=26000,604 d=26000,604
X854 a_11499_29984 a_10639_30440 Vdd.t818 Vdd.t817 pfet_03v3
**devattr s=52800,1376 d=31200,704
X855 a_23865_30170.t2 adc_PISO_0.2inmux_4.OUT.t3 Vdd.t97 Vdd.t96 pfet_03v3
**devattr s=26000,604 d=44000,1176
X856 adc_PISO_0.B1.t2 SARlogic_0.dffrs_4.Qb.t8 Vdd.t177 Vdd.t176 pfet_03v3
**devattr s=44000,1176 d=26000,604
X857 Vss.t277 comparator_no_offsetcal_0.x5.out comparator_no_offsetcal_0.x2.Vout2 Vss.t276 nfet_03v3
**devattr s=17600,576 d=17600,576
X858 a_18743_30440 inv2_0.out.t27 a_18555_31160.t1 Vss.t589 nfet_03v3
**devattr s=17600,576 d=10400,304
X859 Vdd.t692 Clk.t29 SARlogic_0.dffrs_3.nand3_8.C.t2 Vdd.t691 pfet_03v3
**devattr s=26000,604 d=26000,604
X860 a_n9429_n2007.t6 Vin1.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t3 Vss.t153 nfet_03v3
**devattr s=15600,404 d=15600,404
X861 Piso_out.t2 Vdd.t474 Vdd.t476 Vdd.t475 pfet_03v3
**devattr s=44000,1176 d=26000,604
X862 a_44479_33720 a_42729_31423.t8 a_44295_33720 Vss.t21 nfet_03v3
**devattr s=10400,304 d=10400,304
X863 a_n2097_11838 SARlogic_0.dffrs_1.nand3_6.C.t9 a_n2281_11838 Vss.t597 nfet_03v3
**devattr s=10400,304 d=10400,304
X864 a_n7625_14043 SARlogic_0.dffrs_0.nand3_8.Z.t7 a_n7809_14043 Vss.t478 nfet_03v3
**devattr s=10400,304 d=10400,304
X865 adc_PISO_0.2inmux_2.Bit.t1 adc_PISO_0.dffrs_0.Qb a_n2881_33719 Vss.t68 nfet_03v3
**devattr s=10400,304 d=17600,576
X866 a_15879_33720 Vdd.t983 Vss.t397 Vss.t396 nfet_03v3
**devattr s=17600,576 d=10400,304
X867 a_23785_29218.t0 a_23865_30170.t7 Vdd.t287 Vdd.t286 pfet_03v3
**devattr s=26000,604 d=44000,1176
X868 a_n4551_30169.t1 adc_PISO_0.2inmux_0.OUT.t3 a_n4367_29309 Vss.t353 nfet_03v3
**devattr s=10400,304 d=17600,576
X869 Vdd.t826 a_4921_30169.t6 a_4841_33627.t3 Vdd.t825 pfet_03v3
**devattr s=26000,604 d=26000,604
X870 Vdd.t664 Reset.t77 SARlogic_0.dffrs_3.nand3_6.C.t3 Vdd.t663 pfet_03v3
**devattr s=26000,604 d=26000,604
X871 Vdd.t473 Vdd.t471 a_42729_31423.t2 Vdd.t472 pfet_03v3
**devattr s=26000,604 d=26000,604
X872 Vdd.t632 SARlogic_0.dffrs_13.nand3_8.C.t7 SARlogic_0.dffrs_13.Qb.t3 Vdd.t631 pfet_03v3
**devattr s=26000,604 d=26000,604
X873 SARlogic_0.dffrs_2.d.t2 SARlogic_0.dffrs_1.Qb.t9 a_n2097_11838 Vss.t38 nfet_03v3
**devattr s=10400,304 d=17600,576
X874 a_n3767_7428 SARlogic_0.dffrs_1.nand3_8.C.t7 Vss.t141 Vss.t140 nfet_03v3
**devattr s=17600,576 d=10400,304
X875 a_4841_33627.t2 Vdd.t468 Vdd.t470 Vdd.t469 pfet_03v3
**devattr s=44000,1176 d=26000,604
X876 SARlogic_0.dffrs_9.nand3_6.C.t1 adc_PISO_0.B2.t11 a_4501_21414 Vss.t499 nfet_03v3
**devattr s=10400,304 d=17600,576
X877 a_5803_21414 SARlogic_0.dffrs_2.Qb.t8 Vss.t381 Vss.t380 nfet_03v3
**devattr s=17600,576 d=10400,304
X878 a_12401_21414 SARlogic_0.dffrs_11.nand3_1.C Vss.t269 Vss.t268 nfet_03v3
**devattr s=17600,576 d=10400,304
X879 a_8543_9633 Clk.t30 a_8359_9633 Vss.t504 nfet_03v3
**devattr s=10400,304 d=10400,304
X880 Vdd.t666 Reset.t78 SARlogic_0.dffrs_10.nand3_6.C.t3 Vdd.t665 pfet_03v3
**devattr s=26000,604 d=26000,604
X881 Vdd.t922 adc_PISO_0.B3.t11 SARlogic_0.dffrs_8.nand3_8.C.t3 Vdd.t921 pfet_03v3
**devattr s=26000,604 d=26000,604
X882 SARlogic_0.dffrs_13.nand3_6.C.t2 Clk.t31 a_n11637_11838 Vss.t518 nfet_03v3
**devattr s=10400,304 d=17600,576
X883 Vdd.t846 a_42809_30170.t7 a_42729_33628.t3 Vdd.t845 pfet_03v3
**devattr s=26000,604 d=26000,604
X884 a_20111_30440 a_18555_31160.t5 Vdd.t467 Vdd.t466 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X885 a_n10335_11838 Reset.t79 Vss.t492 Vss.t491 nfet_03v3
**devattr s=17600,576 d=10400,304
X886 a_n6693_1497 a_n6893_1405 Vdd.t463 Vdd.t462 pfet_03v3
**devattr s=10400,304 d=17600,576
X887 a_n6323_19213 adc_PISO_0.B6.t8 Vss.t576 Vss.t575 nfet_03v3
**devattr s=17600,576 d=10400,304
X888 a_9845_9634 SARlogic_0.dffrs_4.Q.t7 Vss.t357 Vss.t356 nfet_03v3
**devattr s=17600,576 d=10400,304
X889 a_37499_31160.t2 inv2_0.out.t28 Vdd.t838 Vdd.t837 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X890 Vss.t91 a_n10567_29019 a_n9673_28099 Vss.t90 nfet_03v3
**devattr s=10400,304 d=17600,576
X891 Vdd.t251 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_1.C Vdd.t250 pfet_03v3
**devattr s=26000,604 d=26000,604
X892 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t9 a_4501_23619 Vss.t635 nfet_03v3
**devattr s=10400,304 d=17600,576
X893 a_12401_23619 SARlogic_0.dffrs_4.Qb.t9 Vss.t157 Vss.t156 nfet_03v3
**devattr s=17600,576 d=10400,304
X894 a_13887_19210 adc_PISO_0.B1.t12 Vss.t322 Vss.t321 nfet_03v3
**devattr s=17600,576 d=10400,304
X895 a_n389_31159.t1 inv2_0.out.t29 a_n201_30439 Vss.t590 nfet_03v3
**devattr s=10400,304 d=17600,576
X896 a_4841_29217.t3 a_4921_30169.t7 a_5105_31514 Vss.t566 nfet_03v3
**devattr s=10400,304 d=17600,576
X897 a_11311_29264.t2 a_10639_28100 Vss.t136 Vss.t135 nfet_03v3
**devattr s=17600,576 d=17600,576
X898 adc_PISO_0.B6.t2 SARlogic_0.dffrs_14.Qb Vdd.t279 Vdd.t278 pfet_03v3
**devattr s=26000,604 d=44000,1176
X899 a_33521_31515 Clk_piso.t22 a_33337_31515 Vss.t387 nfet_03v3
**devattr s=10400,304 d=10400,304
X900 adc_PISO_0.dffrs_5.Qb Piso_out.t5 Vdd.t449 Vdd.t448 pfet_03v3
**devattr s=44000,1176 d=26000,604
X901 a_44479_31516 a_42729_29218.t7 a_44295_31516 Vss.t294 nfet_03v3
**devattr s=10400,304 d=10400,304
X902 Vdd.t626 a_n4551_30169.t7 a_n4631_33627.t3 Vdd.t625 pfet_03v3
**devattr s=26000,604 d=26000,604
X903 a_4841_31422.t2 Clk_piso.t23 a_5105_33719 Vss.t472 nfet_03v3
**devattr s=10400,304 d=17600,576
X904 a_6407_33719 Vdd.t984 Vss.t395 Vss.t394 nfet_03v3
**devattr s=17600,576 d=10400,304
X905 a_15879_31516 adc_PISO_0.dffrs_2.Q.t7 Vss.t637 Vss.t636 nfet_03v3
**devattr s=17600,576 d=10400,304
X906 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t16 a_n9933_n1136 a_n10021_n1044 Vss.t228 nfet_03v3
**devattr s=26400,776 d=15600,404
X907 adc_PISO_0.2inmux_0.OUT.t0 a_n7633_29263.t5 Vss.t338 Vss.t337 nfet_03v3
**devattr s=17600,576 d=17600,576
X908 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t10 a_12585_17004 Vss.t310 nfet_03v3
**devattr s=10400,304 d=17600,576
X909 a_36793_29020 inv2_0.out.t30 Vss.t592 Vss.t591 nfet_03v3
**devattr s=17600,576 d=17600,576
X910 Vdd.t295 a_n10831_4320 Comp_out.t4 Vdd.t294 pfet_03v3
**devattr s=18700,450 d=18700,450
X911 SARlogic_0.dffrs_4.nand3_1.C.t2 SARlogic_0.dffrs_4.nand3_6.C.t9 a_8543_14043 Vss.t371 nfet_03v3
**devattr s=10400,304 d=17600,576
X912 a_42809_30170.t2 adc_PISO_0.2inmux_1.OUT.t3 a_42993_29310 Vss.t352 nfet_03v3
**devattr s=10400,304 d=17600,576
X913 a_14577_29310 Vdd.t985 a_14393_29310 Vss.t393 nfet_03v3
**devattr s=10400,304 d=10400,304
X914 SARlogic_0.dffrs_11.nand3_8.C.t0 SARlogic_0.dffrs_11.nand3_8.Z a_12585_19209 Vss.t151 nfet_03v3
**devattr s=10400,304 d=17600,576
X915 a_4317_21414 SARlogic_0.dffrs_9.nand3_1.C Vss.t302 Vss.t301 nfet_03v3
**devattr s=17600,576 d=10400,304
X916 SARlogic_0.dffrs_0.d.t1 SARlogic_0.dffrs_13.Qb.t9 a_n10151_11838 Vss.t165 nfet_03v3
**devattr s=10400,304 d=17600,576
X917 a_39055_30440 a_37499_31160.t5 Vdd.t165 Vdd.t164 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X918 Vdd.t141 a_29583_30440 a_30443_29984 Vdd.t140 pfet_03v3
**devattr s=31200,704 d=52800,1376
X919 a_4501_17004 Reset.t80 a_4317_17004 Vss.t493 nfet_03v3
**devattr s=10400,304 d=10400,304
X920 a_18555_28820.t1 adc_PISO_0.B3.t12 a_18743_28100 Vss.t661 nfet_03v3
**devattr s=10400,304 d=17600,576
X921 SARlogic_0.dffrs_14.Qb Reset.t81 a_n6139_19213 Vss.t523 nfet_03v3
**devattr s=10400,304 d=17600,576
X922 a_n11821_9633 SARlogic_0.dffrs_13.nand3_6.C.t9 Vss.t599 Vss.t598 nfet_03v3
**devattr s=17600,576 d=10400,304
X923 SARlogic_0.dffrs_5.nand3_1.C.t2 SARlogic_0.dffrs_5.nand3_6.C.t8 Vdd.t167 Vdd.t166 pfet_03v3
**devattr s=26000,604 d=44000,1176
X924 a_4317_23619 SARlogic_0.dffrs_2.Qb.t9 Vss.t383 Vss.t382 nfet_03v3
**devattr s=17600,576 d=10400,304
X925 adc_PISO_0.2inmux_1.Bit.t2 adc_PISO_0.dffrs_4.Qb Vdd.t938 Vdd.t937 pfet_03v3
**devattr s=26000,604 d=44000,1176
X926 a_n9673_30439 inv2_0.out.t31 a_n9861_31159.t1 Vss.t593 nfet_03v3
**devattr s=17600,576 d=10400,304
X927 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t17 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t5 Vss.t210 nfet_03v3
**devattr s=20800,504 d=20800,504
X928 a_4501_19209 adc_PISO_0.B2.t12 a_4317_19209 Vss.t500 nfet_03v3
**devattr s=10400,304 d=10400,304
X929 SARlogic_0.dffrs_5.Q.t1 SARlogic_0.dffrs_5.Qb.t9 a_14071_11838 Vss.t29 nfet_03v3
**devattr s=10400,304 d=17600,576
X930 a_n3767_11838 SARlogic_0.dffrs_1.nand3_1.C.t5 Vss.t54 Vss.t53 nfet_03v3
**devattr s=17600,576 d=10400,304
X931 Vdd.t65 SARlogic_0.dffrs_3.nand3_8.Z.t7 SARlogic_0.dffrs_3.nand3_1.C.t0 Vdd.t64 pfet_03v3
**devattr s=26000,604 d=26000,604
X932 a_42809_31515 a_42729_31423.t9 Vss.t23 Vss.t22 nfet_03v3
**devattr s=17600,576 d=10400,304
X933 a_14071_11838 SARlogic_0.dffrs_5.nand3_6.C.t9 a_13887_11838 Vss.t147 nfet_03v3
**devattr s=10400,304 d=10400,304
X934 Vss.t639 adc_PISO_0.dffrs_2.Q.t8 a_18743_30440 Vss.t638 nfet_03v3
**devattr s=10400,304 d=17600,576
X935 a_5105_29309 Vdd.t986 a_4921_29309 Vss.t392 nfet_03v3
**devattr s=10400,304 d=10400,304
X936 Vdd.t870 SARlogic_0.dffrs_12.nand3_6.C.t9 SARlogic_0.dffrs_12.Q.t3 Vdd.t869 pfet_03v3
**devattr s=26000,604 d=26000,604
X937 SARlogic_0.dffrs_13.nand3_8.Z.t1 Vss.t680 Vdd.t768 Vdd.t767 pfet_03v3
**devattr s=26000,604 d=44000,1176
X938 a_8359_14043 Vdd.t987 Vss.t391 Vss.t390 nfet_03v3
**devattr s=17600,576 d=10400,304
X939 a_4921_29309 a_4841_29217.t7 Vss.t365 Vss.t364 nfet_03v3
**devattr s=17600,576 d=10400,304
X940 SARlogic_0.dffrs_12.nand3_6.C.t2 Vss.t681 Vdd.t770 Vdd.t769 pfet_03v3
**devattr s=26000,604 d=44000,1176
X941 a_4501_9633 Clk.t32 a_4317_9633 Vss.t519 nfet_03v3
**devattr s=10400,304 d=10400,304
X942 a_9083_28820.t2 adc_PISO_0.B4.t12 Vdd.t83 Vdd.t82 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X943 Vdd.t127 adc_PISO_0.B5.t12 SARlogic_0.dffrs_14.nand3_8.C.t0 Vdd.t126 pfet_03v3
**devattr s=26000,604 d=26000,604
X944 Vdd.t898 adc_PISO_0.dffrs_1.Q.t8 a_9083_31160.t0 Vdd.t897 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X945 Vss.t123 Vss.t121 a_n9673_30439 Vss.t122 nfet_03v3
**devattr s=10400,304 d=17600,576
X946 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t11 Vdd.t327 Vdd.t326 pfet_03v3
**devattr s=26000,604 d=44000,1176
R0 adc_PISO_0.B4.n3 adc_PISO_0.B4.t8 41.0041
R1 adc_PISO_0.B4.n4 adc_PISO_0.B4.t4 40.8177
R2 adc_PISO_0.B4.n7 adc_PISO_0.B4.t7 40.6313
R3 adc_PISO_0.B4.n1 adc_PISO_0.B4.t12 34.2529
R4 adc_PISO_0.B4.n6 SARlogic_0.dffrs_7.clk 33.3108
R5 adc_PISO_0.B4.n7 adc_PISO_0.B4.t5 27.3166
R6 adc_PISO_0.B4.n4 adc_PISO_0.B4.t10 27.1302
R7 adc_PISO_0.B4.n3 adc_PISO_0.B4.t9 26.9438
R8 adc_PISO_0.B4.n0 adc_PISO_0.B4.t6 19.673
R9 adc_PISO_0.B4.n0 adc_PISO_0.B4.t11 19.4007
R10 adc_PISO_0.B4.n9 adc_PISO_0.B4.n8 14.0582
R11 adc_PISO_0.B4.n9 adc_PISO_0.B4.n6 11.1633
R12 SARlogic_0.d3 adc_PISO_0.B4.n2 10.6816
R13 adc_PISO_0.B4.n12 adc_PISO_0.B4.t1 10.0473
R14 adc_PISO_0.B4.n2 adc_PISO_0.B4.n1 8.05164
R15 adc_PISO_0.B4.n11 adc_PISO_0.B4.t0 6.51042
R16 adc_PISO_0.B4.n11 adc_PISO_0.B4.n10 6.04952
R17 SARlogic_0.dffrs_7.nand3_1.A adc_PISO_0.B4.n3 5.7755
R18 SARlogic_0.dffrs_7.nand3_6.B adc_PISO_0.B4.n4 5.47979
R19 adc_PISO_0.B4.n8 adc_PISO_0.B4.n7 5.13907
R20 SARlogic_0.dffrs_8.nand3_2.Z adc_PISO_0.B4.n12 4.72925
R21 adc_PISO_0.B4.n5 SARlogic_0.dffrs_7.nand3_6.B 2.17818
R22 adc_PISO_0.B4.n6 SARlogic_0.d3 1.54657
R23 adc_PISO_0.B4.n5 SARlogic_0.dffrs_7.nand3_1.A 1.34729
R24 adc_PISO_0.B4.n12 adc_PISO_0.B4.n11 0.732092
R25 adc_PISO_0.B4.n10 adc_PISO_0.B4.t2 0.7285
R26 adc_PISO_0.B4.n10 adc_PISO_0.B4.t3 0.7285
R27 SARlogic_0.dffrs_7.clk adc_PISO_0.B4.n5 0.610571
R28 SARlogic_0.dffrs_8.nand3_2.Z adc_PISO_0.B4.n9 0.166901
R29 adc_PISO_0.B4.n1 adc_PISO_0.B4.n0 0.106438
R30 adc_PISO_0.B4.n8 SARlogic_0.dffrs_8.nand3_7.C 0.0455
R31 adc_PISO_0.B4.n2 adc_PISO_0.2inmux_3.In 0.0455
R32 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t6 40.8177
R33 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t5 40.6313
R34 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t7 27.3166
R35 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t4 27.1302
R36 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_8.C.n2 14.119
R37 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.t1 10.0473
R38 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.t0 6.51042
R39 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.n4 6.04952
R40 SARlogic_0.dffrs_7.nand3_7.B SARlogic_0.dffrs_7.nand3_8.C.n0 5.47979
R41 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C.n1 5.13907
R42 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n6 4.72925
R43 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.n5 0.732092
R44 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t2 0.7285
R45 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t3 0.7285
R46 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_7.B 0.438233
R47 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n3 0.166901
R48 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C 0.0455
R49 Vdd.n1018 Vdd.t651 869.717
R50 Vdd.n1007 Vdd.t234 869.717
R51 Vdd.t230 Vdd.t462 490.324
R52 Vdd.t232 Vdd.t230 490.324
R53 Vdd.t685 Vdd.t232 490.324
R54 Vdd.t649 Vdd.t685 490.324
R55 Vdd.t314 Vdd.t649 490.324
R56 Vdd.t228 Vdd.t314 490.324
R57 Vdd.t713 Vdd.t228 490.324
R58 Vdd.t715 Vdd.t713 490.324
R59 Vdd.t24 Vdd.t715 490.324
R60 Vdd.t462 Vdd.n1054 467.743
R61 Vdd.n1056 Vdd.t24 467.743
R62 Vdd.n1057 Vdd.t735 398.652
R63 Vdd.n1039 Vdd.t719 398.652
R64 Vdd.t735 Vdd.n1056 389.878
R65 Vdd.n1054 Vdd.t719 389.878
R66 Vdd.t112 Vdd.n1011 372.543
R67 Vdd.n1014 Vdd.t66 372.543
R68 Vdd.n1013 Vdd.t112 370.969
R69 Vdd.t66 Vdd.n1013 370.969
R70 Vdd.n1034 Vdd.n1032 287.351
R71 Vdd.n1035 Vdd.n1033 287.351
R72 Vdd.t296 Vdd.t294 265.625
R73 Vdd.t190 Vdd.n4 250.9
R74 Vdd.n5 Vdd.t538 250.9
R75 Vdd.t404 Vdd.n1093 250.9
R76 Vdd.n1094 Vdd.t653 250.9
R77 Vdd.t268 Vdd.n9 250.9
R78 Vdd.n10 Vdd.t559 250.9
R79 Vdd.t286 Vdd.n1081 250.9
R80 Vdd.n1082 Vdd.t931 250.9
R81 Vdd.t532 Vdd.n1087 250.9
R82 Vdd.n1088 Vdd.t655 250.9
R83 Vdd.t96 Vdd.n1074 250.9
R84 Vdd.n1075 Vdd.t98 250.9
R85 Vdd.t280 Vdd.n51 250.9
R86 Vdd.n52 Vdd.t586 250.9
R87 Vdd.t611 Vdd.n62 250.9
R88 Vdd.n63 Vdd.t829 250.9
R89 Vdd.t320 Vdd.n57 250.9
R90 Vdd.n58 Vdd.t475 250.9
R91 Vdd.t835 Vdd.n74 250.9
R92 Vdd.n75 Vdd.t284 250.9
R93 Vdd.t514 Vdd.n68 250.9
R94 Vdd.n69 Vdd.t448 250.9
R95 Vdd.t426 Vdd.n85 250.9
R96 Vdd.n86 Vdd.t410 250.9
R97 Vdd.t236 Vdd.n124 250.9
R98 Vdd.n125 Vdd.t565 250.9
R99 Vdd.t641 Vdd.n135 250.9
R100 Vdd.n136 Vdd.t216 250.9
R101 Vdd.t937 Vdd.n130 250.9
R102 Vdd.n131 Vdd.t577 250.9
R103 Vdd.t889 Vdd.n147 250.9
R104 Vdd.n148 Vdd.t240 250.9
R105 Vdd.t601 Vdd.n141 250.9
R106 Vdd.n142 Vdd.t919 250.9
R107 Vdd.t12 Vdd.n158 250.9
R108 Vdd.n159 Vdd.t28 250.9
R109 Vdd.t460 Vdd.n204 250.9
R110 Vdd.n205 Vdd.t496 250.9
R111 Vdd.t517 Vdd.n209 250.9
R112 Vdd.n210 Vdd.t32 250.9
R113 Vdd.t865 Vdd.n198 250.9
R114 Vdd.n199 Vdd.t102 250.9
R115 Vdd.t769 Vdd.n999 250.9
R116 Vdd.n1000 Vdd.t46 250.9
R117 Vdd.t158 Vdd.n982 250.9
R118 Vdd.n983 Vdd.t36 250.9
R119 Vdd.t20 Vdd.n987 250.9
R120 Vdd.n988 Vdd.t867 250.9
R121 Vdd.t743 Vdd.n993 250.9
R122 Vdd.n994 Vdd.t793 250.9
R123 Vdd.t761 Vdd.n975 250.9
R124 Vdd.n976 Vdd.t883 250.9
R125 Vdd.t851 Vdd.n503 250.9
R126 Vdd.n504 Vdd.t481 250.9
R127 Vdd.t635 Vdd.n509 250.9
R128 Vdd.n510 Vdd.t266 250.9
R129 Vdd.t935 Vdd.n515 250.9
R130 Vdd.n516 Vdd.t879 250.9
R131 Vdd.t450 Vdd.n966 250.9
R132 Vdd.n967 Vdd.t813 250.9
R133 Vdd.t775 Vdd.n752 250.9
R134 Vdd.n753 Vdd.t368 250.9
R135 Vdd.t56 Vdd.n791 250.9
R136 Vdd.n792 Vdd.t264 250.9
R137 Vdd.t218 Vdd.n829 250.9
R138 Vdd.n830 Vdd.t272 250.9
R139 Vdd.t901 Vdd.n867 250.9
R140 Vdd.n868 Vdd.t747 250.9
R141 Vdd.t370 Vdd.n906 250.9
R142 Vdd.n907 Vdd.t212 250.9
R143 Vdd.t202 Vdd.n944 250.9
R144 Vdd.n945 Vdd.t911 250.9
R145 Vdd.t458 Vdd.n670 250.9
R146 Vdd.n671 Vdd.t394 250.9
R147 Vdd.t278 Vdd.n763 250.9
R148 Vdd.n764 Vdd.t186 250.9
R149 Vdd.t84 Vdd.n398 250.9
R150 Vdd.n399 Vdd.t124 250.9
R151 Vdd.t887 Vdd.n802 250.9
R152 Vdd.n803 Vdd.t42 250.9
R153 Vdd.t925 Vdd.n368 250.9
R154 Vdd.n369 Vdd.t50 250.9
R155 Vdd.t76 Vdd.n840 250.9
R156 Vdd.n841 Vdd.t270 250.9
R157 Vdd.t683 Vdd.n338 250.9
R158 Vdd.n339 Vdd.t366 250.9
R159 Vdd.t128 Vdd.n879 250.9
R160 Vdd.n880 Vdd.t745 250.9
R161 Vdd.t795 Vdd.n302 250.9
R162 Vdd.n303 Vdd.t290 250.9
R163 Vdd.t434 Vdd.n917 250.9
R164 Vdd.n918 Vdd.t210 250.9
R165 Vdd.t791 Vdd.n272 250.9
R166 Vdd.n273 Vdd.t312 250.9
R167 Vdd.t168 Vdd.n955 250.9
R168 Vdd.n956 Vdd.t176 250.9
R169 Vdd.t781 Vdd.n747 250.9
R170 Vdd.n748 Vdd.t777 250.9
R171 Vdd.t669 Vdd.n660 250.9
R172 Vdd.n661 Vdd.t929 250.9
R173 Vdd.t72 Vdd.n786 250.9
R174 Vdd.n787 Vdd.t148 250.9
R175 Vdd.t356 Vdd.n388 250.9
R176 Vdd.n389 Vdd.t174 250.9
R177 Vdd.t4 Vdd.n824 250.9
R178 Vdd.n825 Vdd.t242 250.9
R179 Vdd.t853 Vdd.n358 250.9
R180 Vdd.n359 Vdd.t86 250.9
R181 Vdd.t607 Vdd.n862 250.9
R182 Vdd.n863 Vdd.t899 250.9
R183 Vdd.t358 Vdd.n322 250.9
R184 Vdd.n323 Vdd.t923 250.9
R185 Vdd.t252 Vdd.n901 250.9
R186 Vdd.n902 Vdd.t200 250.9
R187 Vdd.t739 Vdd.n292 250.9
R188 Vdd.n293 Vdd.t681 250.9
R189 Vdd.t172 Vdd.n939 250.9
R190 Vdd.n940 Vdd.t372 250.9
R191 Vdd.t344 Vdd.n262 250.9
R192 Vdd.n263 Vdd.t797 250.9
R193 Vdd.t326 Vdd.n675 250.9
R194 Vdd.n676 Vdd.t787 250.9
R195 Vdd.t382 Vdd.n403 250.9
R196 Vdd.n404 Vdd.t907 250.9
R197 Vdd.t276 Vdd.n373 250.9
R198 Vdd.n374 Vdd.t322 250.9
R199 Vdd.t378 Vdd.n343 250.9
R200 Vdd.n344 Vdd.t258 250.9
R201 Vdd.t274 Vdd.n307 250.9
R202 Vdd.n308 Vdd.t849 250.9
R203 Vdd.t376 Vdd.n277 250.9
R204 Vdd.n278 Vdd.t226 250.9
R205 Vdd.t420 Vdd.n742 250.9
R206 Vdd.n743 Vdd.t571 250.9
R207 Vdd.t725 Vdd.n680 250.9
R208 Vdd.n681 Vdd.t318 250.9
R209 Vdd.t843 Vdd.n781 250.9
R210 Vdd.n782 Vdd.t478 250.9
R211 Vdd.t44 Vdd.n758 250.9
R212 Vdd.n759 Vdd.t562 250.9
R213 Vdd.t723 Vdd.n408 250.9
R214 Vdd.n409 Vdd.t0 250.9
R215 Vdd.t388 Vdd.n819 250.9
R216 Vdd.n820 Vdd.t526 250.9
R217 Vdd.t48 Vdd.n797 250.9
R218 Vdd.n798 Vdd.t520 250.9
R219 Vdd.t697 Vdd.n378 250.9
R220 Vdd.n379 Vdd.t913 250.9
R221 Vdd.t831 Vdd.n857 250.9
R222 Vdd.n858 Vdd.t574 250.9
R223 Vdd.t811 Vdd.n835 250.9
R224 Vdd.n836 Vdd.t544 250.9
R225 Vdd.t701 Vdd.n348 250.9
R226 Vdd.n349 Vdd.t40 250.9
R227 Vdd.t424 Vdd.n896 250.9
R228 Vdd.n897 Vdd.t535 250.9
R229 Vdd.t214 Vdd.n874 250.9
R230 Vdd.n875 Vdd.t592 250.9
R231 Vdd.t733 Vdd.n312 250.9
R232 Vdd.n313 Vdd.t871 250.9
R233 Vdd.t166 Vdd.n934 250.9
R234 Vdd.n935 Vdd.t580 250.9
R235 Vdd.t909 Vdd.n912 250.9
R236 Vdd.n913 Vdd.t541 250.9
R237 Vdd.t689 Vdd.n282 250.9
R238 Vdd.n283 Vdd.t188 250.9
R239 Vdd.t38 Vdd.n950 250.9
R240 Vdd.n951 Vdd.t556 250.9
R241 Vdd.t891 Vdd.n737 250.9
R242 Vdd.n738 Vdd.t418 250.9
R243 Vdd.t362 Vdd.n665 250.9
R244 Vdd.n666 Vdd.t412 250.9
R245 Vdd.t619 Vdd.n776 250.9
R246 Vdd.n777 Vdd.t841 250.9
R247 Vdd.t861 Vdd.n393 250.9
R248 Vdd.n394 Vdd.t428 250.9
R249 Vdd.t452 Vdd.n814 250.9
R250 Vdd.n815 Vdd.t384 250.9
R251 Vdd.t346 Vdd.n363 250.9
R252 Vdd.n364 Vdd.t821 250.9
R253 Vdd.t62 Vdd.n852 250.9
R254 Vdd.n853 Vdd.t693 250.9
R255 Vdd.t334 Vdd.n327 250.9
R256 Vdd.n328 Vdd.t877 250.9
R257 Vdd.t400 Vdd.n891 250.9
R258 Vdd.n892 Vdd.t422 250.9
R259 Vdd.t342 Vdd.n297 250.9
R260 Vdd.n298 Vdd.t432 250.9
R261 Vdd.t34 Vdd.n929 250.9
R262 Vdd.n930 Vdd.t254 250.9
R263 Vdd.t857 Vdd.n267 250.9
R264 Vdd.n268 Vdd.t18 250.9
R265 Vdd.t180 Vdd.n685 250.9
R266 Vdd.n686 Vdd.t246 250.9
R267 Vdd.t464 Vdd.n413 250.9
R268 Vdd.n414 Vdd.t146 250.9
R269 Vdd.t454 Vdd.n383 250.9
R270 Vdd.n384 Vdd.t222 250.9
R271 Vdd.t398 Vdd.n353 250.9
R272 Vdd.n354 Vdd.t160 250.9
R273 Vdd.t875 Vdd.n317 250.9
R274 Vdd.n318 Vdd.t637 250.9
R275 Vdd.t438 Vdd.n287 250.9
R276 Vdd.n288 Vdd.t60 250.9
R277 Vdd.t629 Vdd.n690 250.9
R278 Vdd.n691 Vdd.t340 250.9
R279 Vdd.t721 Vdd.n706 250.9
R280 Vdd.n707 Vdd.t615 250.9
R281 Vdd.t184 Vdd.n701 250.9
R282 Vdd.n702 Vdd.t338 250.9
R283 Vdd.t136 Vdd.n724 250.9
R284 Vdd.n725 Vdd.t627 250.9
R285 Vdd.t589 Vdd.n730 250.9
R286 Vdd.n731 Vdd.t178 250.9
R287 Vdd.t767 Vdd.n718 250.9
R288 Vdd.n719 Vdd.t364 250.9
R289 Vdd.t182 Vdd.n623 250.9
R290 Vdd.n624 Vdd.t484 250.9
R291 Vdd.t609 Vdd.n634 250.9
R292 Vdd.n635 Vdd.t414 250.9
R293 Vdd.t80 Vdd.n629 250.9
R294 Vdd.n630 Vdd.t523 250.9
R295 Vdd.t623 Vdd.n646 250.9
R296 Vdd.n647 Vdd.t328 250.9
R297 Vdd.t598 Vdd.n640 250.9
R298 Vdd.n641 Vdd.t941 250.9
R299 Vdd.t613 Vdd.n653 250.9
R300 Vdd.n654 Vdd.t873 250.9
R301 Vdd.t306 Vdd.n554 250.9
R302 Vdd.n555 Vdd.t469 250.9
R303 Vdd.t446 Vdd.n565 250.9
R304 Vdd.n566 Vdd.t915 250.9
R305 Vdd.t14 Vdd.n560 250.9
R306 Vdd.n561 Vdd.t490 250.9
R307 Vdd.t823 Vdd.n577 250.9
R308 Vdd.n578 Vdd.t310 250.9
R309 Vdd.t499 Vdd.n571 250.9
R310 Vdd.n572 Vdd.t106 250.9
R311 Vdd.t8 Vdd.n584 250.9
R312 Vdd.n585 Vdd.t440 250.9
R313 Vdd.n1025 Vdd.t114 242.189
R314 Vdd.n186 Vdd.t90 236.083
R315 Vdd.t118 Vdd.n183 236.083
R316 Vdd.t749 Vdd.n166 236.083
R317 Vdd.n172 Vdd.t771 236.083
R318 Vdd.n113 Vdd.t164 236.083
R319 Vdd.t837 Vdd.n110 236.083
R320 Vdd.t603 Vdd.n93 236.083
R321 Vdd.n99 Vdd.t799 236.083
R322 Vdd.n45 Vdd.t939 236.083
R323 Vdd.n39 Vdd.t707 236.083
R324 Vdd.n29 Vdd.t204 236.083
R325 Vdd.n23 Vdd.t142 236.083
R326 Vdd.t436 Vdd.n231 236.083
R327 Vdd.n237 Vdd.t927 236.083
R328 Vdd.n612 Vdd.t380 236.083
R329 Vdd.t134 Vdd.n609 236.083
R330 Vdd.t316 Vdd.n592 236.083
R331 Vdd.n598 Vdd.t456 236.083
R332 Vdd.n543 Vdd.t92 236.083
R333 Vdd.t116 Vdd.n540 236.083
R334 Vdd.t895 Vdd.n523 236.083
R335 Vdd.n529 Vdd.t82 236.083
R336 Vdd.n497 Vdd.t430 236.083
R337 Vdd.n491 Vdd.t817 236.083
R338 Vdd.n481 Vdd.t705 236.083
R339 Vdd.n475 Vdd.t304 236.083
R340 Vdd.t74 Vdd.n451 236.083
R341 Vdd.n457 Vdd.t827 236.083
R342 Vdd.t224 Vdd.n435 236.083
R343 Vdd.n443 Vdd.t759 236.083
R344 Vdd.t402 Vdd.n422 236.083
R345 Vdd.n433 Vdd.t54 236.083
R346 Vdd.t466 Vdd.n247 236.083
R347 Vdd.n251 Vdd.t753 236.083
R348 Vdd.t244 Vdd.n221 236.083
R349 Vdd.n223 Vdd.t154 236.083
R350 Vdd.t90 Vdd.n185 235.294
R351 Vdd.n185 Vdd.t118 235.294
R352 Vdd.n171 Vdd.t749 235.294
R353 Vdd.t771 Vdd.n171 235.294
R354 Vdd.t164 Vdd.n112 235.294
R355 Vdd.n112 Vdd.t837 235.294
R356 Vdd.n98 Vdd.t603 235.294
R357 Vdd.t799 Vdd.n98 235.294
R358 Vdd.t939 Vdd.n44 235.294
R359 Vdd.n44 Vdd.t261 235.294
R360 Vdd.t260 Vdd.n42 235.294
R361 Vdd.n42 Vdd.t709 235.294
R362 Vdd.t204 Vdd.n28 235.294
R363 Vdd.n28 Vdd.t11 235.294
R364 Vdd.t10 Vdd.n26 235.294
R365 Vdd.n26 Vdd.t140 235.294
R366 Vdd.n236 Vdd.t436 235.294
R367 Vdd.t927 Vdd.n236 235.294
R368 Vdd.t380 Vdd.n611 235.294
R369 Vdd.n611 Vdd.t134 235.294
R370 Vdd.n597 Vdd.t316 235.294
R371 Vdd.t456 Vdd.n597 235.294
R372 Vdd.t92 Vdd.n542 235.294
R373 Vdd.n542 Vdd.t116 235.294
R374 Vdd.n528 Vdd.t895 235.294
R375 Vdd.t82 Vdd.n528 235.294
R376 Vdd.t430 Vdd.n496 235.294
R377 Vdd.n496 Vdd.t152 235.294
R378 Vdd.t153 Vdd.n494 235.294
R379 Vdd.n494 Vdd.t819 235.294
R380 Vdd.t705 Vdd.n480 235.294
R381 Vdd.n480 Vdd.t109 235.294
R382 Vdd.t108 Vdd.n478 235.294
R383 Vdd.n478 Vdd.t302 235.294
R384 Vdd.n456 Vdd.t74 235.294
R385 Vdd.t827 Vdd.n456 235.294
R386 Vdd.n442 Vdd.t224 235.294
R387 Vdd.t759 Vdd.n442 235.294
R388 Vdd.n430 Vdd.t402 235.294
R389 Vdd.t123 Vdd.n430 235.294
R390 Vdd.n432 Vdd.t122 235.294
R391 Vdd.t52 Vdd.n432 235.294
R392 Vdd.n250 Vdd.t466 235.294
R393 Vdd.t753 Vdd.n250 235.294
R394 Vdd.n227 Vdd.t244 235.294
R395 Vdd.n227 Vdd.t288 235.294
R396 Vdd.t289 Vdd.n226 235.294
R397 Vdd.n226 Vdd.t156 235.294
R398 Vdd.t933 Vdd.t190 200
R399 Vdd.t538 Vdd.t933 200
R400 Vdd.t529 Vdd.t404 200
R401 Vdd.t653 Vdd.t529 200
R402 Vdd.t192 Vdd.t268 200
R403 Vdd.t559 Vdd.t192 200
R404 Vdd.t643 Vdd.t286 200
R405 Vdd.t931 Vdd.t643 200
R406 Vdd.t100 Vdd.t532 200
R407 Vdd.t655 Vdd.t100 200
R408 Vdd.t568 Vdd.t96 200
R409 Vdd.t98 Vdd.t568 200
R410 Vdd.t845 Vdd.t280 200
R411 Vdd.t586 Vdd.t845 200
R412 Vdd.t472 Vdd.t611 200
R413 Vdd.t829 Vdd.t472 200
R414 Vdd.t282 Vdd.t320 200
R415 Vdd.t475 Vdd.t282 200
R416 Vdd.t647 Vdd.t835 200
R417 Vdd.t284 Vdd.t647 200
R418 Vdd.t408 Vdd.t514 200
R419 Vdd.t448 Vdd.t408 200
R420 Vdd.t508 Vdd.t426 200
R421 Vdd.t410 Vdd.t508 200
R422 Vdd.t261 Vdd.t260 200
R423 Vdd.t707 Vdd.t709 200
R424 Vdd.t885 Vdd.t236 200
R425 Vdd.t565 Vdd.t885 200
R426 Vdd.t595 Vdd.t641 200
R427 Vdd.t216 Vdd.t595 200
R428 Vdd.t238 Vdd.t937 200
R429 Vdd.t577 Vdd.t238 200
R430 Vdd.t444 Vdd.t889 200
R431 Vdd.t240 Vdd.t444 200
R432 Vdd.t262 Vdd.t601 200
R433 Vdd.t919 Vdd.t262 200
R434 Vdd.t493 Vdd.t12 200
R435 Vdd.t28 Vdd.t493 200
R436 Vdd.t11 Vdd.t10 200
R437 Vdd.t142 Vdd.t140 200
R438 Vdd.t881 Vdd.t460 200
R439 Vdd.t496 Vdd.t881 200
R440 Vdd.t815 Vdd.t517 200
R441 Vdd.t32 Vdd.t815 200
R442 Vdd.t22 Vdd.t865 200
R443 Vdd.t102 Vdd.t22 200
R444 Vdd.t805 Vdd.t769 200
R445 Vdd.t46 Vdd.t805 200
R446 Vdd.t869 Vdd.t158 200
R447 Vdd.t36 Vdd.t869 200
R448 Vdd.t765 Vdd.t20 200
R449 Vdd.t867 Vdd.t765 200
R450 Vdd.t94 Vdd.t743 200
R451 Vdd.t793 Vdd.t94 200
R452 Vdd.t809 Vdd.t761 200
R453 Vdd.t883 Vdd.t809 200
R454 Vdd.t104 Vdd.t851 200
R455 Vdd.t481 Vdd.t104 200
R456 Vdd.t511 Vdd.t635 200
R457 Vdd.t266 Vdd.t511 200
R458 Vdd.t406 Vdd.t935 200
R459 Vdd.t879 Vdd.t406 200
R460 Vdd.t553 Vdd.t450 200
R461 Vdd.t813 Vdd.t553 200
R462 Vdd.t783 Vdd.t775 200
R463 Vdd.t368 Vdd.t783 200
R464 Vdd.t70 Vdd.t56 200
R465 Vdd.t264 Vdd.t70 200
R466 Vdd.t6 Vdd.t218 200
R467 Vdd.t272 Vdd.t6 200
R468 Vdd.t605 Vdd.t901 200
R469 Vdd.t747 Vdd.t605 200
R470 Vdd.t250 Vdd.t370 200
R471 Vdd.t212 Vdd.t250 200
R472 Vdd.t170 Vdd.t202 200
R473 Vdd.t911 Vdd.t170 200
R474 Vdd.t392 Vdd.t458 200
R475 Vdd.t394 Vdd.t392 200
R476 Vdd.t773 Vdd.t278 200
R477 Vdd.t186 Vdd.t773 200
R478 Vdd.t673 Vdd.t84 200
R479 Vdd.t124 Vdd.t673 200
R480 Vdd.t150 Vdd.t887 200
R481 Vdd.t42 Vdd.t150 200
R482 Vdd.t807 Vdd.t925 200
R483 Vdd.t50 Vdd.t807 200
R484 Vdd.t220 Vdd.t76 200
R485 Vdd.t270 Vdd.t220 200
R486 Vdd.t348 Vdd.t683 200
R487 Vdd.t366 Vdd.t348 200
R488 Vdd.t903 Vdd.t128 200
R489 Vdd.t745 Vdd.t903 200
R490 Vdd.t665 Vdd.t795 200
R491 Vdd.t290 Vdd.t665 200
R492 Vdd.t198 Vdd.t434 200
R493 Vdd.t210 Vdd.t198 200
R494 Vdd.t332 Vdd.t791 200
R495 Vdd.t312 Vdd.t332 200
R496 Vdd.t374 Vdd.t168 200
R497 Vdd.t176 Vdd.t374 200
R498 Vdd.t126 Vdd.t781 200
R499 Vdd.t777 Vdd.t126 200
R500 Vdd.t785 Vdd.t669 200
R501 Vdd.t929 Vdd.t785 200
R502 Vdd.t88 Vdd.t72 200
R503 Vdd.t148 Vdd.t88 200
R504 Vdd.t905 Vdd.t356 200
R505 Vdd.t174 Vdd.t905 200
R506 Vdd.t921 Vdd.t4 200
R507 Vdd.t242 Vdd.t921 200
R508 Vdd.t324 Vdd.t853 200
R509 Vdd.t86 Vdd.t324 200
R510 Vdd.t679 Vdd.t607 200
R511 Vdd.t899 Vdd.t679 200
R512 Vdd.t208 Vdd.t358 200
R513 Vdd.t923 Vdd.t208 200
R514 Vdd.t390 Vdd.t252 200
R515 Vdd.t200 Vdd.t390 200
R516 Vdd.t847 Vdd.t739 200
R517 Vdd.t681 Vdd.t847 200
R518 Vdd.t789 Vdd.t172 200
R519 Vdd.t372 Vdd.t789 200
R520 Vdd.t779 Vdd.t344 200
R521 Vdd.t797 Vdd.t779 200
R522 Vdd.t859 Vdd.t326 200
R523 Vdd.t787 Vdd.t859 200
R524 Vdd.t741 Vdd.t382 200
R525 Vdd.t907 Vdd.t741 200
R526 Vdd.t677 Vdd.t276 200
R527 Vdd.t322 Vdd.t677 200
R528 Vdd.t354 Vdd.t378 200
R529 Vdd.t258 Vdd.t354 200
R530 Vdd.t863 Vdd.t274 200
R531 Vdd.t849 Vdd.t863 200
R532 Vdd.t661 Vdd.t376 200
R533 Vdd.t226 Vdd.t661 200
R534 Vdd.t893 Vdd.t420 200
R535 Vdd.t571 Vdd.t893 200
R536 Vdd.t675 Vdd.t725 200
R537 Vdd.t318 Vdd.t675 200
R538 Vdd.t396 Vdd.t843 200
R539 Vdd.t478 Vdd.t396 200
R540 Vdd.t206 Vdd.t44 200
R541 Vdd.t562 Vdd.t206 200
R542 Vdd.t352 Vdd.t723 200
R543 Vdd.t0 Vdd.t352 200
R544 Vdd.t633 Vdd.t388 200
R545 Vdd.t526 Vdd.t633 200
R546 Vdd.t839 Vdd.t48 200
R547 Vdd.t520 Vdd.t839 200
R548 Vdd.t360 Vdd.t697 200
R549 Vdd.t913 Vdd.t360 200
R550 Vdd.t64 Vdd.t831 200
R551 Vdd.t574 Vdd.t64 200
R552 Vdd.t386 Vdd.t811 200
R553 Vdd.t544 Vdd.t386 200
R554 Vdd.t663 Vdd.t701 200
R555 Vdd.t40 Vdd.t663 200
R556 Vdd.t711 Vdd.t424 200
R557 Vdd.t535 Vdd.t711 200
R558 Vdd.t833 Vdd.t214 200
R559 Vdd.t592 Vdd.t833 200
R560 Vdd.t667 Vdd.t733 200
R561 Vdd.t871 Vdd.t667 200
R562 Vdd.t2 Vdd.t166 200
R563 Vdd.t580 Vdd.t2 200
R564 Vdd.t617 Vdd.t909 200
R565 Vdd.t541 Vdd.t617 200
R566 Vdd.t803 Vdd.t689 200
R567 Vdd.t188 Vdd.t803 200
R568 Vdd.t256 Vdd.t38 200
R569 Vdd.t556 Vdd.t256 200
R570 Vdd.t729 Vdd.t891 200
R571 Vdd.t418 Vdd.t729 200
R572 Vdd.t248 Vdd.t362 200
R573 Vdd.t412 Vdd.t248 200
R574 Vdd.t717 Vdd.t619 200
R575 Vdd.t841 Vdd.t717 200
R576 Vdd.t144 Vdd.t861 200
R577 Vdd.t428 Vdd.t144 200
R578 Vdd.t699 Vdd.t452 200
R579 Vdd.t384 Vdd.t699 200
R580 Vdd.t196 Vdd.t346 200
R581 Vdd.t821 Vdd.t196 200
R582 Vdd.t691 Vdd.t62 200
R583 Vdd.t693 Vdd.t691 200
R584 Vdd.t162 Vdd.t334 200
R585 Vdd.t877 Vdd.t162 200
R586 Vdd.t727 Vdd.t400 200
R587 Vdd.t422 Vdd.t727 200
R588 Vdd.t639 Vdd.t342 200
R589 Vdd.t432 Vdd.t639 200
R590 Vdd.t703 Vdd.t34 200
R591 Vdd.t254 Vdd.t703 200
R592 Vdd.t58 Vdd.t857 200
R593 Vdd.t18 Vdd.t58 200
R594 Vdd.t671 Vdd.t180 200
R595 Vdd.t246 Vdd.t671 200
R596 Vdd.t350 Vdd.t464 200
R597 Vdd.t146 Vdd.t350 200
R598 Vdd.t659 Vdd.t454 200
R599 Vdd.t222 Vdd.t659 200
R600 Vdd.t855 Vdd.t398 200
R601 Vdd.t160 Vdd.t855 200
R602 Vdd.t737 Vdd.t875 200
R603 Vdd.t637 Vdd.t737 200
R604 Vdd.t336 Vdd.t438 200
R605 Vdd.t60 Vdd.t336 200
R606 Vdd.t138 Vdd.t629 200
R607 Vdd.t340 Vdd.t138 200
R608 Vdd.t487 Vdd.t721 200
R609 Vdd.t615 Vdd.t487 200
R610 Vdd.t621 Vdd.t184 200
R611 Vdd.t338 Vdd.t621 200
R612 Vdd.t687 Vdd.t136 200
R613 Vdd.t627 Vdd.t687 200
R614 Vdd.t631 Vdd.t589 200
R615 Vdd.t178 Vdd.t631 200
R616 Vdd.t583 Vdd.t767 200
R617 Vdd.t364 Vdd.t583 200
R618 Vdd.t625 Vdd.t182 200
R619 Vdd.t484 Vdd.t625 200
R620 Vdd.t502 Vdd.t609 200
R621 Vdd.t414 Vdd.t502 200
R622 Vdd.t330 Vdd.t80 200
R623 Vdd.t523 Vdd.t330 200
R624 Vdd.t416 Vdd.t623 200
R625 Vdd.t328 Vdd.t416 200
R626 Vdd.t292 Vdd.t598 200
R627 Vdd.t941 Vdd.t292 200
R628 Vdd.t547 Vdd.t613 200
R629 Vdd.t873 Vdd.t547 200
R630 Vdd.t825 Vdd.t306 200
R631 Vdd.t469 Vdd.t825 200
R632 Vdd.t505 Vdd.t446 200
R633 Vdd.t915 Vdd.t505 200
R634 Vdd.t308 Vdd.t14 200
R635 Vdd.t490 Vdd.t308 200
R636 Vdd.t645 Vdd.t823 200
R637 Vdd.t310 Vdd.t645 200
R638 Vdd.t442 Vdd.t499 200
R639 Vdd.t106 Vdd.t442 200
R640 Vdd.t550 Vdd.t8 200
R641 Vdd.t440 Vdd.t550 200
R642 Vdd.t152 Vdd.t153 200
R643 Vdd.t817 Vdd.t819 200
R644 Vdd.t109 Vdd.t108 200
R645 Vdd.t304 Vdd.t302 200
R646 Vdd.t122 Vdd.t123 200
R647 Vdd.t54 Vdd.t52 200
R648 Vdd.t288 Vdd.t289 200
R649 Vdd.t154 Vdd.t156 200
R650 Vdd.t300 Vdd.n1027 195.312
R651 Vdd.n1061 Vdd.t695 190.464
R652 Vdd.n1037 Vdd.t731 190.464
R653 Vdd.n1028 Vdd.t300 179.689
R654 Vdd.t114 Vdd.n1024 145.413
R655 Vdd.n15 Vdd.t657 131.589
R656 Vdd.n174 Vdd.t801 131.589
R657 Vdd.n31 Vdd.t917 131.589
R658 Vdd.n101 Vdd.t68 131.589
R659 Vdd.n239 Vdd.t78 131.589
R660 Vdd.n253 Vdd.t30 131.589
R661 Vdd.n467 Vdd.t26 131.589
R662 Vdd.n600 Vdd.t16 131.589
R663 Vdd.n483 Vdd.t897 131.589
R664 Vdd.n531 Vdd.t194 131.589
R665 Vdd.n459 Vdd.t110 131.589
R666 Vdd.n445 Vdd.t763 131.589
R667 Vdd.n1004 Vdd.n259 130.231
R668 Vdd.n1004 Vdd.n980 121.085
R669 Vdd.n117 Vdd.t132 118.543
R670 Vdd.n190 Vdd.t757 118.543
R671 Vdd.n547 Vdd.t120 118.543
R672 Vdd.n616 Vdd.t755 118.543
R673 Vdd.n437 Vdd.t751 118.543
R674 Vdd.n255 Vdd.t130 118.543
R675 Vdd.n259 Vdd.n258 117.481
R676 Vdd.n39 Vdd.n38 96.0755
R677 Vdd.n40 Vdd.n39 96.0755
R678 Vdd.n23 Vdd.n22 96.0755
R679 Vdd.n24 Vdd.n23 96.0755
R680 Vdd.n491 Vdd.n490 96.0755
R681 Vdd.n492 Vdd.n491 96.0755
R682 Vdd.n475 Vdd.n474 96.0755
R683 Vdd.n476 Vdd.n475 96.0755
R684 Vdd.n433 Vdd.n425 96.0755
R685 Vdd.n433 Vdd.n426 96.0755
R686 Vdd.n223 Vdd.n222 96.0755
R687 Vdd.n224 Vdd.n223 96.0755
R688 Vdd.n1028 Vdd.t296 85.938
R689 Vdd.n168 Vdd.n166 78.2255
R690 Vdd.n172 Vdd.n168 78.2255
R691 Vdd.n172 Vdd.n169 78.2255
R692 Vdd.n169 Vdd.n166 78.2255
R693 Vdd.n95 Vdd.n93 78.2255
R694 Vdd.n99 Vdd.n95 78.2255
R695 Vdd.n99 Vdd.n96 78.2255
R696 Vdd.n96 Vdd.n93 78.2255
R697 Vdd.n45 Vdd.n36 78.2255
R698 Vdd.n45 Vdd.n37 78.2255
R699 Vdd.n113 Vdd.n108 78.2255
R700 Vdd.n113 Vdd.n109 78.2255
R701 Vdd.n110 Vdd.n108 78.2255
R702 Vdd.n110 Vdd.n109 78.2255
R703 Vdd.n29 Vdd.n20 78.2255
R704 Vdd.n29 Vdd.n21 78.2255
R705 Vdd.n186 Vdd.n181 78.2255
R706 Vdd.n186 Vdd.n182 78.2255
R707 Vdd.n183 Vdd.n181 78.2255
R708 Vdd.n183 Vdd.n182 78.2255
R709 Vdd.n233 Vdd.n231 78.2255
R710 Vdd.n237 Vdd.n233 78.2255
R711 Vdd.n237 Vdd.n234 78.2255
R712 Vdd.n234 Vdd.n231 78.2255
R713 Vdd.n594 Vdd.n592 78.2255
R714 Vdd.n598 Vdd.n594 78.2255
R715 Vdd.n598 Vdd.n595 78.2255
R716 Vdd.n595 Vdd.n592 78.2255
R717 Vdd.n525 Vdd.n523 78.2255
R718 Vdd.n529 Vdd.n525 78.2255
R719 Vdd.n529 Vdd.n526 78.2255
R720 Vdd.n526 Vdd.n523 78.2255
R721 Vdd.n497 Vdd.n488 78.2255
R722 Vdd.n497 Vdd.n489 78.2255
R723 Vdd.n543 Vdd.n538 78.2255
R724 Vdd.n543 Vdd.n539 78.2255
R725 Vdd.n540 Vdd.n538 78.2255
R726 Vdd.n540 Vdd.n539 78.2255
R727 Vdd.n481 Vdd.n472 78.2255
R728 Vdd.n481 Vdd.n473 78.2255
R729 Vdd.n612 Vdd.n607 78.2255
R730 Vdd.n612 Vdd.n608 78.2255
R731 Vdd.n609 Vdd.n607 78.2255
R732 Vdd.n609 Vdd.n608 78.2255
R733 Vdd.n453 Vdd.n451 78.2255
R734 Vdd.n457 Vdd.n453 78.2255
R735 Vdd.n457 Vdd.n454 78.2255
R736 Vdd.n454 Vdd.n451 78.2255
R737 Vdd.n439 Vdd.n435 78.2255
R738 Vdd.n443 Vdd.n439 78.2255
R739 Vdd.n443 Vdd.n440 78.2255
R740 Vdd.n440 Vdd.n435 78.2255
R741 Vdd.n427 Vdd.n422 78.2255
R742 Vdd.n428 Vdd.n422 78.2255
R743 Vdd.n247 Vdd.n215 78.2255
R744 Vdd.n251 Vdd.n215 78.2255
R745 Vdd.n251 Vdd.n216 78.2255
R746 Vdd.n247 Vdd.n216 78.2255
R747 Vdd.n221 Vdd.n219 78.2255
R748 Vdd.n221 Vdd.n220 78.2255
R749 Vdd.n1027 Vdd.t298 70.313
R750 Vdd.n5 Vdd.n4 68.0765
R751 Vdd.n1094 Vdd.n1093 68.0765
R752 Vdd.n10 Vdd.n9 68.0765
R753 Vdd.n1082 Vdd.n1081 68.0765
R754 Vdd.n1088 Vdd.n1087 68.0765
R755 Vdd.n1075 Vdd.n1074 68.0765
R756 Vdd.n52 Vdd.n51 68.0765
R757 Vdd.n63 Vdd.n62 68.0765
R758 Vdd.n58 Vdd.n57 68.0765
R759 Vdd.n75 Vdd.n74 68.0765
R760 Vdd.n69 Vdd.n68 68.0765
R761 Vdd.n86 Vdd.n85 68.0765
R762 Vdd.n125 Vdd.n124 68.0765
R763 Vdd.n136 Vdd.n135 68.0765
R764 Vdd.n131 Vdd.n130 68.0765
R765 Vdd.n148 Vdd.n147 68.0765
R766 Vdd.n142 Vdd.n141 68.0765
R767 Vdd.n159 Vdd.n158 68.0765
R768 Vdd.n205 Vdd.n204 68.0765
R769 Vdd.n210 Vdd.n209 68.0765
R770 Vdd.n199 Vdd.n198 68.0765
R771 Vdd.n1000 Vdd.n999 68.0765
R772 Vdd.n983 Vdd.n982 68.0765
R773 Vdd.n988 Vdd.n987 68.0765
R774 Vdd.n994 Vdd.n993 68.0765
R775 Vdd.n976 Vdd.n975 68.0765
R776 Vdd.n504 Vdd.n503 68.0765
R777 Vdd.n510 Vdd.n509 68.0765
R778 Vdd.n516 Vdd.n515 68.0765
R779 Vdd.n967 Vdd.n966 68.0765
R780 Vdd.n753 Vdd.n752 68.0765
R781 Vdd.n792 Vdd.n791 68.0765
R782 Vdd.n830 Vdd.n829 68.0765
R783 Vdd.n868 Vdd.n867 68.0765
R784 Vdd.n907 Vdd.n906 68.0765
R785 Vdd.n945 Vdd.n944 68.0765
R786 Vdd.n671 Vdd.n670 68.0765
R787 Vdd.n764 Vdd.n763 68.0765
R788 Vdd.n399 Vdd.n398 68.0765
R789 Vdd.n803 Vdd.n802 68.0765
R790 Vdd.n369 Vdd.n368 68.0765
R791 Vdd.n841 Vdd.n840 68.0765
R792 Vdd.n339 Vdd.n338 68.0765
R793 Vdd.n880 Vdd.n879 68.0765
R794 Vdd.n303 Vdd.n302 68.0765
R795 Vdd.n918 Vdd.n917 68.0765
R796 Vdd.n273 Vdd.n272 68.0765
R797 Vdd.n956 Vdd.n955 68.0765
R798 Vdd.n748 Vdd.n747 68.0765
R799 Vdd.n661 Vdd.n660 68.0765
R800 Vdd.n787 Vdd.n786 68.0765
R801 Vdd.n389 Vdd.n388 68.0765
R802 Vdd.n825 Vdd.n824 68.0765
R803 Vdd.n359 Vdd.n358 68.0765
R804 Vdd.n863 Vdd.n862 68.0765
R805 Vdd.n323 Vdd.n322 68.0765
R806 Vdd.n902 Vdd.n901 68.0765
R807 Vdd.n293 Vdd.n292 68.0765
R808 Vdd.n940 Vdd.n939 68.0765
R809 Vdd.n263 Vdd.n262 68.0765
R810 Vdd.n676 Vdd.n675 68.0765
R811 Vdd.n404 Vdd.n403 68.0765
R812 Vdd.n374 Vdd.n373 68.0765
R813 Vdd.n344 Vdd.n343 68.0765
R814 Vdd.n308 Vdd.n307 68.0765
R815 Vdd.n278 Vdd.n277 68.0765
R816 Vdd.n743 Vdd.n742 68.0765
R817 Vdd.n681 Vdd.n680 68.0765
R818 Vdd.n782 Vdd.n781 68.0765
R819 Vdd.n759 Vdd.n758 68.0765
R820 Vdd.n409 Vdd.n408 68.0765
R821 Vdd.n820 Vdd.n819 68.0765
R822 Vdd.n798 Vdd.n797 68.0765
R823 Vdd.n379 Vdd.n378 68.0765
R824 Vdd.n858 Vdd.n857 68.0765
R825 Vdd.n836 Vdd.n835 68.0765
R826 Vdd.n349 Vdd.n348 68.0765
R827 Vdd.n897 Vdd.n896 68.0765
R828 Vdd.n875 Vdd.n874 68.0765
R829 Vdd.n313 Vdd.n312 68.0765
R830 Vdd.n935 Vdd.n934 68.0765
R831 Vdd.n913 Vdd.n912 68.0765
R832 Vdd.n283 Vdd.n282 68.0765
R833 Vdd.n951 Vdd.n950 68.0765
R834 Vdd.n738 Vdd.n737 68.0765
R835 Vdd.n666 Vdd.n665 68.0765
R836 Vdd.n777 Vdd.n776 68.0765
R837 Vdd.n394 Vdd.n393 68.0765
R838 Vdd.n815 Vdd.n814 68.0765
R839 Vdd.n364 Vdd.n363 68.0765
R840 Vdd.n853 Vdd.n852 68.0765
R841 Vdd.n328 Vdd.n327 68.0765
R842 Vdd.n892 Vdd.n891 68.0765
R843 Vdd.n298 Vdd.n297 68.0765
R844 Vdd.n930 Vdd.n929 68.0765
R845 Vdd.n268 Vdd.n267 68.0765
R846 Vdd.n686 Vdd.n685 68.0765
R847 Vdd.n414 Vdd.n413 68.0765
R848 Vdd.n384 Vdd.n383 68.0765
R849 Vdd.n354 Vdd.n353 68.0765
R850 Vdd.n318 Vdd.n317 68.0765
R851 Vdd.n288 Vdd.n287 68.0765
R852 Vdd.n691 Vdd.n690 68.0765
R853 Vdd.n707 Vdd.n706 68.0765
R854 Vdd.n702 Vdd.n701 68.0765
R855 Vdd.n725 Vdd.n724 68.0765
R856 Vdd.n731 Vdd.n730 68.0765
R857 Vdd.n719 Vdd.n718 68.0765
R858 Vdd.n624 Vdd.n623 68.0765
R859 Vdd.n635 Vdd.n634 68.0765
R860 Vdd.n630 Vdd.n629 68.0765
R861 Vdd.n647 Vdd.n646 68.0765
R862 Vdd.n641 Vdd.n640 68.0765
R863 Vdd.n654 Vdd.n653 68.0765
R864 Vdd.n555 Vdd.n554 68.0765
R865 Vdd.n566 Vdd.n565 68.0765
R866 Vdd.n561 Vdd.n560 68.0765
R867 Vdd.n578 Vdd.n577 68.0765
R868 Vdd.n572 Vdd.n571 68.0765
R869 Vdd.n585 Vdd.n584 68.0765
R870 Vdd.n38 Vdd.n36 59.8505
R871 Vdd.n40 Vdd.n37 59.8505
R872 Vdd.n22 Vdd.n20 59.8505
R873 Vdd.n24 Vdd.n21 59.8505
R874 Vdd.n490 Vdd.n488 59.8505
R875 Vdd.n492 Vdd.n489 59.8505
R876 Vdd.n474 Vdd.n472 59.8505
R877 Vdd.n476 Vdd.n473 59.8505
R878 Vdd.n427 Vdd.n425 59.8505
R879 Vdd.n428 Vdd.n426 59.8505
R880 Vdd.n222 Vdd.n219 59.8505
R881 Vdd.n224 Vdd.n220 59.8505
R882 Vdd.n1011 Vdd.n1009 58.9755
R883 Vdd.n1014 Vdd.n1009 58.9755
R884 Vdd.n1014 Vdd.n1010 58.9755
R885 Vdd.n1011 Vdd.n1010 58.9755
R886 Vdd.n1057 Vdd.n1032 54.0755
R887 Vdd.n1039 Vdd.n1034 54.0755
R888 Vdd.n1039 Vdd.n1035 54.0755
R889 Vdd.n1057 Vdd.n1033 54.0755
R890 Vdd.n192 Vdd.t531 41.0041
R891 Vdd.n79 Vdd.t513 41.0041
R892 Vdd.n152 Vdd.t600 41.0041
R893 Vdd.n960 Vdd.t516 41.0041
R894 Vdd.n711 Vdd.t588 41.0041
R895 Vdd.n417 Vdd.t597 41.0041
R896 Vdd.n331 Vdd.t498 41.0041
R897 Vdd.n194 Vdd.t567 40.8177
R898 Vdd.n193 Vdd.t528 40.8177
R899 Vdd.n81 Vdd.t507 40.8177
R900 Vdd.n80 Vdd.t471 40.8177
R901 Vdd.n154 Vdd.t492 40.8177
R902 Vdd.n153 Vdd.t594 40.8177
R903 Vdd.n962 Vdd.t552 40.8177
R904 Vdd.n961 Vdd.t510 40.8177
R905 Vdd.n714 Vdd.t582 40.8177
R906 Vdd.n713 Vdd.t486 40.8177
R907 Vdd.n419 Vdd.t546 40.8177
R908 Vdd.n418 Vdd.t501 40.8177
R909 Vdd.n333 Vdd.t549 40.8177
R910 Vdd.n332 Vdd.t504 40.8177
R911 Vdd.n47 Vdd.t585 40.6313
R912 Vdd.n46 Vdd.t474 40.6313
R913 Vdd.n120 Vdd.t564 40.6313
R914 Vdd.n119 Vdd.t576 40.6313
R915 Vdd.n499 Vdd.t480 40.6313
R916 Vdd.n498 Vdd.t495 40.6313
R917 Vdd.n771 Vdd.t477 40.6313
R918 Vdd.n769 Vdd.t519 40.6313
R919 Vdd.n809 Vdd.t525 40.6313
R920 Vdd.n807 Vdd.t543 40.6313
R921 Vdd.n847 Vdd.t573 40.6313
R922 Vdd.n845 Vdd.t591 40.6313
R923 Vdd.n886 Vdd.t534 40.6313
R924 Vdd.n884 Vdd.t540 40.6313
R925 Vdd.n924 Vdd.t579 40.6313
R926 Vdd.n922 Vdd.t555 40.6313
R927 Vdd.n696 Vdd.t570 40.6313
R928 Vdd.n694 Vdd.t561 40.6313
R929 Vdd.n550 Vdd.t468 40.6313
R930 Vdd.n549 Vdd.t489 40.6313
R931 Vdd.n619 Vdd.t483 40.6313
R932 Vdd.n618 Vdd.t522 40.6313
R933 Vdd.n1 Vdd.t537 40.6313
R934 Vdd.n0 Vdd.t558 40.6313
R935 Vdd.n170 Vdd.n168 36.2255
R936 Vdd.n170 Vdd.n169 36.2255
R937 Vdd.n97 Vdd.n95 36.2255
R938 Vdd.n97 Vdd.n96 36.2255
R939 Vdd.n41 Vdd.n38 36.2255
R940 Vdd.n41 Vdd.n40 36.2255
R941 Vdd.n43 Vdd.n36 36.2255
R942 Vdd.n43 Vdd.n37 36.2255
R943 Vdd.n111 Vdd.n108 36.2255
R944 Vdd.n111 Vdd.n109 36.2255
R945 Vdd.n25 Vdd.n22 36.2255
R946 Vdd.n25 Vdd.n24 36.2255
R947 Vdd.n27 Vdd.n20 36.2255
R948 Vdd.n27 Vdd.n21 36.2255
R949 Vdd.n184 Vdd.n181 36.2255
R950 Vdd.n184 Vdd.n182 36.2255
R951 Vdd.n235 Vdd.n233 36.2255
R952 Vdd.n235 Vdd.n234 36.2255
R953 Vdd.n596 Vdd.n594 36.2255
R954 Vdd.n596 Vdd.n595 36.2255
R955 Vdd.n527 Vdd.n525 36.2255
R956 Vdd.n527 Vdd.n526 36.2255
R957 Vdd.n493 Vdd.n490 36.2255
R958 Vdd.n493 Vdd.n492 36.2255
R959 Vdd.n495 Vdd.n488 36.2255
R960 Vdd.n495 Vdd.n489 36.2255
R961 Vdd.n541 Vdd.n538 36.2255
R962 Vdd.n541 Vdd.n539 36.2255
R963 Vdd.n477 Vdd.n474 36.2255
R964 Vdd.n477 Vdd.n476 36.2255
R965 Vdd.n479 Vdd.n472 36.2255
R966 Vdd.n479 Vdd.n473 36.2255
R967 Vdd.n610 Vdd.n607 36.2255
R968 Vdd.n610 Vdd.n608 36.2255
R969 Vdd.n455 Vdd.n453 36.2255
R970 Vdd.n455 Vdd.n454 36.2255
R971 Vdd.n441 Vdd.n439 36.2255
R972 Vdd.n441 Vdd.n440 36.2255
R973 Vdd.n431 Vdd.n425 36.2255
R974 Vdd.n431 Vdd.n426 36.2255
R975 Vdd.n429 Vdd.n427 36.2255
R976 Vdd.n429 Vdd.n428 36.2255
R977 Vdd.n249 Vdd.n215 36.2255
R978 Vdd.n249 Vdd.n216 36.2255
R979 Vdd.n225 Vdd.n222 36.2255
R980 Vdd.n225 Vdd.n224 36.2255
R981 Vdd.n228 Vdd.n219 36.2255
R982 Vdd.n228 Vdd.n220 36.2255
R983 Vdd.n768 Vdd.n658 32.646
R984 Vdd.n1061 Vdd.n1060 29.3622
R985 Vdd.n1038 Vdd.n1037 29.3622
R986 Vdd.n47 Vdd.t956 27.3166
R987 Vdd.n46 Vdd.t948 27.3166
R988 Vdd.n120 Vdd.t961 27.3166
R989 Vdd.n119 Vdd.t959 27.3166
R990 Vdd.n499 Vdd.t947 27.3166
R991 Vdd.n498 Vdd.t983 27.3166
R992 Vdd.n771 Vdd.t958 27.3166
R993 Vdd.n769 Vdd.t974 27.3166
R994 Vdd.n809 Vdd.t946 27.3166
R995 Vdd.n807 Vdd.t965 27.3166
R996 Vdd.n847 Vdd.t969 27.3166
R997 Vdd.n845 Vdd.t954 27.3166
R998 Vdd.n886 Vdd.t987 27.3166
R999 Vdd.n884 Vdd.t966 27.3166
R1000 Vdd.n924 Vdd.t968 27.3166
R1001 Vdd.n922 Vdd.t964 27.3166
R1002 Vdd.n696 Vdd.t970 27.3166
R1003 Vdd.n694 Vdd.t962 27.3166
R1004 Vdd.n550 Vdd.t950 27.3166
R1005 Vdd.n549 Vdd.t984 27.3166
R1006 Vdd.n619 Vdd.t945 27.3166
R1007 Vdd.n618 Vdd.t973 27.3166
R1008 Vdd.n1 Vdd.t967 27.3166
R1009 Vdd.n0 Vdd.t963 27.3166
R1010 Vdd.n194 Vdd.t980 27.1302
R1011 Vdd.n193 Vdd.t972 27.1302
R1012 Vdd.n81 Vdd.t955 27.1302
R1013 Vdd.n80 Vdd.t949 27.1302
R1014 Vdd.n154 Vdd.t960 27.1302
R1015 Vdd.n153 Vdd.t953 27.1302
R1016 Vdd.n962 Vdd.t985 27.1302
R1017 Vdd.n961 Vdd.t977 27.1302
R1018 Vdd.n714 Vdd.t957 27.1302
R1019 Vdd.n713 Vdd.t944 27.1302
R1020 Vdd.n419 Vdd.t943 27.1302
R1021 Vdd.n418 Vdd.t981 27.1302
R1022 Vdd.n333 Vdd.t986 27.1302
R1023 Vdd.n332 Vdd.t978 27.1302
R1024 Vdd.n192 Vdd.t971 26.9438
R1025 Vdd.n79 Vdd.t976 26.9438
R1026 Vdd.n152 Vdd.t951 26.9438
R1027 Vdd.n960 Vdd.t975 26.9438
R1028 Vdd.n711 Vdd.t979 26.9438
R1029 Vdd.n417 Vdd.t952 26.9438
R1030 Vdd.n331 Vdd.t982 26.9438
R1031 Vdd.t294 Vdd.n1025 23.438
R1032 Vdd.n1053 Vdd.n1034 20.1255
R1033 Vdd.n1053 Vdd.n1035 20.1255
R1034 Vdd.n1055 Vdd.n1032 20.1255
R1035 Vdd.n1055 Vdd.n1033 20.1255
R1036 Vdd.n1062 Vdd.n1061 19.9167
R1037 Vdd.n1037 Vdd.n1036 19.9167
R1038 Vdd.n1012 Vdd.n1009 18.7255
R1039 Vdd.n1012 Vdd.n1010 18.7255
R1040 Vdd.n722 SARlogic_0.dffrs_13.resetb 18.2673
R1041 Vdd.n89 adc_PISO_0.dffrs_5.resetb 18.2415
R1042 Vdd.n162 adc_PISO_0.dffrs_4.resetb 18.2415
R1043 Vdd.n1072 adc_PISO_0.dffrs_3.resetb 18.2061
R1044 Vdd.n971 adc_PISO_0.dffrs_2.resetb 18.2061
R1045 Vdd.n658 adc_PISO_0.dffrs_0.resetb 18.2061
R1046 Vdd.n336 adc_PISO_0.dffrs_1.resetb 18.2061
R1047 Vdd.n55 Vdd.n49 18.0418
R1048 Vdd.n128 Vdd.n122 18.0418
R1049 Vdd.n507 Vdd.n501 18.0418
R1050 Vdd.n558 Vdd.n552 18.0418
R1051 Vdd.n627 Vdd.n621 18.0418
R1052 Vdd.n1099 Vdd.n1098 18.0418
R1053 Vdd.n774 Vdd.n773 18.0005
R1054 Vdd.n812 Vdd.n811 18.0005
R1055 Vdd.n850 Vdd.n849 18.0005
R1056 Vdd.n889 Vdd.n888 18.0005
R1057 Vdd.n927 Vdd.n926 18.0005
R1058 Vdd.n699 Vdd.n698 18.0005
R1059 Vdd.n195 Vdd.n193 17.6364
R1060 Vdd.n82 Vdd.n80 17.6364
R1061 Vdd.n155 Vdd.n153 17.6364
R1062 Vdd.n963 Vdd.n961 17.6364
R1063 Vdd.n420 Vdd.n418 17.6364
R1064 Vdd.n334 Vdd.n332 17.6364
R1065 Vdd.n1064 Vdd.n1063 14.6602
R1066 Vdd.n48 Vdd.n46 14.3609
R1067 Vdd.n121 Vdd.n119 14.3609
R1068 Vdd.n500 Vdd.n498 14.3609
R1069 Vdd.n551 Vdd.n549 14.3609
R1070 Vdd.n620 Vdd.n618 14.3609
R1071 Vdd.n2 Vdd.n0 14.3609
R1072 Vdd.n213 Vdd.n207 13.5842
R1073 Vdd.n507 Vdd.n506 13.5431
R1074 Vdd.n1098 Vdd.n7 13.5174
R1075 Vdd.n55 Vdd.n54 13.5174
R1076 Vdd.n128 Vdd.n127 13.5174
R1077 Vdd.n627 Vdd.n626 13.5174
R1078 Vdd.n558 Vdd.n557 13.5174
R1079 Vdd.n699 Vdd.n693 13.5152
R1080 Vdd.n1097 Vdd.n1096 13.5005
R1081 Vdd.n1097 Vdd.n12 13.5005
R1082 Vdd.n1085 Vdd.n1084 13.5005
R1083 Vdd.n1091 Vdd.n1090 13.5005
R1084 Vdd.n1078 Vdd.n1077 13.5005
R1085 Vdd.n66 Vdd.n65 13.5005
R1086 Vdd.n66 Vdd.n60 13.5005
R1087 Vdd.n78 Vdd.n77 13.5005
R1088 Vdd.n72 Vdd.n71 13.5005
R1089 Vdd.n89 Vdd.n88 13.5005
R1090 Vdd.n139 Vdd.n138 13.5005
R1091 Vdd.n139 Vdd.n133 13.5005
R1092 Vdd.n151 Vdd.n150 13.5005
R1093 Vdd.n145 Vdd.n144 13.5005
R1094 Vdd.n162 Vdd.n161 13.5005
R1095 Vdd.n213 Vdd.n212 13.5005
R1096 Vdd.n202 Vdd.n201 13.5005
R1097 Vdd.n1003 Vdd.n1002 13.5005
R1098 Vdd.n1003 Vdd.n985 13.5005
R1099 Vdd.n991 Vdd.n990 13.5005
R1100 Vdd.n997 Vdd.n996 13.5005
R1101 Vdd.n979 Vdd.n978 13.5005
R1102 Vdd.n513 Vdd.n512 13.5005
R1103 Vdd.n519 Vdd.n518 13.5005
R1104 Vdd.n970 Vdd.n969 13.5005
R1105 Vdd.n756 Vdd.n755 13.5005
R1106 Vdd.n795 Vdd.n794 13.5005
R1107 Vdd.n833 Vdd.n832 13.5005
R1108 Vdd.n871 Vdd.n870 13.5005
R1109 Vdd.n910 Vdd.n909 13.5005
R1110 Vdd.n948 Vdd.n947 13.5005
R1111 Vdd.n756 Vdd.n673 13.5005
R1112 Vdd.n767 Vdd.n766 13.5005
R1113 Vdd.n795 Vdd.n401 13.5005
R1114 Vdd.n806 Vdd.n805 13.5005
R1115 Vdd.n833 Vdd.n371 13.5005
R1116 Vdd.n844 Vdd.n843 13.5005
R1117 Vdd.n871 Vdd.n341 13.5005
R1118 Vdd.n883 Vdd.n882 13.5005
R1119 Vdd.n910 Vdd.n305 13.5005
R1120 Vdd.n921 Vdd.n920 13.5005
R1121 Vdd.n948 Vdd.n275 13.5005
R1122 Vdd.n959 Vdd.n958 13.5005
R1123 Vdd.n756 Vdd.n750 13.5005
R1124 Vdd.n767 Vdd.n663 13.5005
R1125 Vdd.n795 Vdd.n789 13.5005
R1126 Vdd.n806 Vdd.n391 13.5005
R1127 Vdd.n833 Vdd.n827 13.5005
R1128 Vdd.n844 Vdd.n361 13.5005
R1129 Vdd.n871 Vdd.n865 13.5005
R1130 Vdd.n883 Vdd.n325 13.5005
R1131 Vdd.n910 Vdd.n904 13.5005
R1132 Vdd.n921 Vdd.n295 13.5005
R1133 Vdd.n948 Vdd.n942 13.5005
R1134 Vdd.n959 Vdd.n265 13.5005
R1135 Vdd.n756 Vdd.n678 13.5005
R1136 Vdd.n795 Vdd.n406 13.5005
R1137 Vdd.n833 Vdd.n376 13.5005
R1138 Vdd.n871 Vdd.n346 13.5005
R1139 Vdd.n910 Vdd.n310 13.5005
R1140 Vdd.n948 Vdd.n280 13.5005
R1141 Vdd.n756 Vdd.n745 13.5005
R1142 Vdd.n756 Vdd.n683 13.5005
R1143 Vdd.n795 Vdd.n784 13.5005
R1144 Vdd.n767 Vdd.n761 13.5005
R1145 Vdd.n795 Vdd.n411 13.5005
R1146 Vdd.n833 Vdd.n822 13.5005
R1147 Vdd.n806 Vdd.n800 13.5005
R1148 Vdd.n833 Vdd.n381 13.5005
R1149 Vdd.n871 Vdd.n860 13.5005
R1150 Vdd.n844 Vdd.n838 13.5005
R1151 Vdd.n871 Vdd.n351 13.5005
R1152 Vdd.n910 Vdd.n899 13.5005
R1153 Vdd.n883 Vdd.n877 13.5005
R1154 Vdd.n910 Vdd.n315 13.5005
R1155 Vdd.n948 Vdd.n937 13.5005
R1156 Vdd.n921 Vdd.n915 13.5005
R1157 Vdd.n948 Vdd.n285 13.5005
R1158 Vdd.n959 Vdd.n953 13.5005
R1159 Vdd.n756 Vdd.n740 13.5005
R1160 Vdd.n767 Vdd.n668 13.5005
R1161 Vdd.n795 Vdd.n779 13.5005
R1162 Vdd.n806 Vdd.n396 13.5005
R1163 Vdd.n833 Vdd.n817 13.5005
R1164 Vdd.n844 Vdd.n366 13.5005
R1165 Vdd.n871 Vdd.n855 13.5005
R1166 Vdd.n883 Vdd.n330 13.5005
R1167 Vdd.n910 Vdd.n894 13.5005
R1168 Vdd.n921 Vdd.n300 13.5005
R1169 Vdd.n948 Vdd.n932 13.5005
R1170 Vdd.n959 Vdd.n270 13.5005
R1171 Vdd.n756 Vdd.n688 13.5005
R1172 Vdd.n795 Vdd.n416 13.5005
R1173 Vdd.n833 Vdd.n386 13.5005
R1174 Vdd.n871 Vdd.n356 13.5005
R1175 Vdd.n910 Vdd.n320 13.5005
R1176 Vdd.n948 Vdd.n290 13.5005
R1177 Vdd.n710 Vdd.n709 13.5005
R1178 Vdd.n710 Vdd.n704 13.5005
R1179 Vdd.n728 Vdd.n727 13.5005
R1180 Vdd.n734 Vdd.n733 13.5005
R1181 Vdd.n722 Vdd.n721 13.5005
R1182 Vdd.n638 Vdd.n637 13.5005
R1183 Vdd.n638 Vdd.n632 13.5005
R1184 Vdd.n650 Vdd.n649 13.5005
R1185 Vdd.n644 Vdd.n643 13.5005
R1186 Vdd.n657 Vdd.n656 13.5005
R1187 Vdd.n569 Vdd.n568 13.5005
R1188 Vdd.n569 Vdd.n563 13.5005
R1189 Vdd.n581 Vdd.n580 13.5005
R1190 Vdd.n575 Vdd.n574 13.5005
R1191 Vdd.n588 Vdd.n587 13.5005
R1192 Vdd.n1069 Vdd.n1006 13.4987
R1193 Vdd.n196 Vdd.n192 13.4839
R1194 Vdd.n83 Vdd.n79 13.4839
R1195 Vdd.n156 Vdd.n152 13.4839
R1196 Vdd.n964 Vdd.n960 13.4839
R1197 Vdd.n421 Vdd.n417 13.4839
R1198 Vdd.n335 Vdd.n331 13.4839
R1199 Vdd.n1025 Vdd.n1019 12.6005
R1200 Vdd.n1029 Vdd.n1028 12.6005
R1201 Vdd.n1027 Vdd.n1026 12.6005
R1202 Vdd.n715 SARlogic_0.dffrs_13.nand3_1.B 12.1571
R1203 Vdd.n1051 Vdd.n1050 12.136
R1204 Vdd.n1049 Vdd.n1048 12.136
R1205 Vdd.n1047 Vdd.n1046 12.136
R1206 Vdd.n1045 Vdd.n1044 12.136
R1207 Vdd.n1043 Vdd.n1042 12.136
R1208 Vdd.n1055 Vdd.n1031 11.111
R1209 Vdd.n1053 Vdd.n1052 11.111
R1210 Vdd.n195 Vdd.n194 10.5752
R1211 Vdd.n82 Vdd.n81 10.5752
R1212 Vdd.n155 Vdd.n154 10.5752
R1213 Vdd.n963 Vdd.n962 10.5752
R1214 Vdd.n420 Vdd.n419 10.5752
R1215 Vdd.n334 Vdd.n333 10.5752
R1216 Vdd.n1036 Vdd.n1006 9.86945
R1217 Vdd.n1041 Vdd.n1040 9.536
R1218 Vdd.n1059 Vdd.n1058 9.536
R1219 Vdd.n1063 Vdd.n1062 9.536
R1220 Vdd.n772 Vdd.n770 9.22229
R1221 Vdd.n810 Vdd.n808 9.22229
R1222 Vdd.n848 Vdd.n846 9.22229
R1223 Vdd.n887 Vdd.n885 9.22229
R1224 Vdd.n925 Vdd.n923 9.22229
R1225 Vdd.n697 Vdd.n695 9.22229
R1226 Vdd.n716 Vdd.n712 7.75389
R1227 Vdd.n1040 Vdd.t720 7.4755
R1228 Vdd.n1058 Vdd.t736 7.4755
R1229 Vdd.n1062 Vdd.t696 7.4755
R1230 Vdd.n1036 Vdd.t732 7.4755
R1231 Vdd.n973 Vdd.n972 6.55364
R1232 Vdd.n7 Vdd.n4 6.4802
R1233 Vdd.n1096 Vdd.n1093 6.4802
R1234 Vdd.n12 Vdd.n9 6.4802
R1235 Vdd.n1084 Vdd.n1081 6.4802
R1236 Vdd.n1090 Vdd.n1087 6.4802
R1237 Vdd.n1077 Vdd.n1074 6.4802
R1238 Vdd.n54 Vdd.n51 6.4802
R1239 Vdd.n65 Vdd.n62 6.4802
R1240 Vdd.n60 Vdd.n57 6.4802
R1241 Vdd.n77 Vdd.n74 6.4802
R1242 Vdd.n71 Vdd.n68 6.4802
R1243 Vdd.n88 Vdd.n85 6.4802
R1244 Vdd.n127 Vdd.n124 6.4802
R1245 Vdd.n138 Vdd.n135 6.4802
R1246 Vdd.n133 Vdd.n130 6.4802
R1247 Vdd.n150 Vdd.n147 6.4802
R1248 Vdd.n144 Vdd.n141 6.4802
R1249 Vdd.n161 Vdd.n158 6.4802
R1250 Vdd.n207 Vdd.n204 6.4802
R1251 Vdd.n212 Vdd.n209 6.4802
R1252 Vdd.n201 Vdd.n198 6.4802
R1253 Vdd.n1002 Vdd.n999 6.4802
R1254 Vdd.n985 Vdd.n982 6.4802
R1255 Vdd.n990 Vdd.n987 6.4802
R1256 Vdd.n996 Vdd.n993 6.4802
R1257 Vdd.n978 Vdd.n975 6.4802
R1258 Vdd.n506 Vdd.n503 6.4802
R1259 Vdd.n512 Vdd.n509 6.4802
R1260 Vdd.n518 Vdd.n515 6.4802
R1261 Vdd.n969 Vdd.n966 6.4802
R1262 Vdd.n755 Vdd.n752 6.4802
R1263 Vdd.n794 Vdd.n791 6.4802
R1264 Vdd.n832 Vdd.n829 6.4802
R1265 Vdd.n870 Vdd.n867 6.4802
R1266 Vdd.n909 Vdd.n906 6.4802
R1267 Vdd.n947 Vdd.n944 6.4802
R1268 Vdd.n673 Vdd.n670 6.4802
R1269 Vdd.n766 Vdd.n763 6.4802
R1270 Vdd.n401 Vdd.n398 6.4802
R1271 Vdd.n805 Vdd.n802 6.4802
R1272 Vdd.n371 Vdd.n368 6.4802
R1273 Vdd.n843 Vdd.n840 6.4802
R1274 Vdd.n341 Vdd.n338 6.4802
R1275 Vdd.n882 Vdd.n879 6.4802
R1276 Vdd.n305 Vdd.n302 6.4802
R1277 Vdd.n920 Vdd.n917 6.4802
R1278 Vdd.n275 Vdd.n272 6.4802
R1279 Vdd.n958 Vdd.n955 6.4802
R1280 Vdd.n750 Vdd.n747 6.4802
R1281 Vdd.n663 Vdd.n660 6.4802
R1282 Vdd.n789 Vdd.n786 6.4802
R1283 Vdd.n391 Vdd.n388 6.4802
R1284 Vdd.n827 Vdd.n824 6.4802
R1285 Vdd.n361 Vdd.n358 6.4802
R1286 Vdd.n865 Vdd.n862 6.4802
R1287 Vdd.n325 Vdd.n322 6.4802
R1288 Vdd.n904 Vdd.n901 6.4802
R1289 Vdd.n295 Vdd.n292 6.4802
R1290 Vdd.n942 Vdd.n939 6.4802
R1291 Vdd.n265 Vdd.n262 6.4802
R1292 Vdd.n678 Vdd.n675 6.4802
R1293 Vdd.n406 Vdd.n403 6.4802
R1294 Vdd.n376 Vdd.n373 6.4802
R1295 Vdd.n346 Vdd.n343 6.4802
R1296 Vdd.n310 Vdd.n307 6.4802
R1297 Vdd.n280 Vdd.n277 6.4802
R1298 Vdd.n745 Vdd.n742 6.4802
R1299 Vdd.n683 Vdd.n680 6.4802
R1300 Vdd.n784 Vdd.n781 6.4802
R1301 Vdd.n761 Vdd.n758 6.4802
R1302 Vdd.n411 Vdd.n408 6.4802
R1303 Vdd.n822 Vdd.n819 6.4802
R1304 Vdd.n800 Vdd.n797 6.4802
R1305 Vdd.n381 Vdd.n378 6.4802
R1306 Vdd.n860 Vdd.n857 6.4802
R1307 Vdd.n838 Vdd.n835 6.4802
R1308 Vdd.n351 Vdd.n348 6.4802
R1309 Vdd.n899 Vdd.n896 6.4802
R1310 Vdd.n877 Vdd.n874 6.4802
R1311 Vdd.n315 Vdd.n312 6.4802
R1312 Vdd.n937 Vdd.n934 6.4802
R1313 Vdd.n915 Vdd.n912 6.4802
R1314 Vdd.n285 Vdd.n282 6.4802
R1315 Vdd.n953 Vdd.n950 6.4802
R1316 Vdd.n740 Vdd.n737 6.4802
R1317 Vdd.n668 Vdd.n665 6.4802
R1318 Vdd.n779 Vdd.n776 6.4802
R1319 Vdd.n396 Vdd.n393 6.4802
R1320 Vdd.n817 Vdd.n814 6.4802
R1321 Vdd.n366 Vdd.n363 6.4802
R1322 Vdd.n855 Vdd.n852 6.4802
R1323 Vdd.n330 Vdd.n327 6.4802
R1324 Vdd.n894 Vdd.n891 6.4802
R1325 Vdd.n300 Vdd.n297 6.4802
R1326 Vdd.n932 Vdd.n929 6.4802
R1327 Vdd.n270 Vdd.n267 6.4802
R1328 Vdd.n688 Vdd.n685 6.4802
R1329 Vdd.n416 Vdd.n413 6.4802
R1330 Vdd.n386 Vdd.n383 6.4802
R1331 Vdd.n356 Vdd.n353 6.4802
R1332 Vdd.n320 Vdd.n317 6.4802
R1333 Vdd.n290 Vdd.n287 6.4802
R1334 Vdd.n693 Vdd.n690 6.4802
R1335 Vdd.n709 Vdd.n706 6.4802
R1336 Vdd.n704 Vdd.n701 6.4802
R1337 Vdd.n727 Vdd.n724 6.4802
R1338 Vdd.n733 Vdd.n730 6.4802
R1339 Vdd.n721 Vdd.n718 6.4802
R1340 Vdd.n626 Vdd.n623 6.4802
R1341 Vdd.n637 Vdd.n634 6.4802
R1342 Vdd.n632 Vdd.n629 6.4802
R1343 Vdd.n649 Vdd.n646 6.4802
R1344 Vdd.n643 Vdd.n640 6.4802
R1345 Vdd.n656 Vdd.n653 6.4802
R1346 Vdd.n557 Vdd.n554 6.4802
R1347 Vdd.n568 Vdd.n565 6.4802
R1348 Vdd.n563 Vdd.n560 6.4802
R1349 Vdd.n580 Vdd.n577 6.4802
R1350 Vdd.n574 Vdd.n571 6.4802
R1351 Vdd.n587 Vdd.n584 6.4802
R1352 Vdd.n7 Vdd.n3 6.25878
R1353 Vdd.n1096 Vdd.n1092 6.25878
R1354 Vdd.n12 Vdd.n8 6.25878
R1355 Vdd.n1084 Vdd.n1080 6.25878
R1356 Vdd.n1090 Vdd.n1086 6.25878
R1357 Vdd.n1077 Vdd.n1073 6.25878
R1358 Vdd.n54 Vdd.n50 6.25878
R1359 Vdd.n65 Vdd.n61 6.25878
R1360 Vdd.n60 Vdd.n56 6.25878
R1361 Vdd.n77 Vdd.n73 6.25878
R1362 Vdd.n71 Vdd.n67 6.25878
R1363 Vdd.n88 Vdd.n84 6.25878
R1364 Vdd.n127 Vdd.n123 6.25878
R1365 Vdd.n138 Vdd.n134 6.25878
R1366 Vdd.n133 Vdd.n129 6.25878
R1367 Vdd.n150 Vdd.n146 6.25878
R1368 Vdd.n144 Vdd.n140 6.25878
R1369 Vdd.n161 Vdd.n157 6.25878
R1370 Vdd.n207 Vdd.n203 6.25878
R1371 Vdd.n212 Vdd.n208 6.25878
R1372 Vdd.n201 Vdd.n197 6.25878
R1373 Vdd.n1002 Vdd.n998 6.25878
R1374 Vdd.n985 Vdd.n981 6.25878
R1375 Vdd.n990 Vdd.n986 6.25878
R1376 Vdd.n996 Vdd.n992 6.25878
R1377 Vdd.n978 Vdd.n974 6.25878
R1378 Vdd.n506 Vdd.n502 6.25878
R1379 Vdd.n512 Vdd.n508 6.25878
R1380 Vdd.n518 Vdd.n514 6.25878
R1381 Vdd.n969 Vdd.n965 6.25878
R1382 Vdd.n755 Vdd.n751 6.25878
R1383 Vdd.n794 Vdd.n790 6.25878
R1384 Vdd.n832 Vdd.n828 6.25878
R1385 Vdd.n870 Vdd.n866 6.25878
R1386 Vdd.n909 Vdd.n905 6.25878
R1387 Vdd.n947 Vdd.n943 6.25878
R1388 Vdd.n673 Vdd.n669 6.25878
R1389 Vdd.n766 Vdd.n762 6.25878
R1390 Vdd.n401 Vdd.n397 6.25878
R1391 Vdd.n805 Vdd.n801 6.25878
R1392 Vdd.n371 Vdd.n367 6.25878
R1393 Vdd.n843 Vdd.n839 6.25878
R1394 Vdd.n341 Vdd.n337 6.25878
R1395 Vdd.n882 Vdd.n878 6.25878
R1396 Vdd.n305 Vdd.n301 6.25878
R1397 Vdd.n920 Vdd.n916 6.25878
R1398 Vdd.n275 Vdd.n271 6.25878
R1399 Vdd.n958 Vdd.n954 6.25878
R1400 Vdd.n750 Vdd.n746 6.25878
R1401 Vdd.n663 Vdd.n659 6.25878
R1402 Vdd.n789 Vdd.n785 6.25878
R1403 Vdd.n391 Vdd.n387 6.25878
R1404 Vdd.n827 Vdd.n823 6.25878
R1405 Vdd.n361 Vdd.n357 6.25878
R1406 Vdd.n865 Vdd.n861 6.25878
R1407 Vdd.n325 Vdd.n321 6.25878
R1408 Vdd.n904 Vdd.n900 6.25878
R1409 Vdd.n295 Vdd.n291 6.25878
R1410 Vdd.n942 Vdd.n938 6.25878
R1411 Vdd.n265 Vdd.n261 6.25878
R1412 Vdd.n678 Vdd.n674 6.25878
R1413 Vdd.n406 Vdd.n402 6.25878
R1414 Vdd.n376 Vdd.n372 6.25878
R1415 Vdd.n346 Vdd.n342 6.25878
R1416 Vdd.n310 Vdd.n306 6.25878
R1417 Vdd.n280 Vdd.n276 6.25878
R1418 Vdd.n745 Vdd.n741 6.25878
R1419 Vdd.n683 Vdd.n679 6.25878
R1420 Vdd.n784 Vdd.n780 6.25878
R1421 Vdd.n761 Vdd.n757 6.25878
R1422 Vdd.n411 Vdd.n407 6.25878
R1423 Vdd.n822 Vdd.n818 6.25878
R1424 Vdd.n800 Vdd.n796 6.25878
R1425 Vdd.n381 Vdd.n377 6.25878
R1426 Vdd.n860 Vdd.n856 6.25878
R1427 Vdd.n838 Vdd.n834 6.25878
R1428 Vdd.n351 Vdd.n347 6.25878
R1429 Vdd.n899 Vdd.n895 6.25878
R1430 Vdd.n877 Vdd.n873 6.25878
R1431 Vdd.n315 Vdd.n311 6.25878
R1432 Vdd.n937 Vdd.n933 6.25878
R1433 Vdd.n915 Vdd.n911 6.25878
R1434 Vdd.n285 Vdd.n281 6.25878
R1435 Vdd.n953 Vdd.n949 6.25878
R1436 Vdd.n740 Vdd.n736 6.25878
R1437 Vdd.n668 Vdd.n664 6.25878
R1438 Vdd.n779 Vdd.n775 6.25878
R1439 Vdd.n396 Vdd.n392 6.25878
R1440 Vdd.n817 Vdd.n813 6.25878
R1441 Vdd.n366 Vdd.n362 6.25878
R1442 Vdd.n855 Vdd.n851 6.25878
R1443 Vdd.n330 Vdd.n326 6.25878
R1444 Vdd.n894 Vdd.n890 6.25878
R1445 Vdd.n300 Vdd.n296 6.25878
R1446 Vdd.n932 Vdd.n928 6.25878
R1447 Vdd.n270 Vdd.n266 6.25878
R1448 Vdd.n688 Vdd.n684 6.25878
R1449 Vdd.n416 Vdd.n412 6.25878
R1450 Vdd.n386 Vdd.n382 6.25878
R1451 Vdd.n356 Vdd.n352 6.25878
R1452 Vdd.n320 Vdd.n316 6.25878
R1453 Vdd.n290 Vdd.n286 6.25878
R1454 Vdd.n693 Vdd.n689 6.25878
R1455 Vdd.n709 Vdd.n705 6.25878
R1456 Vdd.n704 Vdd.n700 6.25878
R1457 Vdd.n727 Vdd.n723 6.25878
R1458 Vdd.n733 Vdd.n729 6.25878
R1459 Vdd.n721 Vdd.n717 6.25878
R1460 Vdd.n626 Vdd.n622 6.25878
R1461 Vdd.n637 Vdd.n633 6.25878
R1462 Vdd.n632 Vdd.n628 6.25878
R1463 Vdd.n649 Vdd.n645 6.25878
R1464 Vdd.n643 Vdd.n639 6.25878
R1465 Vdd.n656 Vdd.n652 6.25878
R1466 Vdd.n557 Vdd.n553 6.25878
R1467 Vdd.n568 Vdd.n564 6.25878
R1468 Vdd.n563 Vdd.n559 6.25878
R1469 Vdd.n580 Vdd.n576 6.25878
R1470 Vdd.n574 Vdd.n570 6.25878
R1471 Vdd.n587 Vdd.n583 6.25878
R1472 Vdd.n196 Vdd.n195 5.93546
R1473 Vdd.n83 Vdd.n82 5.93546
R1474 Vdd.n156 Vdd.n155 5.93546
R1475 Vdd.n964 Vdd.n963 5.93546
R1476 Vdd.n716 Vdd.n715 5.93546
R1477 Vdd.n421 Vdd.n420 5.93546
R1478 Vdd.n335 Vdd.n334 5.93546
R1479 Vdd.n712 Vdd.n711 5.7305
R1480 SARlogic_0.dffrs_13.nand3_8.B Vdd.n714 5.47979
R1481 SARlogic_0.dffrs_13.nand3_1.B Vdd.n713 5.47979
R1482 Vdd.n7 Vdd.n6 5.44497
R1483 Vdd.n1096 Vdd.n1095 5.44497
R1484 Vdd.n12 Vdd.n11 5.44497
R1485 Vdd.n1084 Vdd.n1083 5.44497
R1486 Vdd.n1090 Vdd.n1089 5.44497
R1487 Vdd.n1077 Vdd.n1076 5.44497
R1488 Vdd.n54 Vdd.n53 5.44497
R1489 Vdd.n65 Vdd.n64 5.44497
R1490 Vdd.n60 Vdd.n59 5.44497
R1491 Vdd.n77 Vdd.n76 5.44497
R1492 Vdd.n71 Vdd.n70 5.44497
R1493 Vdd.n88 Vdd.n87 5.44497
R1494 Vdd.n127 Vdd.n126 5.44497
R1495 Vdd.n138 Vdd.n137 5.44497
R1496 Vdd.n133 Vdd.n132 5.44497
R1497 Vdd.n150 Vdd.n149 5.44497
R1498 Vdd.n144 Vdd.n143 5.44497
R1499 Vdd.n161 Vdd.n160 5.44497
R1500 Vdd.n207 Vdd.n206 5.44497
R1501 Vdd.n212 Vdd.n211 5.44497
R1502 Vdd.n201 Vdd.n200 5.44497
R1503 Vdd.n1002 Vdd.n1001 5.44497
R1504 Vdd.n985 Vdd.n984 5.44497
R1505 Vdd.n990 Vdd.n989 5.44497
R1506 Vdd.n996 Vdd.n995 5.44497
R1507 Vdd.n978 Vdd.n977 5.44497
R1508 Vdd.n506 Vdd.n505 5.44497
R1509 Vdd.n512 Vdd.n511 5.44497
R1510 Vdd.n518 Vdd.n517 5.44497
R1511 Vdd.n969 Vdd.n968 5.44497
R1512 Vdd.n755 Vdd.n754 5.44497
R1513 Vdd.n794 Vdd.n793 5.44497
R1514 Vdd.n832 Vdd.n831 5.44497
R1515 Vdd.n870 Vdd.n869 5.44497
R1516 Vdd.n909 Vdd.n908 5.44497
R1517 Vdd.n947 Vdd.n946 5.44497
R1518 Vdd.n673 Vdd.n672 5.44497
R1519 Vdd.n766 Vdd.n765 5.44497
R1520 Vdd.n401 Vdd.n400 5.44497
R1521 Vdd.n805 Vdd.n804 5.44497
R1522 Vdd.n371 Vdd.n370 5.44497
R1523 Vdd.n843 Vdd.n842 5.44497
R1524 Vdd.n341 Vdd.n340 5.44497
R1525 Vdd.n882 Vdd.n881 5.44497
R1526 Vdd.n305 Vdd.n304 5.44497
R1527 Vdd.n920 Vdd.n919 5.44497
R1528 Vdd.n275 Vdd.n274 5.44497
R1529 Vdd.n958 Vdd.n957 5.44497
R1530 Vdd.n750 Vdd.n749 5.44497
R1531 Vdd.n663 Vdd.n662 5.44497
R1532 Vdd.n789 Vdd.n788 5.44497
R1533 Vdd.n391 Vdd.n390 5.44497
R1534 Vdd.n827 Vdd.n826 5.44497
R1535 Vdd.n361 Vdd.n360 5.44497
R1536 Vdd.n865 Vdd.n864 5.44497
R1537 Vdd.n325 Vdd.n324 5.44497
R1538 Vdd.n904 Vdd.n903 5.44497
R1539 Vdd.n295 Vdd.n294 5.44497
R1540 Vdd.n942 Vdd.n941 5.44497
R1541 Vdd.n265 Vdd.n264 5.44497
R1542 Vdd.n678 Vdd.n677 5.44497
R1543 Vdd.n406 Vdd.n405 5.44497
R1544 Vdd.n376 Vdd.n375 5.44497
R1545 Vdd.n346 Vdd.n345 5.44497
R1546 Vdd.n310 Vdd.n309 5.44497
R1547 Vdd.n280 Vdd.n279 5.44497
R1548 Vdd.n745 Vdd.n744 5.44497
R1549 Vdd.n683 Vdd.n682 5.44497
R1550 Vdd.n784 Vdd.n783 5.44497
R1551 Vdd.n761 Vdd.n760 5.44497
R1552 Vdd.n411 Vdd.n410 5.44497
R1553 Vdd.n822 Vdd.n821 5.44497
R1554 Vdd.n800 Vdd.n799 5.44497
R1555 Vdd.n381 Vdd.n380 5.44497
R1556 Vdd.n860 Vdd.n859 5.44497
R1557 Vdd.n838 Vdd.n837 5.44497
R1558 Vdd.n351 Vdd.n350 5.44497
R1559 Vdd.n899 Vdd.n898 5.44497
R1560 Vdd.n877 Vdd.n876 5.44497
R1561 Vdd.n315 Vdd.n314 5.44497
R1562 Vdd.n937 Vdd.n936 5.44497
R1563 Vdd.n915 Vdd.n914 5.44497
R1564 Vdd.n285 Vdd.n284 5.44497
R1565 Vdd.n953 Vdd.n952 5.44497
R1566 Vdd.n740 Vdd.n739 5.44497
R1567 Vdd.n668 Vdd.n667 5.44497
R1568 Vdd.n779 Vdd.n778 5.44497
R1569 Vdd.n396 Vdd.n395 5.44497
R1570 Vdd.n817 Vdd.n816 5.44497
R1571 Vdd.n366 Vdd.n365 5.44497
R1572 Vdd.n855 Vdd.n854 5.44497
R1573 Vdd.n330 Vdd.n329 5.44497
R1574 Vdd.n894 Vdd.n893 5.44497
R1575 Vdd.n300 Vdd.n299 5.44497
R1576 Vdd.n932 Vdd.n931 5.44497
R1577 Vdd.n270 Vdd.n269 5.44497
R1578 Vdd.n688 Vdd.n687 5.44497
R1579 Vdd.n416 Vdd.n415 5.44497
R1580 Vdd.n386 Vdd.n385 5.44497
R1581 Vdd.n356 Vdd.n355 5.44497
R1582 Vdd.n320 Vdd.n319 5.44497
R1583 Vdd.n290 Vdd.n289 5.44497
R1584 Vdd.n693 Vdd.n692 5.44497
R1585 Vdd.n709 Vdd.n708 5.44497
R1586 Vdd.n704 Vdd.n703 5.44497
R1587 Vdd.n727 Vdd.n726 5.44497
R1588 Vdd.n733 Vdd.n732 5.44497
R1589 Vdd.n721 Vdd.n720 5.44497
R1590 Vdd.n626 Vdd.n625 5.44497
R1591 Vdd.n637 Vdd.n636 5.44497
R1592 Vdd.n632 Vdd.n631 5.44497
R1593 Vdd.n649 Vdd.n648 5.44497
R1594 Vdd.n643 Vdd.n642 5.44497
R1595 Vdd.n656 Vdd.n655 5.44497
R1596 Vdd.n557 Vdd.n556 5.44497
R1597 Vdd.n568 Vdd.n567 5.44497
R1598 Vdd.n563 Vdd.n562 5.44497
R1599 Vdd.n580 Vdd.n579 5.44497
R1600 Vdd.n574 Vdd.n573 5.44497
R1601 Vdd.n587 Vdd.n586 5.44497
R1602 Vdd.n48 Vdd.n47 5.14711
R1603 Vdd.n121 Vdd.n120 5.14711
R1604 Vdd.n500 Vdd.n499 5.14711
R1605 Vdd.n772 Vdd.n771 5.14711
R1606 Vdd.n810 Vdd.n809 5.14711
R1607 Vdd.n848 Vdd.n847 5.14711
R1608 Vdd.n887 Vdd.n886 5.14711
R1609 Vdd.n925 Vdd.n924 5.14711
R1610 Vdd.n697 Vdd.n696 5.14711
R1611 Vdd.n551 Vdd.n550 5.14711
R1612 Vdd.n620 Vdd.n619 5.14711
R1613 Vdd.n2 Vdd.n1 5.14711
R1614 Vdd.n770 Vdd.n769 5.13907
R1615 Vdd.n808 Vdd.n807 5.13907
R1616 Vdd.n846 Vdd.n845 5.13907
R1617 Vdd.n885 Vdd.n884 5.13907
R1618 Vdd.n923 Vdd.n922 5.13907
R1619 Vdd.n695 Vdd.n694 5.13907
R1620 Vdd.n715 SARlogic_0.dffrs_13.nand3_8.B 5.09593
R1621 Vdd.n1070 Vdd.n1069 4.98176
R1622 Vdd.n1015 Vdd.t67 4.4205
R1623 Vdd.n1008 Vdd.t113 4.4205
R1624 Vdd.n973 Vdd.n260 4.3905
R1625 Vdd.n1026 Vdd.t299 3.38176
R1626 Vdd.n178 Vdd.n177 2.49936
R1627 Vdd.n105 Vdd.n104 2.49936
R1628 Vdd.n243 Vdd.n242 2.49936
R1629 Vdd.n604 Vdd.n603 2.49936
R1630 Vdd.n535 Vdd.n534 2.49936
R1631 Vdd.n463 Vdd.n462 2.49936
R1632 Vdd.n1040 Vdd.n1039 2.1905
R1633 Vdd.n1058 Vdd.n1057 2.1905
R1634 Vdd.n1021 Vdd.n1020 2.16583
R1635 Vdd.n1023 Vdd.n1022 2.16583
R1636 Vdd.n1007 Vdd.t235 1.99236
R1637 Vdd.n177 Vdd.n166 1.93883
R1638 Vdd.n104 Vdd.n93 1.93883
R1639 Vdd.n242 Vdd.n231 1.93883
R1640 Vdd.n603 Vdd.n592 1.93883
R1641 Vdd.n534 Vdd.n523 1.93883
R1642 Vdd.n462 Vdd.n451 1.93883
R1643 Vdd.n1017 Vdd.t652 1.91107
R1644 Vdd.n979 Vdd.n973 1.89424
R1645 Vdd.n6 Vdd.t539 1.85637
R1646 Vdd.n1095 Vdd.t654 1.85637
R1647 Vdd.n11 Vdd.t560 1.85637
R1648 Vdd.n1083 Vdd.t932 1.85637
R1649 Vdd.n1089 Vdd.t656 1.85637
R1650 Vdd.n1076 Vdd.t99 1.85637
R1651 Vdd.n53 Vdd.t587 1.85637
R1652 Vdd.n64 Vdd.t830 1.85637
R1653 Vdd.n59 Vdd.t476 1.85637
R1654 Vdd.n76 Vdd.t285 1.85637
R1655 Vdd.n70 Vdd.t449 1.85637
R1656 Vdd.n87 Vdd.t411 1.85637
R1657 Vdd.n126 Vdd.t566 1.85637
R1658 Vdd.n137 Vdd.t217 1.85637
R1659 Vdd.n132 Vdd.t578 1.85637
R1660 Vdd.n149 Vdd.t241 1.85637
R1661 Vdd.n143 Vdd.t920 1.85637
R1662 Vdd.n160 Vdd.t29 1.85637
R1663 Vdd.n206 Vdd.t497 1.85637
R1664 Vdd.n211 Vdd.t33 1.85637
R1665 Vdd.n200 Vdd.t103 1.85637
R1666 Vdd.n1001 Vdd.t47 1.85637
R1667 Vdd.n984 Vdd.t37 1.85637
R1668 Vdd.n989 Vdd.t868 1.85637
R1669 Vdd.n995 Vdd.t794 1.85637
R1670 Vdd.n977 Vdd.t884 1.85637
R1671 Vdd.n505 Vdd.t482 1.85637
R1672 Vdd.n511 Vdd.t267 1.85637
R1673 Vdd.n517 Vdd.t880 1.85637
R1674 Vdd.n968 Vdd.t814 1.85637
R1675 Vdd.n754 Vdd.t369 1.85637
R1676 Vdd.n793 Vdd.t265 1.85637
R1677 Vdd.n831 Vdd.t273 1.85637
R1678 Vdd.n869 Vdd.t748 1.85637
R1679 Vdd.n908 Vdd.t213 1.85637
R1680 Vdd.n946 Vdd.t912 1.85637
R1681 Vdd.n672 Vdd.t395 1.85637
R1682 Vdd.n765 Vdd.t187 1.85637
R1683 Vdd.n400 Vdd.t125 1.85637
R1684 Vdd.n804 Vdd.t43 1.85637
R1685 Vdd.n370 Vdd.t51 1.85637
R1686 Vdd.n842 Vdd.t271 1.85637
R1687 Vdd.n340 Vdd.t367 1.85637
R1688 Vdd.n881 Vdd.t746 1.85637
R1689 Vdd.n304 Vdd.t291 1.85637
R1690 Vdd.n919 Vdd.t211 1.85637
R1691 Vdd.n274 Vdd.t313 1.85637
R1692 Vdd.n957 Vdd.t177 1.85637
R1693 Vdd.n749 Vdd.t778 1.85637
R1694 Vdd.n662 Vdd.t930 1.85637
R1695 Vdd.n788 Vdd.t149 1.85637
R1696 Vdd.n390 Vdd.t175 1.85637
R1697 Vdd.n826 Vdd.t243 1.85637
R1698 Vdd.n360 Vdd.t87 1.85637
R1699 Vdd.n864 Vdd.t900 1.85637
R1700 Vdd.n324 Vdd.t924 1.85637
R1701 Vdd.n903 Vdd.t201 1.85637
R1702 Vdd.n294 Vdd.t682 1.85637
R1703 Vdd.n941 Vdd.t373 1.85637
R1704 Vdd.n264 Vdd.t798 1.85637
R1705 Vdd.n677 Vdd.t788 1.85637
R1706 Vdd.n405 Vdd.t908 1.85637
R1707 Vdd.n375 Vdd.t323 1.85637
R1708 Vdd.n345 Vdd.t259 1.85637
R1709 Vdd.n309 Vdd.t850 1.85637
R1710 Vdd.n279 Vdd.t227 1.85637
R1711 Vdd.n744 Vdd.t572 1.85637
R1712 Vdd.n682 Vdd.t319 1.85637
R1713 Vdd.n783 Vdd.t479 1.85637
R1714 Vdd.n760 Vdd.t563 1.85637
R1715 Vdd.n410 Vdd.t1 1.85637
R1716 Vdd.n821 Vdd.t527 1.85637
R1717 Vdd.n799 Vdd.t521 1.85637
R1718 Vdd.n380 Vdd.t914 1.85637
R1719 Vdd.n859 Vdd.t575 1.85637
R1720 Vdd.n837 Vdd.t545 1.85637
R1721 Vdd.n350 Vdd.t41 1.85637
R1722 Vdd.n898 Vdd.t536 1.85637
R1723 Vdd.n876 Vdd.t593 1.85637
R1724 Vdd.n314 Vdd.t872 1.85637
R1725 Vdd.n936 Vdd.t581 1.85637
R1726 Vdd.n914 Vdd.t542 1.85637
R1727 Vdd.n284 Vdd.t189 1.85637
R1728 Vdd.n952 Vdd.t557 1.85637
R1729 Vdd.n739 Vdd.t419 1.85637
R1730 Vdd.n667 Vdd.t413 1.85637
R1731 Vdd.n778 Vdd.t842 1.85637
R1732 Vdd.n395 Vdd.t429 1.85637
R1733 Vdd.n816 Vdd.t385 1.85637
R1734 Vdd.n365 Vdd.t822 1.85637
R1735 Vdd.n854 Vdd.t694 1.85637
R1736 Vdd.n329 Vdd.t878 1.85637
R1737 Vdd.n893 Vdd.t423 1.85637
R1738 Vdd.n299 Vdd.t433 1.85637
R1739 Vdd.n931 Vdd.t255 1.85637
R1740 Vdd.n269 Vdd.t19 1.85637
R1741 Vdd.n687 Vdd.t247 1.85637
R1742 Vdd.n415 Vdd.t147 1.85637
R1743 Vdd.n385 Vdd.t223 1.85637
R1744 Vdd.n355 Vdd.t161 1.85637
R1745 Vdd.n319 Vdd.t638 1.85637
R1746 Vdd.n289 Vdd.t61 1.85637
R1747 Vdd.n692 Vdd.t341 1.85637
R1748 Vdd.n708 Vdd.t616 1.85637
R1749 Vdd.n703 Vdd.t339 1.85637
R1750 Vdd.n726 Vdd.t628 1.85637
R1751 Vdd.n732 Vdd.t179 1.85637
R1752 Vdd.n720 Vdd.t365 1.85637
R1753 Vdd.n625 Vdd.t485 1.85637
R1754 Vdd.n636 Vdd.t415 1.85637
R1755 Vdd.n631 Vdd.t524 1.85637
R1756 Vdd.n648 Vdd.t329 1.85637
R1757 Vdd.n642 Vdd.t942 1.85637
R1758 Vdd.n655 Vdd.t874 1.85637
R1759 Vdd.n556 Vdd.t470 1.85637
R1760 Vdd.n567 Vdd.t916 1.85637
R1761 Vdd.n562 Vdd.t491 1.85637
R1762 Vdd.n579 Vdd.t311 1.85637
R1763 Vdd.n573 Vdd.t107 1.85637
R1764 Vdd.n586 Vdd.t441 1.85637
R1765 Vdd.n1066 Vdd.n1018 1.83762
R1766 Vdd.n1068 Vdd.n1007 1.83762
R1767 Vdd.n1050 Vdd.t463 1.8205
R1768 Vdd.n1050 Vdd.t231 1.8205
R1769 Vdd.n1048 Vdd.t233 1.8205
R1770 Vdd.n1048 Vdd.t686 1.8205
R1771 Vdd.n1046 Vdd.t650 1.8205
R1772 Vdd.n1046 Vdd.t315 1.8205
R1773 Vdd.n1044 Vdd.t229 1.8205
R1774 Vdd.n1044 Vdd.t714 1.8205
R1775 Vdd.n1042 Vdd.t716 1.8205
R1776 Vdd.n1042 Vdd.t25 1.8205
R1777 Vdd.n91 Vdd.n45 1.80479
R1778 Vdd.n164 Vdd.n29 1.80479
R1779 Vdd.n521 Vdd.n497 1.80479
R1780 Vdd.n590 Vdd.n481 1.80479
R1781 Vdd.n465 Vdd.n422 1.80479
R1782 Vdd.n221 Vdd.n13 1.80479
R1783 Vdd.n114 Vdd.n113 1.78583
R1784 Vdd.n187 Vdd.n186 1.78583
R1785 Vdd.n544 Vdd.n543 1.78583
R1786 Vdd.n613 Vdd.n612 1.78583
R1787 Vdd.n448 Vdd.n435 1.78583
R1788 Vdd.n247 Vdd.n246 1.78583
R1789 Vdd.n117 Vdd.t133 1.74654
R1790 Vdd.n190 Vdd.t758 1.74654
R1791 Vdd.n547 Vdd.t121 1.74654
R1792 Vdd.n616 Vdd.t756 1.74654
R1793 Vdd.n437 Vdd.t752 1.74654
R1794 Vdd.n255 Vdd.t131 1.74654
R1795 Vdd.n1013 Vdd.n1012 1.5755
R1796 Vdd.n1015 Vdd.n1014 1.5755
R1797 Vdd.n1011 Vdd.n1008 1.5755
R1798 Vdd.n1054 Vdd.n1053 1.5755
R1799 Vdd.n1056 Vdd.n1055 1.5755
R1800 Vdd.n15 Vdd.t658 1.49467
R1801 Vdd.n174 Vdd.t802 1.49467
R1802 Vdd.n173 Vdd.t772 1.49467
R1803 Vdd.n31 Vdd.t918 1.49467
R1804 Vdd.n101 Vdd.t69 1.49467
R1805 Vdd.n100 Vdd.t800 1.49467
R1806 Vdd.n30 Vdd.t838 1.49467
R1807 Vdd.n14 Vdd.t119 1.49467
R1808 Vdd.n239 Vdd.t79 1.49467
R1809 Vdd.n238 Vdd.t928 1.49467
R1810 Vdd.n253 Vdd.t31 1.49467
R1811 Vdd.n252 Vdd.t754 1.49467
R1812 Vdd.n467 Vdd.t27 1.49467
R1813 Vdd.n600 Vdd.t17 1.49467
R1814 Vdd.n599 Vdd.t457 1.49467
R1815 Vdd.n483 Vdd.t898 1.49467
R1816 Vdd.n531 Vdd.t195 1.49467
R1817 Vdd.n530 Vdd.t83 1.49467
R1818 Vdd.n482 Vdd.t117 1.49467
R1819 Vdd.n466 Vdd.t135 1.49467
R1820 Vdd.n459 Vdd.t111 1.49467
R1821 Vdd.n458 Vdd.t828 1.49467
R1822 Vdd.n445 Vdd.t764 1.49467
R1823 Vdd.n444 Vdd.t760 1.49467
R1824 Vdd.n167 Vdd.t750 1.47383
R1825 Vdd.n94 Vdd.t604 1.47383
R1826 Vdd.n33 Vdd.t708 1.47383
R1827 Vdd.n34 Vdd.t710 1.47383
R1828 Vdd.n35 Vdd.t940 1.47383
R1829 Vdd.n32 Vdd.t165 1.47383
R1830 Vdd.n17 Vdd.t143 1.47383
R1831 Vdd.n18 Vdd.t141 1.47383
R1832 Vdd.n19 Vdd.t205 1.47383
R1833 Vdd.n16 Vdd.t91 1.47383
R1834 Vdd.n232 Vdd.t437 1.47383
R1835 Vdd.n593 Vdd.t317 1.47383
R1836 Vdd.n524 Vdd.t896 1.47383
R1837 Vdd.n485 Vdd.t818 1.47383
R1838 Vdd.n486 Vdd.t820 1.47383
R1839 Vdd.n487 Vdd.t431 1.47383
R1840 Vdd.n484 Vdd.t93 1.47383
R1841 Vdd.n469 Vdd.t305 1.47383
R1842 Vdd.n470 Vdd.t303 1.47383
R1843 Vdd.n471 Vdd.t706 1.47383
R1844 Vdd.n468 Vdd.t381 1.47383
R1845 Vdd.n452 Vdd.t75 1.47383
R1846 Vdd.n436 Vdd.t225 1.47383
R1847 Vdd.n434 Vdd.t55 1.47383
R1848 Vdd.n424 Vdd.t53 1.47383
R1849 Vdd.n423 Vdd.t403 1.47383
R1850 Vdd.n248 Vdd.t467 1.47383
R1851 Vdd.n217 Vdd.t155 1.47383
R1852 Vdd.n218 Vdd.t157 1.47383
R1853 Vdd.n229 Vdd.t245 1.47383
R1854 Vdd.n163 Vdd.n118 1.19311
R1855 Vdd.n1079 Vdd.n191 1.19311
R1856 Vdd.n582 Vdd.n548 1.19311
R1857 Vdd.n651 Vdd.n617 1.19311
R1858 Vdd.n257 Vdd.n256 1.19311
R1859 Vdd.n1020 Vdd.t297 1.13285
R1860 Vdd.n1020 Vdd.t301 1.13285
R1861 Vdd.n1022 Vdd.t115 1.13285
R1862 Vdd.n1022 Vdd.t295 1.13285
R1863 Vdd.n1067 Vdd.n1016 1.058
R1864 Vdd.n6 Vdd.n5 1.04105
R1865 Vdd.n1095 Vdd.n1094 1.04105
R1866 Vdd.n11 Vdd.n10 1.04105
R1867 Vdd.n1083 Vdd.n1082 1.04105
R1868 Vdd.n1089 Vdd.n1088 1.04105
R1869 Vdd.n1076 Vdd.n1075 1.04105
R1870 Vdd.n53 Vdd.n52 1.04105
R1871 Vdd.n64 Vdd.n63 1.04105
R1872 Vdd.n59 Vdd.n58 1.04105
R1873 Vdd.n76 Vdd.n75 1.04105
R1874 Vdd.n70 Vdd.n69 1.04105
R1875 Vdd.n87 Vdd.n86 1.04105
R1876 Vdd.n126 Vdd.n125 1.04105
R1877 Vdd.n137 Vdd.n136 1.04105
R1878 Vdd.n132 Vdd.n131 1.04105
R1879 Vdd.n149 Vdd.n148 1.04105
R1880 Vdd.n143 Vdd.n142 1.04105
R1881 Vdd.n160 Vdd.n159 1.04105
R1882 Vdd.n206 Vdd.n205 1.04105
R1883 Vdd.n211 Vdd.n210 1.04105
R1884 Vdd.n200 Vdd.n199 1.04105
R1885 Vdd.n1001 Vdd.n1000 1.04105
R1886 Vdd.n984 Vdd.n983 1.04105
R1887 Vdd.n989 Vdd.n988 1.04105
R1888 Vdd.n995 Vdd.n994 1.04105
R1889 Vdd.n977 Vdd.n976 1.04105
R1890 Vdd.n505 Vdd.n504 1.04105
R1891 Vdd.n511 Vdd.n510 1.04105
R1892 Vdd.n517 Vdd.n516 1.04105
R1893 Vdd.n968 Vdd.n967 1.04105
R1894 Vdd.n754 Vdd.n753 1.04105
R1895 Vdd.n793 Vdd.n792 1.04105
R1896 Vdd.n831 Vdd.n830 1.04105
R1897 Vdd.n869 Vdd.n868 1.04105
R1898 Vdd.n908 Vdd.n907 1.04105
R1899 Vdd.n946 Vdd.n945 1.04105
R1900 Vdd.n672 Vdd.n671 1.04105
R1901 Vdd.n765 Vdd.n764 1.04105
R1902 Vdd.n400 Vdd.n399 1.04105
R1903 Vdd.n804 Vdd.n803 1.04105
R1904 Vdd.n370 Vdd.n369 1.04105
R1905 Vdd.n842 Vdd.n841 1.04105
R1906 Vdd.n340 Vdd.n339 1.04105
R1907 Vdd.n881 Vdd.n880 1.04105
R1908 Vdd.n304 Vdd.n303 1.04105
R1909 Vdd.n919 Vdd.n918 1.04105
R1910 Vdd.n274 Vdd.n273 1.04105
R1911 Vdd.n957 Vdd.n956 1.04105
R1912 Vdd.n749 Vdd.n748 1.04105
R1913 Vdd.n662 Vdd.n661 1.04105
R1914 Vdd.n788 Vdd.n787 1.04105
R1915 Vdd.n390 Vdd.n389 1.04105
R1916 Vdd.n826 Vdd.n825 1.04105
R1917 Vdd.n360 Vdd.n359 1.04105
R1918 Vdd.n864 Vdd.n863 1.04105
R1919 Vdd.n324 Vdd.n323 1.04105
R1920 Vdd.n903 Vdd.n902 1.04105
R1921 Vdd.n294 Vdd.n293 1.04105
R1922 Vdd.n941 Vdd.n940 1.04105
R1923 Vdd.n264 Vdd.n263 1.04105
R1924 Vdd.n677 Vdd.n676 1.04105
R1925 Vdd.n405 Vdd.n404 1.04105
R1926 Vdd.n375 Vdd.n374 1.04105
R1927 Vdd.n345 Vdd.n344 1.04105
R1928 Vdd.n309 Vdd.n308 1.04105
R1929 Vdd.n279 Vdd.n278 1.04105
R1930 Vdd.n744 Vdd.n743 1.04105
R1931 Vdd.n682 Vdd.n681 1.04105
R1932 Vdd.n783 Vdd.n782 1.04105
R1933 Vdd.n760 Vdd.n759 1.04105
R1934 Vdd.n410 Vdd.n409 1.04105
R1935 Vdd.n821 Vdd.n820 1.04105
R1936 Vdd.n799 Vdd.n798 1.04105
R1937 Vdd.n380 Vdd.n379 1.04105
R1938 Vdd.n859 Vdd.n858 1.04105
R1939 Vdd.n837 Vdd.n836 1.04105
R1940 Vdd.n350 Vdd.n349 1.04105
R1941 Vdd.n898 Vdd.n897 1.04105
R1942 Vdd.n876 Vdd.n875 1.04105
R1943 Vdd.n314 Vdd.n313 1.04105
R1944 Vdd.n936 Vdd.n935 1.04105
R1945 Vdd.n914 Vdd.n913 1.04105
R1946 Vdd.n284 Vdd.n283 1.04105
R1947 Vdd.n952 Vdd.n951 1.04105
R1948 Vdd.n739 Vdd.n738 1.04105
R1949 Vdd.n667 Vdd.n666 1.04105
R1950 Vdd.n778 Vdd.n777 1.04105
R1951 Vdd.n395 Vdd.n394 1.04105
R1952 Vdd.n816 Vdd.n815 1.04105
R1953 Vdd.n365 Vdd.n364 1.04105
R1954 Vdd.n854 Vdd.n853 1.04105
R1955 Vdd.n329 Vdd.n328 1.04105
R1956 Vdd.n893 Vdd.n892 1.04105
R1957 Vdd.n299 Vdd.n298 1.04105
R1958 Vdd.n931 Vdd.n930 1.04105
R1959 Vdd.n269 Vdd.n268 1.04105
R1960 Vdd.n687 Vdd.n686 1.04105
R1961 Vdd.n415 Vdd.n414 1.04105
R1962 Vdd.n385 Vdd.n384 1.04105
R1963 Vdd.n355 Vdd.n354 1.04105
R1964 Vdd.n319 Vdd.n318 1.04105
R1965 Vdd.n289 Vdd.n288 1.04105
R1966 Vdd.n692 Vdd.n691 1.04105
R1967 Vdd.n708 Vdd.n707 1.04105
R1968 Vdd.n703 Vdd.n702 1.04105
R1969 Vdd.n726 Vdd.n725 1.04105
R1970 Vdd.n732 Vdd.n731 1.04105
R1971 Vdd.n720 Vdd.n719 1.04105
R1972 Vdd.n625 Vdd.n624 1.04105
R1973 Vdd.n636 Vdd.n635 1.04105
R1974 Vdd.n631 Vdd.n630 1.04105
R1975 Vdd.n648 Vdd.n647 1.04105
R1976 Vdd.n642 Vdd.n641 1.04105
R1977 Vdd.n655 Vdd.n654 1.04105
R1978 Vdd.n556 Vdd.n555 1.04105
R1979 Vdd.n567 Vdd.n566 1.04105
R1980 Vdd.n562 Vdd.n561 1.04105
R1981 Vdd.n579 Vdd.n578 1.04105
R1982 Vdd.n573 Vdd.n572 1.04105
R1983 Vdd.n586 Vdd.n585 1.04105
R1984 Vdd.n1016 Vdd.n1008 1.01373
R1985 Vdd.n1016 Vdd.n1015 0.979984
R1986 Vdd.n91 Vdd.n90 0.809622
R1987 Vdd.n164 Vdd.n163 0.809622
R1988 Vdd.n521 Vdd.n520 0.809622
R1989 Vdd.n590 Vdd.n589 0.809622
R1990 Vdd.n651 Vdd.n465 0.809622
R1991 Vdd.n1079 Vdd.n13 0.809622
R1992 Vdd.n170 Vdd.n167 0.788
R1993 Vdd.n171 Vdd.n170 0.788
R1994 Vdd.n173 Vdd.n172 0.788
R1995 Vdd.n97 Vdd.n94 0.788
R1996 Vdd.n98 Vdd.n97 0.788
R1997 Vdd.n100 Vdd.n99 0.788
R1998 Vdd.n41 Vdd.n34 0.788
R1999 Vdd.n42 Vdd.n41 0.788
R2000 Vdd.n43 Vdd.n35 0.788
R2001 Vdd.n44 Vdd.n43 0.788
R2002 Vdd.n39 Vdd.n33 0.788
R2003 Vdd.n111 Vdd.n32 0.788
R2004 Vdd.n112 Vdd.n111 0.788
R2005 Vdd.n110 Vdd.n30 0.788
R2006 Vdd.n25 Vdd.n18 0.788
R2007 Vdd.n26 Vdd.n25 0.788
R2008 Vdd.n27 Vdd.n19 0.788
R2009 Vdd.n28 Vdd.n27 0.788
R2010 Vdd.n23 Vdd.n17 0.788
R2011 Vdd.n184 Vdd.n16 0.788
R2012 Vdd.n185 Vdd.n184 0.788
R2013 Vdd.n183 Vdd.n14 0.788
R2014 Vdd.n235 Vdd.n232 0.788
R2015 Vdd.n236 Vdd.n235 0.788
R2016 Vdd.n238 Vdd.n237 0.788
R2017 Vdd.n596 Vdd.n593 0.788
R2018 Vdd.n597 Vdd.n596 0.788
R2019 Vdd.n599 Vdd.n598 0.788
R2020 Vdd.n527 Vdd.n524 0.788
R2021 Vdd.n528 Vdd.n527 0.788
R2022 Vdd.n530 Vdd.n529 0.788
R2023 Vdd.n493 Vdd.n486 0.788
R2024 Vdd.n494 Vdd.n493 0.788
R2025 Vdd.n495 Vdd.n487 0.788
R2026 Vdd.n496 Vdd.n495 0.788
R2027 Vdd.n491 Vdd.n485 0.788
R2028 Vdd.n541 Vdd.n484 0.788
R2029 Vdd.n542 Vdd.n541 0.788
R2030 Vdd.n540 Vdd.n482 0.788
R2031 Vdd.n477 Vdd.n470 0.788
R2032 Vdd.n478 Vdd.n477 0.788
R2033 Vdd.n479 Vdd.n471 0.788
R2034 Vdd.n480 Vdd.n479 0.788
R2035 Vdd.n475 Vdd.n469 0.788
R2036 Vdd.n610 Vdd.n468 0.788
R2037 Vdd.n611 Vdd.n610 0.788
R2038 Vdd.n609 Vdd.n466 0.788
R2039 Vdd.n455 Vdd.n452 0.788
R2040 Vdd.n456 Vdd.n455 0.788
R2041 Vdd.n458 Vdd.n457 0.788
R2042 Vdd.n441 Vdd.n436 0.788
R2043 Vdd.n442 Vdd.n441 0.788
R2044 Vdd.n444 Vdd.n443 0.788
R2045 Vdd.n431 Vdd.n424 0.788
R2046 Vdd.n432 Vdd.n431 0.788
R2047 Vdd.n429 Vdd.n423 0.788
R2048 Vdd.n430 Vdd.n429 0.788
R2049 Vdd.n434 Vdd.n433 0.788
R2050 Vdd.n249 Vdd.n248 0.788
R2051 Vdd.n250 Vdd.n249 0.788
R2052 Vdd.n252 Vdd.n251 0.788
R2053 Vdd.n225 Vdd.n218 0.788
R2054 Vdd.n226 Vdd.n225 0.788
R2055 Vdd.n229 Vdd.n228 0.788
R2056 Vdd.n228 Vdd.n227 0.788
R2057 Vdd.n223 Vdd.n217 0.788
R2058 Vdd.n49 Vdd.n48 0.754571
R2059 Vdd.n122 Vdd.n121 0.754571
R2060 Vdd.n501 Vdd.n500 0.754571
R2061 Vdd.n552 Vdd.n551 0.754571
R2062 Vdd.n621 Vdd.n620 0.754571
R2063 Vdd.n1099 Vdd.n2 0.754571
R2064 Vdd.n1065 Vdd.n1030 0.750875
R2065 Vdd.n3 Vdd.t191 0.7285
R2066 Vdd.n3 Vdd.t934 0.7285
R2067 Vdd.n1092 Vdd.t405 0.7285
R2068 Vdd.n1092 Vdd.t530 0.7285
R2069 Vdd.n8 Vdd.t269 0.7285
R2070 Vdd.n8 Vdd.t193 0.7285
R2071 Vdd.n1080 Vdd.t287 0.7285
R2072 Vdd.n1080 Vdd.t644 0.7285
R2073 Vdd.n1086 Vdd.t533 0.7285
R2074 Vdd.n1086 Vdd.t101 0.7285
R2075 Vdd.n1073 Vdd.t97 0.7285
R2076 Vdd.n1073 Vdd.t569 0.7285
R2077 Vdd.n50 Vdd.t281 0.7285
R2078 Vdd.n50 Vdd.t846 0.7285
R2079 Vdd.n61 Vdd.t612 0.7285
R2080 Vdd.n61 Vdd.t473 0.7285
R2081 Vdd.n56 Vdd.t321 0.7285
R2082 Vdd.n56 Vdd.t283 0.7285
R2083 Vdd.n73 Vdd.t836 0.7285
R2084 Vdd.n73 Vdd.t648 0.7285
R2085 Vdd.n67 Vdd.t515 0.7285
R2086 Vdd.n67 Vdd.t409 0.7285
R2087 Vdd.n84 Vdd.t427 0.7285
R2088 Vdd.n84 Vdd.t509 0.7285
R2089 Vdd.n123 Vdd.t237 0.7285
R2090 Vdd.n123 Vdd.t886 0.7285
R2091 Vdd.n134 Vdd.t642 0.7285
R2092 Vdd.n134 Vdd.t596 0.7285
R2093 Vdd.n129 Vdd.t938 0.7285
R2094 Vdd.n129 Vdd.t239 0.7285
R2095 Vdd.n146 Vdd.t890 0.7285
R2096 Vdd.n146 Vdd.t445 0.7285
R2097 Vdd.n140 Vdd.t602 0.7285
R2098 Vdd.n140 Vdd.t263 0.7285
R2099 Vdd.n157 Vdd.t13 0.7285
R2100 Vdd.n157 Vdd.t494 0.7285
R2101 Vdd.n203 Vdd.t461 0.7285
R2102 Vdd.n203 Vdd.t882 0.7285
R2103 Vdd.n208 Vdd.t518 0.7285
R2104 Vdd.n208 Vdd.t816 0.7285
R2105 Vdd.n197 Vdd.t866 0.7285
R2106 Vdd.n197 Vdd.t23 0.7285
R2107 Vdd.n998 Vdd.t770 0.7285
R2108 Vdd.n998 Vdd.t806 0.7285
R2109 Vdd.n981 Vdd.t159 0.7285
R2110 Vdd.n981 Vdd.t870 0.7285
R2111 Vdd.n986 Vdd.t21 0.7285
R2112 Vdd.n986 Vdd.t766 0.7285
R2113 Vdd.n992 Vdd.t744 0.7285
R2114 Vdd.n992 Vdd.t95 0.7285
R2115 Vdd.n974 Vdd.t762 0.7285
R2116 Vdd.n974 Vdd.t810 0.7285
R2117 Vdd.n502 Vdd.t852 0.7285
R2118 Vdd.n502 Vdd.t105 0.7285
R2119 Vdd.n508 Vdd.t636 0.7285
R2120 Vdd.n508 Vdd.t512 0.7285
R2121 Vdd.n514 Vdd.t936 0.7285
R2122 Vdd.n514 Vdd.t407 0.7285
R2123 Vdd.n965 Vdd.t451 0.7285
R2124 Vdd.n965 Vdd.t554 0.7285
R2125 Vdd.n751 Vdd.t776 0.7285
R2126 Vdd.n751 Vdd.t784 0.7285
R2127 Vdd.n790 Vdd.t57 0.7285
R2128 Vdd.n790 Vdd.t71 0.7285
R2129 Vdd.n828 Vdd.t219 0.7285
R2130 Vdd.n828 Vdd.t7 0.7285
R2131 Vdd.n866 Vdd.t902 0.7285
R2132 Vdd.n866 Vdd.t606 0.7285
R2133 Vdd.n905 Vdd.t371 0.7285
R2134 Vdd.n905 Vdd.t251 0.7285
R2135 Vdd.n943 Vdd.t203 0.7285
R2136 Vdd.n943 Vdd.t171 0.7285
R2137 Vdd.n669 Vdd.t459 0.7285
R2138 Vdd.n669 Vdd.t393 0.7285
R2139 Vdd.n762 Vdd.t279 0.7285
R2140 Vdd.n762 Vdd.t774 0.7285
R2141 Vdd.n397 Vdd.t85 0.7285
R2142 Vdd.n397 Vdd.t674 0.7285
R2143 Vdd.n801 Vdd.t888 0.7285
R2144 Vdd.n801 Vdd.t151 0.7285
R2145 Vdd.n367 Vdd.t926 0.7285
R2146 Vdd.n367 Vdd.t808 0.7285
R2147 Vdd.n839 Vdd.t77 0.7285
R2148 Vdd.n839 Vdd.t221 0.7285
R2149 Vdd.n337 Vdd.t684 0.7285
R2150 Vdd.n337 Vdd.t349 0.7285
R2151 Vdd.n878 Vdd.t129 0.7285
R2152 Vdd.n878 Vdd.t904 0.7285
R2153 Vdd.n301 Vdd.t796 0.7285
R2154 Vdd.n301 Vdd.t666 0.7285
R2155 Vdd.n916 Vdd.t435 0.7285
R2156 Vdd.n916 Vdd.t199 0.7285
R2157 Vdd.n271 Vdd.t792 0.7285
R2158 Vdd.n271 Vdd.t333 0.7285
R2159 Vdd.n954 Vdd.t169 0.7285
R2160 Vdd.n954 Vdd.t375 0.7285
R2161 Vdd.n746 Vdd.t782 0.7285
R2162 Vdd.n746 Vdd.t127 0.7285
R2163 Vdd.n659 Vdd.t670 0.7285
R2164 Vdd.n659 Vdd.t786 0.7285
R2165 Vdd.n785 Vdd.t73 0.7285
R2166 Vdd.n785 Vdd.t89 0.7285
R2167 Vdd.n387 Vdd.t357 0.7285
R2168 Vdd.n387 Vdd.t906 0.7285
R2169 Vdd.n823 Vdd.t5 0.7285
R2170 Vdd.n823 Vdd.t922 0.7285
R2171 Vdd.n357 Vdd.t854 0.7285
R2172 Vdd.n357 Vdd.t325 0.7285
R2173 Vdd.n861 Vdd.t608 0.7285
R2174 Vdd.n861 Vdd.t680 0.7285
R2175 Vdd.n321 Vdd.t359 0.7285
R2176 Vdd.n321 Vdd.t209 0.7285
R2177 Vdd.n900 Vdd.t253 0.7285
R2178 Vdd.n900 Vdd.t391 0.7285
R2179 Vdd.n291 Vdd.t740 0.7285
R2180 Vdd.n291 Vdd.t848 0.7285
R2181 Vdd.n938 Vdd.t173 0.7285
R2182 Vdd.n938 Vdd.t790 0.7285
R2183 Vdd.n261 Vdd.t345 0.7285
R2184 Vdd.n261 Vdd.t780 0.7285
R2185 Vdd.n674 Vdd.t327 0.7285
R2186 Vdd.n674 Vdd.t860 0.7285
R2187 Vdd.n402 Vdd.t383 0.7285
R2188 Vdd.n402 Vdd.t742 0.7285
R2189 Vdd.n372 Vdd.t277 0.7285
R2190 Vdd.n372 Vdd.t678 0.7285
R2191 Vdd.n342 Vdd.t379 0.7285
R2192 Vdd.n342 Vdd.t355 0.7285
R2193 Vdd.n306 Vdd.t275 0.7285
R2194 Vdd.n306 Vdd.t864 0.7285
R2195 Vdd.n276 Vdd.t377 0.7285
R2196 Vdd.n276 Vdd.t662 0.7285
R2197 Vdd.n741 Vdd.t421 0.7285
R2198 Vdd.n741 Vdd.t894 0.7285
R2199 Vdd.n679 Vdd.t726 0.7285
R2200 Vdd.n679 Vdd.t676 0.7285
R2201 Vdd.n780 Vdd.t844 0.7285
R2202 Vdd.n780 Vdd.t397 0.7285
R2203 Vdd.n757 Vdd.t45 0.7285
R2204 Vdd.n757 Vdd.t207 0.7285
R2205 Vdd.n407 Vdd.t724 0.7285
R2206 Vdd.n407 Vdd.t353 0.7285
R2207 Vdd.n818 Vdd.t389 0.7285
R2208 Vdd.n818 Vdd.t634 0.7285
R2209 Vdd.n796 Vdd.t49 0.7285
R2210 Vdd.n796 Vdd.t840 0.7285
R2211 Vdd.n377 Vdd.t698 0.7285
R2212 Vdd.n377 Vdd.t361 0.7285
R2213 Vdd.n856 Vdd.t832 0.7285
R2214 Vdd.n856 Vdd.t65 0.7285
R2215 Vdd.n834 Vdd.t812 0.7285
R2216 Vdd.n834 Vdd.t387 0.7285
R2217 Vdd.n347 Vdd.t702 0.7285
R2218 Vdd.n347 Vdd.t664 0.7285
R2219 Vdd.n895 Vdd.t425 0.7285
R2220 Vdd.n895 Vdd.t712 0.7285
R2221 Vdd.n873 Vdd.t215 0.7285
R2222 Vdd.n873 Vdd.t834 0.7285
R2223 Vdd.n311 Vdd.t734 0.7285
R2224 Vdd.n311 Vdd.t668 0.7285
R2225 Vdd.n933 Vdd.t167 0.7285
R2226 Vdd.n933 Vdd.t3 0.7285
R2227 Vdd.n911 Vdd.t910 0.7285
R2228 Vdd.n911 Vdd.t618 0.7285
R2229 Vdd.n281 Vdd.t690 0.7285
R2230 Vdd.n281 Vdd.t804 0.7285
R2231 Vdd.n949 Vdd.t39 0.7285
R2232 Vdd.n949 Vdd.t257 0.7285
R2233 Vdd.n736 Vdd.t892 0.7285
R2234 Vdd.n736 Vdd.t730 0.7285
R2235 Vdd.n664 Vdd.t363 0.7285
R2236 Vdd.n664 Vdd.t249 0.7285
R2237 Vdd.n775 Vdd.t620 0.7285
R2238 Vdd.n775 Vdd.t718 0.7285
R2239 Vdd.n392 Vdd.t862 0.7285
R2240 Vdd.n392 Vdd.t145 0.7285
R2241 Vdd.n813 Vdd.t453 0.7285
R2242 Vdd.n813 Vdd.t700 0.7285
R2243 Vdd.n362 Vdd.t347 0.7285
R2244 Vdd.n362 Vdd.t197 0.7285
R2245 Vdd.n851 Vdd.t63 0.7285
R2246 Vdd.n851 Vdd.t692 0.7285
R2247 Vdd.n326 Vdd.t335 0.7285
R2248 Vdd.n326 Vdd.t163 0.7285
R2249 Vdd.n890 Vdd.t401 0.7285
R2250 Vdd.n890 Vdd.t728 0.7285
R2251 Vdd.n296 Vdd.t343 0.7285
R2252 Vdd.n296 Vdd.t640 0.7285
R2253 Vdd.n928 Vdd.t35 0.7285
R2254 Vdd.n928 Vdd.t704 0.7285
R2255 Vdd.n266 Vdd.t858 0.7285
R2256 Vdd.n266 Vdd.t59 0.7285
R2257 Vdd.n684 Vdd.t181 0.7285
R2258 Vdd.n684 Vdd.t672 0.7285
R2259 Vdd.n412 Vdd.t465 0.7285
R2260 Vdd.n412 Vdd.t351 0.7285
R2261 Vdd.n382 Vdd.t455 0.7285
R2262 Vdd.n382 Vdd.t660 0.7285
R2263 Vdd.n352 Vdd.t399 0.7285
R2264 Vdd.n352 Vdd.t856 0.7285
R2265 Vdd.n316 Vdd.t876 0.7285
R2266 Vdd.n316 Vdd.t738 0.7285
R2267 Vdd.n286 Vdd.t439 0.7285
R2268 Vdd.n286 Vdd.t337 0.7285
R2269 Vdd.n689 Vdd.t630 0.7285
R2270 Vdd.n689 Vdd.t139 0.7285
R2271 Vdd.n705 Vdd.t722 0.7285
R2272 Vdd.n705 Vdd.t488 0.7285
R2273 Vdd.n700 Vdd.t185 0.7285
R2274 Vdd.n700 Vdd.t622 0.7285
R2275 Vdd.n723 Vdd.t137 0.7285
R2276 Vdd.n723 Vdd.t688 0.7285
R2277 Vdd.n729 Vdd.t590 0.7285
R2278 Vdd.n729 Vdd.t632 0.7285
R2279 Vdd.n717 Vdd.t768 0.7285
R2280 Vdd.n717 Vdd.t584 0.7285
R2281 Vdd.n622 Vdd.t183 0.7285
R2282 Vdd.n622 Vdd.t626 0.7285
R2283 Vdd.n633 Vdd.t610 0.7285
R2284 Vdd.n633 Vdd.t503 0.7285
R2285 Vdd.n628 Vdd.t81 0.7285
R2286 Vdd.n628 Vdd.t331 0.7285
R2287 Vdd.n645 Vdd.t624 0.7285
R2288 Vdd.n645 Vdd.t417 0.7285
R2289 Vdd.n639 Vdd.t599 0.7285
R2290 Vdd.n639 Vdd.t293 0.7285
R2291 Vdd.n652 Vdd.t614 0.7285
R2292 Vdd.n652 Vdd.t548 0.7285
R2293 Vdd.n553 Vdd.t307 0.7285
R2294 Vdd.n553 Vdd.t826 0.7285
R2295 Vdd.n564 Vdd.t447 0.7285
R2296 Vdd.n564 Vdd.t506 0.7285
R2297 Vdd.n559 Vdd.t15 0.7285
R2298 Vdd.n559 Vdd.t309 0.7285
R2299 Vdd.n576 Vdd.t824 0.7285
R2300 Vdd.n576 Vdd.t646 0.7285
R2301 Vdd.n570 Vdd.t500 0.7285
R2302 Vdd.n570 Vdd.t443 0.7285
R2303 Vdd.n583 Vdd.t9 0.7285
R2304 Vdd.n583 Vdd.t551 0.7285
R2305 Vdd.n773 SARlogic_0.dffrs_1.nand3_0.C 0.717607
R2306 Vdd.n811 SARlogic_0.dffrs_2.nand3_0.C 0.717607
R2307 Vdd.n849 SARlogic_0.dffrs_3.nand3_0.C 0.717607
R2308 Vdd.n888 SARlogic_0.dffrs_4.nand3_0.C 0.717607
R2309 Vdd.n926 SARlogic_0.dffrs_5.nand3_0.C 0.717607
R2310 Vdd.n698 SARlogic_0.dffrs_0.nand3_0.C 0.717607
R2311 Vdd.n1045 Vdd.n1043 0.667
R2312 Vdd.n1051 Vdd.n1049 0.662
R2313 Vdd.n1047 Vdd.n1045 0.643429
R2314 Vdd.n1049 Vdd.n1047 0.638429
R2315 Vdd.n1060 Vdd.n1059 0.58325
R2316 Vdd.n1041 Vdd.n1038 0.58325
R2317 Vdd.n176 Vdd.n167 0.561043
R2318 Vdd.n103 Vdd.n94 0.561043
R2319 Vdd.n107 Vdd.n33 0.561043
R2320 Vdd.n106 Vdd.n34 0.561043
R2321 Vdd.n92 Vdd.n35 0.561043
R2322 Vdd.n115 Vdd.n32 0.561043
R2323 Vdd.n180 Vdd.n17 0.561043
R2324 Vdd.n179 Vdd.n18 0.561043
R2325 Vdd.n165 Vdd.n19 0.561043
R2326 Vdd.n188 Vdd.n16 0.561043
R2327 Vdd.n241 Vdd.n232 0.561043
R2328 Vdd.n602 Vdd.n593 0.561043
R2329 Vdd.n533 Vdd.n524 0.561043
R2330 Vdd.n537 Vdd.n485 0.561043
R2331 Vdd.n536 Vdd.n486 0.561043
R2332 Vdd.n522 Vdd.n487 0.561043
R2333 Vdd.n545 Vdd.n484 0.561043
R2334 Vdd.n606 Vdd.n469 0.561043
R2335 Vdd.n605 Vdd.n470 0.561043
R2336 Vdd.n591 Vdd.n471 0.561043
R2337 Vdd.n614 Vdd.n468 0.561043
R2338 Vdd.n461 Vdd.n452 0.561043
R2339 Vdd.n447 Vdd.n436 0.561043
R2340 Vdd.n449 Vdd.n434 0.561043
R2341 Vdd.n450 Vdd.n424 0.561043
R2342 Vdd.n464 Vdd.n423 0.561043
R2343 Vdd.n248 Vdd.n214 0.561043
R2344 Vdd.n245 Vdd.n217 0.561043
R2345 Vdd.n244 Vdd.n218 0.561043
R2346 Vdd.n230 Vdd.n229 0.561043
R2347 Vdd.n438 Vdd.n437 0.510024
R2348 Vdd.n118 Vdd.n116 0.490037
R2349 Vdd.n191 Vdd.n189 0.490037
R2350 Vdd.n548 Vdd.n546 0.490037
R2351 Vdd.n617 Vdd.n615 0.490037
R2352 Vdd.n256 Vdd.n254 0.490037
R2353 Vdd.n1043 Vdd.n1031 0.47525
R2354 Vdd.n1052 Vdd.n1051 0.47525
R2355 Vdd.n118 Vdd.n117 0.436534
R2356 Vdd.n191 Vdd.n190 0.436534
R2357 Vdd.n548 Vdd.n547 0.436534
R2358 Vdd.n617 Vdd.n616 0.436534
R2359 Vdd.n256 Vdd.n255 0.436534
R2360 Vdd.n446 Vdd.n438 0.415037
R2361 Vdd.n756 Vdd.n735 0.403945
R2362 Vdd.n1065 Vdd.n1064 0.381816
R2363 Vdd.n1063 Vdd.n1060 0.34025
R2364 Vdd.n1059 Vdd.n1031 0.34025
R2365 Vdd.n1052 Vdd.n1041 0.34025
R2366 Vdd.n1069 Vdd.n1068 0.313132
R2367 Vdd.n1068 Vdd.n1067 0.289447
R2368 Vdd.n1067 Vdd.n1066 0.279974
R2369 Vdd.n1071 Vdd.n1070 0.265225
R2370 Vdd.n1066 Vdd.n1065 0.256289
R2371 Vdd.n176 Vdd.n175 0.255737
R2372 Vdd.n103 Vdd.n102 0.255737
R2373 Vdd.n116 Vdd.n115 0.255737
R2374 Vdd.n189 Vdd.n188 0.255737
R2375 Vdd.n241 Vdd.n240 0.255737
R2376 Vdd.n602 Vdd.n601 0.255737
R2377 Vdd.n533 Vdd.n532 0.255737
R2378 Vdd.n546 Vdd.n545 0.255737
R2379 Vdd.n615 Vdd.n614 0.255737
R2380 Vdd.n461 Vdd.n460 0.255737
R2381 Vdd.n447 Vdd.n446 0.255737
R2382 Vdd.n254 Vdd.n214 0.255737
R2383 Vdd.n258 Vdd.n202 0.236406
R2384 Vdd.n115 Vdd.n114 0.2165
R2385 Vdd.n188 Vdd.n187 0.2165
R2386 Vdd.n545 Vdd.n544 0.2165
R2387 Vdd.n614 Vdd.n613 0.2165
R2388 Vdd.n448 Vdd.n447 0.2165
R2389 Vdd.n246 Vdd.n214 0.2165
R2390 Vdd.n1017 comparator_no_offsetcal_0.x3.avdd 0.207699
R2391 Vdd.n972 Vdd.n971 0.165959
R2392 Vdd.n1070 Vdd 0.162037
R2393 Vdd.n114 Vdd.n107 0.148424
R2394 Vdd.n187 Vdd.n180 0.148424
R2395 Vdd.n544 Vdd.n537 0.148424
R2396 Vdd.n613 Vdd.n606 0.148424
R2397 Vdd.n449 Vdd.n448 0.148424
R2398 Vdd.n246 Vdd.n245 0.148424
R2399 adc_PISO_0.dffrs_3.resetb Vdd.n196 0.136036
R2400 adc_PISO_0.dffrs_5.resetb Vdd.n83 0.136036
R2401 adc_PISO_0.dffrs_4.resetb Vdd.n156 0.136036
R2402 adc_PISO_0.dffrs_2.resetb Vdd.n964 0.136036
R2403 SARlogic_0.dffrs_13.resetb Vdd.n716 0.136036
R2404 adc_PISO_0.dffrs_0.resetb Vdd.n421 0.136036
R2405 adc_PISO_0.dffrs_1.resetb Vdd.n335 0.136036
R2406 Vdd.n1026 Vdd.n1021 0.1355
R2407 Vdd.n1024 Vdd.n1023 0.109786
R2408 Vdd.n1030 Vdd.n1019 0.103357
R2409 Vdd.n519 Vdd.n513 0.101647
R2410 Vdd.n1071 Vdd.n1005 0.0967961
R2411 Vdd.n1018 Vdd.n1017 0.0965492
R2412 Vdd.n1064 comparator_no_offsetcal_0.VDD 0.0942895
R2413 Vdd.n971 Vdd.n970 0.0898578
R2414 Vdd.n973 Vdd.n259 0.0817571
R2415 Vdd.n520 Vdd.n519 0.0720596
R2416 Vdd.n1072 Vdd.n1071 0.0680047
R2417 Vdd.n872 Vdd.n336 0.0660636
R2418 Vdd.n177 Vdd.n176 0.0635
R2419 Vdd.n104 Vdd.n103 0.0635
R2420 Vdd.n242 Vdd.n241 0.0635
R2421 Vdd.n603 Vdd.n602 0.0635
R2422 Vdd.n534 Vdd.n533 0.0635
R2423 Vdd.n462 Vdd.n461 0.0635
R2424 Vdd.n257 Vdd.n213 0.0597785
R2425 Vdd.n513 Vdd.n507 0.0590321
R2426 Vdd.n1030 Vdd.n1029 0.0519286
R2427 Vdd.n1023 Vdd.n1019 0.0455
R2428 Vdd.n770 SARlogic_0.dffrs_1.nand3_2.C 0.0455
R2429 Vdd.n808 SARlogic_0.dffrs_2.nand3_2.C 0.0455
R2430 Vdd.n846 SARlogic_0.dffrs_3.nand3_2.C 0.0455
R2431 Vdd.n885 SARlogic_0.dffrs_4.nand3_2.C 0.0455
R2432 Vdd.n923 SARlogic_0.dffrs_5.nand3_2.C 0.0455
R2433 Vdd.n695 SARlogic_0.dffrs_0.nand3_2.C 0.0455
R2434 Vdd.n712 SARlogic_0.dffrs_13.nand3_7.A 0.0455
R2435 Vdd.n107 Vdd.n106 0.0452384
R2436 Vdd.n180 Vdd.n179 0.0452384
R2437 Vdd.n537 Vdd.n536 0.0452384
R2438 Vdd.n606 Vdd.n605 0.0452384
R2439 Vdd.n450 Vdd.n449 0.0452384
R2440 Vdd.n245 Vdd.n244 0.0452384
R2441 Vdd.n72 Vdd.n66 0.0405727
R2442 Vdd.n145 Vdd.n139 0.0405727
R2443 Vdd.n575 Vdd.n569 0.0405727
R2444 Vdd.n644 Vdd.n638 0.0405727
R2445 Vdd.n1097 Vdd.n1091 0.0405727
R2446 SARlogic_0.dffrs_1.nand3_0.C Vdd.n772 0.0374643
R2447 SARlogic_0.dffrs_2.nand3_0.C Vdd.n810 0.0374643
R2448 SARlogic_0.dffrs_3.nand3_0.C Vdd.n848 0.0374643
R2449 SARlogic_0.dffrs_4.nand3_0.C Vdd.n887 0.0374643
R2450 SARlogic_0.dffrs_5.nand3_0.C Vdd.n925 0.0374643
R2451 SARlogic_0.dffrs_0.nand3_0.C Vdd.n697 0.0374643
R2452 Vdd.n1003 Vdd.n997 0.0373206
R2453 Vdd.n588 Vdd.n336 0.0359182
R2454 Vdd.n658 Vdd.n657 0.0359182
R2455 Vdd.n1078 Vdd.n1072 0.0359182
R2456 Vdd.n728 Vdd.n722 0.0339767
R2457 Vdd.n49 adc_PISO_0.dffrs_5.setb 0.032
R2458 Vdd.n122 adc_PISO_0.dffrs_4.setb 0.032
R2459 Vdd.n501 adc_PISO_0.dffrs_2.setb 0.032
R2460 Vdd.n773 SARlogic_0.dffrs_1.setb 0.032
R2461 Vdd.n811 SARlogic_0.dffrs_2.setb 0.032
R2462 Vdd.n849 SARlogic_0.dffrs_3.setb 0.032
R2463 Vdd.n888 SARlogic_0.dffrs_4.setb 0.032
R2464 Vdd.n926 SARlogic_0.dffrs_5.setb 0.032
R2465 Vdd.n698 SARlogic_0.dffrs_0.setb 0.032
R2466 Vdd.n552 adc_PISO_0.dffrs_1.setb 0.032
R2467 Vdd.n621 adc_PISO_0.dffrs_0.setb 0.032
R2468 adc_PISO_0.dffrs_3.setb Vdd.n1099 0.032
R2469 Vdd.n735 Vdd.n710 0.0316083
R2470 Vdd.n175 Vdd.n173 0.0313054
R2471 Vdd.n175 Vdd.n174 0.0313054
R2472 Vdd.n102 Vdd.n100 0.0313054
R2473 Vdd.n102 Vdd.n101 0.0313054
R2474 Vdd.n116 Vdd.n30 0.0313054
R2475 Vdd.n116 Vdd.n31 0.0313054
R2476 Vdd.n189 Vdd.n14 0.0313054
R2477 Vdd.n189 Vdd.n15 0.0313054
R2478 Vdd.n240 Vdd.n238 0.0313054
R2479 Vdd.n240 Vdd.n239 0.0313054
R2480 Vdd.n601 Vdd.n599 0.0313054
R2481 Vdd.n601 Vdd.n600 0.0313054
R2482 Vdd.n532 Vdd.n530 0.0313054
R2483 Vdd.n532 Vdd.n531 0.0313054
R2484 Vdd.n546 Vdd.n482 0.0313054
R2485 Vdd.n546 Vdd.n483 0.0313054
R2486 Vdd.n615 Vdd.n466 0.0313054
R2487 Vdd.n615 Vdd.n467 0.0313054
R2488 Vdd.n460 Vdd.n458 0.0313054
R2489 Vdd.n460 Vdd.n459 0.0313054
R2490 Vdd.n446 Vdd.n444 0.0313054
R2491 Vdd.n446 Vdd.n445 0.0313054
R2492 Vdd.n254 Vdd.n252 0.0313054
R2493 Vdd.n254 Vdd.n253 0.0313054
R2494 Vdd.n105 Vdd.n92 0.0295407
R2495 Vdd.n178 Vdd.n165 0.0295407
R2496 Vdd.n535 Vdd.n522 0.0295407
R2497 Vdd.n604 Vdd.n591 0.0295407
R2498 Vdd.n464 Vdd.n463 0.0295407
R2499 Vdd.n243 Vdd.n230 0.0295407
R2500 Vdd.n90 Vdd.n78 0.0288636
R2501 Vdd.n163 Vdd.n151 0.0288636
R2502 Vdd.n651 Vdd.n650 0.0288636
R2503 Vdd.n1085 Vdd.n1079 0.0288636
R2504 Vdd.n582 Vdd.n581 0.0288455
R2505 Vdd.n991 Vdd.n980 0.0286958
R2506 Vdd.n970 Vdd.n260 0.0279312
R2507 Vdd.n1005 Vdd.n202 0.0273926
R2508 Vdd.n66 Vdd.n55 0.0237
R2509 Vdd.n139 Vdd.n128 0.0237
R2510 Vdd.n569 Vdd.n558 0.0237
R2511 Vdd.n638 Vdd.n627 0.0237
R2512 Vdd.n1098 Vdd.n1097 0.0237
R2513 Vdd.n1029 Vdd.n1021 0.0197857
R2514 Vdd.n710 Vdd.n699 0.0192652
R2515 Vdd.n106 Vdd.n105 0.0161977
R2516 Vdd.n179 Vdd.n178 0.0161977
R2517 Vdd.n536 Vdd.n535 0.0161977
R2518 Vdd.n605 Vdd.n604 0.0161977
R2519 Vdd.n463 Vdd.n450 0.0161977
R2520 Vdd.n244 Vdd.n243 0.0161977
R2521 Vdd.n92 Vdd.n91 0.0129273
R2522 Vdd.n165 Vdd.n164 0.0129273
R2523 Vdd.n522 Vdd.n521 0.0129273
R2524 Vdd.n591 Vdd.n590 0.0129273
R2525 Vdd.n465 Vdd.n464 0.0129273
R2526 Vdd.n230 Vdd.n13 0.0129273
R2527 Vdd.n438 adc_PISO_0.avdd 0.0128676
R2528 Vdd.n90 Vdd.n89 0.0122273
R2529 Vdd.n163 Vdd.n162 0.0122273
R2530 Vdd.n589 Vdd.n588 0.0122273
R2531 Vdd.n657 Vdd.n651 0.0122273
R2532 Vdd.n1079 Vdd.n1078 0.0122273
R2533 Vdd.n980 Vdd.n979 0.0113078
R2534 Vdd.n1038 Vdd.n1006 0.0068
R2535 Vdd.n1005 Vdd.n1004 0.00613636
R2536 Vdd.n927 Vdd.n921 0.00505026
R2537 Vdd.n889 Vdd.n883 0.00505026
R2538 Vdd.n850 Vdd.n844 0.00505026
R2539 Vdd.n812 Vdd.n806 0.00505026
R2540 Vdd.n1004 Vdd.n1003 0.00441736
R2541 Vdd.n948 Vdd.n927 0.00430496
R2542 Vdd.n910 Vdd.n889 0.00430496
R2543 Vdd.n871 Vdd.n850 0.00430496
R2544 Vdd.n833 Vdd.n812 0.00430496
R2545 Vdd.n795 Vdd.n774 0.00430496
R2546 Vdd.n1024 comparator_no_offsetcal_0.x4.VDD 0.00371429
R2547 SARlogic_0.dffrs_5.vdd Vdd.n948 0.00349428
R2548 SARlogic_0.dffrs_4.vdd Vdd.n910 0.00349428
R2549 SARlogic_0.dffrs_3.vdd Vdd.n871 0.00349428
R2550 SARlogic_0.dffrs_2.vdd Vdd.n833 0.00349428
R2551 SARlogic_0.dffrs_1.vdd Vdd.n795 0.00349428
R2552 SARlogic_0.dffrs_0.vdd Vdd.n756 0.00349428
R2553 Vdd.n768 Vdd.n767 0.00291569
R2554 Vdd.n735 Vdd.n734 0.00285324
R2555 Vdd.n520 Vdd.n260 0.00265596
R2556 Vdd.n774 Vdd.n768 0.00263457
R2557 Vdd.n959 SARlogic_0.dffrs_5.vdd 0.00236325
R2558 Vdd.n921 SARlogic_0.dffrs_4.vdd 0.00236325
R2559 Vdd.n844 SARlogic_0.dffrs_2.vdd 0.00236325
R2560 Vdd.n806 SARlogic_0.dffrs_1.vdd 0.00236325
R2561 Vdd.n767 SARlogic_0.dffrs_0.vdd 0.00236325
R2562 Vdd.n258 Vdd.n257 0.00228481
R2563 Vdd.n883 Vdd.n872 0.0014349
R2564 Vdd.n872 SARlogic_0.dffrs_3.vdd 0.00142836
R2565 Vdd.n972 Vdd.n959 0.0008465
R2566 Vdd.n78 Vdd.n72 0.000518182
R2567 Vdd.n151 Vdd.n145 0.000518182
R2568 Vdd.n581 Vdd.n575 0.000518182
R2569 Vdd.n589 Vdd.n582 0.000518182
R2570 Vdd.n650 Vdd.n644 0.000518182
R2571 Vdd.n1091 Vdd.n1085 0.000518182
R2572 Vdd.n997 Vdd.n991 0.000517689
R2573 Vdd.n734 Vdd.n728 0.000515182
R2574 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t6 41.0041
R2575 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t5 40.6313
R2576 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t4 27.3166
R2577 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t7 26.9438
R2578 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d 17.5382
R2579 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d.n2 14.0582
R2580 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.t0 10.0473
R2581 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.t1 6.51042
R2582 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.n4 6.04952
R2583 SARlogic_0.dffrs_4.nand3_8.A SARlogic_0.dffrs_4.d.n0 5.7755
R2584 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_4.d.n1 5.13907
R2585 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n6 4.72925
R2586 SARlogic_0.dffrs_4.d SARlogic_0.dffrs_4.nand3_8.A 0.784786
R2587 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.n5 0.732092
R2588 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t3 0.7285
R2589 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t2 0.7285
R2590 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n3 0.166901
R2591 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_3.nand3_7.C 0.0455
R2592 Vss.n1474 Vss.n1473 1.11127e+06
R2593 Vss.n1508 Vss.n252 1.11127e+06
R2594 Vss.n1452 Vss.n1451 1.03768e+06
R2595 Vss.n1470 Vss.n1469 653018
R2596 Vss.n1468 Vss.n1467 533628
R2597 Vss.n1472 Vss.n1471 511643
R2598 Vss.n1777 Vss.n1776 149960
R2599 Vss.n1452 Vss.n289 136500
R2600 Vss.n1469 Vss.n1468 106786
R2601 Vss.n1471 Vss.n1470 106786
R2602 Vss.n190 Vss.n188 106554
R2603 Vss.n850 Vss.n849 50714
R2604 Vss.n1362 Vss.n1230 50260.2
R2605 Vss.n1660 Vss.n167 47256
R2606 Vss.n1467 Vss.n1466 42535.5
R2607 Vss.n1669 Vss.n1668 41697.6
R2608 Vss.n1454 Vss.n278 32884
R2609 Vss.n646 Vss.n518 32356.2
R2610 Vss.n1668 Vss.n1667 26779.4
R2611 Vss.n1064 Vss.n1063 24208.9
R2612 Vss.n24 Vss.n16 22665.9
R2613 Vss.n581 Vss.n580 22665.9
R2614 Vss.t129 Vss.n107 18167.5
R2615 Vss.n327 Vss.n278 17319
R2616 Vss.n847 Vss.n835 17088.9
R2617 Vss.n1063 Vss.n369 16547
R2618 Vss.n646 Vss.n645 16547
R2619 Vss.n252 Vss.n70 16020.5
R2620 Vss.n1504 Vss.n252 16020.5
R2621 Vss.n582 Vss.n581 15733.7
R2622 Vss.n1867 Vss.n24 15733.7
R2623 Vss.n1041 Vss.n390 15356.8
R2624 Vss.n1466 Vss.n278 14805.6
R2625 Vss.n834 Vss.n833 13656.9
R2626 Vss.n1165 Vss.n1144 13507.5
R2627 Vss.n1118 Vss.n1117 13264.1
R2628 Vss.n391 Vss.n369 12982.5
R2629 Vss.n1193 Vss.n1180 11672.3
R2630 Vss.n1880 Vss.n13 11672.3
R2631 Vss.n1072 Vss.n1071 11670.6
R2632 Vss.n682 Vss.n679 11510.4
R2633 Vss.n1071 Vss.n366 11510.4
R2634 Vss.n1288 Vss.n1129 11510.4
R2635 Vss.n1371 Vss.n1370 11510.4
R2636 Vss.n1180 Vss.n1176 11510.4
R2637 Vss.n709 Vss.n13 11510.4
R2638 Vss.n848 Vss.n847 11510.4
R2639 Vss.n679 Vss.n678 11510.4
R2640 Vss.n1038 Vss.n395 10562.5
R2641 Vss.n1668 Vss.n167 10357.6
R2642 Vss.n1660 Vss.t94 10202.1
R2643 Vss.t207 Vss.n1605 9747.75
R2644 Vss.n1471 Vss.n273 9694.18
R2645 Vss.n270 Vss.n70 9694.18
R2646 Vss.n1471 Vss.n270 9687.98
R2647 Vss.n1506 Vss.n1504 9687.98
R2648 Vss.n834 Vss.n392 9486.49
R2649 Vss.n857 Vss.n491 9213.04
R2650 Vss.n716 Vss.n499 9213.04
R2651 Vss.n1228 Vss.n1227 8696.91
R2652 Vss.n1195 Vss.n1117 7467.21
R2653 Vss.n317 Vss.n288 7154.22
R2654 Vss.n549 Vss.n534 7143.16
R2655 Vss.n797 Vss.n796 7143.16
R2656 Vss.n833 Vss.n798 7143.16
R2657 Vss.n581 Vss.n498 7082.44
R2658 Vss.n490 Vss.n24 7082.44
R2659 Vss.n351 Vss.n350 6961.73
R2660 Vss.n1164 Vss.n1142 6961.73
R2661 Vss.n832 Vss.n389 6961.73
R2662 Vss.n794 Vss.n793 6961.73
R2663 Vss.n560 Vss.n559 6961.73
R2664 Vss.n621 Vss.n601 6925.27
R2665 Vss.n1193 Vss.n1192 6921.73
R2666 Vss.n1880 Vss.n14 6921.73
R2667 Vss.n698 Vss.n697 6921.73
R2668 Vss.n1670 Vss.n188 6841.13
R2669 Vss.n1454 Vss.n277 6737.81
R2670 Vss.n1227 Vss.n1131 6393.51
R2671 Vss.n1368 Vss.n1362 6375
R2672 Vss.n1467 Vss.n277 6373.63
R2673 Vss.n1661 Vss.n1660 6317.73
R2674 Vss.n755 Vss.n392 6190.48
R2675 Vss.n1072 Vss.n315 6190.48
R2676 Vss.n1392 Vss.n1116 6157.34
R2677 Vss.n1041 Vss.n1040 5894.95
R2678 Vss.n1779 Vss.n1778 5751.62
R2679 Vss.n1036 Vss.n397 5557.62
R2680 Vss.n1008 Vss.n1006 5557.62
R2681 Vss.n1005 Vss.n208 5557.62
R2682 Vss.n128 Vss.n101 5557.62
R2683 Vss.n1807 Vss.n83 5557.62
R2684 Vss.n1806 Vss.n85 5557.62
R2685 Vss.n1404 Vss.n60 5557.62
R2686 Vss.n1831 Vss.n61 5557.62
R2687 Vss.n1348 Vss.n124 5557.62
R2688 Vss.n1347 Vss.n1346 5557.62
R2689 Vss.n939 Vss.n448 5557.62
R2690 Vss.n902 Vss.n393 5557.62
R2691 Vss.n623 Vss.n622 5557.62
R2692 Vss.n560 Vss.n547 5551.58
R2693 Vss.n793 Vss.n762 5551.58
R2694 Vss.n959 Vss.n448 5551.58
R2695 Vss.n1762 Vss.n124 5551.58
R2696 Vss.n1559 Vss.n208 5551.58
R2697 Vss.n1581 Vss.n61 5551.58
R2698 Vss.n1006 Vss.n1005 5551.58
R2699 Vss.n1202 Vss.n1142 5551.58
R2700 Vss.n351 Vss.n338 5551.58
R2701 Vss.n1051 Vss.n389 5551.58
R2702 Vss.n1749 Vss.n128 5551.58
R2703 Vss.n1684 Vss.n85 5551.58
R2704 Vss.n1807 Vss.n1806 5551.58
R2705 Vss.n1831 Vss.n60 5551.58
R2706 Vss.n1348 Vss.n1347 5551.58
R2707 Vss.n939 Vss.n397 5551.58
R2708 Vss.n903 Vss.n902 5551.58
R2709 Vss.n623 Vss.n524 5551.58
R2710 Vss.n1072 Vss.n365 5418.32
R2711 Vss.n1193 Vss.n289 5416.67
R2712 Vss.n1880 Vss.n11 5416.67
R2713 Vss.n834 Vss.n390 5243.79
R2714 Vss.n1780 Vss.n1779 4925
R2715 Vss.n1633 Vss.n189 4797.83
R2716 Vss.n1779 Vss.n107 4745.41
R2717 Vss.n1038 Vss.n1037 4485.19
R2718 Vss.n920 Vss.n449 4456.62
R2719 Vss.n1331 Vss.n1120 4448.54
R2720 Vss.n678 Vss.n677 4366.67
R2721 Vss.n395 Vss.n370 4316.58
R2722 Vss.n533 Vss.n532 4273.71
R2723 Vss.n1040 Vss.n392 4229.5
R2724 Vss.n1229 Vss.n1118 4107.2
R2725 Vss.n1605 Vss.n189 3983.8
R2726 Vss.n395 Vss.n391 3889.63
R2727 Vss.n1040 Vss.n1039 3784.25
R2728 Vss.n865 Vss.n864 3765.76
R2729 Vss.n722 Vss.n721 3765.76
R2730 Vss.n622 Vss.n533 3568.02
R2731 Vss.n1652 Vss.t515 3463.67
R2732 Vss.n1791 Vss.n100 3217.05
R2733 Vss.n159 Vss.n158 3214.99
R2734 Vss.n1369 Vss.n1229 3201.53
R2735 Vss.n1369 Vss.n1368 3178.74
R2736 Vss.n1531 Vss.n1529 3157.03
R2737 Vss.n1546 Vss.n217 3157.03
R2738 Vss.n1021 Vss.n1020 3157.03
R2739 Vss.n1818 Vss.n73 3157.03
R2740 Vss.n1394 Vss.n75 3157.03
R2741 Vss.n1426 Vss.n1425 3157.03
R2742 Vss.n1844 Vss.n1843 3157.03
R2743 Vss.n1481 Vss.n251 3157.03
R2744 Vss.n1728 Vss.n170 3157.03
R2745 Vss.n921 Vss.n396 3157.03
R2746 Vss.n1565 Vss.n206 3155.01
R2747 Vss.n1548 Vss.n1547 3155.01
R2748 Vss.n1022 Vss.n217 3155.01
R2749 Vss.n1699 Vss.n1698 3155.01
R2750 Vss.n1818 Vss.n1817 3155.01
R2751 Vss.n1481 Vss.n268 3155.01
R2752 Vss.n1531 Vss.n48 3155.01
R2753 Vss.n1593 Vss.n195 3155.01
R2754 Vss.n1730 Vss.n1729 3155.01
R2755 Vss.n1330 Vss.n170 3148.94
R2756 Vss.n1391 Vss.n1119 3122.83
R2757 Vss.n650 Vss.n648 2945.66
R2758 Vss.n364 Vss.n363 2944.88
R2759 Vss.n1167 Vss.n1166 2944.88
R2760 Vss.n795 Vss.n15 2944.88
R2761 Vss.n600 Vss.n599 2944.88
R2762 Vss.n1668 Vss.n1605 2850.36
R2763 Vss.n1670 Vss.n1669 2846.85
R2764 Vss.n1507 Vss.n188 2814.38
R2765 Vss.n1009 Vss.n383 2720.84
R2766 Vss.t207 Vss.n1614 2698.96
R2767 Vss.t515 Vss.n1614 2698.96
R2768 Vss.n364 Vss.n317 2677.48
R2769 Vss.n363 Vss.n316 2677.48
R2770 Vss.n1166 Vss.n1165 2677.48
R2771 Vss.n1194 Vss.n1167 2677.48
R2772 Vss.n796 Vss.n795 2677.48
R2773 Vss.n1879 Vss.n15 2677.48
R2774 Vss.n600 Vss.n534 2677.48
R2775 Vss.n599 Vss.n505 2677.48
R2776 Vss.n1373 Vss.n1372 2575.98
R2777 Vss.n1368 Vss.t204 2437.5
R2778 Vss.n350 Vss.n317 2353.3
R2779 Vss.n1165 Vss.n1164 2353.3
R2780 Vss.n833 Vss.n832 2353.3
R2781 Vss.n796 Vss.n794 2353.3
R2782 Vss.n559 Vss.n534 2353.3
R2783 Vss.n1391 Vss.n1118 2306.19
R2784 Vss.n1144 Vss.n1131 2303.4
R2785 Vss.n1455 Vss.n1453 2267.8
R2786 Vss.n820 Vss.n368 2257.8
R2787 Vss.n583 Vss.n569 2257.8
R2788 Vss.n1868 Vss.n23 2257.8
R2789 Vss.n1392 Vss.n1391 2253.62
R2790 Vss.n1370 Vss.n107 2145.4
R2791 Vss.n328 Vss.n316 2028.48
R2792 Vss.n1196 Vss.n1194 2027.23
R2793 Vss.n1879 Vss.n1878 2027.23
R2794 Vss.n575 Vss.n505 2027.23
R2795 Vss.n1697 Vss.n181 1972.34
R2796 Vss.n1697 Vss.n1696 1972.34
R2797 Vss.n1733 Vss.n1732 1972.34
R2798 Vss.n1742 Vss.n160 1953.93
R2799 Vss.n1742 Vss.n1741 1953.93
R2800 Vss.t122 Vss.n1371 1950
R2801 Vss.n1072 Vss.n316 1891.48
R2802 Vss.n1194 Vss.n1193 1890.32
R2803 Vss.n1880 Vss.n1879 1890.32
R2804 Vss.n697 Vss.n505 1890.32
R2805 Vss.n1019 Vss.n1008 1883.67
R2806 Vss.n1393 Vss.n83 1883.67
R2807 Vss.n1470 Vss.n274 1883.67
R2808 Vss.n1404 Vss.n47 1883.67
R2809 Vss.n1037 Vss.n1036 1883.67
R2810 Vss.n1790 Vss.n101 1861.56
R2811 Vss.n383 Vss.n382 1775.77
R2812 Vss.n835 Vss.n834 1732.36
R2813 Vss.n1732 Vss.n167 1726.87
R2814 Vss.n820 Vss.n365 1659.81
R2815 Vss.n569 Vss.n11 1659.81
R2816 Vss.n835 Vss.n23 1659.81
R2817 Vss.t129 Vss.t122 1657.5
R2818 Vss.n1392 Vss.n1117 1579.08
R2819 Vss.n1212 Vss.n1117 1476.63
R2820 Vss.n1393 Vss.n1392 1450.15
R2821 Vss.n1451 Vss.n277 1392.86
R2822 Vss.n888 Vss.n396 1336.79
R2823 Vss.n1020 Vss.n406 1336.79
R2824 Vss.n1845 Vss.n1844 1336.79
R2825 Vss.n1427 Vss.n1426 1336.79
R2826 Vss.n1395 Vss.n1394 1336.79
R2827 Vss.n1549 Vss.n1548 1336.25
R2828 Vss.n1565 Vss.n1564 1336.25
R2829 Vss.n1730 Vss.n168 1336.25
R2830 Vss.n1698 Vss.n179 1336.25
R2831 Vss.n1792 Vss.n1791 1314.68
R2832 Vss.n159 Vss.n129 1314.15
R2833 Vss.n1652 Vss.n108 1303.34
R2834 Vss.n1618 Vss.n108 1223
R2835 Vss.n609 Vss.n533 1212.42
R2836 Vss.n1452 Vss.n288 1205.38
R2837 Vss.n311 Vss.n47 1201.62
R2838 Vss.n1062 Vss.n383 1200.6
R2839 Vss.n1370 Vss.n1369 1153.88
R2840 Vss.n1020 Vss.n1019 1095.12
R2841 Vss.n1791 Vss.n1790 1095.12
R2842 Vss.n1394 Vss.n1393 1095.12
R2843 Vss.n1844 Vss.n47 1095.12
R2844 Vss.n1037 Vss.n396 1095.12
R2845 Vss.n1568 Vss.n1565 1094.63
R2846 Vss.n1548 Vss.n215 1094.63
R2847 Vss.n1742 Vss.n159 1094.63
R2848 Vss.n1698 Vss.n1697 1094.63
R2849 Vss.n1732 Vss.n1730 1094.63
R2850 Vss.n600 Vss.n504 1086.49
R2851 Vss.n1453 Vss.n1452 1062.42
R2852 Vss.n1393 Vss.n1115 1055.77
R2853 Vss.n697 Vss.n504 1048.57
R2854 Vss.n1040 Vss.n391 996.898
R2855 Vss.n1391 Vss.n1120 933.769
R2856 Vss.n1776 Vss.n109 928.572
R2857 Vss.n953 Vss.n449 927.706
R2858 Vss.n622 Vss.n621 897.806
R2859 Vss.n1508 Vss.n1507 885.807
R2860 Vss.n1064 Vss.n367 873.918
R2861 Vss.n677 Vss.n671 873.918
R2862 Vss.n1372 Vss.t111 857.144
R2863 Vss.n1781 Vss.t111 857.144
R2864 Vss.t137 Vss.n30 849.126
R2865 Vss.n733 Vss.t116 849.126
R2866 Vss.t204 Vss.n1363 847.827
R2867 Vss.t122 Vss.n1129 847.827
R2868 Vss.n1373 Vss.t129 847.827
R2869 Vss.n1192 Vss.t99 847.827
R2870 Vss.t99 Vss.n1116 847.827
R2871 Vss.t101 Vss.n14 847.827
R2872 Vss.n491 Vss.t101 847.827
R2873 Vss.t215 Vss.n865 847.827
R2874 Vss.n874 Vss.t215 847.827
R2875 Vss.n873 Vss.t251 847.827
R2876 Vss.n870 Vss.t251 847.827
R2877 Vss.n869 Vss.t137 847.827
R2878 Vss.n698 Vss.t591 847.827
R2879 Vss.t591 Vss.n499 847.827
R2880 Vss.n722 Vss.t183 847.827
R2881 Vss.n725 Vss.t183 847.827
R2882 Vss.t3 Vss.n726 847.827
R2883 Vss.n731 Vss.t3 847.827
R2884 Vss.t116 Vss.n732 847.827
R2885 Vss.n451 Vss.n448 832.22
R2886 Vss.n232 Vss.n61 832.22
R2887 Vss.n218 Vss.n208 832.22
R2888 Vss.n1006 Vss.n412 832.22
R2889 Vss.n351 Vss.n339 832.22
R2890 Vss.n149 Vss.n128 832.22
R2891 Vss.n1153 Vss.n1142 832.22
R2892 Vss.n1707 Vss.n85 832.22
R2893 Vss.n1808 Vss.n1807 832.22
R2894 Vss.n60 Vss.n59 832.22
R2895 Vss.n171 Vss.n124 832.22
R2896 Vss.n1347 Vss.n1282 832.22
R2897 Vss.n922 Vss.n397 832.22
R2898 Vss.n810 Vss.n389 832.22
R2899 Vss.n902 Vss.n900 832.22
R2900 Vss.n793 Vss.n763 832.22
R2901 Vss.n560 Vss.n548 832.22
R2902 Vss.n623 Vss.n531 832.22
R2903 Vss.n448 Vss.n447 832.101
R2904 Vss.n1514 Vss.n61 832.101
R2905 Vss.n236 Vss.n208 832.101
R2906 Vss.n1006 Vss.n422 832.101
R2907 Vss.n352 Vss.n351 832.101
R2908 Vss.n128 Vss.n127 832.101
R2909 Vss.n1142 Vss.n1141 832.101
R2910 Vss.n1714 Vss.n85 832.101
R2911 Vss.n1807 Vss.n84 832.101
R2912 Vss.n1410 Vss.n60 832.101
R2913 Vss.n130 Vss.n124 832.101
R2914 Vss.n1347 Vss.n1283 832.101
R2915 Vss.n404 Vss.n397 832.101
R2916 Vss.n819 Vss.n389 832.101
R2917 Vss.n902 Vss.n901 832.101
R2918 Vss.n793 Vss.n792 832.101
R2919 Vss.n561 Vss.n560 832.101
R2920 Vss.n624 Vss.n623 832.101
R2921 Vss.n1037 Vss.n383 829.364
R2922 Vss.n1506 Vss.n1505 814.398
R2923 Vss.n270 Vss.n269 814.398
R2924 Vss.n1212 Vss.t353 812.5
R2925 Vss.t255 Vss.n1119 812.5
R2926 Vss.n857 Vss.t83 812.5
R2927 Vss.n716 Vss.t489 812.5
R2928 Vss.n1465 Vss.n279 798.088
R2929 Vss.n647 Vss.n646 767.827
R2930 Vss.n1371 Vss.n1130 755.625
R2931 Vss.n280 Vss.n47 750.922
R2932 Vss.n1455 Vss.n1454 748.735
R2933 Vss.t129 Vss.t122 720.653
R2934 Vss.n874 Vss.n873 720.653
R2935 Vss.n870 Vss.n869 720.653
R2936 Vss.n726 Vss.n725 720.653
R2937 Vss.n732 Vss.n731 720.653
R2938 Vss.n1669 Vss.n1604 702.332
R2939 Vss.n1426 Vss.n274 698.639
R2940 Vss.n338 Vss.n337 693.082
R2941 Vss.n585 Vss.n547 692.747
R2942 Vss.n1203 Vss.n1202 692.747
R2943 Vss.n762 Vss.n761 692.747
R2944 Vss.n1667 Vss.t276 676.471
R2945 Vss.n1614 Vss.t276 676.471
R2946 Vss.n1614 Vss.t148 676.471
R2947 Vss.n1661 Vss.t148 676.471
R2948 Vss.n382 Vss.t325 670.104
R2949 Vss.t325 Vss.n381 670.104
R2950 Vss.n378 Vss.t135 670.104
R2951 Vss.n375 Vss.t135 670.104
R2952 Vss.n374 Vss.t569 670.104
R2953 Vss.t569 Vss.n367 670.104
R2954 Vss.n648 Vss.t671 670.104
R2955 Vss.n662 Vss.t671 670.104
R2956 Vss.n663 Vss.t229 670.104
R2957 Vss.n667 Vss.t229 670.104
R2958 Vss.t512 Vss.n670 670.104
R2959 Vss.n671 Vss.t512 670.104
R2960 Vss.n1064 Vss.n368 665.564
R2961 Vss.n583 Vss.n582 665.564
R2962 Vss.n1868 Vss.n1867 665.564
R2963 Vss.n1473 Vss.n270 662.646
R2964 Vss.n338 Vss.n336 662.074
R2965 Vss.n1202 Vss.n1201 661.665
R2966 Vss.n762 Vss.n760 661.665
R2967 Vss.n579 Vss.n547 661.665
R2968 Vss.t353 Vss.t458 650
R2969 Vss.t458 Vss.t255 650
R2970 Vss.t400 Vss.t86 650
R2971 Vss.t432 Vss.t235 650
R2972 Vss.t567 Vss.n1062 642.183
R2973 Vss.t352 Vss.n647 642.183
R2974 Vss.n651 Vss.t340 642.183
R2975 Vss.n1781 Vss.n1780 607.144
R2976 Vss.n798 Vss.n365 597.985
R2977 Vss.n549 Vss.n11 597.985
R2978 Vss.n835 Vss.n797 597.985
R2979 Vss.n1229 Vss.n1228 596.029
R2980 Vss.n1367 Vss.t103 590.91
R2981 Vss.t204 Vss.n1367 590.91
R2982 Vss.t77 Vss.n1065 590.909
R2983 Vss.n1069 Vss.t77 590.909
R2984 Vss.t232 Vss.n1069 590.909
R2985 Vss.n1071 Vss.t98 590.909
R2986 Vss.n1071 Vss.t629 590.909
R2987 Vss.n1073 Vss.t631 590.909
R2988 Vss.n1450 Vss.t311 590.909
R2989 Vss.n1179 Vss.t311 590.909
R2990 Vss.t590 Vss.n1179 590.909
R2991 Vss.n1180 Vss.t114 590.909
R2992 Vss.t675 Vss.n1180 590.909
R2993 Vss.n1188 Vss.t19 590.909
R2994 Vss.n574 Vss.t75 590.909
R2995 Vss.t75 Vss.n573 590.909
R2996 Vss.n573 Vss.t233 590.909
R2997 Vss.t528 Vss.n13 590.909
R2998 Vss.n13 Vss.t225 590.909
R2999 Vss.n1881 Vss.t474 590.909
R3000 Vss.n1866 Vss.t388 590.909
R3001 Vss.n838 Vss.t388 590.909
R3002 Vss.t113 Vss.n838 590.909
R3003 Vss.n847 Vss.t589 590.909
R3004 Vss.n847 Vss.t638 590.909
R3005 Vss.t245 Vss.n846 590.909
R3006 Vss.n676 Vss.t649 590.909
R3007 Vss.t649 Vss.n675 590.909
R3008 Vss.n675 Vss.t529 590.909
R3009 Vss.n679 Vss.t231 590.909
R3010 Vss.n679 Vss.t653 590.909
R3011 Vss.n696 Vss.t657 590.909
R3012 Vss.n1528 Vss.t194 582.165
R3013 Vss.n232 Vss.t441 582.165
R3014 Vss.n1545 Vss.t648 582.165
R3015 Vss.n218 Vss.t420 582.165
R3016 Vss.t358 Vss.n405 582.165
R3017 Vss.n412 Vss.t195 582.165
R3018 Vss.n362 Vss.t5 582.165
R3019 Vss.n339 Vss.t394 582.165
R3020 Vss.n150 Vss.t165 582.165
R3021 Vss.t491 Vss.n149 582.165
R3022 Vss.t68 Vss.n1143 582.165
R3023 Vss.n1153 Vss.t408 582.165
R3024 Vss.n1708 Vss.t38 582.165
R3025 Vss.t406 Vss.n1707 582.165
R3026 Vss.n1809 Vss.t625 582.165
R3027 Vss.t237 Vss.n1808 582.165
R3028 Vss.n1424 Vss.t63 582.165
R3029 Vss.t34 Vss.n271 582.165
R3030 Vss.n1842 Vss.t108 582.165
R3031 Vss.n59 Vss.t380 582.165
R3032 Vss.n1510 Vss.t565 582.165
R3033 Vss.t422 Vss.n1509 582.165
R3034 Vss.n1727 Vss.t239 582.165
R3035 Vss.n171 Vss.t428 582.165
R3036 Vss.n1332 Vss.t248 582.165
R3037 Vss.t305 Vss.n1282 582.165
R3038 Vss.n923 Vss.t150 582.165
R3039 Vss.t192 Vss.n922 582.165
R3040 Vss.n458 Vss.t29 582.165
R3041 Vss.n451 Vss.t424 582.165
R3042 Vss.t384 Vss.n809 582.165
R3043 Vss.n810 Vss.t396 582.165
R3044 Vss.n757 Vss.t139 582.165
R3045 Vss.n900 Vss.t27 582.165
R3046 Vss.n774 Vss.t244 582.165
R3047 Vss.t426 Vss.n763 582.165
R3048 Vss.n598 Vss.t670 582.165
R3049 Vss.n548 Vss.t433 582.165
R3050 Vss.n609 Vss.t274 582.165
R3051 Vss.t449 Vss.n531 582.165
R3052 Vss.n585 Vss.t624 581.712
R3053 Vss.t145 Vss.n584 581.712
R3054 Vss.t618 Vss.n394 581.712
R3055 Vss.n888 Vss.t25 581.712
R3056 Vss.n1035 Vss.t182 581.712
R3057 Vss.n406 Vss.t156 581.712
R3058 Vss.n996 Vss.t220 581.712
R3059 Vss.t179 Vss.n230 581.712
R3060 Vss.n1534 Vss.t371 581.712
R3061 Vss.t390 Vss.n1533 581.712
R3062 Vss.n941 Vss.t151 581.712
R3063 Vss.t307 Vss.n431 581.712
R3064 Vss.n440 Vss.t24 581.712
R3065 Vss.n1549 Vss.t222 581.712
R3066 Vss.n933 Vss.t224 581.712
R3067 Vss.n978 Vss.t416 581.712
R3068 Vss.n447 Vss.t510 581.712
R3069 Vss.t303 Vss.n216 581.712
R3070 Vss.n1582 Vss.t48 581.712
R3071 Vss.t581 Vss.n194 581.712
R3072 Vss.n1560 Vss.t514 581.712
R3073 Vss.n1564 Vss.t466 581.712
R3074 Vss.t522 Vss.n1514 581.712
R3075 Vss.n1515 Vss.t30 581.712
R3076 Vss.t508 Vss.n236 581.712
R3077 Vss.n237 Vss.t621 581.712
R3078 Vss.n422 Vss.t553 581.712
R3079 Vss.n414 Vss.t253 581.712
R3080 Vss.n1007 Vss.t177 581.712
R3081 Vss.n1845 Vss.t197 581.712
R3082 Vss.t635 Vss.n1405 581.712
R3083 Vss.n1427 Vss.t382 581.712
R3084 Vss.n1163 Vss.t278 581.712
R3085 Vss.n1145 Vss.t455 581.712
R3086 Vss.n352 Vss.t472 581.712
R3087 Vss.t651 Vss.n287 581.712
R3088 Vss.n349 Vss.t267 581.712
R3089 Vss.n340 Vss.t446 581.712
R3090 Vss.n337 Vss.t566 581.712
R3091 Vss.n1456 Vss.t51 581.712
R3092 Vss.t669 Vss.n1052 581.712
R3093 Vss.n1053 Vss.t551 581.712
R3094 Vss.n1276 Vss.t540 581.712
R3095 Vss.t535 Vss.n1233 581.712
R3096 Vss.n1793 Vss.t188 581.712
R3097 Vss.t412 Vss.n1792 581.712
R3098 Vss.n1761 Vss.t477 581.712
R3099 Vss.n129 Vss.t348 581.712
R3100 Vss.n1750 Vss.t115 581.712
R3101 Vss.t598 Vss.n110 581.712
R3102 Vss.n136 Vss.t469 581.712
R3103 Vss.t495 Vss.n111 581.712
R3104 Vss.n127 Vss.t518 581.712
R3105 Vss.n1775 Vss.t463 581.712
R3106 Vss.n1141 Vss.t81 581.712
R3107 Vss.n1226 Vss.t345 581.712
R3108 Vss.n1203 Vss.t470 581.712
R3109 Vss.t279 Vss.n1132 581.712
R3110 Vss.n1316 Vss.t44 581.712
R3111 Vss.t240 Vss.n1315 581.712
R3112 Vss.t202 Vss.n272 581.712
R3113 Vss.n1395 Vss.t36 581.712
R3114 Vss.t61 Vss.n87 581.712
R3115 Vss.n1268 Vss.t548 581.712
R3116 Vss.t596 Vss.n88 581.712
R3117 Vss.n1265 Vss.t435 581.712
R3118 Vss.n1821 Vss.t1 581.712
R3119 Vss.t213 Vss.n1820 581.712
R3120 Vss.n1503 Vss.t316 581.712
R3121 Vss.t453 Vss.n71 581.712
R3122 Vss.n1685 Vss.t468 581.712
R3123 Vss.t594 Vss.n168 581.712
R3124 Vss.n1505 Vss.t521 581.712
R3125 Vss.n1700 Vss.t119 581.712
R3126 Vss.n1671 Vss.t473 581.712
R3127 Vss.t317 Vss.n179 581.712
R3128 Vss.n1714 Vss.t509 581.712
R3129 Vss.t53 Vss.n169 581.712
R3130 Vss.t71 Vss.n84 581.712
R3131 Vss.n1329 Vss.t106 581.712
R3132 Vss.n269 Vss.t662 581.712
R3133 Vss.n1816 Vss.t39 581.712
R3134 Vss.t499 Vss.n1410 581.712
R3135 Vss.n1411 Vss.t301 581.712
R3136 Vss.n1829 Vss.t462 581.712
R3137 Vss.n261 Vss.t633 581.712
R3138 Vss.t580 Vss.n63 581.712
R3139 Vss.n267 Vss.t414 581.712
R3140 Vss.n130 Vss.t507 581.712
R3141 Vss.n157 Vss.t272 581.712
R3142 Vss.n1283 Vss.t298 581.712
R3143 Vss.n1361 Vss.t323 581.712
R3144 Vss.n1343 Vss.t534 581.712
R3145 Vss.t163 Vss.n1234 581.712
R3146 Vss.t465 Vss.n404 581.712
R3147 Vss.n1023 Vss.t268 581.712
R3148 Vss.n480 Vss.t12 581.712
R3149 Vss.n474 Vss.t619 581.712
R3150 Vss.n831 Vss.t550 581.712
R3151 Vss.n799 Vss.t451 581.712
R3152 Vss.t347 Vss.n819 581.712
R3153 Vss.n821 Vss.t242 581.712
R3154 Vss.n901 Vss.t132 581.712
R3155 Vss.n919 Vss.t32 581.712
R3156 Vss.n759 Vss.t169 581.712
R3157 Vss.t418 Vss.n758 581.712
R3158 Vss.n792 Vss.t354 581.712
R3159 Vss.n764 Vss.t484 581.712
R3160 Vss.n561 Vss.t339 581.712
R3161 Vss.n568 Vss.t199 581.712
R3162 Vss.n558 Vss.t211 581.712
R3163 Vss.n550 Vss.t430 581.712
R3164 Vss.n636 Vss.t586 581.712
R3165 Vss.t22 Vss.n635 581.712
R3166 Vss.n761 Vss.t668 581.712
R3167 Vss.n1869 Vss.t167 581.712
R3168 Vss.t82 Vss.n624 581.712
R3169 Vss.n625 Vss.t577 581.712
R3170 Vss.n620 Vss.t249 581.712
R3171 Vss.n602 Vss.t438 581.712
R3172 Vss.n381 Vss.n378 569.588
R3173 Vss.n375 Vss.n374 569.588
R3174 Vss.n663 Vss.n662 569.588
R3175 Vss.n670 Vss.n667 569.588
R3176 Vss.n1369 Vss.n1131 565.155
R3177 Vss.t86 Vss.n490 561.686
R3178 Vss.t235 Vss.n498 561.686
R3179 Vss.n1036 Vss.n1035 548.236
R3180 Vss.n1008 Vss.n1007 548.236
R3181 Vss.n1405 Vss.n1404 548.236
R3182 Vss.n136 Vss.n101 548.236
R3183 Vss.n1316 Vss.n83 548.236
R3184 Vss.n1582 Vss.n1581 548.058
R3185 Vss.n1560 Vss.n1559 548.058
R3186 Vss.n1052 Vss.n1051 548.058
R3187 Vss.n1762 Vss.n1761 548.058
R3188 Vss.n1750 Vss.n1749 548.058
R3189 Vss.n1685 Vss.n1684 548.058
R3190 Vss.n636 Vss.n524 548.058
R3191 Vss.t374 Vss.t393 513.746
R3192 Vss.t393 Vss.t567 513.746
R3193 Vss.t440 Vss.t352 513.746
R3194 Vss.t340 Vss.t440 513.746
R3195 Vss.t98 Vss.t232 502.274
R3196 Vss.t629 Vss.t631 502.274
R3197 Vss.t103 Vss.t593 502.274
R3198 Vss.t114 Vss.t590 502.274
R3199 Vss.t19 Vss.t675 502.274
R3200 Vss.t233 Vss.t528 502.274
R3201 Vss.t225 Vss.t474 502.274
R3202 Vss.t589 Vss.t113 502.274
R3203 Vss.t638 Vss.t245 502.274
R3204 Vss.t529 Vss.t231 502.274
R3205 Vss.t653 Vss.t657 502.274
R3206 Vss.n1581 Vss.n1580 484.702
R3207 Vss.n1559 Vss.n1558 484.702
R3208 Vss.n1051 Vss.n1050 484.702
R3209 Vss.n1749 Vss.n1748 484.702
R3210 Vss.n1684 Vss.n1683 484.702
R3211 Vss.n1763 Vss.n1762 484.702
R3212 Vss.n644 Vss.n524 484.702
R3213 Vss.t579 Vss.t194 465.733
R3214 Vss.t441 Vss.t579 465.733
R3215 Vss.t370 Vss.t648 465.733
R3216 Vss.t420 Vss.t370 465.733
R3217 Vss.t178 Vss.t358 465.733
R3218 Vss.t195 Vss.t178 465.733
R3219 Vss.t50 Vss.t5 465.733
R3220 Vss.t394 Vss.t50 465.733
R3221 Vss.t165 Vss.t471 465.733
R3222 Vss.t471 Vss.t491 465.733
R3223 Vss.t158 Vss.t68 465.733
R3224 Vss.t408 Vss.t158 465.733
R3225 Vss.t38 Vss.t597 465.733
R3226 Vss.t597 Vss.t406 465.733
R3227 Vss.t625 Vss.t43 465.733
R3228 Vss.t43 Vss.t237 465.733
R3229 Vss.t63 Vss.t203 465.733
R3230 Vss.t203 Vss.t34 465.733
R3231 Vss.t644 Vss.t108 465.733
R3232 Vss.t380 Vss.t644 465.733
R3233 Vss.t565 Vss.t319 465.733
R3234 Vss.t319 Vss.t422 465.733
R3235 Vss.t187 Vss.t239 465.733
R3236 Vss.t428 Vss.t187 465.733
R3237 Vss.t248 Vss.t533 465.733
R3238 Vss.t533 Vss.t305 465.733
R3239 Vss.t150 Vss.t181 465.733
R3240 Vss.t181 Vss.t192 465.733
R3241 Vss.t147 Vss.t29 465.733
R3242 Vss.t424 Vss.t147 465.733
R3243 Vss.t603 Vss.t384 465.733
R3244 Vss.t396 Vss.t603 465.733
R3245 Vss.t139 Vss.t617 465.733
R3246 Vss.t617 Vss.t27 465.733
R3247 Vss.t244 Vss.t366 465.733
R3248 Vss.t366 Vss.t426 465.733
R3249 Vss.t212 Vss.t670 465.733
R3250 Vss.t433 Vss.t212 465.733
R3251 Vss.t274 Vss.t21 465.733
R3252 Vss.t21 Vss.t449 465.733
R3253 Vss.t624 Vss.t387 465.37
R3254 Vss.t387 Vss.t145 465.37
R3255 Vss.t13 Vss.t618 465.37
R3256 Vss.t25 Vss.t13 465.37
R3257 Vss.t152 Vss.t182 465.37
R3258 Vss.t156 Vss.t152 465.37
R3259 Vss.t220 Vss.t554 465.37
R3260 Vss.t554 Vss.t179 465.37
R3261 Vss.t371 Vss.t335 465.37
R3262 Vss.t335 Vss.t390 465.37
R3263 Vss.t151 Vss.t336 465.37
R3264 Vss.t336 Vss.t307 465.37
R3265 Vss.t24 Vss.t505 465.37
R3266 Vss.t505 Vss.t222 465.37
R3267 Vss.t224 Vss.t0 465.37
R3268 Vss.t0 Vss.t416 465.37
R3269 Vss.t510 Vss.t524 465.37
R3270 Vss.t524 Vss.t303 465.37
R3271 Vss.t48 Vss.t519 465.37
R3272 Vss.t519 Vss.t581 465.37
R3273 Vss.t514 Vss.t504 465.37
R3274 Vss.t504 Vss.t466 465.37
R3275 Vss.t561 Vss.t522 465.37
R3276 Vss.t30 Vss.t561 465.37
R3277 Vss.t607 Vss.t508 465.37
R3278 Vss.t621 Vss.t607 465.37
R3279 Vss.t562 Vss.t553 465.37
R3280 Vss.t253 Vss.t562 465.37
R3281 Vss.t177 Vss.t221 465.37
R3282 Vss.t221 Vss.t197 465.37
R3283 Vss.t461 Vss.t635 465.37
R3284 Vss.t382 Vss.t461 465.37
R3285 Vss.t330 Vss.t278 465.37
R3286 Vss.t455 Vss.t330 465.37
R3287 Vss.t472 Vss.t402 465.37
R3288 Vss.t402 Vss.t651 465.37
R3289 Vss.t572 Vss.t267 465.37
R3290 Vss.t446 Vss.t572 465.37
R3291 Vss.t566 Vss.t331 465.37
R3292 Vss.t331 Vss.t51 465.37
R3293 Vss.t355 Vss.t669 465.37
R3294 Vss.t551 Vss.t355 465.37
R3295 Vss.t540 Vss.t155 465.37
R3296 Vss.t155 Vss.t535 465.37
R3297 Vss.t188 Vss.t478 465.37
R3298 Vss.t478 Vss.t412 465.37
R3299 Vss.t501 Vss.t477 465.37
R3300 Vss.t348 Vss.t501 465.37
R3301 Vss.t115 Vss.t520 465.37
R3302 Vss.t520 Vss.t598 465.37
R3303 Vss.t469 Vss.t281 465.37
R3304 Vss.t281 Vss.t495 465.37
R3305 Vss.t518 Vss.t457 465.37
R3306 Vss.t457 Vss.t463 465.37
R3307 Vss.t81 Vss.t399 465.37
R3308 Vss.t399 Vss.t345 465.37
R3309 Vss.t470 Vss.t386 465.37
R3310 Vss.t386 Vss.t279 465.37
R3311 Vss.t44 Vss.t62 465.37
R3312 Vss.t62 Vss.t240 465.37
R3313 Vss.t2 Vss.t202 465.37
R3314 Vss.t36 Vss.t2 465.37
R3315 Vss.t70 Vss.t61 465.37
R3316 Vss.t548 Vss.t70 465.37
R3317 Vss.t329 Vss.t596 465.37
R3318 Vss.t435 Vss.t329 465.37
R3319 Vss.t1 Vss.t664 465.37
R3320 Vss.t664 Vss.t213 465.37
R3321 Vss.t316 Vss.t375 465.37
R3322 Vss.t375 Vss.t453 465.37
R3323 Vss.t468 Vss.t511 465.37
R3324 Vss.t511 Vss.t594 465.37
R3325 Vss.t521 Vss.t282 465.37
R3326 Vss.t282 Vss.t119 465.37
R3327 Vss.t473 Vss.t506 465.37
R3328 Vss.t506 Vss.t317 465.37
R3329 Vss.t509 Vss.t490 465.37
R3330 Vss.t490 Vss.t53 465.37
R3331 Vss.t292 Vss.t71 465.37
R3332 Vss.t106 Vss.t292 465.37
R3333 Vss.t662 Vss.t606 465.37
R3334 Vss.t606 Vss.t39 465.37
R3335 Vss.t283 Vss.t499 465.37
R3336 Vss.t301 Vss.t283 465.37
R3337 Vss.t500 Vss.t462 465.37
R3338 Vss.t633 Vss.t500 465.37
R3339 Vss.t49 Vss.t580 465.37
R3340 Vss.t414 Vss.t49 465.37
R3341 Vss.t507 Vss.t293 465.37
R3342 Vss.t293 Vss.t272 465.37
R3343 Vss.t298 Vss.t494 465.37
R3344 Vss.t494 Vss.t323 465.37
R3345 Vss.t534 Vss.t541 465.37
R3346 Vss.t541 Vss.t163 465.37
R3347 Vss.t616 Vss.t465 465.37
R3348 Vss.t268 Vss.t616 465.37
R3349 Vss.t125 Vss.t12 465.37
R3350 Vss.t619 Vss.t125 465.37
R3351 Vss.t84 Vss.t550 465.37
R3352 Vss.t451 Vss.t84 465.37
R3353 Vss.t403 Vss.t347 465.37
R3354 Vss.t242 Vss.t403 465.37
R3355 Vss.t132 Vss.t525 465.37
R3356 Vss.t525 Vss.t32 465.37
R3357 Vss.t169 Vss.t250 465.37
R3358 Vss.t250 Vss.t418 465.37
R3359 Vss.t410 Vss.t354 465.37
R3360 Vss.t484 Vss.t410 465.37
R3361 Vss.t339 Vss.t443 465.37
R3362 Vss.t443 Vss.t199 465.37
R3363 Vss.t626 Vss.t211 465.37
R3364 Vss.t430 Vss.t626 465.37
R3365 Vss.t586 Vss.t332 465.37
R3366 Vss.t332 Vss.t22 465.37
R3367 Vss.t668 Vss.t476 465.37
R3368 Vss.t476 Vss.t167 465.37
R3369 Vss.t448 Vss.t82 465.37
R3370 Vss.t577 Vss.t448 465.37
R3371 Vss.t585 Vss.t249 465.37
R3372 Vss.t438 Vss.t585 465.37
R3373 Vss.n336 Vss.t627 462.849
R3374 Vss.n1201 Vss.t17 462.562
R3375 Vss.n760 Vss.t487 462.562
R3376 Vss.t655 Vss.n579 462.562
R3377 Vss.n961 Vss.n215 443.358
R3378 Vss.n215 Vss.n213 443.358
R3379 Vss.n1569 Vss.n1568 443.358
R3380 Vss.n1568 Vss.n1567 443.358
R3381 Vss.n423 Vss.n217 435.214
R3382 Vss.n1818 Vss.n74 435.214
R3383 Vss.n1531 Vss.n1530 435.214
R3384 Vss.n1481 Vss.n1480 435.214
R3385 Vss.n1281 Vss.n170 435.012
R3386 Vss.n1646 Vss.n1617 414.478
R3387 Vss.n979 Vss.n217 404.991
R3388 Vss.n1819 Vss.n1818 404.991
R3389 Vss.n1532 Vss.n1531 404.991
R3390 Vss.n1482 Vss.n1481 404.991
R3391 Vss.n1267 Vss.n170 404.803
R3392 Vss.n1063 Vss.n370 402.062
R3393 Vss.t261 Vss.t259 384.214
R3394 Vss.n715 Vss.n707 383.418
R3395 Vss.n715 Vss.n714 383.418
R3396 Vss.n856 Vss.n746 383.418
R3397 Vss.n856 Vss.n855 383.418
R3398 Vss.t398 Vss.t486 370.279
R3399 Vss.t486 Vss.t627 370.279
R3400 Vss.t444 Vss.t623 370.05
R3401 Vss.t623 Vss.t17 370.05
R3402 Vss.t85 Vss.t411 370.05
R3403 Vss.t487 Vss.t85 370.05
R3404 Vss.t445 Vss.t234 370.05
R3405 Vss.t234 Vss.t655 370.05
R3406 Vss.n856 Vss.t400 367.392
R3407 Vss.n715 Vss.t432 367.392
R3408 Vss.n328 Vss.n327 366.255
R3409 Vss.n988 Vss.t314 366.243
R3410 Vss.t601 Vss.n231 366.243
R3411 Vss.n932 Vss.t310 366.243
R3412 Vss.n980 Vss.t537 366.243
R3413 Vss.n1804 Vss.t309 366.243
R3414 Vss.n1266 Vss.t645 366.243
R3415 Vss.n1490 Vss.t315 366.243
R3416 Vss.t665 Vss.n72 366.243
R3417 Vss.t247 Vss.n62 366.243
R3418 Vss.n1483 Vss.t189 366.243
R3419 Vss.n1196 Vss.n1195 366.027
R3420 Vss.n1878 Vss.n16 366.027
R3421 Vss.n580 Vss.n575 366.027
R3422 Vss.n1243 Vss.t313 365.705
R3423 Vss.t543 Vss.n1232 365.705
R3424 Vss.t593 Vss.n1130 361.933
R3425 Vss.t94 Vss.n1609 350.313
R3426 Vss.n1566 Vss.t609 338.849
R3427 Vss.n1580 Vss.t15 338.849
R3428 Vss.n214 Vss.t290 338.849
R3429 Vss.n1558 Vss.t356 338.849
R3430 Vss.n1042 Vss.t405 338.849
R3431 Vss.n1743 Vss.t401 338.849
R3432 Vss.n1748 Vss.t640 338.849
R3433 Vss.t610 Vss.n180 338.849
R3434 Vss.n1683 Vss.t377 338.849
R3435 Vss.n1731 Vss.t611 338.849
R3436 Vss.n1763 Vss.t343 338.849
R3437 Vss.n532 Vss.t404 338.849
R3438 Vss.t368 Vss.n644 338.849
R3439 Vss.n650 Vss.n649 330.211
R3440 Vss.n1130 Vss.n1129 328.534
R3441 Vss.n601 Vss.n600 307.176
R3442 Vss.t314 Vss.t497 292.995
R3443 Vss.t497 Vss.t601 292.995
R3444 Vss.t310 Vss.t563 292.995
R3445 Vss.t563 Vss.t537 292.995
R3446 Vss.t287 Vss.t309 292.995
R3447 Vss.t645 Vss.t287 292.995
R3448 Vss.t315 Vss.t288 292.995
R3449 Vss.t288 Vss.t665 292.995
R3450 Vss.t493 Vss.t247 292.995
R3451 Vss.t189 Vss.t493 292.995
R3452 Vss.t313 Vss.t527 292.565
R3453 Vss.t527 Vss.t543 292.565
R3454 Vss.t83 Vss.n856 282.61
R3455 Vss.t489 Vss.n715 282.61
R3456 Vss.t257 Vss.n1654 282.512
R3457 Vss.n1604 Vss.t376 282.289
R3458 Vss.t174 Vss.n181 282.289
R3459 Vss.n1696 Vss.t342 282.289
R3460 Vss.n182 Vss.t140 282.289
R3461 Vss.n1733 Vss.t642 282.289
R3462 Vss.t218 Vss.n160 282.289
R3463 Vss.n1741 Vss.t134 282.289
R3464 Vss.n112 Vss.t296 282.289
R3465 Vss.t609 Vss.t142 271.079
R3466 Vss.t142 Vss.t15 271.079
R3467 Vss.t290 Vss.t479 271.079
R3468 Vss.t479 Vss.t356 271.079
R3469 Vss.t405 Vss.t667 271.079
R3470 Vss.t667 Vss.t636 271.079
R3471 Vss.t401 Vss.t295 271.079
R3472 Vss.t295 Vss.t640 271.079
R3473 Vss.t118 Vss.t610 271.079
R3474 Vss.t377 Vss.t118 271.079
R3475 Vss.t611 Vss.t217 271.079
R3476 Vss.t217 Vss.t343 271.079
R3477 Vss.t294 Vss.t368 271.079
R3478 Vss.n1789 Vss.n102 266.082
R3479 Vss.n1655 Vss.t257 259.911
R3480 Vss.n1776 Vss.n102 250.827
R3481 Vss.n864 Vss.n490 250.815
R3482 Vss.n721 Vss.n498 250.815
R3483 Vss.n953 Vss.n952 247.475
R3484 Vss.t94 Vss.n1659 246.108
R3485 Vss.n182 Vss.n167 245.469
R3486 Vss.n1063 Vss.t374 240.12
R3487 Vss.n1473 Vss.n1472 232.143
R3488 Vss.n1474 Vss.n252 232.143
R3489 Vss.n1468 Vss.n276 229.095
R3490 Vss.n1170 Vss.t270 228.071
R3491 Vss.n1170 Vss.t379 228.071
R3492 Vss.n1176 Vss.t154 228.071
R3493 Vss.n1176 Vss.t6 228.071
R3494 Vss.t8 Vss.n1115 228.071
R3495 Vss.t59 Vss.n1009 228.004
R3496 Vss.n1018 Vss.t69 228.004
R3497 Vss.t72 Vss.n366 228.004
R3498 Vss.t172 Vss.n366 228.004
R3499 Vss.n1013 Vss.t170 228.004
R3500 Vss.t263 Vss.n1652 226.008
R3501 Vss.t376 Vss.t614 225.832
R3502 Vss.t614 Vss.t174 225.832
R3503 Vss.t284 Vss.t342 225.832
R3504 Vss.t140 Vss.t284 225.832
R3505 Vss.t642 Vss.t608 225.832
R3506 Vss.t608 Vss.t218 225.832
R3507 Vss.t296 Vss.t437 225.832
R3508 Vss.n1362 Vss.n1231 225.304
R3509 Vss.n645 Vss.t294 220.988
R3510 Vss.n1050 Vss.n369 213.623
R3511 Vss.n1363 Vss.n1362 211.958
R3512 Vss.n1636 Vss.n1622 205.139
R3513 Vss.n1622 Vss.n1616 205.139
R3514 Vss.n1637 Vss.n1616 205.139
R3515 Vss.n1637 Vss.n1636 205.139
R3516 Vss.n1593 Vss.n1592 200.773
R3517 Vss.t379 Vss.t154 193.861
R3518 Vss.t6 Vss.t8 193.861
R3519 Vss.t69 Vss.t72 193.804
R3520 Vss.t170 Vss.t172 193.804
R3521 Vss.n1635 Vss.n1633 193.476
R3522 Vss.n1639 Vss.n1618 193.476
R3523 Vss.n275 Vss.n273 191.959
R3524 Vss.n1594 Vss.n1593 186.831
R3525 Vss.n314 Vss.t109 179.683
R3526 Vss.n311 Vss.t109 179.683
R3527 Vss.t673 Vss.n279 179.683
R3528 Vss.n1092 Vss.t673 179.683
R3529 Vss.n1097 Vss.t88 179.683
R3530 Vss.n1098 Vss.t265 179.683
R3531 Vss.t265 Vss.n276 179.683
R3532 Vss.n1568 Vss.n1566 178.264
R3533 Vss.n215 Vss.n214 178.264
R3534 Vss.n1697 Vss.n180 178.264
R3535 Vss.n1732 Vss.n1731 178.264
R3536 Vss.n280 Vss.t97 172.196
R3537 Vss.n1300 Vss.t41 170.268
R3538 Vss.t41 Vss.n1231 170.268
R3539 Vss.n1013 Vss.n315 167.056
R3540 Vss.n1631 Vss.n1624 166.989
R3541 Vss.n1644 Vss.n1619 166.989
R3542 Vss.n1019 Vss.n1018 166.254
R3543 Vss.n1005 Vss.n1004 165.725
R3544 Vss.n1806 Vss.n86 165.725
R3545 Vss.n1832 Vss.n1831 165.725
R3546 Vss.n939 Vss.n938 165.725
R3547 Vss.n1349 Vss.n1348 165.648
R3548 Vss.n1166 Vss.n289 161.839
R3549 Vss.n795 Vss.n11 161.839
R3550 Vss.n365 Vss.n364 160.189
R3551 Vss.n1743 Vss.n1742 156.166
R3552 Vss.n315 Vss.n314 154.976
R3553 Vss.n1093 Vss.n1092 152.731
R3554 Vss.n1098 Vss.n1097 152.731
R3555 Vss.n1529 Vss.n1528 151.869
R3556 Vss.n1546 Vss.n1545 151.869
R3557 Vss.n1021 Vss.n405 151.869
R3558 Vss.n363 Vss.n362 151.869
R3559 Vss.n150 Vss.n100 151.869
R3560 Vss.n1167 Vss.n1143 151.869
R3561 Vss.n1708 Vss.n73 151.869
R3562 Vss.n1809 Vss.n75 151.869
R3563 Vss.n1425 Vss.n1424 151.869
R3564 Vss.n1472 Vss.n271 151.869
R3565 Vss.n1843 Vss.n1842 151.869
R3566 Vss.n1510 Vss.n251 151.869
R3567 Vss.n1509 Vss.n1508 151.869
R3568 Vss.n1728 Vss.n1727 151.869
R3569 Vss.n1332 Vss.n1331 151.869
R3570 Vss.n923 Vss.n921 151.869
R3571 Vss.n953 Vss.n458 151.869
R3572 Vss.n809 Vss.n390 151.869
R3573 Vss.n849 Vss.n757 151.869
R3574 Vss.n774 Vss.n15 151.869
R3575 Vss.n599 Vss.n598 151.869
R3576 Vss.n584 Vss.n583 151.751
R3577 Vss.n1038 Vss.n394 151.751
R3578 Vss.n996 Vss.n229 151.751
R3579 Vss.n1532 Vss.n230 151.751
R3580 Vss.n1534 Vss.n229 151.751
R3581 Vss.n1533 Vss.n1532 151.751
R3582 Vss.n941 Vss.n940 151.751
R3583 Vss.n979 Vss.n431 151.751
R3584 Vss.n960 Vss.n440 151.751
R3585 Vss.n940 Vss.n933 151.751
R3586 Vss.n979 Vss.n978 151.751
R3587 Vss.n1547 Vss.n216 151.751
R3588 Vss.n1594 Vss.n194 151.751
R3589 Vss.n1515 Vss.n195 151.751
R3590 Vss.n237 Vss.n206 151.751
R3591 Vss.n414 Vss.n48 151.751
R3592 Vss.n1164 Vss.n1163 151.751
R3593 Vss.n1145 Vss.n1144 151.751
R3594 Vss.n1453 Vss.n287 151.751
R3595 Vss.n350 Vss.n349 151.751
R3596 Vss.n340 Vss.n288 151.751
R3597 Vss.n1456 Vss.n1455 151.751
R3598 Vss.n1053 Vss.n368 151.751
R3599 Vss.n1276 Vss.n99 151.751
R3600 Vss.n1362 Vss.n1233 151.751
R3601 Vss.n1793 Vss.n99 151.751
R3602 Vss.n1776 Vss.n110 151.751
R3603 Vss.n1776 Vss.n111 151.751
R3604 Vss.n1776 Vss.n1775 151.751
R3605 Vss.n1227 Vss.n1226 151.751
R3606 Vss.n1228 Vss.n1132 151.751
R3607 Vss.n1315 Vss.n1120 151.751
R3608 Vss.n1471 Vss.n272 151.751
R3609 Vss.n1805 Vss.n87 151.751
R3610 Vss.n1268 Vss.n1267 151.751
R3611 Vss.n1805 Vss.n88 151.751
R3612 Vss.n1267 Vss.n1265 151.751
R3613 Vss.n1821 Vss.n70 151.751
R3614 Vss.n1820 Vss.n1819 151.751
R3615 Vss.n1504 Vss.n1503 151.751
R3616 Vss.n1819 Vss.n71 151.751
R3617 Vss.n1700 Vss.n1699 151.751
R3618 Vss.n1671 Vss.n1670 151.751
R3619 Vss.n1729 Vss.n169 151.751
R3620 Vss.n1330 Vss.n1329 151.751
R3621 Vss.n1817 Vss.n1816 151.751
R3622 Vss.n1411 Vss.n268 151.751
R3623 Vss.n1830 Vss.n1829 151.751
R3624 Vss.n1482 Vss.n261 151.751
R3625 Vss.n1830 Vss.n63 151.751
R3626 Vss.n1482 Vss.n267 151.751
R3627 Vss.n158 Vss.n157 151.751
R3628 Vss.n1362 Vss.n1361 151.751
R3629 Vss.n1344 Vss.n1343 151.751
R3630 Vss.n1362 Vss.n1234 151.751
R3631 Vss.n1023 Vss.n1022 151.751
R3632 Vss.n482 Vss.n480 151.751
R3633 Vss.n474 Vss.n449 151.751
R3634 Vss.n832 Vss.n831 151.751
R3635 Vss.n799 Vss.n798 151.751
R3636 Vss.n821 Vss.n820 151.751
R3637 Vss.n920 Vss.n919 151.751
R3638 Vss.n794 Vss.n759 151.751
R3639 Vss.n797 Vss.n758 151.751
R3640 Vss.n764 Vss.n23 151.751
R3641 Vss.n569 Vss.n568 151.751
R3642 Vss.n559 Vss.n558 151.751
R3643 Vss.n550 Vss.n549 151.751
R3644 Vss.n635 Vss.n503 151.751
R3645 Vss.n1869 Vss.n1868 151.751
R3646 Vss.n625 Vss.n504 151.751
R3647 Vss.n621 Vss.n620 151.751
R3648 Vss.n602 Vss.n601 151.751
R3649 Vss.n1065 Vss.n1064 147.727
R3650 Vss.n1073 Vss.n1072 147.727
R3651 Vss.n1451 Vss.n1450 147.727
R3652 Vss.n1193 Vss.n1188 147.727
R3653 Vss.n582 Vss.n574 147.727
R3654 Vss.n1881 Vss.n1880 147.727
R3655 Vss.n1867 Vss.n1866 147.727
R3656 Vss.n846 Vss.n392 147.727
R3657 Vss.n677 Vss.n676 147.727
R3658 Vss.n697 Vss.n696 147.727
R3659 Vss.n1093 Vss.n274 143.746
R3660 Vss.t97 Vss.t392 137.756
R3661 Vss.t392 Vss.t364 137.756
R3662 Vss.n1005 Vss.n229 135.501
R3663 Vss.n1806 Vss.n1805 135.501
R3664 Vss.n1831 Vss.n1830 135.501
R3665 Vss.n940 Vss.n939 135.501
R3666 Vss.n1348 Vss.n99 135.439
R3667 Vss.n1367 Vss.n1366 129.76
R3668 Vss.t636 Vss.n369 125.228
R3669 Vss.n1655 Vss.t261 124.305
R3670 Vss.t134 Vss.n109 120.279
R3671 Vss.n754 Vss.t587 119.157
R3672 Vss.n751 Vss.t587 119.157
R3673 Vss.n1641 Vss.n1621 118.222
R3674 Vss.n423 Vss.t613 115.856
R3675 Vss.n1004 Vss.t530 115.856
R3676 Vss.t526 Vss.n74 115.856
R3677 Vss.n86 Vss.t299 115.856
R3678 Vss.n1530 Vss.t564 115.856
R3679 Vss.n1832 Vss.t659 115.856
R3680 Vss.n1480 Vss.t560 115.856
R3681 Vss.n1475 Vss.t73 115.856
R3682 Vss.t605 Vss.n450 115.856
R3683 Vss.n938 Vss.t321 115.856
R3684 Vss.t523 Vss.n1281 115.802
R3685 Vss.n1349 Vss.t575 115.802
R3686 Vss.n1390 Vss.t337 114.944
R3687 Vss.t337 Vss.n1389 114.944
R3688 Vss.n1386 Vss.t104 114.944
R3689 Vss.n1466 Vss.t364 113.799
R3690 Vss.n751 Vss.n393 113.695
R3691 Vss.n1039 Vss.n1038 108.731
R3692 Vss.t385 Vss.t96 108.138
R3693 Vss.t166 Vss.t483 108.138
R3694 Vss.t159 Vss.t482 108.138
R3695 Vss.t363 Vss.t517 108.138
R3696 Vss.t206 Vss.t372 108.138
R3697 Vss.t210 Vss.t160 108.138
R3698 Vss.t209 Vss.t362 108.138
R3699 Vss.t545 Vss.t228 108.138
R3700 Vss.t437 Vss.n109 105.552
R3701 Vss.n755 Vss.n754 102.773
R3702 Vss.n1654 Vss.t263 101.704
R3703 Vss.t502 Vss.t373 99.0183
R3704 Vss.t153 Vss.t502 99.0183
R3705 Vss.n1389 Vss.n1386 97.7016
R3706 Vss.n327 Vss.t398 96.5949
R3707 Vss.n1195 Vss.t444 96.5352
R3708 Vss.t411 Vss.n16 96.5352
R3709 Vss.n580 Vss.t445 96.5352
R3710 Vss.n988 Vss.n229 95.5419
R3711 Vss.n1532 Vss.n231 95.5419
R3712 Vss.n940 Vss.n932 95.5419
R3713 Vss.n980 Vss.n979 95.5419
R3714 Vss.n1805 Vss.n1804 95.5419
R3715 Vss.n1267 Vss.n1266 95.5419
R3716 Vss.n1490 Vss.n252 95.5419
R3717 Vss.n1819 Vss.n72 95.5419
R3718 Vss.n1830 Vss.n62 95.5419
R3719 Vss.n1483 Vss.n1482 95.5419
R3720 Vss.n1243 Vss.n99 95.4017
R3721 Vss.n1362 Vss.n1232 95.4017
R3722 Vss.t613 Vss.t600 92.6849
R3723 Vss.t600 Vss.t530 92.6849
R3724 Vss.t647 Vss.t526 92.6849
R3725 Vss.t299 Vss.t647 92.6849
R3726 Vss.t564 Vss.t191 92.6849
R3727 Vss.t191 Vss.t659 92.6849
R3728 Vss.t275 Vss.t560 92.6849
R3729 Vss.t73 Vss.t275 92.6849
R3730 Vss.t539 Vss.t605 92.6849
R3731 Vss.t321 Vss.t539 92.6849
R3732 Vss.t542 Vss.t523 92.6419
R3733 Vss.t575 Vss.t542 92.6419
R3734 Vss.t96 Vss.t166 89.8983
R3735 Vss.t483 Vss.t159 89.8983
R3736 Vss.t482 Vss.t363 89.8983
R3737 Vss.t517 Vss.t161 89.8983
R3738 Vss.t162 Vss.t206 89.8983
R3739 Vss.t372 Vss.t210 89.8983
R3740 Vss.t160 Vss.t209 89.8983
R3741 Vss.t362 Vss.t545 89.8983
R3742 Vss.n1042 Vss.n1041 88.3958
R3743 Vss.n695 Vss.n506 87.3061
R3744 Vss.n695 Vss.n507 87.3061
R3745 Vss.n745 Vss.n492 87.3061
R3746 Vss.n745 Vss.n493 87.3061
R3747 Vss.n706 Vss.n500 87.3061
R3748 Vss.n706 Vss.n501 87.3061
R3749 Vss.n845 Vss.n840 87.3061
R3750 Vss.n845 Vss.n841 87.3061
R3751 Vss.n1882 Vss.n9 87.3061
R3752 Vss.n1882 Vss.n10 87.3061
R3753 Vss.n1014 Vss.n1012 87.3061
R3754 Vss.n1015 Vss.n1014 87.3061
R3755 Vss.n1173 Vss.n1168 87.3061
R3756 Vss.n1174 Vss.n1173 87.3061
R3757 Vss.n1187 Vss.n1181 87.3061
R3758 Vss.n1187 Vss.n1182 87.3061
R3759 Vss.n1074 Vss.n308 87.3061
R3760 Vss.n1074 Vss.n309 87.3061
R3761 Vss.n850 Vss.n749 87.3061
R3762 Vss.n851 Vss.n850 87.3061
R3763 Vss.n1374 Vss.n1126 87.3061
R3764 Vss.n1374 Vss.n1127 87.3061
R3765 Vss.n1788 Vss.n103 87.3061
R3766 Vss.n1788 Vss.n104 87.3061
R3767 Vss.n1391 Vss.n1390 86.8248
R3768 Vss.n1635 Vss.t385 80.7782
R3769 Vss.n1634 Vss.t227 80.7782
R3770 Vss.n1640 Vss.t367 80.7782
R3771 Vss.t228 Vss.n1639 80.7782
R3772 Vss.n1624 Vss.n1619 80.5005
R3773 Vss.n959 Vss.n958 76.452
R3774 Vss.n1776 Vss.n112 73.641
R3775 Vss.n849 Vss.n755 72.984
R3776 Vss.t227 Vss.t201 69.0524
R3777 Vss.t367 Vss.t583 69.0524
R3778 Vss.n672 Vss.n510 67.4727
R3779 Vss.n673 Vss.n510 67.4727
R3780 Vss.n710 Vss.n496 67.4727
R3781 Vss.n711 Vss.n496 67.4727
R3782 Vss.n515 Vss.n514 67.4727
R3783 Vss.n516 Vss.n514 67.4727
R3784 Vss.n1865 Vss.n25 67.4727
R3785 Vss.n1865 Vss.n26 67.4727
R3786 Vss.n570 Vss.n6 67.4727
R3787 Vss.n571 Vss.n6 67.4727
R3788 Vss.n1010 Vss.n301 67.4727
R3789 Vss.n1016 Vss.n301 67.4727
R3790 Vss.n1169 Vss.n1101 67.4727
R3791 Vss.n1172 Vss.n1101 67.4727
R3792 Vss.n1449 Vss.n290 67.4727
R3793 Vss.n1449 Vss.n291 67.4727
R3794 Vss.n1066 Vss.n305 67.4727
R3795 Vss.n1067 Vss.n305 67.4727
R3796 Vss.n747 Vss.n31 67.4727
R3797 Vss.n852 Vss.n31 67.4727
R3798 Vss.n1364 Vss.n1123 67.4727
R3799 Vss.n1365 Vss.n1123 67.4727
R3800 Vss.n1284 Vss.n1230 67.4727
R3801 Vss.n1285 Vss.n1230 67.4727
R3802 Vss.n1345 Vss.n1344 67.0503
R3803 Vss.n672 Vss.n506 66.5005
R3804 Vss.n673 Vss.n507 66.5005
R3805 Vss.n710 Vss.n492 66.5005
R3806 Vss.n711 Vss.n493 66.5005
R3807 Vss.n515 Vss.n500 66.5005
R3808 Vss.n516 Vss.n501 66.5005
R3809 Vss.n840 Vss.n25 66.5005
R3810 Vss.n841 Vss.n26 66.5005
R3811 Vss.n570 Vss.n9 66.5005
R3812 Vss.n571 Vss.n10 66.5005
R3813 Vss.n1012 Vss.n1010 66.5005
R3814 Vss.n1016 Vss.n1015 66.5005
R3815 Vss.n1169 Vss.n1168 66.5005
R3816 Vss.n1174 Vss.n1172 66.5005
R3817 Vss.n1181 Vss.n290 66.5005
R3818 Vss.n1182 Vss.n291 66.5005
R3819 Vss.n1066 Vss.n308 66.5005
R3820 Vss.n1067 Vss.n309 66.5005
R3821 Vss.n749 Vss.n747 66.5005
R3822 Vss.n852 Vss.n851 66.5005
R3823 Vss.n1364 Vss.n1126 66.5005
R3824 Vss.n1365 Vss.n1127 66.5005
R3825 Vss.n1284 Vss.n103 66.5005
R3826 Vss.n1285 Vss.n104 66.5005
R3827 Vss.n1666 Vss.n1606 65.5283
R3828 Vss.n1662 Vss.n1606 65.5283
R3829 Vss.n1662 Vss.n1607 65.5283
R3830 Vss.n1666 Vss.n1607 65.5283
R3831 Vss.n962 Vss.t361 63.4555
R3832 Vss.t45 Vss.n961 63.4555
R3833 Vss.n213 Vss.t14 63.4555
R3834 Vss.n1569 Vss.t480 63.4555
R3835 Vss.n1567 Vss.t571 63.4555
R3836 Vss.n1595 Vss.t143 63.4555
R3837 Vss.n960 Vss.n959 62.5094
R3838 Vss.n1346 Vss.n1345 61.7821
R3839 Vss.n1019 Vss.t59 61.7514
R3840 Vss.n1550 Vss.n212 61.0571
R3841 Vss.n977 Vss.n432 61.0571
R3842 Vss.n446 Vss.n441 61.0571
R3843 Vss.n1162 Vss.n1146 61.0571
R3844 Vss.n348 Vss.n341 61.0571
R3845 Vss.n1049 Vss.n1043 61.0571
R3846 Vss.n1752 Vss.n1751 61.0571
R3847 Vss.n138 Vss.n137 61.0571
R3848 Vss.n1815 Vss.n76 61.0571
R3849 Vss.n1342 Vss.n1301 61.0571
R3850 Vss.n830 Vss.n800 61.0571
R3851 Vss.n899 Vss.n483 61.0571
R3852 Vss.n783 Vss.n782 61.0571
R3853 Vss.n557 Vss.n551 61.0571
R3854 Vss.n619 Vss.n603 61.0571
R3855 Vss.n626 Vss.n530 61.0561
R3856 Vss.n578 Vss.n576 61.0561
R3857 Vss.n720 Vss.n717 61.0561
R3858 Vss.n1870 Vss.n21 61.0561
R3859 Vss.n1877 Vss.n17 61.0561
R3860 Vss.n863 Vss.n858 61.0561
R3861 Vss.n567 Vss.n562 61.0561
R3862 Vss.n586 Vss.n546 61.0561
R3863 Vss.n791 Vss.n765 61.0561
R3864 Vss.n775 Vss.n773 61.0561
R3865 Vss.n918 Vss.n468 61.0561
R3866 Vss.n822 Vss.n818 61.0561
R3867 Vss.n811 Vss.n808 61.0561
R3868 Vss.n1061 Vss.n384 61.0561
R3869 Vss.n890 Vss.n889 61.0561
R3870 Vss.n951 Vss.n459 61.0561
R3871 Vss.n457 Vss.n452 61.0561
R3872 Vss.n957 Vss.n955 61.0561
R3873 Vss.n937 Vss.n934 61.0561
R3874 Vss.n1024 Vss.n403 61.0561
R3875 Vss.n924 Vss.n467 61.0561
R3876 Vss.n1360 Vss.n1235 61.0561
R3877 Vss.n1334 Vss.n1333 61.0561
R3878 Vss.n1350 Vss.n1280 61.0561
R3879 Vss.n156 Vss.n131 61.0561
R3880 Vss.n1726 Vss.n172 61.0561
R3881 Vss.n1764 Vss.n123 61.0561
R3882 Vss.n1740 Vss.n161 61.0561
R3883 Vss.n1735 Vss.n1734 61.0561
R3884 Vss.n1695 Vss.n183 61.0561
R3885 Vss.n1603 Vss.n191 61.0561
R3886 Vss.n1591 Vss.n197 61.0561
R3887 Vss.n1511 Vss.n250 61.0561
R3888 Vss.n1479 Vss.n1476 61.0561
R3889 Vss.n1484 Vss.n260 61.0561
R3890 Vss.n266 Vss.n262 61.0561
R3891 Vss.n1828 Vss.n64 61.0561
R3892 Vss.n1833 Vss.n58 61.0561
R3893 Vss.n1412 Vss.n1409 61.0561
R3894 Vss.n1841 Vss.n49 61.0561
R3895 Vss.n1846 Vss.n46 61.0561
R3896 Vss.n1034 Vss.n398 61.0561
R3897 Vss.n1003 Vss.n424 61.0561
R3898 Vss.n989 Vss.n987 61.0561
R3899 Vss.n1535 Vss.n228 61.0561
R3900 Vss.n997 Vss.n995 61.0561
R3901 Vss.n981 Vss.n430 61.0561
R3902 Vss.n942 Vss.n931 61.0561
R3903 Vss.n238 Vss.n235 61.0561
R3904 Vss.n1544 Vss.n219 61.0561
R3905 Vss.n1557 Vss.n209 61.0561
R3906 Vss.n1596 Vss.n193 61.0561
R3907 Vss.n1570 Vss.n205 61.0561
R3908 Vss.n963 Vss.n439 61.0561
R3909 Vss.n1579 Vss.n200 61.0561
R3910 Vss.n1584 Vss.n1583 61.0561
R3911 Vss.n1563 Vss.n1561 61.0561
R3912 Vss.n1516 Vss.n246 61.0561
R3913 Vss.n1527 Vss.n233 61.0561
R3914 Vss.n421 Vss.n415 61.0561
R3915 Vss.n411 Vss.n407 61.0561
R3916 Vss.n1464 Vss.n281 61.0561
R3917 Vss.n1428 Vss.n1403 61.0561
R3918 Vss.n1423 Vss.n1406 61.0561
R3919 Vss.n1214 Vss.n1213 61.0561
R3920 Vss.n1205 Vss.n1204 61.0561
R3921 Vss.n1200 Vss.n1197 61.0561
R3922 Vss.n1225 Vss.n1133 61.0561
R3923 Vss.n1155 Vss.n1154 61.0561
R3924 Vss.n335 Vss.n329 61.0561
R3925 Vss.n1457 Vss.n286 61.0561
R3926 Vss.n353 Vss.n326 61.0561
R3927 Vss.n361 Vss.n318 61.0561
R3928 Vss.n1054 Vss.n388 61.0561
R3929 Vss.n1277 Vss.n1275 61.0561
R3930 Vss.n1245 Vss.n1244 61.0561
R3931 Vss.n1794 Vss.n98 61.0561
R3932 Vss.n1747 Vss.n1744 61.0561
R3933 Vss.n1760 Vss.n125 61.0561
R3934 Vss.n1774 Vss.n113 61.0561
R3935 Vss.n151 Vss.n148 61.0561
R3936 Vss.n1317 Vss.n1314 61.0561
R3937 Vss.n1397 Vss.n1396 61.0561
R3938 Vss.n1251 Vss.n1250 61.0561
R3939 Vss.n1803 Vss.n89 61.0561
R3940 Vss.n1264 Vss.n1260 61.0561
R3941 Vss.n1269 Vss.n1259 61.0561
R3942 Vss.n1491 Vss.n1489 61.0561
R3943 Vss.n1502 Vss.n253 61.0561
R3944 Vss.n1822 Vss.n69 61.0561
R3945 Vss.n1716 Vss.n1715 61.0561
R3946 Vss.n1709 Vss.n1706 61.0561
R3947 Vss.n1682 Vss.n1679 61.0561
R3948 Vss.n1686 Vss.n1678 61.0561
R3949 Vss.n1673 Vss.n1672 61.0561
R3950 Vss.n1701 Vss.n178 61.0561
R3951 Vss.n1328 Vss.n1307 61.0561
R3952 Vss.n1810 Vss.n82 61.0561
R3953 Vss.n479 Vss.n475 61.0561
R3954 Vss.n905 Vss.n473 61.0561
R3955 Vss.n597 Vss.n535 61.0561
R3956 Vss.n652 Vss.n523 61.0561
R3957 Vss.n643 Vss.n525 61.0561
R3958 Vss.n637 Vss.n634 61.0561
R3959 Vss.n611 Vss.n610 61.0561
R3960 Vss.n1289 Vss.t327 60.019
R3961 Vss.n1289 Vss.t573 60.019
R3962 Vss.t574 Vss.n1288 60.019
R3963 Vss.n1288 Vss.t90 60.019
R3964 Vss.t92 Vss.n1789 60.019
R3965 Vss.n1466 Vss.n1465 58.3972
R3966 Vss.n1469 Vss.n275 57.018
R3967 Vss.n1362 Vss.t327 54.0171
R3968 Vss.n1592 Vss.t285 53.4468
R3969 Vss.n196 Vss.t333 53.4468
R3970 Vss.n954 Vss.t604 53.4468
R3971 Vss.n958 Vss.t10 53.4468
R3972 Vss.n1346 Vss.t104 53.1614
R3973 Vss.t573 Vss.t574 51.0162
R3974 Vss.t361 Vss.t612 50.7645
R3975 Vss.t612 Vss.t45 50.7645
R3976 Vss.t14 Vss.t289 50.7645
R3977 Vss.t289 Vss.t480 50.7645
R3978 Vss.t571 Vss.t286 50.7645
R3979 Vss.t286 Vss.t143 50.7645
R3980 Vss.n645 Vss.t404 50.0912
R3981 Vss.n1344 Vss.n1300 45.4054
R3982 Vss.n904 Vss.n903 45.3808
R3983 Vss.n1299 Vss.n1295 44.1404
R3984 Vss.n666 Vss.n664 44.1404
R3985 Vss.n669 Vss.n513 44.1404
R3986 Vss.n733 Vss.n497 44.1394
R3987 Vss.n730 Vss.n4 44.1394
R3988 Vss.n724 Vss.n723 44.1394
R3989 Vss.n700 Vss.n699 44.1394
R3990 Vss.n868 Vss.n30 44.1394
R3991 Vss.n872 Vss.n871 44.1394
R3992 Vss.n875 Vss.n489 44.1394
R3993 Vss.n740 Vss.n739 44.1394
R3994 Vss.n753 Vss.n752 44.1394
R3995 Vss.n373 Vss.n302 44.1394
R3996 Vss.n377 Vss.n376 44.1394
R3997 Vss.n380 Vss.n36 44.1394
R3998 Vss.n1385 Vss.n1121 44.1394
R3999 Vss.n1388 Vss.n1106 44.1394
R4000 Vss.n1100 Vss.n1099 44.1394
R4001 Vss.n1096 Vss.n1094 44.1394
R4002 Vss.n1091 Vss.n296 44.1394
R4003 Vss.n313 Vss.n312 44.1394
R4004 Vss.n1191 Vss.n1190 44.1394
R4005 Vss.n1782 Vss.n106 44.1394
R4006 Vss.n661 Vss.n519 44.1394
R4007 Vss.t176 Vss.t285 42.7575
R4008 Vss.t333 Vss.t176 42.7575
R4009 Vss.t604 Vss.t47 42.7575
R4010 Vss.t47 Vss.t10 42.7575
R4011 Vss.n678 Vss.n518 42.4436
R4012 Vss.n911 Vss.t681 41.0041
R4013 Vss.n947 Vss.t677 41.0041
R4014 Vss.n163 Vss.t680 41.0041
R4015 Vss.n912 Vss.t679 40.8177
R4016 Vss.n1790 Vss.t90 38.0122
R4017 Vss.n903 Vss.n482 37.1047
R4018 Vss.t270 Vss.n273 36.1116
R4019 Vss.t88 Vss.n274 35.9369
R4020 Vss.n481 Vss.t127 35.0024
R4021 Vss.n952 Vss.t79 35.0024
R4022 Vss.n1377 Vss.t678 34.1066
R4023 Vss.t259 Vss.n1609 33.9022
R4024 Vss.n756 Vss.t615 31.7253
R4025 Vss.n904 Vss.t546 31.7253
R4026 Vss.n651 Vss.n650 30.7136
R4027 Vss.n1638 Vss.n1622 30.5283
R4028 Vss.n1638 Vss.n1637 30.5283
R4029 Vss.n1475 Vss.n1474 30.2237
R4030 Vss.n953 Vss.n450 30.2237
R4031 Vss.n1656 Vss.n1655 29.4859
R4032 Vss.t127 Vss.t291 28.002
R4033 Vss.t291 Vss.t79 28.002
R4034 Vss.n1654 Vss.n1653 27.3737
R4035 Vss.t161 Vss.n1634 27.3607
R4036 Vss.n1640 Vss.t162 27.3607
R4037 Vss.n912 Vss.t124 27.1302
R4038 Vss.n911 Vss.t131 26.9438
R4039 Vss.n947 Vss.t126 26.9438
R4040 Vss.n163 Vss.t133 26.9438
R4041 Vss.t615 Vss.t643 25.3804
R4042 Vss.t643 Vss.t546 25.3804
R4043 Vss.n1778 Vss.t350 24.9198
R4044 Vss.n1039 Vss.n393 24.8248
R4045 Vss.n649 Vss.t459 24.1401
R4046 Vss.n683 Vss.t459 24.1401
R4047 Vss.n683 Vss.t555 24.1401
R4048 Vss.t320 Vss.n682 24.1401
R4049 Vss.n682 Vss.t55 24.1401
R4050 Vss.n707 Vss.t57 24.1401
R4051 Vss.n714 Vss.t185 24.1401
R4052 Vss.t185 Vss.n713 24.1401
R4053 Vss.n713 Vss.t498 24.1401
R4054 Vss.t532 Vss.n709 24.1401
R4055 Vss.n709 Vss.t558 24.1401
R4056 Vss.n746 Vss.t556 24.1401
R4057 Vss.n855 Vss.t359 24.1401
R4058 Vss.t359 Vss.n854 24.1401
R4059 Vss.n854 Vss.t661 24.1401
R4060 Vss.n848 Vss.t663 24.1401
R4061 Vss.t64 Vss.n848 24.1401
R4062 Vss.t201 Vss.t373 20.8464
R4063 Vss.t583 Vss.t153 20.8464
R4064 Vss.n517 Vss.n506 20.8061
R4065 Vss.n517 Vss.n507 20.8061
R4066 Vss.n674 Vss.n672 20.8061
R4067 Vss.n674 Vss.n673 20.8061
R4068 Vss.n708 Vss.n492 20.8061
R4069 Vss.n708 Vss.n493 20.8061
R4070 Vss.n712 Vss.n710 20.8061
R4071 Vss.n712 Vss.n711 20.8061
R4072 Vss.n681 Vss.n500 20.8061
R4073 Vss.n681 Vss.n501 20.8061
R4074 Vss.n684 Vss.n515 20.8061
R4075 Vss.n684 Vss.n516 20.8061
R4076 Vss.n840 Vss.n839 20.8061
R4077 Vss.n841 Vss.n839 20.8061
R4078 Vss.n837 Vss.n25 20.8061
R4079 Vss.n837 Vss.n26 20.8061
R4080 Vss.n12 Vss.n9 20.8061
R4081 Vss.n12 Vss.n10 20.8061
R4082 Vss.n572 Vss.n570 20.8061
R4083 Vss.n572 Vss.n571 20.8061
R4084 Vss.n1012 Vss.n1011 20.8061
R4085 Vss.n1015 Vss.n1011 20.8061
R4086 Vss.n1017 Vss.n1010 20.8061
R4087 Vss.n1017 Vss.n1016 20.8061
R4088 Vss.n1175 Vss.n1168 20.8061
R4089 Vss.n1175 Vss.n1174 20.8061
R4090 Vss.n1171 Vss.n1169 20.8061
R4091 Vss.n1172 Vss.n1171 20.8061
R4092 Vss.n1183 Vss.n1181 20.8061
R4093 Vss.n1183 Vss.n1182 20.8061
R4094 Vss.n1178 Vss.n290 20.8061
R4095 Vss.n1178 Vss.n291 20.8061
R4096 Vss.n1068 Vss.n1066 20.8061
R4097 Vss.n1068 Vss.n1067 20.8061
R4098 Vss.n1070 Vss.n308 20.8061
R4099 Vss.n1070 Vss.n309 20.8061
R4100 Vss.n853 Vss.n747 20.8061
R4101 Vss.n853 Vss.n852 20.8061
R4102 Vss.n749 Vss.n748 20.8061
R4103 Vss.n851 Vss.n748 20.8061
R4104 Vss.n1128 Vss.n1126 20.8061
R4105 Vss.n1128 Vss.n1127 20.8061
R4106 Vss.n1366 Vss.n1364 20.8061
R4107 Vss.n1366 Vss.n1365 20.8061
R4108 Vss.n1613 Vss.n1606 20.8061
R4109 Vss.n1613 Vss.n1607 20.8061
R4110 Vss.n1287 Vss.n103 20.8061
R4111 Vss.n1287 Vss.n104 20.8061
R4112 Vss.n1290 Vss.n1284 20.8061
R4113 Vss.n1290 Vss.n1285 20.8061
R4114 Vss.t555 Vss.t320 20.5192
R4115 Vss.t55 Vss.t57 20.5192
R4116 Vss.t498 Vss.t532 20.5192
R4117 Vss.t558 Vss.t556 20.5192
R4118 Vss.t663 Vss.t661 20.5192
R4119 Vss.t66 Vss.t64 20.5192
R4120 Vss.n1669 Vss.n189 19.8869
R4121 Vss.n1376 Vss.t121 19.673
R4122 Vss.n1376 Vss.t128 19.4007
R4123 Vss.n1641 Vss.n1619 18.8616
R4124 Vss.n1624 Vss.n1621 18.8616
R4125 Vss.n1776 Vss.t350 18.5862
R4126 Vss.n518 Vss.n503 18.022
R4127 comparator_no_offsetcal_0.x3.avss Vss.n1649 17.8218
R4128 Vss.n1657 Vss.n1609 17.4164
R4129 Vss.n1628 comparator_no_offsetcal_0.x5.avss 16.7565
R4130 Vss.n962 Vss.n960 16.554
R4131 Vss.n1595 Vss.n1594 16.554
R4132 Vss.n1780 Vss.n102 16.1938
R4133 Vss.n196 Vss.n190 15.5696
R4134 Vss.n849 Vss.t66 14.6854
R4135 Vss.n1379 Vss.n1378 14.6135
R4136 Vss.n954 Vss.n953 13.943
R4137 Vss.n164 SARlogic_0.dffrs_13.d 13.7563
R4138 Vss.n914 SARlogic_0.dffrs_12.clk 13.599
R4139 Vss.n948 SARlogic_0.dffrs_12.d 13.599
R4140 Vss.n1790 Vss.t92 13.0045
R4141 Vss.n1642 Vss.n1620 11.0305
R4142 Vss.n482 Vss.n481 9.13142
R4143 Vss.n1628 Vss.n1625 9.05474
R4144 Vss.n165 Vss.n164 9.04466
R4145 Vss.n949 Vss.n948 9.04027
R4146 Vss.n965 Vss.n964 9.03475
R4147 Vss.n461 Vss.n460 9.03475
R4148 Vss.n544 Vss.n541 9.0005
R4149 Vss.n790 Vss.n789 9.0005
R4150 Vss.n859 Vss.n20 9.0005
R4151 Vss.n1874 Vss.n1873 9.0005
R4152 Vss.n817 Vss.n816 9.0005
R4153 Vss.n892 Vss.n891 9.0005
R4154 Vss.n1026 Vss.n401 9.0005
R4155 Vss.n263 Vss.n257 9.0005
R4156 Vss.n966 Vss.n211 9.0005
R4157 Vss.n973 Vss.n972 9.0005
R4158 Vss.n445 Vss.n444 9.0005
R4159 Vss.n456 Vss.n434 9.0005
R4160 Vss.n455 Vss.n453 9.0005
R4161 Vss.n1520 Vss.n1519 9.0005
R4162 Vss.n1525 Vss.n1523 9.0005
R4163 Vss.n420 Vss.n419 9.0005
R4164 Vss.n45 Vss.n42 9.0005
R4165 Vss.n409 Vss.n400 9.0005
R4166 Vss.n1408 Vss.n1407 9.0005
R4167 Vss.n53 Vss.n51 9.0005
R4168 Vss.n1402 Vss.n1111 9.0005
R4169 Vss.n1135 Vss.n1134 9.0005
R4170 Vss.n1161 Vss.n1160 9.0005
R4171 Vss.n1148 Vss.n1136 9.0005
R4172 Vss.n330 Vss.n282 9.0005
R4173 Vss.n347 Vss.n346 9.0005
R4174 Vss.n345 Vss.n343 9.0005
R4175 Vss.n360 Vss.n319 9.0005
R4176 Vss.n359 Vss.n357 9.0005
R4177 Vss.n355 Vss.n354 9.0005
R4178 Vss.n324 Vss.n323 9.0005
R4179 Vss.n1462 Vss.n1461 9.0005
R4180 Vss.n331 Vss.n285 9.0005
R4181 Vss.n1460 Vss.n1459 9.0005
R4182 Vss.n1044 Vss.n385 9.0005
R4183 Vss.n1045 Vss.n387 9.0005
R4184 Vss.n1057 Vss.n1056 9.0005
R4185 Vss.n1059 Vss.n1058 9.0005
R4186 Vss.n115 Vss.n114 9.0005
R4187 Vss.n1754 Vss.n117 9.0005
R4188 Vss.n142 Vss.n141 9.0005
R4189 Vss.n140 Vss.n116 9.0005
R4190 Vss.n1772 Vss.n1771 9.0005
R4191 Vss.n146 Vss.n145 9.0005
R4192 Vss.n1211 Vss.n1210 9.0005
R4193 Vss.n1209 Vss.n1208 9.0005
R4194 Vss.n1207 Vss.n1139 9.0005
R4195 Vss.n1217 Vss.n1216 9.0005
R4196 Vss.n1223 Vss.n1222 9.0005
R4197 Vss.n1157 Vss.n1156 9.0005
R4198 Vss.n1151 Vss.n1150 9.0005
R4199 Vss.n1261 Vss.n92 9.0005
R4200 Vss.n1720 Vss.n1719 9.0005
R4201 Vss.n1704 Vss.n175 9.0005
R4202 Vss.n1417 Vss.n77 9.0005
R4203 Vss.n1421 Vss.n1419 9.0005
R4204 Vss.n1341 Vss.n1340 9.0005
R4205 Vss.n1303 Vss.n1238 9.0005
R4206 Vss.n1337 Vss.n1336 9.0005
R4207 Vss.n1237 Vss.n1236 9.0005
R4208 Vss.n1358 Vss.n1357 9.0005
R4209 Vss.n1273 Vss.n1239 9.0005
R4210 Vss.n1248 Vss.n1247 9.0005
R4211 Vss.n154 Vss.n153 9.0005
R4212 Vss.n153 Vss.n152 9.0005
R4213 Vss.n133 Vss.n96 9.0005
R4214 Vss.n1738 Vss.n1737 9.0005
R4215 Vss.n1739 Vss.n1738 9.0005
R4216 Vss.n1758 Vss.n1756 9.0005
R4217 Vss.n1756 Vss.n1755 9.0005
R4218 Vss.n1693 Vss.n1691 9.0005
R4219 Vss.n1691 Vss.n166 9.0005
R4220 Vss.n1676 Vss.n122 9.0005
R4221 Vss.n1759 Vss.n122 9.0005
R4222 Vss.n1718 Vss.n173 9.0005
R4223 Vss.n1725 Vss.n173 9.0005
R4224 Vss.n1262 Vss.n93 9.0005
R4225 Vss.n1724 Vss.n1722 9.0005
R4226 Vss.n134 Vss.n132 9.0005
R4227 Vss.n1796 Vss.n1795 9.0005
R4228 Vss.n1801 Vss.n1799 9.0005
R4229 Vss.n1242 Vss.n91 9.0005
R4230 Vss.n1272 Vss.n1271 9.0005
R4231 Vss.n1279 Vss.n1278 9.0005
R4232 Vss.n1326 Vss.n1325 9.0005
R4233 Vss.n1324 Vss.n1306 9.0005
R4234 Vss.n1312 Vss.n1311 9.0005
R4235 Vss.n1309 Vss.n80 9.0005
R4236 Vss.n1322 Vss.n1308 9.0005
R4237 Vss.n1319 Vss.n1318 9.0005
R4238 Vss.n1399 Vss.n1398 9.0005
R4239 Vss.n1813 Vss.n1812 9.0005
R4240 Vss.n1812 Vss.n1811 9.0005
R4241 Vss.n1113 Vss.n1112 9.0005
R4242 Vss.n1487 Vss.n90 9.0005
R4243 Vss.n1802 Vss.n90 9.0005
R4244 Vss.n1257 Vss.n67 9.0005
R4245 Vss.n1258 Vss.n1257 9.0005
R4246 Vss.n1711 Vss.n1703 9.0005
R4247 Vss.n1711 Vss.n1710 9.0005
R4248 Vss.n1500 Vss.n1498 9.0005
R4249 Vss.n1601 Vss.n184 9.0005
R4250 Vss.n1694 Vss.n184 9.0005
R4251 Vss.n1688 Vss.n1675 9.0005
R4252 Vss.n1688 Vss.n1687 9.0005
R4253 Vss.n1599 Vss.n1598 9.0005
R4254 Vss.n1602 Vss.n1599 9.0005
R4255 Vss.n1587 Vss.n1586 9.0005
R4256 Vss.n1587 Vss.n187 9.0005
R4257 Vss.n1518 Vss.n1513 9.0005
R4258 Vss.n1513 Vss.n1512 9.0005
R4259 Vss.n264 Vss.n258 9.0005
R4260 Vss.n254 Vss.n248 9.0005
R4261 Vss.n255 Vss.n177 9.0005
R4262 Vss.n1501 Vss.n1496 9.0005
R4263 Vss.n1493 Vss.n1486 9.0005
R4264 Vss.n1493 Vss.n1492 9.0005
R4265 Vss.n1826 Vss.n1824 9.0005
R4266 Vss.n1824 Vss.n1823 9.0005
R4267 Vss.n1415 Vss.n1414 9.0005
R4268 Vss.n1422 Vss.n1415 9.0005
R4269 Vss.n1431 Vss.n1430 9.0005
R4270 Vss.n1839 Vss.n52 9.0005
R4271 Vss.n1840 Vss.n1839 9.0005
R4272 Vss.n1849 Vss.n1848 9.0005
R4273 Vss.n985 Vss.n984 9.0005
R4274 Vss.n984 Vss.n259 9.0005
R4275 Vss.n993 Vss.n57 9.0005
R4276 Vss.n1827 Vss.n57 9.0005
R4277 Vss.n241 Vss.n240 9.0005
R4278 Vss.n1526 Vss.n241 9.0005
R4279 Vss.n242 Vss.n226 9.0005
R4280 Vss.n1573 Vss.n1572 9.0005
R4281 Vss.n1573 Vss.n192 9.0005
R4282 Vss.n1575 Vss.n202 9.0005
R4283 Vss.n1575 Vss.n199 9.0005
R4284 Vss.n437 Vss.n436 9.0005
R4285 Vss.n436 Vss.n204 9.0005
R4286 Vss.n1553 Vss.n1552 9.0005
R4287 Vss.n1553 Vss.n207 9.0005
R4288 Vss.n443 Vss.n220 9.0005
R4289 Vss.n1543 Vss.n220 9.0005
R4290 Vss.n975 Vss.n974 9.0005
R4291 Vss.n1542 Vss.n1540 9.0005
R4292 Vss.n234 Vss.n223 9.0005
R4293 Vss.n1537 Vss.n1536 9.0005
R4294 Vss.n991 Vss.n983 9.0005
R4295 Vss.n991 Vss.n990 9.0005
R4296 Vss.n999 Vss.n425 9.0005
R4297 Vss.n999 Vss.n998 9.0005
R4298 Vss.n408 Vss.n401 9.0005
R4299 Vss.n1032 Vss.n1030 9.0005
R4300 Vss.n1033 Vss.n399 9.0005
R4301 Vss.n1028 Vss.n1027 9.0005
R4302 Vss.n465 Vss.n464 9.0005
R4303 Vss.n829 Vss.n828 9.0005
R4304 Vss.n827 Vss.n802 9.0005
R4305 Vss.n825 Vss.n824 9.0005
R4306 Vss.n807 Vss.n806 9.0005
R4307 Vss.n814 Vss.n813 9.0005
R4308 Vss.n485 Vss.n484 9.0005
R4309 Vss.n897 Vss.n896 9.0005
R4310 Vss.n894 Vss.n469 9.0005
R4311 Vss.n478 Vss.n472 9.0005
R4312 Vss.n477 Vss.n462 9.0005
R4313 Vss.n916 Vss.n915 9.0005
R4314 Vss.n886 Vss.n885 9.0005
R4315 Vss.n429 Vss.n428 9.0005
R4316 Vss.n944 Vss.n943 9.0005
R4317 Vss.n926 Vss.n925 9.0005
R4318 Vss.n861 Vss.n860 9.0005
R4319 Vss.n1872 Vss.n22 9.0005
R4320 Vss.n781 Vss.n780 9.0005
R4321 Vss.n786 Vss.n785 9.0005
R4322 Vss.n788 Vss.n767 9.0005
R4323 Vss.n777 Vss.n776 9.0005
R4324 Vss.n771 Vss.n770 9.0005
R4325 Vss.n556 Vss.n555 9.0005
R4326 Vss.n554 Vss.n553 9.0005
R4327 Vss.n596 Vss.n536 9.0005
R4328 Vss.n595 Vss.n593 9.0005
R4329 Vss.n563 Vss.n538 9.0005
R4330 Vss.n565 Vss.n564 9.0005
R4331 Vss.n588 Vss.n587 9.0005
R4332 Vss.n639 Vss.n638 9.0005
R4333 Vss.n618 Vss.n617 9.0005
R4334 Vss.n605 Vss.n527 9.0005
R4335 Vss.n608 Vss.n607 9.0005
R4336 Vss.n614 Vss.n613 9.0005
R4337 Vss.n529 Vss.n528 9.0005
R4338 Vss.n629 Vss.n628 9.0005
R4339 Vss.n632 Vss.n521 9.0005
R4340 Vss.n522 Vss.n520 9.0005
R4341 Vss.n655 Vss.n654 9.0005
R4342 Vss.n1653 Vss.t264 8.70131
R4343 Vss.n849 Vss.n756 8.27654
R4344 Vss.n1331 Vss.n1330 8.08508
R4345 Vss.n1304 Vss.n1108 8.05717
R4346 Vss.n1648 Vss.n1647 7.7564
R4347 Vss.n1629 Vss.n1623 7.59387
R4348 Vss.n1507 Vss.n1506 7.29099
R4349 Vss.n576 Vss.n542 6.9012
R4350 Vss.n1877 Vss.n1876 6.9012
R4351 Vss.n935 Vss.n934 6.9012
R4352 Vss.n1352 Vss.n1280 6.9012
R4353 Vss.n1766 Vss.n123 6.9012
R4354 Vss.n1591 Vss.n1590 6.9012
R4355 Vss.n1479 Vss.n1478 6.9012
R4356 Vss.n1835 Vss.n58 6.9012
R4357 Vss.n1001 Vss.n424 6.9012
R4358 Vss.n1555 Vss.n209 6.9012
R4359 Vss.n955 Vss.n435 6.9012
R4360 Vss.n1577 Vss.n200 6.9012
R4361 Vss.n333 Vss.n329 6.9012
R4362 Vss.n1047 Vss.n1043 6.9012
R4363 Vss.n1745 Vss.n1744 6.9012
R4364 Vss.n1198 Vss.n1197 6.9012
R4365 Vss.n1253 Vss.n1250 6.9012
R4366 Vss.n1680 Vss.n1679 6.9012
R4367 Vss.n907 Vss.n473 6.9012
R4368 Vss.n641 Vss.n525 6.9012
R4369 Vss.n718 Vss.n717 6.90005
R4370 Vss.n1631 Vss.n1630 6.64904
R4371 Vss.n1658 Vss.n1610 6.5795
R4372 Vss.n1612 Vss.n1611 6.5795
R4373 Vss.n530 Vss.n529 6.46296
R4374 Vss.n563 Vss.n562 6.46296
R4375 Vss.n587 Vss.n586 6.46296
R4376 Vss.n791 Vss.n790 6.46296
R4377 Vss.n1873 Vss.n21 6.46296
R4378 Vss.n469 Vss.n468 6.46296
R4379 Vss.n818 Vss.n817 6.46296
R4380 Vss.n1027 Vss.n403 6.46296
R4381 Vss.n1236 Vss.n1235 6.46296
R4382 Vss.n1333 Vss.n1306 6.46296
R4383 Vss.n132 Vss.n131 6.46296
R4384 Vss.n1726 Vss.n1725 6.46296
R4385 Vss.n1512 Vss.n1511 6.46296
R4386 Vss.n1828 Vss.n1827 6.46296
R4387 Vss.n998 Vss.n997 6.46296
R4388 Vss.n943 Vss.n942 6.46296
R4389 Vss.n235 Vss.n234 6.46296
R4390 Vss.n1544 Vss.n1543 6.46296
R4391 Vss.n212 Vss.n211 6.46296
R4392 Vss.n446 Vss.n445 6.46296
R4393 Vss.n457 Vss.n456 6.46296
R4394 Vss.n1583 Vss.n199 6.46296
R4395 Vss.n1561 Vss.n207 6.46296
R4396 Vss.n1519 Vss.n246 6.46296
R4397 Vss.n1527 Vss.n1526 6.46296
R4398 Vss.n421 Vss.n420 6.46296
R4399 Vss.n408 Vss.n407 6.46296
R4400 Vss.n1409 Vss.n1408 6.46296
R4401 Vss.n1841 Vss.n1840 6.46296
R4402 Vss.n1134 Vss.n1133 6.46296
R4403 Vss.n354 Vss.n353 6.46296
R4404 Vss.n361 Vss.n360 6.46296
R4405 Vss.n286 Vss.n285 6.46296
R4406 Vss.n388 Vss.n387 6.46296
R4407 Vss.n1278 Vss.n1277 6.46296
R4408 Vss.n1760 Vss.n1759 6.46296
R4409 Vss.n114 Vss.n113 6.46296
R4410 Vss.n1755 Vss.n1751 6.46296
R4411 Vss.n152 Vss.n151 6.46296
R4412 Vss.n1208 Vss.n1204 6.46296
R4413 Vss.n1156 Vss.n1155 6.46296
R4414 Vss.n1259 Vss.n1258 6.46296
R4415 Vss.n1823 Vss.n1822 6.46296
R4416 Vss.n1719 Vss.n1715 6.46296
R4417 Vss.n1710 Vss.n1709 6.46296
R4418 Vss.n1687 Vss.n1686 6.46296
R4419 Vss.n1672 Vss.n187 6.46296
R4420 Vss.n178 Vss.n177 6.46296
R4421 Vss.n1308 Vss.n1307 6.46296
R4422 Vss.n1811 Vss.n1810 6.46296
R4423 Vss.n77 Vss.n76 6.46296
R4424 Vss.n1423 Vss.n1422 6.46296
R4425 Vss.n925 Vss.n924 6.46296
R4426 Vss.n479 Vss.n478 6.46296
R4427 Vss.n808 Vss.n807 6.46296
R4428 Vss.n484 Vss.n483 6.46296
R4429 Vss.n776 Vss.n775 6.46296
R4430 Vss.n597 Vss.n596 6.46296
R4431 Vss.n638 Vss.n637 6.46296
R4432 Vss.n610 Vss.n608 6.46296
R4433 Vss.n859 Vss.n858 6.4618
R4434 Vss.n891 Vss.n890 6.4618
R4435 Vss.n460 Vss.n459 6.4618
R4436 Vss.n1734 Vss.n166 6.4618
R4437 Vss.n1695 Vss.n1694 6.4618
R4438 Vss.n1603 Vss.n1602 6.4618
R4439 Vss.n260 Vss.n259 6.4618
R4440 Vss.n263 Vss.n262 6.4618
R4441 Vss.n1034 Vss.n1033 6.4618
R4442 Vss.n990 Vss.n989 6.4618
R4443 Vss.n1536 Vss.n1535 6.4618
R4444 Vss.n430 Vss.n429 6.4618
R4445 Vss.n193 Vss.n192 6.4618
R4446 Vss.n205 Vss.n204 6.4618
R4447 Vss.n973 Vss.n432 6.4618
R4448 Vss.n964 Vss.n963 6.4618
R4449 Vss.n46 Vss.n45 6.4618
R4450 Vss.n1403 Vss.n1402 6.4618
R4451 Vss.n1162 Vss.n1161 6.4618
R4452 Vss.n282 Vss.n281 6.4618
R4453 Vss.n348 Vss.n347 6.4618
R4454 Vss.n385 Vss.n384 6.4618
R4455 Vss.n1244 Vss.n1242 6.4618
R4456 Vss.n1795 Vss.n1794 6.4618
R4457 Vss.n1740 Vss.n1739 6.4618
R4458 Vss.n141 Vss.n137 6.4618
R4459 Vss.n1213 Vss.n1211 6.4618
R4460 Vss.n1318 Vss.n1317 6.4618
R4461 Vss.n1398 Vss.n1397 6.4618
R4462 Vss.n1803 Vss.n1802 6.4618
R4463 Vss.n1261 Vss.n1260 6.4618
R4464 Vss.n1492 Vss.n1491 6.4618
R4465 Vss.n1502 Vss.n1501 6.4618
R4466 Vss.n1342 Vss.n1341 6.4618
R4467 Vss.n830 Vss.n829 6.4618
R4468 Vss.n782 Vss.n781 6.4618
R4469 Vss.n557 Vss.n556 6.4618
R4470 Vss.n523 Vss.n522 6.4618
R4471 Vss.n619 Vss.n618 6.4618
R4472 Vss.n1647 Vss.n1616 6.33584
R4473 Vss.n1636 Vss.n1623 6.32806
R4474 Vss.n1642 Vss.n1641 6.23383
R4475 SARlogic_0.dffrs_12.nand3_1.A Vss.n911 5.7755
R4476 SARlogic_0.dffrs_12.nand3_8.A Vss.n947 5.7755
R4477 SARlogic_0.dffrs_13.nand3_8.A Vss.n163 5.7755
R4478 SARlogic_0.dffrs_12.nand3_6.B Vss.n912 5.47979
R4479 Vss.n1876 Vss.n18 5.47239
R4480 Vss.n936 Vss.n935 5.47239
R4481 Vss.n1352 Vss.n1351 5.47239
R4482 Vss.n1766 Vss.n1765 5.47239
R4483 Vss.n1590 Vss.n1589 5.47239
R4484 Vss.n1478 Vss.n1477 5.47239
R4485 Vss.n1835 Vss.n1834 5.47239
R4486 Vss.n1002 Vss.n1001 5.47239
R4487 Vss.n1556 Vss.n1555 5.47239
R4488 Vss.n956 Vss.n435 5.47239
R4489 Vss.n1578 Vss.n1577 5.47239
R4490 Vss.n334 Vss.n333 5.47239
R4491 Vss.n1048 Vss.n1047 5.47239
R4492 Vss.n1746 Vss.n1745 5.47239
R4493 Vss.n1199 Vss.n1198 5.47239
R4494 Vss.n1253 Vss.n1252 5.47239
R4495 Vss.n1681 Vss.n1680 5.47239
R4496 Vss.n907 Vss.n906 5.47239
R4497 Vss.n577 Vss.n542 5.47239
R4498 Vss.n719 Vss.n718 5.47239
R4499 Vss.n642 Vss.n641 5.47239
R4500 Vss.n1378 Vss.n1377 5.18044
R4501 Vss.n628 Vss.n627 5.03414
R4502 Vss.n566 Vss.n565 5.03414
R4503 Vss.n545 Vss.n544 5.03414
R4504 Vss.n772 Vss.n771 5.03414
R4505 Vss.n767 Vss.n766 5.03414
R4506 Vss.n862 Vss.n861 5.03414
R4507 Vss.n1872 Vss.n1871 5.03414
R4508 Vss.n917 Vss.n916 5.03414
R4509 Vss.n813 Vss.n812 5.03414
R4510 Vss.n824 Vss.n823 5.03414
R4511 Vss.n887 Vss.n886 5.03414
R4512 Vss.n950 Vss.n949 5.03414
R4513 Vss.n466 Vss.n465 5.03414
R4514 Vss.n1026 Vss.n1025 5.03414
R4515 Vss.n1359 Vss.n1358 5.03414
R4516 Vss.n1336 Vss.n1335 5.03414
R4517 Vss.n155 Vss.n154 5.03414
R4518 Vss.n1724 Vss.n1723 5.03414
R4519 Vss.n1737 Vss.n1736 5.03414
R4520 Vss.n1693 Vss.n1692 5.03414
R4521 Vss.n1601 Vss.n1600 5.03414
R4522 Vss.n249 Vss.n248 5.03414
R4523 Vss.n1486 Vss.n1485 5.03414
R4524 Vss.n265 Vss.n264 5.03414
R4525 Vss.n1826 Vss.n1825 5.03414
R4526 Vss.n1032 Vss.n1031 5.03414
R4527 Vss.n986 Vss.n985 5.03414
R4528 Vss.n227 Vss.n226 5.03414
R4529 Vss.n994 Vss.n993 5.03414
R4530 Vss.n983 Vss.n982 5.03414
R4531 Vss.n930 Vss.n425 5.03414
R4532 Vss.n240 Vss.n239 5.03414
R4533 Vss.n1542 Vss.n1541 5.03414
R4534 Vss.n1598 Vss.n1597 5.03414
R4535 Vss.n1572 Vss.n1571 5.03414
R4536 Vss.n438 Vss.n437 5.03414
R4537 Vss.n1552 Vss.n1551 5.03414
R4538 Vss.n976 Vss.n975 5.03414
R4539 Vss.n443 Vss.n442 5.03414
R4540 Vss.n455 Vss.n454 5.03414
R4541 Vss.n1586 Vss.n1585 5.03414
R4542 Vss.n1562 Vss.n202 5.03414
R4543 Vss.n1525 Vss.n1524 5.03414
R4544 Vss.n1518 Vss.n1517 5.03414
R4545 Vss.n410 Vss.n409 5.03414
R4546 Vss.n413 Vss.n52 5.03414
R4547 Vss.n1848 Vss.n1847 5.03414
R4548 Vss.n1430 Vss.n1429 5.03414
R4549 Vss.n1414 Vss.n1413 5.03414
R4550 Vss.n51 Vss.n50 5.03414
R4551 Vss.n1421 Vss.n1420 5.03414
R4552 Vss.n1152 Vss.n1151 5.03414
R4553 Vss.n1224 Vss.n1223 5.03414
R4554 Vss.n1148 Vss.n1147 5.03414
R4555 Vss.n1459 Vss.n1458 5.03414
R4556 Vss.n1463 Vss.n1462 5.03414
R4557 Vss.n325 Vss.n324 5.03414
R4558 Vss.n359 Vss.n358 5.03414
R4559 Vss.n343 Vss.n342 5.03414
R4560 Vss.n1060 Vss.n1059 5.03414
R4561 Vss.n1056 Vss.n1055 5.03414
R4562 Vss.n1274 Vss.n1273 5.03414
R4563 Vss.n1247 Vss.n1246 5.03414
R4564 Vss.n97 Vss.n96 5.03414
R4565 Vss.n1758 Vss.n1757 5.03414
R4566 Vss.n147 Vss.n146 5.03414
R4567 Vss.n1773 Vss.n1772 5.03414
R4568 Vss.n1754 Vss.n1753 5.03414
R4569 Vss.n165 Vss.n162 5.03414
R4570 Vss.n140 Vss.n139 5.03414
R4571 Vss.n1216 Vss.n1215 5.03414
R4572 Vss.n1207 Vss.n1206 5.03414
R4573 Vss.n1313 Vss.n1312 5.03414
R4574 Vss.n1114 Vss.n1113 5.03414
R4575 Vss.n1801 Vss.n1800 5.03414
R4576 Vss.n1263 Vss.n1262 5.03414
R4577 Vss.n1271 Vss.n1270 5.03414
R4578 Vss.n1488 Vss.n1487 5.03414
R4579 Vss.n1500 Vss.n1499 5.03414
R4580 Vss.n68 Vss.n67 5.03414
R4581 Vss.n1705 Vss.n1704 5.03414
R4582 Vss.n1718 Vss.n1717 5.03414
R4583 Vss.n1677 Vss.n1676 5.03414
R4584 Vss.n1675 Vss.n1674 5.03414
R4585 Vss.n1703 Vss.n1702 5.03414
R4586 Vss.n1327 Vss.n1326 5.03414
R4587 Vss.n81 Vss.n80 5.03414
R4588 Vss.n1814 Vss.n1813 5.03414
R4589 Vss.n1303 Vss.n1302 5.03414
R4590 Vss.n477 Vss.n476 5.03414
R4591 Vss.n802 Vss.n801 5.03414
R4592 Vss.n898 Vss.n897 5.03414
R4593 Vss.n785 Vss.n784 5.03414
R4594 Vss.n595 Vss.n594 5.03414
R4595 Vss.n553 Vss.n552 5.03414
R4596 Vss.n654 Vss.n653 5.03414
R4597 Vss.n633 Vss.n632 5.03414
R4598 Vss.n613 Vss.n612 5.03414
R4599 Vss.n605 Vss.n604 5.03414
R4600 Vss.n1777 Vss.t351 4.8595
R4601 Vss.n867 Vss.t138 4.84702
R4602 Vss.n866 Vss.t252 4.84702
R4603 Vss.n372 Vss.t570 4.84702
R4604 Vss.n371 Vss.t136 4.84702
R4605 Vss.n295 Vss.t266 4.84702
R4606 Vss.n1095 Vss.t89 4.84702
R4607 Vss.n1298 Vss.t42 4.84702
R4608 Vss.n1296 Vss.t105 4.84702
R4609 Vss.n668 Vss.t513 4.84702
R4610 Vss.n665 Vss.t230 4.84702
R4611 Vss.n727 Vss.t117 4.84702
R4612 Vss.n729 Vss.t4 4.84702
R4613 Vss.n1776 Vss.n108 4.79462
R4614 Vss.n627 Vss.t578 4.7885
R4615 Vss.n738 Vss.t102 4.7885
R4616 Vss.n719 Vss.t236 4.7885
R4617 Vss.n577 Vss.t656 4.7885
R4618 Vss.n566 Vss.t200 4.7885
R4619 Vss.n545 Vss.t146 4.7885
R4620 Vss.n7 Vss.t76 4.7885
R4621 Vss.n8 Vss.t226 4.7885
R4622 Vss.n1883 Vss.t475 4.7885
R4623 Vss.n772 Vss.t427 4.7885
R4624 Vss.n766 Vss.t485 4.7885
R4625 Vss.n862 Vss.t87 4.7885
R4626 Vss.n1871 Vss.t168 4.7885
R4627 Vss.n18 Vss.t488 4.7885
R4628 Vss.n917 Vss.t33 4.7885
R4629 Vss.n812 Vss.t397 4.7885
R4630 Vss.n823 Vss.t243 4.7885
R4631 Vss.n887 Vss.t26 4.7885
R4632 Vss.n950 Vss.t80 4.7885
R4633 Vss.n936 Vss.t322 4.7885
R4634 Vss.n466 Vss.t193 4.7885
R4635 Vss.n1025 Vss.t269 4.7885
R4636 Vss.n1359 Vss.t324 4.7885
R4637 Vss.n1335 Vss.t306 4.7885
R4638 Vss.n1351 Vss.t576 4.7885
R4639 Vss.n155 Vss.t273 4.7885
R4640 Vss.n1723 Vss.t429 4.7885
R4641 Vss.n1765 Vss.t344 4.7885
R4642 Vss.n1736 Vss.t219 4.7885
R4643 Vss.n1692 Vss.t141 4.7885
R4644 Vss.n1600 Vss.t175 4.7885
R4645 Vss.n1589 Vss.t334 4.7885
R4646 Vss.n249 Vss.t423 4.7885
R4647 Vss.n1477 Vss.t74 4.7885
R4648 Vss.n1485 Vss.t190 4.7885
R4649 Vss.n265 Vss.t415 4.7885
R4650 Vss.n1825 Vss.t634 4.7885
R4651 Vss.n1834 Vss.t660 4.7885
R4652 Vss.n1031 Vss.t157 4.7885
R4653 Vss.n1002 Vss.t531 4.7885
R4654 Vss.n986 Vss.t602 4.7885
R4655 Vss.n227 Vss.t391 4.7885
R4656 Vss.n994 Vss.t180 4.7885
R4657 Vss.n982 Vss.t538 4.7885
R4658 Vss.n930 Vss.t308 4.7885
R4659 Vss.n239 Vss.t622 4.7885
R4660 Vss.n1541 Vss.t421 4.7885
R4661 Vss.n1556 Vss.t357 4.7885
R4662 Vss.n1597 Vss.t144 4.7885
R4663 Vss.n1571 Vss.t481 4.7885
R4664 Vss.n438 Vss.t46 4.7885
R4665 Vss.n1551 Vss.t223 4.7885
R4666 Vss.n956 Vss.t11 4.7885
R4667 Vss.n976 Vss.t417 4.7885
R4668 Vss.n442 Vss.t304 4.7885
R4669 Vss.n454 Vss.t425 4.7885
R4670 Vss.n1578 Vss.t16 4.7885
R4671 Vss.n1585 Vss.t582 4.7885
R4672 Vss.n1562 Vss.t467 4.7885
R4673 Vss.n1524 Vss.t442 4.7885
R4674 Vss.n1517 Vss.t31 4.7885
R4675 Vss.n410 Vss.t196 4.7885
R4676 Vss.n413 Vss.t254 4.7885
R4677 Vss.n1847 Vss.t198 4.7885
R4678 Vss.n1429 Vss.t383 4.7885
R4679 Vss.n1413 Vss.t302 4.7885
R4680 Vss.n50 Vss.t381 4.7885
R4681 Vss.n1420 Vss.t35 4.7885
R4682 Vss.n1152 Vss.t409 4.7885
R4683 Vss.n1224 Vss.t346 4.7885
R4684 Vss.n1147 Vss.t456 4.7885
R4685 Vss.n1177 Vss.t312 4.7885
R4686 Vss.n1184 Vss.t676 4.7885
R4687 Vss.n1186 Vss.t20 4.7885
R4688 Vss.n307 Vss.t630 4.7885
R4689 Vss.n306 Vss.t78 4.7885
R4690 Vss.n1458 Vss.t52 4.7885
R4691 Vss.n334 Vss.t628 4.7885
R4692 Vss.n1463 Vss.t365 4.7885
R4693 Vss.n325 Vss.t652 4.7885
R4694 Vss.n358 Vss.t395 4.7885
R4695 Vss.n342 Vss.t447 4.7885
R4696 Vss.n1075 Vss.t632 4.7885
R4697 Vss.n1060 Vss.t568 4.7885
R4698 Vss.n1055 Vss.t552 4.7885
R4699 Vss.n1048 Vss.t637 4.7885
R4700 Vss.n836 Vss.t389 4.7885
R4701 Vss.n842 Vss.t639 4.7885
R4702 Vss.n844 Vss.t246 4.7885
R4703 Vss.n876 Vss.t216 4.7885
R4704 Vss.n32 Vss.t360 4.7885
R4705 Vss.n33 Vss.t65 4.7885
R4706 Vss.n34 Vss.t67 4.7885
R4707 Vss.n750 Vss.t588 4.7885
R4708 Vss.n379 Vss.t326 4.7885
R4709 Vss.n300 Vss.t60 4.7885
R4710 Vss.n299 Vss.t173 4.7885
R4711 Vss.n298 Vss.t171 4.7885
R4712 Vss.n310 Vss.t110 4.7885
R4713 Vss.n1090 Vss.t674 4.7885
R4714 Vss.n1102 Vss.t271 4.7885
R4715 Vss.n1103 Vss.t7 4.7885
R4716 Vss.n1104 Vss.t9 4.7885
R4717 Vss.n1189 Vss.t100 4.7885
R4718 Vss.n1387 Vss.t338 4.7885
R4719 Vss.n1124 Vss.t205 4.7885
R4720 Vss.n1125 Vss.t123 4.7885
R4721 Vss.n1375 Vss.t130 4.7885
R4722 Vss.n1665 Vss.t277 4.7885
R4723 Vss.n1663 Vss.t149 4.7885
R4724 Vss.n1274 Vss.t536 4.7885
R4725 Vss.n1246 Vss.t544 4.7885
R4726 Vss.n1783 Vss.t112 4.7885
R4727 Vss.n1291 Vss.t328 4.7885
R4728 Vss.n1286 Vss.t91 4.7885
R4729 Vss.n1787 Vss.t93 4.7885
R4730 Vss.n97 Vss.t413 4.7885
R4731 Vss.n1746 Vss.t641 4.7885
R4732 Vss.n1757 Vss.t349 4.7885
R4733 Vss.n147 Vss.t492 4.7885
R4734 Vss.n1773 Vss.t464 4.7885
R4735 Vss.n1753 Vss.t599 4.7885
R4736 Vss.n162 Vss.t297 4.7885
R4737 Vss.n139 Vss.t496 4.7885
R4738 Vss.n1215 Vss.t256 4.7885
R4739 Vss.n1206 Vss.t280 4.7885
R4740 Vss.n1199 Vss.t18 4.7885
R4741 Vss.n1313 Vss.t241 4.7885
R4742 Vss.n1114 Vss.t37 4.7885
R4743 Vss.n1252 Vss.t300 4.7885
R4744 Vss.n1800 Vss.t646 4.7885
R4745 Vss.n1263 Vss.t436 4.7885
R4746 Vss.n1270 Vss.t549 4.7885
R4747 Vss.n1488 Vss.t666 4.7885
R4748 Vss.n1499 Vss.t454 4.7885
R4749 Vss.n68 Vss.t214 4.7885
R4750 Vss.n1705 Vss.t407 4.7885
R4751 Vss.n1717 Vss.t54 4.7885
R4752 Vss.n1681 Vss.t378 4.7885
R4753 Vss.n1677 Vss.t595 4.7885
R4754 Vss.n1674 Vss.t318 4.7885
R4755 Vss.n1702 Vss.t120 4.7885
R4756 Vss.n1327 Vss.t107 4.7885
R4757 Vss.n81 Vss.t238 4.7885
R4758 Vss.n1814 Vss.t40 4.7885
R4759 Vss.n1302 Vss.t164 4.7885
R4760 Vss.n476 Vss.t620 4.7885
R4761 Vss.n906 Vss.t547 4.7885
R4762 Vss.n801 Vss.t452 4.7885
R4763 Vss.n898 Vss.t28 4.7885
R4764 Vss.n784 Vss.t419 4.7885
R4765 Vss.n594 Vss.t434 4.7885
R4766 Vss.n552 Vss.t431 4.7885
R4767 Vss.n509 Vss.t650 4.7885
R4768 Vss.n508 Vss.t654 4.7885
R4769 Vss.n694 Vss.t658 4.7885
R4770 Vss.n660 Vss.t672 4.7885
R4771 Vss.n653 Vss.t341 4.7885
R4772 Vss.n633 Vss.t23 4.7885
R4773 Vss.n642 Vss.t369 4.7885
R4774 Vss.n685 Vss.t460 4.7885
R4775 Vss.n680 Vss.t56 4.7885
R4776 Vss.n705 Vss.t58 4.7885
R4777 Vss.n701 Vss.t592 4.7885
R4778 Vss.n3 Vss.t184 4.7885
R4779 Vss.n495 Vss.t186 4.7885
R4780 Vss.n494 Vss.t559 4.7885
R4781 Vss.n744 Vss.t557 4.7885
R4782 Vss.n612 Vss.t450 4.7885
R4783 Vss.n604 Vss.t439 4.7885
R4784 Vss.n718 Vss.n0 4.28213
R4785 Vss.n589 Vss.n542 4.28213
R4786 Vss.n1876 Vss.n1875 4.28213
R4787 Vss.n967 Vss.n435 4.28213
R4788 Vss.n333 Vss.n332 4.28213
R4789 Vss.n1047 Vss.n1046 4.28213
R4790 Vss.n1198 Vss.n1138 4.28213
R4791 Vss.n1745 Vss.n119 4.28213
R4792 Vss.n1767 Vss.n1766 4.28213
R4793 Vss.n1353 Vss.n1352 4.28213
R4794 Vss.n1254 Vss.n1253 4.28213
R4795 Vss.n1680 Vss.n186 4.28213
R4796 Vss.n1590 Vss.n1588 4.28213
R4797 Vss.n1478 Vss.n65 4.28213
R4798 Vss.n1836 Vss.n1835 4.28213
R4799 Vss.n1577 Vss.n1576 4.28213
R4800 Vss.n1555 Vss.n1554 4.28213
R4801 Vss.n1001 Vss.n1000 4.28213
R4802 Vss.n908 Vss.n907 4.28213
R4803 Vss.n935 Vss.n929 4.28213
R4804 Vss.n641 Vss.n640 4.28213
R4805 Vss.n1644 Vss.n1643 3.8722
R4806 Vss.n1623 Vss.n1617 3.52248
R4807 Vss.n1647 Vss.n1646 3.51469
R4808 Vss.n1448 Vss.n1447 3.51467
R4809 Vss.n1079 Vss.n1078 3.51467
R4810 Vss.n1864 Vss.n1863 3.51467
R4811 Vss.n1383 Vss.n1382 3.51467
R4812 Vss.n691 Vss.n690 3.51467
R4813 Vss.n1887 Vss.n1886 3.51467
R4814 Vss.n1626 Vss.t207 3.46717
R4815 Vss.t515 Vss.n1651 3.46717
R4816 Vss.n1627 Vss.t208 2.9111
R4817 Vss.n1650 Vss.t516 2.9111
R4818 Vss.n1778 Vss.n1777 2.49629
R4819 Vss.n1220 Vss.n1219 2.45741
R4820 Vss.n1219 Vss.n1109 2.21573
R4821 Vss.n913 SARlogic_0.dffrs_12.nand3_6.B 2.17818
R4822 Vss.n158 Vss.n100 2.06007
R4823 Vss.n1886 Vss.n6 2.06002
R4824 Vss.n1449 Vss.n1448 2.06002
R4825 Vss.n1078 Vss.n305 2.06002
R4826 Vss.n1865 Vss.n1864 2.06002
R4827 Vss.n1382 Vss.n1123 2.06002
R4828 Vss.n691 Vss.n510 2.06002
R4829 Vss.n1620 Vss.t503 2.048
R4830 Vss.n1620 Vss.t584 2.048
R4831 Vss.n1610 Vss.t95 2.03874
R4832 Vss.n1610 Vss.t260 2.03874
R4833 Vss.n1611 Vss.t262 2.03874
R4834 Vss.n1611 Vss.t258 2.03874
R4835 Vss.n1529 Vss.n206 2.02164
R4836 Vss.n1547 Vss.n1546 2.02164
R4837 Vss.n1022 Vss.n1021 2.02164
R4838 Vss.n1699 Vss.n73 2.02164
R4839 Vss.n1817 Vss.n75 2.02164
R4840 Vss.n1425 Vss.n268 2.02164
R4841 Vss.n1843 Vss.n48 2.02164
R4842 Vss.n251 Vss.n195 2.02164
R4843 Vss.n1729 Vss.n1728 2.02164
R4844 Vss.n921 Vss.n920 2.02164
R4845 Vss.n658 Vss.n519 1.92616
R4846 Vss.n489 Vss.n488 1.90702
R4847 Vss.n872 Vss.n28 1.90702
R4848 Vss.n1861 Vss.n30 1.90702
R4849 Vss.n1860 Vss.n31 1.90702
R4850 Vss.n753 Vss.n35 1.90702
R4851 Vss.n1855 Vss.n36 1.90702
R4852 Vss.n377 Vss.n304 1.90702
R4853 Vss.n1081 Vss.n302 1.90702
R4854 Vss.n1082 Vss.n301 1.90702
R4855 Vss.n313 Vss.n297 1.90702
R4856 Vss.n1087 Vss.n296 1.90702
R4857 Vss.n1094 Vss.n293 1.90702
R4858 Vss.n1445 Vss.n1100 1.90702
R4859 Vss.n1444 Vss.n1101 1.90702
R4860 Vss.n1191 Vss.n1105 1.90702
R4861 Vss.n1439 Vss.n1106 1.90702
R4862 Vss.n1385 Vss.n1384 1.90702
R4863 Vss.n1784 Vss.n106 1.90702
R4864 Vss.n1293 Vss.n1230 1.90702
R4865 Vss.n1295 Vss.n1294 1.90702
R4866 Vss.n664 Vss.n511 1.90702
R4867 Vss.n688 Vss.n513 1.90702
R4868 Vss.n687 Vss.n514 1.90702
R4869 Vss.n702 Vss.n699 1.90702
R4870 Vss.n723 Vss.n2 1.90702
R4871 Vss.n1888 Vss.n4 1.90702
R4872 Vss.n734 Vss.n733 1.90702
R4873 Vss.n735 Vss.n496 1.90702
R4874 Vss.n741 Vss.n740 1.90702
R4875 Vss.n1634 Vss.n1621 1.73383
R4876 Vss.n1641 Vss.n1640 1.73383
R4877 Vss.n1626 Vss.n1608 1.70279
R4878 Vss.n1651 Vss.n1608 1.62925
R4879 Vss.n1669 Vss.n190 1.62713
R4880 Vss.n1378 adc_PISO_0.2inmux_0.Bit 1.54251
R4881 Vss.n913 SARlogic_0.dffrs_12.nand3_1.A 1.34729
R4882 Vss.n586 Vss.n585 1.3005
R4883 Vss.n546 Vss.n545 1.3005
R4884 Vss.n584 Vss.n546 1.3005
R4885 Vss.n890 Vss.n394 1.3005
R4886 Vss.n889 Vss.n887 1.3005
R4887 Vss.n889 Vss.n888 1.3005
R4888 Vss.n1035 Vss.n1034 1.3005
R4889 Vss.n1031 Vss.n398 1.3005
R4890 Vss.n406 Vss.n398 1.3005
R4891 Vss.n997 Vss.n996 1.3005
R4892 Vss.n995 Vss.n994 1.3005
R4893 Vss.n995 Vss.n230 1.3005
R4894 Vss.n1535 Vss.n1534 1.3005
R4895 Vss.n228 Vss.n227 1.3005
R4896 Vss.n1533 Vss.n228 1.3005
R4897 Vss.n989 Vss.n988 1.3005
R4898 Vss.n987 Vss.n986 1.3005
R4899 Vss.n987 Vss.n231 1.3005
R4900 Vss.n942 Vss.n941 1.3005
R4901 Vss.n931 Vss.n930 1.3005
R4902 Vss.n931 Vss.n431 1.3005
R4903 Vss.n932 Vss.n430 1.3005
R4904 Vss.n982 Vss.n981 1.3005
R4905 Vss.n981 Vss.n980 1.3005
R4906 Vss.n1551 Vss.n1550 1.3005
R4907 Vss.n1550 Vss.n1549 1.3005
R4908 Vss.n440 Vss.n212 1.3005
R4909 Vss.n977 Vss.n976 1.3005
R4910 Vss.n978 Vss.n977 1.3005
R4911 Vss.n933 Vss.n432 1.3005
R4912 Vss.n442 Vss.n441 1.3005
R4913 Vss.n441 Vss.n216 1.3005
R4914 Vss.n447 Vss.n446 1.3005
R4915 Vss.n1583 Vss.n1582 1.3005
R4916 Vss.n1585 Vss.n1584 1.3005
R4917 Vss.n1584 Vss.n194 1.3005
R4918 Vss.n1561 Vss.n1560 1.3005
R4919 Vss.n1563 Vss.n1562 1.3005
R4920 Vss.n1564 Vss.n1563 1.3005
R4921 Vss.n1528 Vss.n1527 1.3005
R4922 Vss.n1524 Vss.n233 1.3005
R4923 Vss.n233 Vss.n232 1.3005
R4924 Vss.n1514 Vss.n246 1.3005
R4925 Vss.n1517 Vss.n1516 1.3005
R4926 Vss.n1516 Vss.n1515 1.3005
R4927 Vss.n1566 Vss.n200 1.3005
R4928 Vss.n1579 Vss.n1578 1.3005
R4929 Vss.n1580 Vss.n1579 1.3005
R4930 Vss.n963 Vss.n962 1.3005
R4931 Vss.n439 Vss.n438 1.3005
R4932 Vss.n961 Vss.n439 1.3005
R4933 Vss.n213 Vss.n205 1.3005
R4934 Vss.n1571 Vss.n1570 1.3005
R4935 Vss.n1570 Vss.n1569 1.3005
R4936 Vss.n1567 Vss.n193 1.3005
R4937 Vss.n1597 Vss.n1596 1.3005
R4938 Vss.n1596 Vss.n1595 1.3005
R4939 Vss.n214 Vss.n209 1.3005
R4940 Vss.n1557 Vss.n1556 1.3005
R4941 Vss.n1558 Vss.n1557 1.3005
R4942 Vss.n1545 Vss.n1544 1.3005
R4943 Vss.n1541 Vss.n219 1.3005
R4944 Vss.n219 Vss.n218 1.3005
R4945 Vss.n236 Vss.n235 1.3005
R4946 Vss.n239 Vss.n238 1.3005
R4947 Vss.n238 Vss.n237 1.3005
R4948 Vss.n407 Vss.n405 1.3005
R4949 Vss.n411 Vss.n410 1.3005
R4950 Vss.n412 Vss.n411 1.3005
R4951 Vss.n422 Vss.n421 1.3005
R4952 Vss.n415 Vss.n413 1.3005
R4953 Vss.n415 Vss.n414 1.3005
R4954 Vss.n424 Vss.n423 1.3005
R4955 Vss.n1003 Vss.n1002 1.3005
R4956 Vss.n1004 Vss.n1003 1.3005
R4957 Vss.n1007 Vss.n46 1.3005
R4958 Vss.n1847 Vss.n1846 1.3005
R4959 Vss.n1846 Vss.n1845 1.3005
R4960 Vss.n1405 Vss.n1403 1.3005
R4961 Vss.n1429 Vss.n1428 1.3005
R4962 Vss.n1428 Vss.n1427 1.3005
R4963 Vss.n1147 Vss.n1146 1.3005
R4964 Vss.n1146 Vss.n1145 1.3005
R4965 Vss.n1163 Vss.n1162 1.3005
R4966 Vss.n362 Vss.n361 1.3005
R4967 Vss.n358 Vss.n318 1.3005
R4968 Vss.n339 Vss.n318 1.3005
R4969 Vss.n353 Vss.n352 1.3005
R4970 Vss.n326 Vss.n325 1.3005
R4971 Vss.n326 Vss.n287 1.3005
R4972 Vss.n342 Vss.n341 1.3005
R4973 Vss.n341 Vss.n340 1.3005
R4974 Vss.n349 Vss.n348 1.3005
R4975 Vss.n337 Vss.n286 1.3005
R4976 Vss.n1458 Vss.n1457 1.3005
R4977 Vss.n1457 Vss.n1456 1.3005
R4978 Vss.n329 Vss.n328 1.3005
R4979 Vss.n335 Vss.n334 1.3005
R4980 Vss.n336 Vss.n335 1.3005
R4981 Vss.n1068 Vss.n306 1.3005
R4982 Vss.n1069 Vss.n1068 1.3005
R4983 Vss.n1065 Vss.n305 1.3005
R4984 Vss.n1070 Vss.n307 1.3005
R4985 Vss.n1071 Vss.n1070 1.3005
R4986 Vss.n1075 Vss.n1074 1.3005
R4987 Vss.n1074 Vss.n1073 1.3005
R4988 Vss.n1052 Vss.n388 1.3005
R4989 Vss.n1055 Vss.n1054 1.3005
R4990 Vss.n1054 Vss.n1053 1.3005
R4991 Vss.n1049 Vss.n1048 1.3005
R4992 Vss.n1050 Vss.n1049 1.3005
R4993 Vss.n1043 Vss.n1042 1.3005
R4994 Vss.n850 Vss.n34 1.3005
R4995 Vss.n1666 Vss.n1665 1.3005
R4996 Vss.n1667 Vss.n1666 1.3005
R4997 Vss.n1614 Vss.n1613 1.3005
R4998 Vss.n1663 Vss.n1662 1.3005
R4999 Vss.n1662 Vss.n1661 1.3005
R5000 Vss.n1244 Vss.n1243 1.3005
R5001 Vss.n1246 Vss.n1245 1.3005
R5002 Vss.n1245 Vss.n1232 1.3005
R5003 Vss.n1277 Vss.n1276 1.3005
R5004 Vss.n1275 Vss.n1274 1.3005
R5005 Vss.n1275 Vss.n1233 1.3005
R5006 Vss.n1794 Vss.n1793 1.3005
R5007 Vss.n98 Vss.n97 1.3005
R5008 Vss.n1792 Vss.n98 1.3005
R5009 Vss.n1761 Vss.n1760 1.3005
R5010 Vss.n1757 Vss.n125 1.3005
R5011 Vss.n129 Vss.n125 1.3005
R5012 Vss.n1753 Vss.n1752 1.3005
R5013 Vss.n1752 Vss.n110 1.3005
R5014 Vss.n1751 Vss.n1750 1.3005
R5015 Vss.n139 Vss.n138 1.3005
R5016 Vss.n138 Vss.n111 1.3005
R5017 Vss.n137 Vss.n136 1.3005
R5018 Vss.n151 Vss.n150 1.3005
R5019 Vss.n148 Vss.n147 1.3005
R5020 Vss.n149 Vss.n148 1.3005
R5021 Vss.n127 Vss.n113 1.3005
R5022 Vss.n1774 Vss.n1773 1.3005
R5023 Vss.n1775 Vss.n1774 1.3005
R5024 Vss.n1744 Vss.n1743 1.3005
R5025 Vss.n1747 Vss.n1746 1.3005
R5026 Vss.n1748 Vss.n1747 1.3005
R5027 Vss.n1291 Vss.n1290 1.3005
R5028 Vss.n1290 Vss.n1289 1.3005
R5029 Vss.n1287 Vss.n1286 1.3005
R5030 Vss.n1288 Vss.n1287 1.3005
R5031 Vss.n1788 Vss.n1787 1.3005
R5032 Vss.n1789 Vss.n1788 1.3005
R5033 Vss.n1372 Vss.n106 1.3005
R5034 Vss.n1783 Vss.n1782 1.3005
R5035 Vss.n1782 Vss.n1781 1.3005
R5036 Vss.n1363 Vss.n1123 1.3005
R5037 Vss.n1366 Vss.n1124 1.3005
R5038 Vss.n1128 Vss.n1125 1.3005
R5039 Vss.n1129 Vss.n1128 1.3005
R5040 Vss.n1375 Vss.n1374 1.3005
R5041 Vss.n1374 Vss.n1373 1.3005
R5042 Vss.n1299 Vss.n1298 1.3005
R5043 Vss.n1300 Vss.n1299 1.3005
R5044 Vss.n1295 Vss.n1231 1.3005
R5045 Vss.n1155 Vss.n1143 1.3005
R5046 Vss.n1154 Vss.n1152 1.3005
R5047 Vss.n1154 Vss.n1153 1.3005
R5048 Vss.n1141 Vss.n1133 1.3005
R5049 Vss.n1225 Vss.n1224 1.3005
R5050 Vss.n1226 Vss.n1225 1.3005
R5051 Vss.n1450 Vss.n1449 1.3005
R5052 Vss.n1178 Vss.n1177 1.3005
R5053 Vss.n1179 Vss.n1178 1.3005
R5054 Vss.n1184 Vss.n1183 1.3005
R5055 Vss.n1183 Vss.n1180 1.3005
R5056 Vss.n1187 Vss.n1186 1.3005
R5057 Vss.n1188 Vss.n1187 1.3005
R5058 Vss.n1197 Vss.n1196 1.3005
R5059 Vss.n1200 Vss.n1199 1.3005
R5060 Vss.n1201 Vss.n1200 1.3005
R5061 Vss.n1204 Vss.n1203 1.3005
R5062 Vss.n1206 Vss.n1205 1.3005
R5063 Vss.n1205 Vss.n1132 1.3005
R5064 Vss.n1192 Vss.n1191 1.3005
R5065 Vss.n1190 Vss.n1189 1.3005
R5066 Vss.n1190 Vss.n1116 1.3005
R5067 Vss.n1213 Vss.n1212 1.3005
R5068 Vss.n1215 Vss.n1214 1.3005
R5069 Vss.n1214 Vss.n1119 1.3005
R5070 Vss.n1317 Vss.n1316 1.3005
R5071 Vss.n1314 Vss.n1313 1.3005
R5072 Vss.n1315 Vss.n1314 1.3005
R5073 Vss.n1397 Vss.n272 1.3005
R5074 Vss.n1396 Vss.n1114 1.3005
R5075 Vss.n1396 Vss.n1395 1.3005
R5076 Vss.n1259 Vss.n87 1.3005
R5077 Vss.n1270 Vss.n1269 1.3005
R5078 Vss.n1269 Vss.n1268 1.3005
R5079 Vss.n1260 Vss.n88 1.3005
R5080 Vss.n1264 Vss.n1263 1.3005
R5081 Vss.n1265 Vss.n1264 1.3005
R5082 Vss.n1804 Vss.n1803 1.3005
R5083 Vss.n1800 Vss.n89 1.3005
R5084 Vss.n1266 Vss.n89 1.3005
R5085 Vss.n1822 Vss.n1821 1.3005
R5086 Vss.n69 Vss.n68 1.3005
R5087 Vss.n1820 Vss.n69 1.3005
R5088 Vss.n1503 Vss.n1502 1.3005
R5089 Vss.n1499 Vss.n253 1.3005
R5090 Vss.n253 Vss.n71 1.3005
R5091 Vss.n1491 Vss.n1490 1.3005
R5092 Vss.n1489 Vss.n1488 1.3005
R5093 Vss.n1489 Vss.n72 1.3005
R5094 Vss.n1686 Vss.n1685 1.3005
R5095 Vss.n1678 Vss.n1677 1.3005
R5096 Vss.n1678 Vss.n168 1.3005
R5097 Vss.n1505 Vss.n178 1.3005
R5098 Vss.n1702 Vss.n1701 1.3005
R5099 Vss.n1701 Vss.n1700 1.3005
R5100 Vss.n1672 Vss.n1671 1.3005
R5101 Vss.n1674 Vss.n1673 1.3005
R5102 Vss.n1673 Vss.n179 1.3005
R5103 Vss.n1679 Vss.n180 1.3005
R5104 Vss.n1682 Vss.n1681 1.3005
R5105 Vss.n1683 Vss.n1682 1.3005
R5106 Vss.n1709 Vss.n1708 1.3005
R5107 Vss.n1706 Vss.n1705 1.3005
R5108 Vss.n1707 Vss.n1706 1.3005
R5109 Vss.n1715 Vss.n1714 1.3005
R5110 Vss.n1717 Vss.n1716 1.3005
R5111 Vss.n1716 Vss.n169 1.3005
R5112 Vss.n1810 Vss.n1809 1.3005
R5113 Vss.n82 Vss.n81 1.3005
R5114 Vss.n1808 Vss.n82 1.3005
R5115 Vss.n1307 Vss.n84 1.3005
R5116 Vss.n1328 Vss.n1327 1.3005
R5117 Vss.n1329 Vss.n1328 1.3005
R5118 Vss.n1250 Vss.n74 1.3005
R5119 Vss.n1252 Vss.n1251 1.3005
R5120 Vss.n1251 Vss.n86 1.3005
R5121 Vss.n1101 Vss.n275 1.3005
R5122 Vss.n1171 Vss.n1102 1.3005
R5123 Vss.n1171 Vss.n1170 1.3005
R5124 Vss.n1175 Vss.n1103 1.3005
R5125 Vss.n1176 Vss.n1175 1.3005
R5126 Vss.n1173 Vss.n1104 1.3005
R5127 Vss.n1173 Vss.n1115 1.3005
R5128 Vss.n1815 Vss.n1814 1.3005
R5129 Vss.n1816 Vss.n1815 1.3005
R5130 Vss.n269 Vss.n76 1.3005
R5131 Vss.n1424 Vss.n1423 1.3005
R5132 Vss.n1420 Vss.n1406 1.3005
R5133 Vss.n1406 Vss.n271 1.3005
R5134 Vss.n314 Vss.n313 1.3005
R5135 Vss.n312 Vss.n310 1.3005
R5136 Vss.n312 Vss.n311 1.3005
R5137 Vss.n281 Vss.n280 1.3005
R5138 Vss.n1464 Vss.n1463 1.3005
R5139 Vss.n1465 Vss.n1464 1.3005
R5140 Vss.n296 Vss.n279 1.3005
R5141 Vss.n1091 Vss.n1090 1.3005
R5142 Vss.n1092 Vss.n1091 1.3005
R5143 Vss.n1094 Vss.n1093 1.3005
R5144 Vss.n1096 Vss.n1095 1.3005
R5145 Vss.n1097 Vss.n1096 1.3005
R5146 Vss.n1099 Vss.n295 1.3005
R5147 Vss.n1099 Vss.n1098 1.3005
R5148 Vss.n1100 Vss.n276 1.3005
R5149 Vss.n1842 Vss.n1841 1.3005
R5150 Vss.n50 Vss.n49 1.3005
R5151 Vss.n59 Vss.n49 1.3005
R5152 Vss.n1410 Vss.n1409 1.3005
R5153 Vss.n1413 Vss.n1412 1.3005
R5154 Vss.n1412 Vss.n1411 1.3005
R5155 Vss.n1530 Vss.n58 1.3005
R5156 Vss.n1834 Vss.n1833 1.3005
R5157 Vss.n1833 Vss.n1832 1.3005
R5158 Vss.n1829 Vss.n1828 1.3005
R5159 Vss.n1825 Vss.n64 1.3005
R5160 Vss.n261 Vss.n64 1.3005
R5161 Vss.n262 Vss.n63 1.3005
R5162 Vss.n266 Vss.n265 1.3005
R5163 Vss.n267 Vss.n266 1.3005
R5164 Vss.n260 Vss.n62 1.3005
R5165 Vss.n1485 Vss.n1484 1.3005
R5166 Vss.n1484 Vss.n1483 1.3005
R5167 Vss.n1480 Vss.n1479 1.3005
R5168 Vss.n1477 Vss.n1476 1.3005
R5169 Vss.n1476 Vss.n1475 1.3005
R5170 Vss.n1511 Vss.n1510 1.3005
R5171 Vss.n250 Vss.n249 1.3005
R5172 Vss.n1509 Vss.n250 1.3005
R5173 Vss.n1592 Vss.n1591 1.3005
R5174 Vss.n1589 Vss.n197 1.3005
R5175 Vss.n197 Vss.n196 1.3005
R5176 Vss.n1604 Vss.n1603 1.3005
R5177 Vss.n1600 Vss.n191 1.3005
R5178 Vss.n191 Vss.n181 1.3005
R5179 Vss.n1696 Vss.n1695 1.3005
R5180 Vss.n1692 Vss.n183 1.3005
R5181 Vss.n183 Vss.n182 1.3005
R5182 Vss.n1734 Vss.n1733 1.3005
R5183 Vss.n1736 Vss.n1735 1.3005
R5184 Vss.n1735 Vss.n160 1.3005
R5185 Vss.n1741 Vss.n1740 1.3005
R5186 Vss.n162 Vss.n161 1.3005
R5187 Vss.n161 Vss.n112 1.3005
R5188 Vss.n1731 Vss.n123 1.3005
R5189 Vss.n1765 Vss.n1764 1.3005
R5190 Vss.n1764 Vss.n1763 1.3005
R5191 Vss.n1727 Vss.n1726 1.3005
R5192 Vss.n1723 Vss.n172 1.3005
R5193 Vss.n172 Vss.n171 1.3005
R5194 Vss.n131 Vss.n130 1.3005
R5195 Vss.n156 Vss.n155 1.3005
R5196 Vss.n157 Vss.n156 1.3005
R5197 Vss.n1281 Vss.n1280 1.3005
R5198 Vss.n1351 Vss.n1350 1.3005
R5199 Vss.n1350 Vss.n1349 1.3005
R5200 Vss.n1333 Vss.n1332 1.3005
R5201 Vss.n1335 Vss.n1334 1.3005
R5202 Vss.n1334 Vss.n1282 1.3005
R5203 Vss.n1283 Vss.n1235 1.3005
R5204 Vss.n1360 Vss.n1359 1.3005
R5205 Vss.n1361 Vss.n1360 1.3005
R5206 Vss.n1390 Vss.n1106 1.3005
R5207 Vss.n1388 Vss.n1387 1.3005
R5208 Vss.n1389 Vss.n1388 1.3005
R5209 Vss.n1386 Vss.n1385 1.3005
R5210 Vss.n1296 Vss.n1121 1.3005
R5211 Vss.n1345 Vss.n1121 1.3005
R5212 Vss.n1302 Vss.n1301 1.3005
R5213 Vss.n1301 Vss.n1234 1.3005
R5214 Vss.n1343 Vss.n1342 1.3005
R5215 Vss.n924 Vss.n923 1.3005
R5216 Vss.n467 Vss.n466 1.3005
R5217 Vss.n922 Vss.n467 1.3005
R5218 Vss.n404 Vss.n403 1.3005
R5219 Vss.n1025 Vss.n1024 1.3005
R5220 Vss.n1024 Vss.n1023 1.3005
R5221 Vss.n934 Vss.n450 1.3005
R5222 Vss.n937 Vss.n936 1.3005
R5223 Vss.n938 Vss.n937 1.3005
R5224 Vss.n955 Vss.n954 1.3005
R5225 Vss.n957 Vss.n956 1.3005
R5226 Vss.n958 Vss.n957 1.3005
R5227 Vss.n458 Vss.n457 1.3005
R5228 Vss.n454 Vss.n452 1.3005
R5229 Vss.n452 Vss.n451 1.3005
R5230 Vss.n480 Vss.n479 1.3005
R5231 Vss.n476 Vss.n475 1.3005
R5232 Vss.n475 Vss.n474 1.3005
R5233 Vss.n756 Vss.n473 1.3005
R5234 Vss.n906 Vss.n905 1.3005
R5235 Vss.n905 Vss.n904 1.3005
R5236 Vss.n481 Vss.n459 1.3005
R5237 Vss.n951 Vss.n950 1.3005
R5238 Vss.n952 Vss.n951 1.3005
R5239 Vss.n1009 Vss.n301 1.3005
R5240 Vss.n1017 Vss.n300 1.3005
R5241 Vss.n1018 Vss.n1017 1.3005
R5242 Vss.n1011 Vss.n299 1.3005
R5243 Vss.n1011 Vss.n366 1.3005
R5244 Vss.n1014 Vss.n298 1.3005
R5245 Vss.n1014 Vss.n1013 1.3005
R5246 Vss.n384 Vss.n370 1.3005
R5247 Vss.n1061 Vss.n1060 1.3005
R5248 Vss.n1062 Vss.n1061 1.3005
R5249 Vss.n382 Vss.n36 1.3005
R5250 Vss.n380 Vss.n379 1.3005
R5251 Vss.n381 Vss.n380 1.3005
R5252 Vss.n378 Vss.n377 1.3005
R5253 Vss.n376 Vss.n371 1.3005
R5254 Vss.n376 Vss.n375 1.3005
R5255 Vss.n373 Vss.n372 1.3005
R5256 Vss.n374 Vss.n373 1.3005
R5257 Vss.n367 Vss.n302 1.3005
R5258 Vss.n801 Vss.n800 1.3005
R5259 Vss.n800 Vss.n799 1.3005
R5260 Vss.n831 Vss.n830 1.3005
R5261 Vss.n809 Vss.n808 1.3005
R5262 Vss.n812 Vss.n811 1.3005
R5263 Vss.n811 Vss.n810 1.3005
R5264 Vss.n819 Vss.n818 1.3005
R5265 Vss.n823 Vss.n822 1.3005
R5266 Vss.n822 Vss.n821 1.3005
R5267 Vss.n754 Vss.n753 1.3005
R5268 Vss.n752 Vss.n750 1.3005
R5269 Vss.n752 Vss.n751 1.3005
R5270 Vss.n901 Vss.n468 1.3005
R5271 Vss.n918 Vss.n917 1.3005
R5272 Vss.n919 Vss.n918 1.3005
R5273 Vss.n899 Vss.n898 1.3005
R5274 Vss.n900 Vss.n899 1.3005
R5275 Vss.n757 Vss.n483 1.3005
R5276 Vss.n784 Vss.n783 1.3005
R5277 Vss.n783 Vss.n758 1.3005
R5278 Vss.n782 Vss.n759 1.3005
R5279 Vss.n775 Vss.n774 1.3005
R5280 Vss.n773 Vss.n772 1.3005
R5281 Vss.n773 Vss.n763 1.3005
R5282 Vss.n792 Vss.n791 1.3005
R5283 Vss.n766 Vss.n765 1.3005
R5284 Vss.n765 Vss.n764 1.3005
R5285 Vss.n574 Vss.n6 1.3005
R5286 Vss.n572 Vss.n7 1.3005
R5287 Vss.n573 Vss.n572 1.3005
R5288 Vss.n12 Vss.n8 1.3005
R5289 Vss.n13 Vss.n12 1.3005
R5290 Vss.n1883 Vss.n1882 1.3005
R5291 Vss.n1882 Vss.n1881 1.3005
R5292 Vss.n598 Vss.n597 1.3005
R5293 Vss.n594 Vss.n535 1.3005
R5294 Vss.n548 Vss.n535 1.3005
R5295 Vss.n562 Vss.n561 1.3005
R5296 Vss.n567 Vss.n566 1.3005
R5297 Vss.n568 Vss.n567 1.3005
R5298 Vss.n552 Vss.n551 1.3005
R5299 Vss.n551 Vss.n550 1.3005
R5300 Vss.n558 Vss.n557 1.3005
R5301 Vss.n637 Vss.n636 1.3005
R5302 Vss.n634 Vss.n633 1.3005
R5303 Vss.n635 Vss.n634 1.3005
R5304 Vss.n532 Vss.n525 1.3005
R5305 Vss.n643 Vss.n642 1.3005
R5306 Vss.n644 Vss.n643 1.3005
R5307 Vss.n647 Vss.n523 1.3005
R5308 Vss.n653 Vss.n652 1.3005
R5309 Vss.n652 Vss.n651 1.3005
R5310 Vss.n648 Vss.n519 1.3005
R5311 Vss.n661 Vss.n660 1.3005
R5312 Vss.n662 Vss.n661 1.3005
R5313 Vss.n664 Vss.n663 1.3005
R5314 Vss.n666 Vss.n665 1.3005
R5315 Vss.n667 Vss.n666 1.3005
R5316 Vss.n669 Vss.n668 1.3005
R5317 Vss.n670 Vss.n669 1.3005
R5318 Vss.n671 Vss.n513 1.3005
R5319 Vss.n740 Vss.n14 1.3005
R5320 Vss.n739 Vss.n738 1.3005
R5321 Vss.n739 Vss.n491 1.3005
R5322 Vss.n858 Vss.n857 1.3005
R5323 Vss.n863 Vss.n862 1.3005
R5324 Vss.n864 Vss.n863 1.3005
R5325 Vss.n865 Vss.n489 1.3005
R5326 Vss.n876 Vss.n875 1.3005
R5327 Vss.n875 Vss.n874 1.3005
R5328 Vss.n873 Vss.n872 1.3005
R5329 Vss.n871 Vss.n866 1.3005
R5330 Vss.n871 Vss.n870 1.3005
R5331 Vss.n868 Vss.n867 1.3005
R5332 Vss.n869 Vss.n868 1.3005
R5333 Vss.n1878 Vss.n1877 1.3005
R5334 Vss.n18 Vss.n17 1.3005
R5335 Vss.n760 Vss.n17 1.3005
R5336 Vss.n761 Vss.n21 1.3005
R5337 Vss.n1871 Vss.n1870 1.3005
R5338 Vss.n1870 Vss.n1869 1.3005
R5339 Vss.n1866 Vss.n1865 1.3005
R5340 Vss.n837 Vss.n836 1.3005
R5341 Vss.n838 Vss.n837 1.3005
R5342 Vss.n842 Vss.n839 1.3005
R5343 Vss.n847 Vss.n839 1.3005
R5344 Vss.n845 Vss.n844 1.3005
R5345 Vss.n846 Vss.n845 1.3005
R5346 Vss.n649 Vss.n514 1.3005
R5347 Vss.n685 Vss.n684 1.3005
R5348 Vss.n684 Vss.n683 1.3005
R5349 Vss.n681 Vss.n680 1.3005
R5350 Vss.n682 Vss.n681 1.3005
R5351 Vss.n706 Vss.n705 1.3005
R5352 Vss.n707 Vss.n706 1.3005
R5353 Vss.n714 Vss.n496 1.3005
R5354 Vss.n712 Vss.n495 1.3005
R5355 Vss.n713 Vss.n712 1.3005
R5356 Vss.n708 Vss.n494 1.3005
R5357 Vss.n709 Vss.n708 1.3005
R5358 Vss.n745 Vss.n744 1.3005
R5359 Vss.n746 Vss.n745 1.3005
R5360 Vss.n855 Vss.n31 1.3005
R5361 Vss.n853 Vss.n32 1.3005
R5362 Vss.n854 Vss.n853 1.3005
R5363 Vss.n748 Vss.n33 1.3005
R5364 Vss.n848 Vss.n748 1.3005
R5365 Vss.n699 Vss.n698 1.3005
R5366 Vss.n701 Vss.n700 1.3005
R5367 Vss.n700 Vss.n499 1.3005
R5368 Vss.n717 Vss.n716 1.3005
R5369 Vss.n720 Vss.n719 1.3005
R5370 Vss.n721 Vss.n720 1.3005
R5371 Vss.n723 Vss.n722 1.3005
R5372 Vss.n724 Vss.n3 1.3005
R5373 Vss.n725 Vss.n724 1.3005
R5374 Vss.n726 Vss.n4 1.3005
R5375 Vss.n730 Vss.n729 1.3005
R5376 Vss.n731 Vss.n730 1.3005
R5377 Vss.n727 Vss.n497 1.3005
R5378 Vss.n732 Vss.n497 1.3005
R5379 Vss.n576 Vss.n575 1.3005
R5380 Vss.n578 Vss.n577 1.3005
R5381 Vss.n579 Vss.n578 1.3005
R5382 Vss.n676 Vss.n510 1.3005
R5383 Vss.n674 Vss.n509 1.3005
R5384 Vss.n675 Vss.n674 1.3005
R5385 Vss.n517 Vss.n508 1.3005
R5386 Vss.n679 Vss.n517 1.3005
R5387 Vss.n695 Vss.n694 1.3005
R5388 Vss.n696 Vss.n695 1.3005
R5389 Vss.n610 Vss.n609 1.3005
R5390 Vss.n612 Vss.n611 1.3005
R5391 Vss.n611 Vss.n531 1.3005
R5392 Vss.n624 Vss.n530 1.3005
R5393 Vss.n627 Vss.n626 1.3005
R5394 Vss.n626 Vss.n625 1.3005
R5395 Vss.n604 Vss.n603 1.3005
R5396 Vss.n603 Vss.n602 1.3005
R5397 Vss.n620 Vss.n619 1.3005
R5398 Vss.n1664 Vss.n1608 1.29323
R5399 Vss.n1665 Vss.n1664 1.00923
R5400 Vss.n1645 Vss.n1644 0.999917
R5401 Vss.n1632 Vss.n1617 0.999917
R5402 Vss.n1632 Vss.n1631 0.999917
R5403 Vss.n1646 Vss.n1645 0.999917
R5404 Vss.n742 Vss.n488 0.990409
R5405 Vss.n1856 Vss.n1855 0.990409
R5406 Vss.n1087 Vss.n1086 0.990409
R5407 Vss.n1440 Vss.n1439 0.990409
R5408 Vss.n703 Vss.n2 0.990409
R5409 Vss.n1664 Vss.n1663 0.984484
R5410 Vss.n1643 Vss.n1615 0.949529
R5411 Vss.n628 Vss.n529 0.92075
R5412 Vss.n565 Vss.n563 0.92075
R5413 Vss.n587 Vss.n544 0.92075
R5414 Vss.n790 Vss.n767 0.92075
R5415 Vss.n861 Vss.n859 0.92075
R5416 Vss.n1873 Vss.n1872 0.92075
R5417 Vss.n916 Vss.n469 0.92075
R5418 Vss.n824 Vss.n817 0.92075
R5419 Vss.n891 Vss.n886 0.92075
R5420 Vss.n949 Vss.n460 0.92075
R5421 Vss.n1027 Vss.n1026 0.92075
R5422 Vss.n1358 Vss.n1236 0.92075
R5423 Vss.n1336 Vss.n1306 0.92075
R5424 Vss.n154 Vss.n132 0.92075
R5425 Vss.n1725 Vss.n1724 0.92075
R5426 Vss.n1737 Vss.n166 0.92075
R5427 Vss.n1694 Vss.n1693 0.92075
R5428 Vss.n1602 Vss.n1601 0.92075
R5429 Vss.n1512 Vss.n248 0.92075
R5430 Vss.n1486 Vss.n259 0.92075
R5431 Vss.n264 Vss.n263 0.92075
R5432 Vss.n1827 Vss.n1826 0.92075
R5433 Vss.n1033 Vss.n1032 0.92075
R5434 Vss.n990 Vss.n985 0.92075
R5435 Vss.n1536 Vss.n226 0.92075
R5436 Vss.n998 Vss.n993 0.92075
R5437 Vss.n983 Vss.n429 0.92075
R5438 Vss.n943 Vss.n425 0.92075
R5439 Vss.n240 Vss.n234 0.92075
R5440 Vss.n1543 Vss.n1542 0.92075
R5441 Vss.n1598 Vss.n192 0.92075
R5442 Vss.n1572 Vss.n204 0.92075
R5443 Vss.n1552 Vss.n211 0.92075
R5444 Vss.n975 Vss.n973 0.92075
R5445 Vss.n445 Vss.n443 0.92075
R5446 Vss.n456 Vss.n455 0.92075
R5447 Vss.n964 Vss.n437 0.92075
R5448 Vss.n1586 Vss.n199 0.92075
R5449 Vss.n207 Vss.n202 0.92075
R5450 Vss.n1519 Vss.n1518 0.92075
R5451 Vss.n1526 Vss.n1525 0.92075
R5452 Vss.n420 Vss.n52 0.92075
R5453 Vss.n1848 Vss.n45 0.92075
R5454 Vss.n409 Vss.n408 0.92075
R5455 Vss.n1414 Vss.n1408 0.92075
R5456 Vss.n1840 Vss.n51 0.92075
R5457 Vss.n1430 Vss.n1402 0.92075
R5458 Vss.n1223 Vss.n1134 0.92075
R5459 Vss.n1161 Vss.n1148 0.92075
R5460 Vss.n1462 Vss.n282 0.92075
R5461 Vss.n354 Vss.n324 0.92075
R5462 Vss.n360 Vss.n359 0.92075
R5463 Vss.n347 Vss.n343 0.92075
R5464 Vss.n1459 Vss.n285 0.92075
R5465 Vss.n1059 Vss.n385 0.92075
R5466 Vss.n1056 Vss.n387 0.92075
R5467 Vss.n1278 Vss.n1273 0.92075
R5468 Vss.n1247 Vss.n1242 0.92075
R5469 Vss.n1795 Vss.n96 0.92075
R5470 Vss.n1759 Vss.n1758 0.92075
R5471 Vss.n1772 Vss.n114 0.92075
R5472 Vss.n1755 Vss.n1754 0.92075
R5473 Vss.n1739 Vss.n165 0.92075
R5474 Vss.n141 Vss.n140 0.92075
R5475 Vss.n152 Vss.n146 0.92075
R5476 Vss.n1216 Vss.n1211 0.92075
R5477 Vss.n1208 Vss.n1207 0.92075
R5478 Vss.n1156 Vss.n1151 0.92075
R5479 Vss.n1318 Vss.n1312 0.92075
R5480 Vss.n1398 Vss.n1113 0.92075
R5481 Vss.n1802 Vss.n1801 0.92075
R5482 Vss.n1262 Vss.n1261 0.92075
R5483 Vss.n1271 Vss.n1258 0.92075
R5484 Vss.n1492 Vss.n1487 0.92075
R5485 Vss.n1501 Vss.n1500 0.92075
R5486 Vss.n1823 Vss.n67 0.92075
R5487 Vss.n1719 Vss.n1718 0.92075
R5488 Vss.n1710 Vss.n1704 0.92075
R5489 Vss.n1687 Vss.n1676 0.92075
R5490 Vss.n1675 Vss.n187 0.92075
R5491 Vss.n1703 Vss.n177 0.92075
R5492 Vss.n1326 Vss.n1308 0.92075
R5493 Vss.n1811 Vss.n80 0.92075
R5494 Vss.n1813 Vss.n77 0.92075
R5495 Vss.n1422 Vss.n1421 0.92075
R5496 Vss.n1341 Vss.n1303 0.92075
R5497 Vss.n925 Vss.n465 0.92075
R5498 Vss.n478 Vss.n477 0.92075
R5499 Vss.n829 Vss.n802 0.92075
R5500 Vss.n813 Vss.n807 0.92075
R5501 Vss.n897 Vss.n484 0.92075
R5502 Vss.n785 Vss.n781 0.92075
R5503 Vss.n776 Vss.n771 0.92075
R5504 Vss.n596 Vss.n595 0.92075
R5505 Vss.n556 Vss.n553 0.92075
R5506 Vss.n654 Vss.n522 0.92075
R5507 Vss.n638 Vss.n632 0.92075
R5508 Vss.n613 Vss.n608 0.92075
R5509 Vss.n618 Vss.n605 0.92075
R5510 Vss.n1630 Vss.n1615 0.907842
R5511 Vss.n1636 Vss.n1635 0.867167
R5512 Vss.t502 Vss.n1638 0.867167
R5513 Vss.n1639 Vss.n1616 0.867167
R5514 SARlogic_0.dffrs_12.d SARlogic_0.dffrs_12.nand3_8.A 0.784786
R5515 SARlogic_0.dffrs_13.d SARlogic_0.dffrs_13.nand3_8.A 0.784786
R5516 Vss.n1248 Vss.n95 0.780467
R5517 Vss.n1884 Vss.n1883 0.771017
R5518 Vss.n1186 Vss.n1185 0.771017
R5519 Vss.n1076 Vss.n1075 0.771017
R5520 Vss.n844 Vss.n843 0.771017
R5521 Vss.n694 Vss.n693 0.771017
R5522 Vss.n1625 Vss.n1 0.714636
R5523 Vss.n1088 Vss.n41 0.669813
R5524 Vss.n1854 Vss.n1853 0.669683
R5525 Vss.n879 Vss.n878 0.669683
R5526 Vss.n1643 comparator_no_offsetcal_0.lvsclean_SAlatch_0.VSS 0.664071
R5527 Vss.n1891 Vss.n1890 0.651683
R5528 Vss.n697 Vss.n503 0.63255
R5529 SARlogic_0.dffrs_12.clk Vss.n913 0.611214
R5530 Vss.n658 Vss.n657 0.601415
R5531 Vss.n1438 Vss.n1437 0.600912
R5532 Vss.n1379 Vss.n1375 0.471317
R5533 Vss.n741 Vss.n738 0.463217
R5534 Vss.n1885 Vss.n7 0.463217
R5535 Vss.n1884 Vss.n8 0.463217
R5536 Vss.n1177 Vss.n292 0.463217
R5537 Vss.n1185 Vss.n1184 0.463217
R5538 Vss.n1076 Vss.n307 0.463217
R5539 Vss.n1077 Vss.n306 0.463217
R5540 Vss.n836 Vss.n27 0.463217
R5541 Vss.n843 Vss.n842 0.463217
R5542 Vss.n877 Vss.n876 0.463217
R5543 Vss.n1859 Vss.n32 0.463217
R5544 Vss.n1858 Vss.n33 0.463217
R5545 Vss.n1857 Vss.n34 0.463217
R5546 Vss.n750 Vss.n35 0.463217
R5547 Vss.n379 Vss.n37 0.463217
R5548 Vss.n1083 Vss.n300 0.463217
R5549 Vss.n1084 Vss.n299 0.463217
R5550 Vss.n1085 Vss.n298 0.463217
R5551 Vss.n310 Vss.n297 0.463217
R5552 Vss.n1090 Vss.n1089 0.463217
R5553 Vss.n1443 Vss.n1102 0.463217
R5554 Vss.n1442 Vss.n1103 0.463217
R5555 Vss.n1441 Vss.n1104 0.463217
R5556 Vss.n1189 Vss.n1105 0.463217
R5557 Vss.n1387 Vss.n1107 0.463217
R5558 Vss.n1381 Vss.n1124 0.463217
R5559 Vss.n1380 Vss.n1125 0.463217
R5560 Vss.n1784 Vss.n1783 0.463217
R5561 Vss.n1292 Vss.n1291 0.463217
R5562 Vss.n1286 Vss.n105 0.463217
R5563 Vss.n1787 Vss.n1786 0.463217
R5564 Vss.n692 Vss.n509 0.463217
R5565 Vss.n693 Vss.n508 0.463217
R5566 Vss.n660 Vss.n659 0.463217
R5567 Vss.n686 Vss.n685 0.463217
R5568 Vss.n680 Vss.n502 0.463217
R5569 Vss.n705 Vss.n704 0.463217
R5570 Vss.n702 Vss.n701 0.463217
R5571 Vss.n1889 Vss.n3 0.463217
R5572 Vss.n736 Vss.n495 0.463217
R5573 Vss.n737 Vss.n494 0.463217
R5574 Vss.n744 Vss.n743 0.463217
R5575 Vss.n883 Vss.n39 0.441453
R5576 Vss.n657 Vss.n1 0.328611
R5577 Vss.n1885 Vss.n1884 0.3083
R5578 Vss.n1185 Vss.n292 0.3083
R5579 Vss.n1077 Vss.n1076 0.3083
R5580 Vss.n843 Vss.n27 0.3083
R5581 Vss.n1859 Vss.n1858 0.3083
R5582 Vss.n1858 Vss.n1857 0.3083
R5583 Vss.n1084 Vss.n1083 0.3083
R5584 Vss.n1085 Vss.n1084 0.3083
R5585 Vss.n1443 Vss.n1442 0.3083
R5586 Vss.n1442 Vss.n1441 0.3083
R5587 Vss.n1381 Vss.n1380 0.3083
R5588 Vss.n1292 Vss.n105 0.3083
R5589 Vss.n1786 Vss.n105 0.3083
R5590 Vss.n693 Vss.n692 0.3083
R5591 Vss.n686 Vss.n502 0.3083
R5592 Vss.n704 Vss.n502 0.3083
R5593 Vss.n737 Vss.n736 0.3083
R5594 Vss.n743 Vss.n737 0.3083
R5595 Vss.n1380 Vss.n1379 0.3002
R5596 Vss.n880 Vss.n879 0.284919
R5597 Vss.n1377 Vss.n1376 0.252687
R5598 Vss.n1649 Vss.n1648 0.238053
R5599 Vss.n1649 comparator_no_offsetcal_0.VSS 0.222184
R5600 Vss.n1860 Vss.n1859 0.2165
R5601 Vss.n1083 Vss.n1082 0.2165
R5602 Vss.n1444 Vss.n1443 0.2165
R5603 Vss.n1293 Vss.n1292 0.2165
R5604 Vss.n687 Vss.n686 0.2165
R5605 Vss.n736 Vss.n735 0.2165
R5606 Vss.n1629 Vss.n1628 0.211763
R5607 Vss.n884 Vss.n883 0.195855
R5608 comparator_no_offsetcal_0.x5.avss Vss.n1627 0.188808
R5609 Vss.n1650 comparator_no_offsetcal_0.x3.avss 0.188808
R5610 Vss.n1857 Vss.n1856 0.1748
R5611 Vss.n1441 Vss.n1440 0.1748
R5612 Vss.n704 Vss.n703 0.1748
R5613 Vss.n743 Vss.n742 0.1748
R5614 Vss.n1086 Vss.n1085 0.17465
R5615 Vss.n1648 Vss.n1615 0.163684
R5616 comparator_no_offsetcal_0.lvsclean_SAlatch_0.VSS Vss.n1642 0.1605
R5617 Vss.n1786 Vss.n1785 0.1598
R5618 Vss.n1657 Vss.n1656 0.154786
R5619 Vss.n1785 Vss.n1784 0.152487
R5620 Vss.n1861 Vss.n1860 0.148459
R5621 Vss.n1082 Vss.n1081 0.148459
R5622 Vss.n1445 Vss.n1444 0.148459
R5623 Vss.n1294 Vss.n1293 0.148459
R5624 Vss.n688 Vss.n687 0.148459
R5625 Vss.n735 Vss.n734 0.148459
R5626 Vss.n1852 Vss.n1851 0.145432
R5627 Vss.n1434 Vss.n1433 0.145432
R5628 Vss.n1249 Vss.n1239 0.143322
R5629 Vss.n884 Vss.n463 0.140365
R5630 Vss.n1086 Vss.n297 0.13865
R5631 Vss.n1856 Vss.n35 0.1385
R5632 Vss.n1440 Vss.n1105 0.1385
R5633 Vss.n703 Vss.n702 0.1385
R5634 Vss.n742 Vss.n741 0.1385
R5635 Vss.n1435 Vss.n1434 0.136253
R5636 Vss.n1653 Vss.n1612 0.1355
R5637 Vss.n1627 Vss.n1626 0.128901
R5638 Vss.n1651 Vss.n1650 0.127885
R5639 Vss.n893 Vss.n486 0.122607
R5640 Vss.n971 Vss.n970 0.122607
R5641 Vss.n1159 Vss.n1158 0.122607
R5642 Vss.n321 Vss.n320 0.122607
R5643 Vss.n805 Vss.n803 0.122607
R5644 Vss.n779 Vss.n778 0.122607
R5645 Vss.n539 Vss.n537 0.122607
R5646 Vss.n616 Vss.n606 0.122607
R5647 Vss.n926 Vss.n463 0.118169
R5648 Vss.n126 Vss.n117 0.115241
R5649 Vss.n1630 Vss.n1629 0.112526
R5650 Vss.n1659 Vss.n1658 0.109786
R5651 Vss.n1851 Vss.n41 0.104592
R5652 Vss.n590 Vss.n540 0.10457
R5653 Vss.n344 Vss.n284 0.10457
R5654 Vss.n826 Vss.n386 0.10457
R5655 Vss.n1770 Vss.n1769 0.10457
R5656 Vss.n1356 Vss.n1355 0.10457
R5657 Vss.n787 Vss.n19 0.10457
R5658 Vss.n631 Vss.n630 0.10457
R5659 SARlogic_0.dffrs_14.vss Vss.n1798 0.102612
R5660 Vss.n1494 SARlogic_0.dffrs_8.vss 0.102537
R5661 SARlogic_0.dffrs_10.vss Vss.n224 0.102537
R5662 Vss.n1497 SARlogic_0.dffrs_7.vss 0.101537
R5663 SARlogic_0.dffrs_9.vss Vss.n225 0.101537
R5664 Vss.n1853 Vss.n1852 0.0911096
R5665 Vss.n914 Vss.n910 0.078611
R5666 Vss.n927 Vss.n926 0.0781858
R5667 Vss.n1434 Vss.n1110 0.0776599
R5668 Vss.n1433 Vss.n1432 0.0776599
R5669 Vss.n1852 Vss.n40 0.0776599
R5670 Vss.n1851 Vss.n1850 0.0776599
R5671 Vss.n1862 Vss.n29 0.073981
R5672 Vss.n1080 Vss.n303 0.073981
R5673 Vss.n1446 Vss.n294 0.073981
R5674 Vss.n1297 Vss.n1122 0.073981
R5675 Vss.n689 Vss.n512 0.073981
R5676 Vss.n728 Vss.n5 0.073981
R5677 Vss.n1874 Vss.n20 0.0679983
R5678 Vss.n331 Vss.n330 0.0679983
R5679 Vss.n1045 Vss.n1044 0.0679983
R5680 Vss.n1210 Vss.n1209 0.0679983
R5681 Vss.n639 Vss.n520 0.0679983
R5682 Vss.n283 Vss.n41 0.0673674
R5683 Vss.n1853 Vss.n38 0.0673025
R5684 Vss.n879 Vss.n487 0.0673025
R5685 Vss.n1221 Vss.n1220 0.0665049
R5686 Vss.n946 Vss.n945 0.0660086
R5687 Vss.n945 Vss.n426 0.0655096
R5688 Vss.n966 Vss.n965 0.0645882
R5689 Vss.n472 Vss.n461 0.0645882
R5690 Vss.n1886 Vss.n1885 0.0635
R5691 Vss.n1448 Vss.n292 0.0635
R5692 Vss.n1078 Vss.n1077 0.0635
R5693 Vss.n1864 Vss.n27 0.0635
R5694 Vss.n1382 Vss.n1381 0.0635
R5695 Vss.n692 Vss.n691 0.0635
R5696 Vss.n135 Vss.n133 0.0625376
R5697 Vss.n606 Vss.n526 0.0622481
R5698 Vss.n778 Vss.n769 0.0622481
R5699 Vss.n970 Vss.n969 0.0622481
R5700 Vss.n322 Vss.n321 0.0622481
R5701 Vss.n805 Vss.n804 0.0622481
R5702 Vss.n1158 Vss.n1137 0.0622481
R5703 Vss.n486 Vss.n471 0.0622481
R5704 Vss.n591 Vss.n539 0.0622481
R5705 Vss.n1721 Vss.n93 0.0616538
R5706 Vss.n1112 Vss.n78 0.0616538
R5707 Vss.n1498 Vss.n176 0.0616538
R5708 Vss.n258 Vss.n245 0.0616538
R5709 Vss.n1431 Vss.n1401 0.0616538
R5710 Vss.n1849 Vss.n44 0.0616538
R5711 Vss.n243 Vss.n242 0.0616538
R5712 Vss.n974 Vss.n221 0.0616538
R5713 Vss.n1030 Vss.n1029 0.0616538
R5714 Vss.n1311 Vss.n1305 0.0615256
R5715 Vss.n1891 Vss.n1 0.0600636
R5716 Vss.n1461 Vss.n1460 0.0568904
R5717 Vss.n1058 Vss.n1057 0.0568904
R5718 Vss.n860 Vss.n22 0.0568904
R5719 Vss.n655 Vss.n521 0.0568904
R5720 Vss.n1220 Vss.n1139 0.0566774
R5721 Vss.n1437 Vss.n1436 0.0561349
R5722 Vss.n881 Vss.n880 0.0551896
R5723 Vss.n884 Vss.n470 0.0551896
R5724 Vss.n590 Vss.n541 0.054837
R5725 Vss.n1460 Vss.n284 0.054837
R5726 Vss.n1057 Vss.n386 0.054837
R5727 Vss.n1769 Vss.n117 0.054837
R5728 Vss.n1355 Vss.n1239 0.054837
R5729 Vss.n22 Vss.n19 0.054837
R5730 Vss.n631 Vss.n521 0.054837
R5731 Vss.n1853 Vss.n39 0.0521009
R5732 Vss.n543 Vss.n541 0.0502328
R5733 Vss.n1437 Vss.n1108 0.0480028
R5734 Vss.n244 Vss.n225 0.0478478
R5735 Vss.n416 Vss.n40 0.0478478
R5736 Vss.n1850 Vss.n43 0.0478478
R5737 Vss.n143 Vss.n95 0.0478478
R5738 Vss.n1497 Vss.n174 0.0478478
R5739 Vss.n1339 Vss.n1304 0.0478478
R5740 Vss.n1798 Vss.n1797 0.0478478
R5741 Vss.n1320 Vss.n1110 0.0478478
R5742 Vss.n1432 Vss.n1400 0.0478478
R5743 Vss.n1495 Vss.n1494 0.0478478
R5744 Vss.n1538 Vss.n224 0.0478478
R5745 Vss.n883 Vss.n882 0.0478478
R5746 Vss.n543 Vss.n0 0.0467
R5747 Vss.n345 Vss.n344 0.0466843
R5748 Vss.n1770 Vss.n116 0.0466843
R5749 Vss.n1356 Vss.n1238 0.0466843
R5750 Vss.n827 Vss.n826 0.0466843
R5751 Vss.n787 Vss.n786 0.0466843
R5752 Vss.n554 Vss.n540 0.0466843
R5753 Vss.n630 Vss.n527 0.0466843
R5754 Vss.n885 Vss.n881 0.0465106
R5755 Vss.n915 Vss.n470 0.0465106
R5756 Vss.n910 Vss.n462 0.0465106
R5757 Vss.n1257 Vss.n1256 0.0465022
R5758 Vss.n1824 Vss.n66 0.0465022
R5759 Vss.n427 Vss.n57 0.0465022
R5760 Vss.n999 Vss.n992 0.0465022
R5761 Vss.n1272 Vss.n1249 0.0464521
R5762 Vss.n1658 Vss.n1657 0.0455
R5763 Vss.n769 Vss.n19 0.0415307
R5764 Vss.n969 Vss.n968 0.0415307
R5765 Vss.n322 Vss.n284 0.0415307
R5766 Vss.n804 Vss.n386 0.0415307
R5767 Vss.n1220 Vss.n1137 0.0415307
R5768 Vss.n909 Vss.n471 0.0415307
R5769 Vss.n591 Vss.n590 0.0415307
R5770 Vss.n631 Vss.n526 0.0415307
R5771 Vss.n1433 Vss.n41 0.0413406
R5772 Vss.n453 Vss.n434 0.0405109
R5773 Vss.n1160 Vss.n1136 0.0405109
R5774 Vss.n346 Vss.n345 0.0405109
R5775 Vss.n357 Vss.n319 0.0405109
R5776 Vss.n355 Vss.n323 0.0405109
R5777 Vss.n142 Vss.n116 0.0405109
R5778 Vss.n1771 Vss.n115 0.0405109
R5779 Vss.n1157 Vss.n1150 0.0405109
R5780 Vss.n1222 Vss.n1135 0.0405109
R5781 Vss.n1340 Vss.n1238 0.0405109
R5782 Vss.n1357 Vss.n1237 0.0405109
R5783 Vss.n828 Vss.n827 0.0405109
R5784 Vss.n814 Vss.n806 0.0405109
R5785 Vss.n825 Vss.n816 0.0405109
R5786 Vss.n896 Vss.n485 0.0405109
R5787 Vss.n786 Vss.n780 0.0405109
R5788 Vss.n777 Vss.n770 0.0405109
R5789 Vss.n789 Vss.n788 0.0405109
R5790 Vss.n555 Vss.n554 0.0405109
R5791 Vss.n593 Vss.n536 0.0405109
R5792 Vss.n564 Vss.n538 0.0405109
R5793 Vss.n617 Vss.n527 0.0405109
R5794 Vss.n614 Vss.n607 0.0405109
R5795 Vss.n629 Vss.n528 0.0405109
R5796 Vss.n928 Vss.n927 0.040346
R5797 Vss.n1862 Vss.n1861 0.0389018
R5798 Vss.n1081 Vss.n1080 0.0389018
R5799 Vss.n1446 Vss.n1445 0.0389018
R5800 Vss.n1294 Vss.n1122 0.0389018
R5801 Vss.n689 Vss.n688 0.0389018
R5802 Vss.n734 Vss.n5 0.0389018
R5803 Vss.n1756 Vss.n126 0.0368083
R5804 Vss.n1690 Vss.n122 0.036505
R5805 Vss.n1689 Vss.n1688 0.036505
R5806 Vss.n1587 Vss.n185 0.036505
R5807 Vss.n1575 Vss.n1574 0.036505
R5808 Vss.n1553 Vss.n203 0.036505
R5809 Vss.n1523 Vss.n243 0.0361576
R5810 Vss.n1029 Vss.n400 0.0361576
R5811 Vss.n53 Vss.n44 0.0361576
R5812 Vss.n145 Vss.n135 0.0361576
R5813 Vss.n176 Vss.n175 0.0361576
R5814 Vss.n1419 Vss.n1401 0.0361576
R5815 Vss.n1337 Vss.n1305 0.0361576
R5816 Vss.n1722 Vss.n1721 0.0361576
R5817 Vss.n1309 Vss.n78 0.0361576
R5818 Vss.n254 Vss.n245 0.0361576
R5819 Vss.n1540 Vss.n221 0.0361576
R5820 Vss.n464 Vss.n463 0.0361576
R5821 Vss.n330 Vss.n283 0.035635
R5822 Vss.n1044 Vss.n38 0.035635
R5823 Vss.n487 Vss.n20 0.035635
R5824 Vss.n656 Vss.n520 0.035635
R5825 Vss.n657 Vss.n656 0.0352182
R5826 Vss.n1875 Vss.n19 0.0349747
R5827 Vss.n968 Vss.n967 0.0349747
R5828 Vss.n332 Vss.n284 0.0349747
R5829 Vss.n1046 Vss.n386 0.0349747
R5830 Vss.n1220 Vss.n1138 0.0349747
R5831 Vss.n909 Vss.n908 0.0349747
R5832 Vss.n590 Vss.n589 0.0349747
R5833 Vss.n640 Vss.n631 0.0349747
R5834 Vss.n1210 Vss.n1140 0.0346145
R5835 Vss.n153 Vss.n135 0.0340549
R5836 Vss.n929 Vss.n928 0.0339793
R5837 Vss.n1721 Vss.n173 0.0335769
R5838 Vss.n1311 Vss.n1310 0.0335769
R5839 Vss.n1112 Vss.n1110 0.0335769
R5840 Vss.n1812 Vss.n78 0.0335769
R5841 Vss.n1711 Vss.n176 0.0335769
R5842 Vss.n1513 Vss.n245 0.0335769
R5843 Vss.n1432 Vss.n1431 0.0335769
R5844 Vss.n1415 Vss.n1401 0.0335769
R5845 Vss.n1850 Vss.n1849 0.0335769
R5846 Vss.n1839 Vss.n44 0.0335769
R5847 Vss.n243 Vss.n241 0.0335769
R5848 Vss.n221 Vss.n220 0.0335769
R5849 Vss.n1030 Vss.n40 0.0335769
R5850 Vss.n1029 Vss.n401 0.0335769
R5851 Vss.n1324 Vss.n1323 0.0334487
R5852 Vss.n769 Vss.n768 0.0322085
R5853 Vss.n895 Vss.n893 0.0322085
R5854 Vss.n1539 Vss.n222 0.0322085
R5855 Vss.n256 Vss.n247 0.0322085
R5856 Vss.n121 Vss.n94 0.0322085
R5857 Vss.n1522 Vss.n244 0.0322085
R5858 Vss.n971 Vss.n433 0.0322085
R5859 Vss.n969 Vss.n433 0.0322085
R5860 Vss.n418 Vss.n416 0.0322085
R5861 Vss.n418 Vss.n417 0.0322085
R5862 Vss.n54 Vss.n43 0.0322085
R5863 Vss.n1159 Vss.n1149 0.0322085
R5864 Vss.n356 Vss.n320 0.0322085
R5865 Vss.n356 Vss.n322 0.0322085
R5866 Vss.n815 Vss.n804 0.0322085
R5867 Vss.n144 Vss.n143 0.0322085
R5868 Vss.n1149 Vss.n1137 0.0322085
R5869 Vss.n1713 Vss.n174 0.0322085
R5870 Vss.n1418 Vss.n1400 0.0322085
R5871 Vss.n1418 Vss.n1416 0.0322085
R5872 Vss.n1339 Vss.n1338 0.0322085
R5873 Vss.n1338 Vss.n1240 0.0322085
R5874 Vss.n144 Vss.n118 0.0322085
R5875 Vss.n1797 Vss.n94 0.0322085
R5876 Vss.n1321 Vss.n1320 0.0322085
R5877 Vss.n1321 Vss.n79 0.0322085
R5878 Vss.n1713 Vss.n1712 0.0322085
R5879 Vss.n1495 Vss.n256 0.0322085
R5880 Vss.n1838 Vss.n54 0.0322085
R5881 Vss.n1522 Vss.n1521 0.0322085
R5882 Vss.n1539 Vss.n1538 0.0322085
R5883 Vss.n882 Vss.n402 0.0322085
R5884 Vss.n927 Vss.n402 0.0322085
R5885 Vss.n815 Vss.n803 0.0322085
R5886 Vss.n895 Vss.n471 0.0322085
R5887 Vss.n779 Vss.n768 0.0322085
R5888 Vss.n592 Vss.n537 0.0322085
R5889 Vss.n592 Vss.n591 0.0322085
R5890 Vss.n616 Vss.n615 0.0322085
R5891 Vss.n615 Vss.n526 0.0322085
R5892 Vss.n1436 Vss.n1109 0.0317776
R5893 Vss.n885 Vss.n884 0.0308765
R5894 Vss.n1436 Vss.n1435 0.0306923
R5895 Vss.n892 Vss.n881 0.0268641
R5896 Vss.n1494 Vss.n257 0.0268641
R5897 Vss.n972 Vss.n224 0.0268641
R5898 Vss.n444 Vss.n221 0.0268641
R5899 Vss.n1520 Vss.n245 0.0268641
R5900 Vss.n1850 Vss.n42 0.0268641
R5901 Vss.n419 Vss.n44 0.0268641
R5902 Vss.n1407 Vss.n1401 0.0268641
R5903 Vss.n1432 Vss.n1111 0.0268641
R5904 Vss.n1798 Vss.n92 0.0268641
R5905 Vss.n1721 Vss.n1720 0.0268641
R5906 Vss.n1417 Vss.n78 0.0268641
R5907 Vss.n135 Vss.n134 0.0268641
R5908 Vss.n1796 Vss.n95 0.0268641
R5909 Vss.n1323 Vss.n1322 0.0268641
R5910 Vss.n1319 Vss.n1310 0.0268641
R5911 Vss.n1399 Vss.n1110 0.0268641
R5912 Vss.n255 Vss.n176 0.0268641
R5913 Vss.n1497 Vss.n1496 0.0268641
R5914 Vss.n243 Vss.n223 0.0268641
R5915 Vss.n1537 Vss.n225 0.0268641
R5916 Vss.n399 Vss.n40 0.0268641
R5917 Vss.n1029 Vss.n1028 0.0268641
R5918 Vss.n894 Vss.n470 0.0268641
R5919 Vss.n1249 Vss.n1248 0.0263346
R5920 Vss.n866 Vss.n29 0.0258591
R5921 Vss.n867 Vss.n29 0.0258591
R5922 Vss.n371 Vss.n303 0.0258591
R5923 Vss.n372 Vss.n303 0.0258591
R5924 Vss.n1095 Vss.n294 0.0258591
R5925 Vss.n295 Vss.n294 0.0258591
R5926 Vss.n1297 Vss.n1296 0.0258591
R5927 Vss.n1298 Vss.n1297 0.0258591
R5928 Vss.n665 Vss.n512 0.0258591
R5929 Vss.n668 Vss.n512 0.0258591
R5930 Vss.n729 Vss.n728 0.0258591
R5931 Vss.n728 Vss.n727 0.0258591
R5932 Vss.n1769 Vss.n118 0.0237454
R5933 Vss.n1768 Vss.n121 0.0235512
R5934 Vss.n1355 Vss.n1240 0.0235512
R5935 Vss.n1241 Vss.n79 0.0235512
R5936 Vss.n1712 Vss.n120 0.0235512
R5937 Vss.n247 Vss.n198 0.0235512
R5938 Vss.n1416 Vss.n56 0.0235512
R5939 Vss.n1838 Vss.n1837 0.0235512
R5940 Vss.n1521 Vss.n201 0.0235512
R5941 Vss.n222 Vss.n210 0.0235512
R5942 Vss.n417 Vss.n55 0.0235512
R5943 Vss.n588 Vss.n543 0.0232899
R5944 Vss.n1863 Vss.n1862 0.023066
R5945 Vss.n1080 Vss.n1079 0.023066
R5946 Vss.n1447 Vss.n1446 0.023066
R5947 Vss.n1383 Vss.n1122 0.023066
R5948 Vss.n690 Vss.n689 0.023066
R5949 Vss.n1887 Vss.n5 0.023066
R5950 Vss.n153 Vss.n118 0.0226532
R5951 Vss.n910 Vss.n909 0.0225109
R5952 Vss.n928 Vss.n55 0.0225109
R5953 Vss.n1837 Vss.n55 0.0225109
R5954 Vss.n1837 Vss.n56 0.0225109
R5955 Vss.n1241 Vss.n56 0.0225109
R5956 Vss.n1354 Vss.n1241 0.0225109
R5957 Vss.n1769 Vss.n1768 0.0225109
R5958 Vss.n1768 Vss.n120 0.0225109
R5959 Vss.n198 Vss.n120 0.0225109
R5960 Vss.n201 Vss.n198 0.0225109
R5961 Vss.n210 Vss.n201 0.0225109
R5962 Vss.n968 Vss.n210 0.0225109
R5963 Vss.n1574 Vss.n203 0.0223682
R5964 Vss.n1574 Vss.n185 0.0223682
R5965 Vss.n1689 Vss.n185 0.0223682
R5966 Vss.n1690 Vss.n1689 0.0223682
R5967 Vss.n1690 Vss.n126 0.0223682
R5968 Vss.n965 Vss.n203 0.0223682
R5969 Vss.n946 Vss.n461 0.0223682
R5970 Vss.n173 Vss.n121 0.0223376
R5971 Vss.n1812 Vss.n79 0.0223376
R5972 Vss.n1712 Vss.n1711 0.0223376
R5973 Vss.n1513 Vss.n247 0.0223376
R5974 Vss.n1416 Vss.n1415 0.0223376
R5975 Vss.n1839 Vss.n1838 0.0223376
R5976 Vss.n1521 Vss.n241 0.0223376
R5977 Vss.n222 Vss.n220 0.0223376
R5978 Vss.n417 Vss.n401 0.0223376
R5979 Vss.n1325 Vss.n1240 0.0222094
R5980 Vss.n1633 Vss.n1632 0.0215413
R5981 Vss.n1645 Vss.n1618 0.0215413
R5982 Vss.n893 Vss.n892 0.0214837
R5983 Vss.n257 Vss.n244 0.0214837
R5984 Vss.n972 Vss.n971 0.0214837
R5985 Vss.n444 Vss.n433 0.0214837
R5986 Vss.n1522 Vss.n1520 0.0214837
R5987 Vss.n416 Vss.n42 0.0214837
R5988 Vss.n419 Vss.n418 0.0214837
R5989 Vss.n1407 Vss.n54 0.0214837
R5990 Vss.n1111 Vss.n43 0.0214837
R5991 Vss.n1160 Vss.n1159 0.0214837
R5992 Vss.n346 Vss.n320 0.0214837
R5993 Vss.n356 Vss.n355 0.0214837
R5994 Vss.n143 Vss.n142 0.0214837
R5995 Vss.n144 Vss.n115 0.0214837
R5996 Vss.n1149 Vss.n1135 0.0214837
R5997 Vss.n174 Vss.n92 0.0214837
R5998 Vss.n1720 Vss.n1713 0.0214837
R5999 Vss.n1418 Vss.n1417 0.0214837
R6000 Vss.n1340 Vss.n1339 0.0214837
R6001 Vss.n1338 Vss.n1237 0.0214837
R6002 Vss.n134 Vss.n94 0.0214837
R6003 Vss.n1797 Vss.n1796 0.0214837
R6004 Vss.n1322 Vss.n1321 0.0214837
R6005 Vss.n1320 Vss.n1319 0.0214837
R6006 Vss.n1400 Vss.n1399 0.0214837
R6007 Vss.n256 Vss.n255 0.0214837
R6008 Vss.n1496 Vss.n1495 0.0214837
R6009 Vss.n1539 Vss.n223 0.0214837
R6010 Vss.n1538 Vss.n1537 0.0214837
R6011 Vss.n882 Vss.n399 0.0214837
R6012 Vss.n1028 Vss.n402 0.0214837
R6013 Vss.n828 Vss.n803 0.0214837
R6014 Vss.n816 Vss.n815 0.0214837
R6015 Vss.n895 Vss.n894 0.0214837
R6016 Vss.n780 Vss.n779 0.0214837
R6017 Vss.n789 Vss.n768 0.0214837
R6018 Vss.n555 Vss.n537 0.0214837
R6019 Vss.n592 Vss.n538 0.0214837
R6020 Vss.n617 Vss.n616 0.0214837
R6021 Vss.n615 Vss.n528 0.0214837
R6022 Vss.n945 Vss.n462 0.0204141
R6023 Vss.n1769 Vss.n119 0.0200312
R6024 Vss.n1738 Vss.n126 0.0199048
R6025 Vss.n1768 Vss.n1767 0.019868
R6026 Vss.n1254 Vss.n1241 0.019868
R6027 Vss.n186 Vss.n120 0.019868
R6028 Vss.n1588 Vss.n198 0.019868
R6029 Vss.n65 Vss.n56 0.019868
R6030 Vss.n1837 Vss.n1836 0.019868
R6031 Vss.n1576 Vss.n201 0.019868
R6032 Vss.n1554 Vss.n210 0.019868
R6033 Vss.n1000 Vss.n55 0.019868
R6034 Vss.n1354 Vss.n1353 0.0197929
R6035 Vss.n1656 Vss.n1612 0.0197857
R6036 Vss.n1691 Vss.n1690 0.0197428
R6037 Vss.n1689 Vss.n184 0.0197428
R6038 Vss.n1599 Vss.n185 0.0197428
R6039 Vss.n1574 Vss.n1573 0.0197428
R6040 Vss.n436 Vss.n203 0.0197428
R6041 Vss.n878 Vss.n488 0.0196349
R6042 Vss.n1855 Vss.n1854 0.0196349
R6043 Vss.n1088 Vss.n1087 0.0196349
R6044 Vss.n1439 Vss.n1438 0.0196349
R6045 Vss.n1890 Vss.n2 0.0196349
R6046 adc_PISO_0.dffrs_4.vss Vss.n1891 0.0170545
R6047 Vss.n428 Vss.n426 0.0164817
R6048 Vss.n1863 Vss.n28 0.0163358
R6049 Vss.n1079 Vss.n304 0.0163358
R6050 Vss.n1447 Vss.n293 0.0163358
R6051 Vss.n1384 Vss.n1383 0.0163358
R6052 Vss.n690 Vss.n511 0.0163358
R6053 Vss.n1888 Vss.n1887 0.0163358
R6054 Vss.n992 Vss.n426 0.0157888
R6055 Vss.n992 Vss.n427 0.0157888
R6056 Vss.n427 Vss.n66 0.0157888
R6057 Vss.n1256 Vss.n66 0.0157888
R6058 Vss.n1256 Vss.n1255 0.0157888
R6059 Vss.n945 Vss.n944 0.0150091
R6060 Vss.n133 Vss.n95 0.0142428
R6061 Vss.n1798 Vss.n93 0.014047
R6062 Vss.n1498 Vss.n1497 0.014047
R6063 Vss.n1494 Vss.n258 0.014047
R6064 Vss.n242 Vss.n225 0.014047
R6065 Vss.n974 Vss.n224 0.014047
R6066 Vss.n877 Vss.n28 0.0139604
R6067 Vss.n304 Vss.n37 0.0139604
R6068 Vss.n1089 Vss.n293 0.0139604
R6069 Vss.n1384 Vss.n1107 0.0139604
R6070 Vss.n659 Vss.n511 0.0139604
R6071 Vss.n1889 Vss.n1888 0.0139604
R6072 Vss.n878 Vss.n877 0.0130367
R6073 Vss.n1854 Vss.n37 0.0130367
R6074 Vss.n1089 Vss.n1088 0.0130367
R6075 Vss.n1438 Vss.n1107 0.0130367
R6076 Vss.n659 Vss.n658 0.0130367
R6077 Vss.n1890 Vss.n1889 0.0130367
R6078 Vss.n453 Vss.n433 0.0121902
R6079 Vss.n1523 Vss.n1522 0.0121902
R6080 Vss.n418 Vss.n400 0.0121902
R6081 Vss.n54 Vss.n53 0.0121902
R6082 Vss.n357 Vss.n356 0.0121902
R6083 Vss.n145 Vss.n144 0.0121902
R6084 Vss.n1150 Vss.n1149 0.0121902
R6085 Vss.n1713 Vss.n175 0.0121902
R6086 Vss.n1419 Vss.n1418 0.0121902
R6087 Vss.n1338 Vss.n1337 0.0121902
R6088 Vss.n1722 Vss.n94 0.0121902
R6089 Vss.n1321 Vss.n1309 0.0121902
R6090 Vss.n256 Vss.n254 0.0121902
R6091 Vss.n1540 Vss.n1539 0.0121902
R6092 Vss.n464 Vss.n402 0.0121902
R6093 Vss.n815 Vss.n814 0.0121902
R6094 Vss.n896 Vss.n895 0.0121902
R6095 Vss.n770 Vss.n768 0.0121902
R6096 Vss.n593 Vss.n592 0.0121902
R6097 Vss.n615 Vss.n614 0.0121902
R6098 Vss.n1785 adc_PISO_0.avss 0.0118245
R6099 Vss.n1218 Vss.n1139 0.0110968
R6100 Vss.n164 Vss.n126 0.0102582
R6101 Vss.n1256 Vss.n90 0.00974555
R6102 Vss.n1493 Vss.n66 0.00974555
R6103 Vss.n984 Vss.n427 0.00974555
R6104 Vss.n992 Vss.n991 0.00974555
R6105 Vss.n1435 Vss.n1108 0.00967928
R6106 Vss.n1255 Vss.n91 0.00967038
R6107 Vss.n970 Vss.n434 0.00915761
R6108 Vss.n321 Vss.n319 0.00915761
R6109 Vss.n1158 Vss.n1157 0.00915761
R6110 Vss.n806 Vss.n805 0.00915761
R6111 Vss.n486 Vss.n485 0.00915761
R6112 Vss.n778 Vss.n777 0.00915761
R6113 Vss.n539 Vss.n536 0.00915761
R6114 Vss.n607 Vss.n606 0.00915761
R6115 Vss.n1140 Vss.n1109 0.00760526
R6116 Vss.n915 Vss.n914 0.00745509
R6117 Vss.n428 SARlogic_0.dffrs_11.vss 0.00734312
R6118 Vss.n344 Vss.n323 0.00720109
R6119 Vss.n1771 Vss.n1770 0.00720109
R6120 Vss.n1357 Vss.n1356 0.00720109
R6121 Vss.n826 Vss.n825 0.00720109
R6122 Vss.n788 Vss.n787 0.00720109
R6123 Vss.n564 Vss.n540 0.00720109
R6124 Vss.n630 Vss.n629 0.00720109
R6125 Vss.n948 Vss.n946 0.00638507
R6126 Vss.n1221 Vss.n1136 0.00617391
R6127 Vss.n1222 Vss.n1221 0.00617391
R6128 Vss.n1217 Vss.n1140 0.00613715
R6129 Vss.n1218 Vss.n1217 0.00613715
R6130 Vss.n1625 Vss 0.00568182
R6131 Vss.n1461 Vss.n283 0.00511663
R6132 Vss.n1058 Vss.n38 0.00511663
R6133 Vss.n860 Vss.n487 0.00511663
R6134 Vss.n656 Vss.n655 0.00511663
R6135 adc_PISO_0.dffrs_4.vss Vss.n0 0.00480909
R6136 Vss.n880 Vss.n39 0.00478552
R6137 SARlogic_0.dffrs_7.vss Vss.n90 0.0044588
R6138 SARlogic_0.dffrs_8.vss Vss.n1493 0.0044588
R6139 Vss.n984 SARlogic_0.dffrs_9.vss 0.0044588
R6140 Vss.n991 SARlogic_0.dffrs_10.vss 0.0044588
R6141 Vss.n1799 SARlogic_0.dffrs_14.vss 0.00438363
R6142 Vss.n1659 comparator_no_offsetcal_0.x4.VSS 0.00371429
R6143 Vss.n1219 Vss.n1218 0.00175057
R6144 Vss.n1323 Vss.n1305 0.000628205
R6145 Vss.n1325 Vss.n1324 0.000628205
R6146 Vss.n1355 Vss.n1354 0.000575167
R6147 Vss.n1279 Vss.n1272 0.000575167
R6148 Vss.n1799 Vss.n91 0.000575167
R6149 Vss.n1255 Vss.n1249 0.000550111
R6150 Vss.n1875 Vss.n1874 0.000544599
R6151 Vss.n967 Vss.n966 0.000544599
R6152 Vss.n332 Vss.n331 0.000544599
R6153 Vss.n1046 Vss.n1045 0.000544599
R6154 Vss.n1209 Vss.n1138 0.000544599
R6155 Vss.n908 Vss.n472 0.000544599
R6156 Vss.n589 Vss.n588 0.000544599
R6157 Vss.n640 Vss.n639 0.000544599
R6158 Vss.n944 Vss.n929 0.000543311
R6159 Vss.n1310 Vss.n1304 0.000542735
R6160 Vss.n1756 Vss.n119 0.000525267
R6161 Vss.n1767 Vss.n122 0.000525056
R6162 Vss.n1353 Vss.n1279 0.000525056
R6163 Vss.n1257 Vss.n1254 0.000525056
R6164 Vss.n1688 Vss.n186 0.000525056
R6165 Vss.n1588 Vss.n1587 0.000525056
R6166 Vss.n1824 Vss.n65 0.000525056
R6167 Vss.n1836 Vss.n57 0.000525056
R6168 Vss.n1576 Vss.n1575 0.000525056
R6169 Vss.n1554 Vss.n1553 0.000525056
R6170 Vss.n1000 Vss.n999 0.000525056
R6171 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t4 41.0041
R6172 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t9 40.8177
R6173 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t8 40.6313
R6174 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t7 27.3166
R6175 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t5 27.1302
R6176 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t6 26.9438
R6177 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.t1 10.0473
R6178 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n4 9.90747
R6179 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n2 9.90116
R6180 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.t2 6.51042
R6181 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.n7 6.04952
R6182 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_6.C.n1 5.7305
R6183 SARlogic_0.dffrs_12.nand3_2.B SARlogic_0.dffrs_12.nand3_6.C.n0 5.47979
R6184 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C.n3 5.13907
R6185 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n9 4.72925
R6186 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_6.C.n5 4.5005
R6187 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.n8 0.732092
R6188 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t3 0.7285
R6189 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t0 0.7285
R6190 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n6 0.449758
R6191 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_2.B 0.166901
R6192 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_0.A 0.0455
R6193 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C 0.0455
R6194 inv2_0.out.n30 inv2_0.out.t25 34.2529
R6195 inv2_0.out.n24 inv2_0.out.t8 34.2529
R6196 inv2_0.out.n18 inv2_0.out.t13 34.2529
R6197 inv2_0.out.n12 inv2_0.out.t21 34.2529
R6198 inv2_0.out.n6 inv2_0.out.t15 34.2529
R6199 inv2_0.out.n1 inv2_0.out.t28 34.2529
R6200 inv2_0.out.n32 inv2_0.out.t20 34.1797
R6201 inv2_0.out.n26 inv2_0.out.t22 34.1797
R6202 inv2_0.out.n20 inv2_0.out.t17 34.1797
R6203 inv2_0.out.n14 inv2_0.out.t5 34.1797
R6204 inv2_0.out.n8 inv2_0.out.t24 34.1797
R6205 inv2_0.out.n3 inv2_0.out.t7 34.1797
R6206 inv2_0.out.n29 inv2_0.out.t31 19.673
R6207 inv2_0.out.n23 inv2_0.out.t11 19.673
R6208 inv2_0.out.n17 inv2_0.out.t12 19.673
R6209 inv2_0.out.n11 inv2_0.out.t27 19.673
R6210 inv2_0.out.n5 inv2_0.out.t19 19.673
R6211 inv2_0.out.n0 inv2_0.out.t2 19.673
R6212 inv2_0.out.n32 inv2_0.out.t9 19.5798
R6213 inv2_0.out.n26 inv2_0.out.t14 19.5798
R6214 inv2_0.out.n20 inv2_0.out.t6 19.5798
R6215 inv2_0.out.n14 inv2_0.out.t26 19.5798
R6216 inv2_0.out.n8 inv2_0.out.t16 19.5798
R6217 inv2_0.out.n3 inv2_0.out.t30 19.5798
R6218 inv2_0.out.n29 inv2_0.out.t18 19.4007
R6219 inv2_0.out.n23 inv2_0.out.t29 19.4007
R6220 inv2_0.out.n17 inv2_0.out.t3 19.4007
R6221 inv2_0.out.n11 inv2_0.out.t10 19.4007
R6222 inv2_0.out.n5 inv2_0.out.t4 19.4007
R6223 inv2_0.out.n0 inv2_0.out.t23 19.4007
R6224 inv2_0.out.n10 inv2_0.out.n4 15.5531
R6225 inv2_0.out.n36 inv2_0.out.t0 9.6935
R6226 inv2_0.out.n34 inv2_0.out.n33 8.46371
R6227 inv2_0.out.n22 inv2_0.out.n21 8.37371
R6228 inv2_0.out.n28 inv2_0.out.n27 8.32871
R6229 inv2_0.out.n16 inv2_0.out.n15 8.32871
R6230 inv2_0.out.n10 inv2_0.out.n9 8.32871
R6231 inv2_0.out.n31 inv2_0.out.n30 7.87164
R6232 inv2_0.out.n25 inv2_0.out.n24 7.87164
R6233 inv2_0.out.n19 inv2_0.out.n18 7.87164
R6234 inv2_0.out.n13 inv2_0.out.n12 7.87164
R6235 inv2_0.out.n7 inv2_0.out.n6 7.87164
R6236 inv2_0.out.n2 inv2_0.out.n1 7.87164
R6237 inv2_0.out.n34 inv2_0.out.n28 7.26762
R6238 inv2_0.out.n16 inv2_0.out.n10 7.22491
R6239 inv2_0.out.n22 inv2_0.out.n16 7.22491
R6240 inv2_0.out.n28 inv2_0.out.n22 7.22491
R6241 inv2_0.out.n33 inv2_0.out.n32 5.00771
R6242 inv2_0.out.n21 inv2_0.out.n20 5.00771
R6243 inv2_0.out.n27 inv2_0.out.n26 4.96432
R6244 inv2_0.out.n15 inv2_0.out.n14 4.96432
R6245 inv2_0.out.n9 inv2_0.out.n8 4.96432
R6246 inv2_0.out.n4 inv2_0.out.n3 4.96432
R6247 inv2_0.out inv2_0.out.n35 4.85086
R6248 inv2_0.out.n36 inv2_0.out.t1 4.35383
R6249 inv2_0.out.n27 inv2_0.out.n25 2.11068
R6250 inv2_0.out.n15 inv2_0.out.n13 2.11068
R6251 inv2_0.out.n9 inv2_0.out.n7 2.11068
R6252 inv2_0.out.n4 inv2_0.out.n2 2.11068
R6253 inv2_0.out.n33 inv2_0.out.n31 2.06729
R6254 inv2_0.out.n21 inv2_0.out.n19 2.06729
R6255 inv2_0.out inv2_0.out.n36 0.254429
R6256 inv2_0.out.n31 adc_PISO_0.2inmux_0.Load 0.2255
R6257 inv2_0.out.n25 adc_PISO_0.2inmux_2.Load 0.2255
R6258 inv2_0.out.n19 adc_PISO_0.2inmux_3.Load 0.2255
R6259 inv2_0.out.n13 adc_PISO_0.2inmux_4.Load 0.2255
R6260 inv2_0.out.n7 adc_PISO_0.2inmux_5.Load 0.2255
R6261 inv2_0.out.n2 adc_PISO_0.2inmux_1.Load 0.2255
R6262 inv2_0.out.n35 inv2_0.out.n34 0.182025
R6263 inv2_0.out.n30 inv2_0.out.n29 0.106438
R6264 inv2_0.out.n24 inv2_0.out.n23 0.106438
R6265 inv2_0.out.n18 inv2_0.out.n17 0.106438
R6266 inv2_0.out.n12 inv2_0.out.n11 0.106438
R6267 inv2_0.out.n6 inv2_0.out.n5 0.106438
R6268 inv2_0.out.n1 inv2_0.out.n0 0.106438
R6269 inv2_0.out.n35 adc_PISO_0.load 0.0294831
R6270 a_37499_31160.n0 a_37499_31160.t5 34.1797
R6271 a_37499_31160.n0 a_37499_31160.t4 19.5798
R6272 a_37499_31160.t1 a_37499_31160.n3 18.7717
R6273 a_37499_31160.n3 a_37499_31160.t0 9.2885
R6274 a_37499_31160.n2 a_37499_31160.n0 4.93379
R6275 a_37499_31160.n1 a_37499_31160.t3 4.23346
R6276 a_37499_31160.n1 a_37499_31160.t2 3.85546
R6277 a_37499_31160.n3 a_37499_31160.n2 0.4055
R6278 a_37499_31160.n2 a_37499_31160.n1 0.352625
R6279 a_n9429_n2007.n12 a_n9429_n2007.n7 11.2899
R6280 a_n9429_n2007.n13 a_n9429_n2007.n12 8.49339
R6281 a_n9429_n2007.n17 a_n9429_n2007.n16 4.89725
R6282 a_n9429_n2007.n9 a_n9429_n2007.n8 4.89725
R6283 a_n9429_n2007.n14 a_n9429_n2007.n5 4.89725
R6284 a_n9429_n2007.n15 a_n9429_n2007.n3 4.89725
R6285 a_n9429_n2007.n2 a_n9429_n2007.n0 4.89725
R6286 a_n9429_n2007.n15 a_n9429_n2007.n4 4.88712
R6287 a_n9429_n2007.n2 a_n9429_n2007.n1 4.88712
R6288 a_n9429_n2007.n18 a_n9429_n2007.n17 4.88712
R6289 a_n9429_n2007.n11 a_n9429_n2007.n10 4.4
R6290 a_n9429_n2007.n13 a_n9429_n2007.n6 4.35275
R6291 a_n9429_n2007.n7 a_n9429_n2007.t10 2.048
R6292 a_n9429_n2007.n7 a_n9429_n2007.t21 2.048
R6293 a_n9429_n2007.n12 a_n9429_n2007.n11 1.95895
R6294 a_n9429_n2007.n16 a_n9429_n2007.t15 1.0925
R6295 a_n9429_n2007.n16 a_n9429_n2007.t6 1.0925
R6296 a_n9429_n2007.n8 a_n9429_n2007.t7 1.0925
R6297 a_n9429_n2007.n8 a_n9429_n2007.t17 1.0925
R6298 a_n9429_n2007.n10 a_n9429_n2007.t2 1.0925
R6299 a_n9429_n2007.n10 a_n9429_n2007.t12 1.0925
R6300 a_n9429_n2007.n5 a_n9429_n2007.t16 1.0925
R6301 a_n9429_n2007.n5 a_n9429_n2007.t1 1.0925
R6302 a_n9429_n2007.n6 a_n9429_n2007.t5 1.0925
R6303 a_n9429_n2007.n6 a_n9429_n2007.t9 1.0925
R6304 a_n9429_n2007.n3 a_n9429_n2007.t18 1.0925
R6305 a_n9429_n2007.n3 a_n9429_n2007.t8 1.0925
R6306 a_n9429_n2007.n4 a_n9429_n2007.t13 1.0925
R6307 a_n9429_n2007.n4 a_n9429_n2007.t3 1.0925
R6308 a_n9429_n2007.n0 a_n9429_n2007.t4 1.0925
R6309 a_n9429_n2007.n0 a_n9429_n2007.t14 1.0925
R6310 a_n9429_n2007.n1 a_n9429_n2007.t11 1.0925
R6311 a_n9429_n2007.n1 a_n9429_n2007.t19 1.0925
R6312 a_n9429_n2007.n18 a_n9429_n2007.t20 1.0925
R6313 a_n9429_n2007.t0 a_n9429_n2007.n18 1.0925
R6314 a_n9429_n2007.n15 a_n9429_n2007.n14 0.849071
R6315 a_n9429_n2007.n9 a_n9429_n2007.n2 0.849071
R6316 a_n9429_n2007.n17 a_n9429_n2007.n2 0.849071
R6317 a_n9429_n2007.n17 a_n9429_n2007.n15 0.849071
R6318 a_n9429_n2007.n14 a_n9429_n2007.n13 0.534875
R6319 a_n9429_n2007.n11 a_n9429_n2007.n9 0.487625
R6320 adc_PISO_0.B2.n3 adc_PISO_0.B2.t9 41.0041
R6321 adc_PISO_0.B2.n4 adc_PISO_0.B2.t7 40.8177
R6322 adc_PISO_0.B2.n7 adc_PISO_0.B2.t8 40.6313
R6323 adc_PISO_0.B2.n1 adc_PISO_0.B2.t4 34.2529
R6324 adc_PISO_0.B2.n6 SARlogic_0.dffrs_9.clk 33.8765
R6325 adc_PISO_0.B2.n7 adc_PISO_0.B2.t5 27.3166
R6326 adc_PISO_0.B2.n4 adc_PISO_0.B2.t12 27.1302
R6327 adc_PISO_0.B2.n3 adc_PISO_0.B2.t11 26.9438
R6328 SARlogic_0.d1 adc_PISO_0.B2 26.2596
R6329 adc_PISO_0.B2.n0 adc_PISO_0.B2.t6 19.673
R6330 adc_PISO_0.B2.n0 adc_PISO_0.B2.t10 19.4007
R6331 adc_PISO_0.B2.n9 adc_PISO_0.B2.n8 14.0582
R6332 adc_PISO_0.B2.n9 adc_PISO_0.B2.n6 11.729
R6333 adc_PISO_0.B2.n12 adc_PISO_0.B2.t2 10.0473
R6334 adc_PISO_0.B2.n2 adc_PISO_0.B2.n1 8.05164
R6335 adc_PISO_0.B2.n11 adc_PISO_0.B2.t3 6.51042
R6336 adc_PISO_0.B2.n11 adc_PISO_0.B2.n10 6.04952
R6337 SARlogic_0.dffrs_9.nand3_1.A adc_PISO_0.B2.n3 5.7755
R6338 SARlogic_0.dffrs_9.nand3_6.B adc_PISO_0.B2.n4 5.47979
R6339 adc_PISO_0.B2.n8 adc_PISO_0.B2.n7 5.13907
R6340 SARlogic_0.dffrs_10.nand3_2.Z adc_PISO_0.B2.n12 4.72925
R6341 adc_PISO_0.B2.n5 SARlogic_0.dffrs_9.nand3_6.B 2.17818
R6342 adc_PISO_0.B2 adc_PISO_0.B2.n2 1.87121
R6343 adc_PISO_0.B2.n5 SARlogic_0.dffrs_9.nand3_1.A 1.34729
R6344 adc_PISO_0.B2.n6 SARlogic_0.d1 0.985679
R6345 adc_PISO_0.B2.n12 adc_PISO_0.B2.n11 0.732092
R6346 adc_PISO_0.B2.n10 adc_PISO_0.B2.t0 0.7285
R6347 adc_PISO_0.B2.n10 adc_PISO_0.B2.t1 0.7285
R6348 SARlogic_0.dffrs_9.clk adc_PISO_0.B2.n5 0.610571
R6349 SARlogic_0.dffrs_10.nand3_2.Z adc_PISO_0.B2.n9 0.166901
R6350 adc_PISO_0.B2.n1 adc_PISO_0.B2.n0 0.106438
R6351 adc_PISO_0.B2.n8 SARlogic_0.dffrs_10.nand3_7.C 0.0455
R6352 adc_PISO_0.B2.n2 adc_PISO_0.2inmux_5.In 0.0455
R6353 a_28027_28820.n0 a_28027_28820.t5 34.1797
R6354 a_28027_28820.n0 a_28027_28820.t4 19.5798
R6355 a_28027_28820.t1 a_28027_28820.n3 18.7717
R6356 a_28027_28820.n3 a_28027_28820.t0 9.2885
R6357 a_28027_28820.n2 a_28027_28820.n0 4.93379
R6358 a_28027_28820.n1 a_28027_28820.t3 4.23346
R6359 a_28027_28820.n1 a_28027_28820.t2 3.85546
R6360 a_28027_28820.n3 a_28027_28820.n2 0.4055
R6361 a_28027_28820.n2 a_28027_28820.n1 0.352625
R6362 Reset.n80 Reset.t25 41.0041
R6363 Reset.n86 Reset.t52 41.0041
R6364 Reset.n66 Reset.t59 41.0041
R6365 Reset.n72 Reset.t1 41.0041
R6366 Reset.n52 Reset.t39 41.0041
R6367 Reset.n58 Reset.t66 41.0041
R6368 Reset.n38 Reset.t48 41.0041
R6369 Reset.n44 Reset.t72 41.0041
R6370 Reset.n24 Reset.t36 41.0041
R6371 Reset.n30 Reset.t64 41.0041
R6372 Reset.n10 Reset.t65 41.0041
R6373 Reset.n16 Reset.t7 41.0041
R6374 Reset.n4 Reset.t38 41.0041
R6375 Reset.n83 Reset.t10 40.8177
R6376 Reset.n82 Reset.t0 40.8177
R6377 Reset.n89 Reset.t26 40.8177
R6378 Reset.n88 Reset.t29 40.8177
R6379 Reset.n69 Reset.t37 40.8177
R6380 Reset.n68 Reset.t28 40.8177
R6381 Reset.n75 Reset.t54 40.8177
R6382 Reset.n74 Reset.t57 40.8177
R6383 Reset.n55 Reset.t30 40.8177
R6384 Reset.n54 Reset.t20 40.8177
R6385 Reset.n61 Reset.t75 40.8177
R6386 Reset.n60 Reset.t51 40.8177
R6387 Reset.n41 Reset.t58 40.8177
R6388 Reset.n40 Reset.t53 40.8177
R6389 Reset.n47 Reset.t42 40.8177
R6390 Reset.n46 Reset.t77 40.8177
R6391 Reset.n27 Reset.t2 40.8177
R6392 Reset.n26 Reset.t78 40.8177
R6393 Reset.n33 Reset.t34 40.8177
R6394 Reset.n32 Reset.t24 40.8177
R6395 Reset.n13 Reset.t76 40.8177
R6396 Reset.n12 Reset.t68 40.8177
R6397 Reset.n19 Reset.t73 40.8177
R6398 Reset.n18 Reset.t13 40.8177
R6399 Reset.n7 Reset.t21 40.8177
R6400 Reset.n6 Reset.t14 40.8177
R6401 Reset.n2 Reset.t63 40.6313
R6402 Reset.n0 Reset.t62 40.6313
R6403 Reset.n2 Reset.t23 27.3166
R6404 Reset.n0 Reset.t79 27.3166
R6405 Reset.n83 Reset.t35 27.1302
R6406 Reset.n82 Reset.t22 27.1302
R6407 Reset.n89 Reset.t45 27.1302
R6408 Reset.n88 Reset.t50 27.1302
R6409 Reset.n69 Reset.t61 27.1302
R6410 Reset.n68 Reset.t49 27.1302
R6411 Reset.n75 Reset.t70 27.1302
R6412 Reset.n74 Reset.t74 27.1302
R6413 Reset.n55 Reset.t55 27.1302
R6414 Reset.n54 Reset.t43 27.1302
R6415 Reset.n61 Reset.t11 27.1302
R6416 Reset.n60 Reset.t67 27.1302
R6417 Reset.n41 Reset.t80 27.1302
R6418 Reset.n40 Reset.t69 27.1302
R6419 Reset.n47 Reset.t60 27.1302
R6420 Reset.n46 Reset.t16 27.1302
R6421 Reset.n27 Reset.t27 27.1302
R6422 Reset.n26 Reset.t17 27.1302
R6423 Reset.n33 Reset.t56 27.1302
R6424 Reset.n32 Reset.t44 27.1302
R6425 Reset.n13 Reset.t18 27.1302
R6426 Reset.n12 Reset.t3 27.1302
R6427 Reset.n19 Reset.t8 27.1302
R6428 Reset.n18 Reset.t31 27.1302
R6429 Reset.n7 Reset.t47 27.1302
R6430 Reset.n6 Reset.t32 27.1302
R6431 Reset.n80 Reset.t81 26.9438
R6432 Reset.n86 Reset.t6 26.9438
R6433 Reset.n66 Reset.t33 26.9438
R6434 Reset.n72 Reset.t5 26.9438
R6435 Reset.n52 Reset.t15 26.9438
R6436 Reset.n58 Reset.t71 26.9438
R6437 Reset.n38 Reset.t19 26.9438
R6438 Reset.n44 Reset.t4 26.9438
R6439 Reset.n24 Reset.t9 26.9438
R6440 Reset.n30 Reset.t46 26.9438
R6441 Reset.n10 Reset.t41 26.9438
R6442 Reset.n16 Reset.t40 26.9438
R6443 Reset.n4 Reset.t12 26.9438
R6444 Reset.n78 SARlogic_0.dffrs_1.resetb 19.0901
R6445 Reset.n64 SARlogic_0.dffrs_2.resetb 19.0901
R6446 Reset.n50 SARlogic_0.dffrs_3.resetb 19.0901
R6447 Reset.n36 SARlogic_0.dffrs_4.resetb 19.0901
R6448 Reset.n22 SARlogic_0.dffrs_5.resetb 19.0901
R6449 Reset.n92 SARlogic_0.dffrs_0.resetb 19.0467
R6450 Reset.n23 SARlogic_0.dffrs_12.resetb 14.0622
R6451 Reset.n84 SARlogic_0.dffrs_14.nand3_1.B 12.1571
R6452 Reset.n90 SARlogic_0.dffrs_0.nand3_1.B 12.1571
R6453 Reset.n70 SARlogic_0.dffrs_7.nand3_1.B 12.1571
R6454 Reset.n76 SARlogic_0.dffrs_1.nand3_1.B 12.1571
R6455 Reset.n56 SARlogic_0.dffrs_8.nand3_1.B 12.1571
R6456 Reset.n62 SARlogic_0.dffrs_2.nand3_1.B 12.1571
R6457 Reset.n42 SARlogic_0.dffrs_9.nand3_1.B 12.1571
R6458 Reset.n48 SARlogic_0.dffrs_3.nand3_1.B 12.1571
R6459 Reset.n28 SARlogic_0.dffrs_10.nand3_1.B 12.1571
R6460 Reset.n34 SARlogic_0.dffrs_4.nand3_1.B 12.1571
R6461 Reset.n14 SARlogic_0.dffrs_11.nand3_1.B 12.1571
R6462 Reset.n20 SARlogic_0.dffrs_5.nand3_1.B 12.1571
R6463 Reset.n8 SARlogic_0.dffrs_12.nand3_1.B 12.1571
R6464 Reset.n3 Reset.n1 9.22229
R6465 Reset.n94 Reset.n93 7.9889
R6466 Reset.n85 Reset.n81 7.75389
R6467 Reset.n91 Reset.n87 7.75389
R6468 Reset.n71 Reset.n67 7.75389
R6469 Reset.n77 Reset.n73 7.75389
R6470 Reset.n57 Reset.n53 7.75389
R6471 Reset.n63 Reset.n59 7.75389
R6472 Reset.n43 Reset.n39 7.75389
R6473 Reset.n49 Reset.n45 7.75389
R6474 Reset.n29 Reset.n25 7.75389
R6475 Reset.n35 Reset.n31 7.75389
R6476 Reset.n15 Reset.n11 7.75389
R6477 Reset.n21 Reset.n17 7.75389
R6478 Reset.n9 Reset.n5 7.75389
R6479 Reset.n94 SARlogic_0.dffrs_13.setb 6.43164
R6480 Reset.n85 Reset.n84 5.93546
R6481 Reset.n91 Reset.n90 5.93546
R6482 Reset.n71 Reset.n70 5.93546
R6483 Reset.n77 Reset.n76 5.93546
R6484 Reset.n57 Reset.n56 5.93546
R6485 Reset.n63 Reset.n62 5.93546
R6486 Reset.n43 Reset.n42 5.93546
R6487 Reset.n49 Reset.n48 5.93546
R6488 Reset.n29 Reset.n28 5.93546
R6489 Reset.n35 Reset.n34 5.93546
R6490 Reset.n15 Reset.n14 5.93546
R6491 Reset.n21 Reset.n20 5.93546
R6492 Reset.n9 Reset.n8 5.93546
R6493 Reset.n78 SARlogic_0.dffrs_7.resetb 5.93246
R6494 Reset.n64 SARlogic_0.dffrs_8.resetb 5.93246
R6495 Reset.n50 SARlogic_0.dffrs_9.resetb 5.93246
R6496 Reset.n36 SARlogic_0.dffrs_10.resetb 5.93246
R6497 Reset.n22 SARlogic_0.dffrs_11.resetb 5.93246
R6498 Reset.n92 SARlogic_0.dffrs_14.resetb 5.88425
R6499 Reset.n81 Reset.n80 5.7305
R6500 Reset.n87 Reset.n86 5.7305
R6501 Reset.n67 Reset.n66 5.7305
R6502 Reset.n73 Reset.n72 5.7305
R6503 Reset.n53 Reset.n52 5.7305
R6504 Reset.n59 Reset.n58 5.7305
R6505 Reset.n39 Reset.n38 5.7305
R6506 Reset.n45 Reset.n44 5.7305
R6507 Reset.n25 Reset.n24 5.7305
R6508 Reset.n31 Reset.n30 5.7305
R6509 Reset.n11 Reset.n10 5.7305
R6510 Reset.n17 Reset.n16 5.7305
R6511 Reset.n5 Reset.n4 5.7305
R6512 SARlogic_0.dffrs_14.nand3_8.B Reset.n83 5.47979
R6513 SARlogic_0.dffrs_14.nand3_1.B Reset.n82 5.47979
R6514 SARlogic_0.dffrs_0.nand3_8.B Reset.n89 5.47979
R6515 SARlogic_0.dffrs_0.nand3_1.B Reset.n88 5.47979
R6516 SARlogic_0.dffrs_7.nand3_8.B Reset.n69 5.47979
R6517 SARlogic_0.dffrs_7.nand3_1.B Reset.n68 5.47979
R6518 SARlogic_0.dffrs_1.nand3_8.B Reset.n75 5.47979
R6519 SARlogic_0.dffrs_1.nand3_1.B Reset.n74 5.47979
R6520 SARlogic_0.dffrs_8.nand3_8.B Reset.n55 5.47979
R6521 SARlogic_0.dffrs_8.nand3_1.B Reset.n54 5.47979
R6522 SARlogic_0.dffrs_2.nand3_8.B Reset.n61 5.47979
R6523 SARlogic_0.dffrs_2.nand3_1.B Reset.n60 5.47979
R6524 SARlogic_0.dffrs_9.nand3_8.B Reset.n41 5.47979
R6525 SARlogic_0.dffrs_9.nand3_1.B Reset.n40 5.47979
R6526 SARlogic_0.dffrs_3.nand3_8.B Reset.n47 5.47979
R6527 SARlogic_0.dffrs_3.nand3_1.B Reset.n46 5.47979
R6528 SARlogic_0.dffrs_10.nand3_8.B Reset.n27 5.47979
R6529 SARlogic_0.dffrs_10.nand3_1.B Reset.n26 5.47979
R6530 SARlogic_0.dffrs_4.nand3_8.B Reset.n33 5.47979
R6531 SARlogic_0.dffrs_4.nand3_1.B Reset.n32 5.47979
R6532 SARlogic_0.dffrs_11.nand3_8.B Reset.n13 5.47979
R6533 SARlogic_0.dffrs_11.nand3_1.B Reset.n12 5.47979
R6534 SARlogic_0.dffrs_5.nand3_8.B Reset.n19 5.47979
R6535 SARlogic_0.dffrs_5.nand3_1.B Reset.n18 5.47979
R6536 SARlogic_0.dffrs_12.nand3_8.B Reset.n7 5.47979
R6537 SARlogic_0.dffrs_12.nand3_1.B Reset.n6 5.47979
R6538 Reset.n3 Reset.n2 5.14711
R6539 Reset.n1 Reset.n0 5.13907
R6540 Reset.n84 SARlogic_0.dffrs_14.nand3_8.B 5.09593
R6541 Reset.n90 SARlogic_0.dffrs_0.nand3_8.B 5.09593
R6542 Reset.n70 SARlogic_0.dffrs_7.nand3_8.B 5.09593
R6543 Reset.n76 SARlogic_0.dffrs_1.nand3_8.B 5.09593
R6544 Reset.n56 SARlogic_0.dffrs_8.nand3_8.B 5.09593
R6545 Reset.n62 SARlogic_0.dffrs_2.nand3_8.B 5.09593
R6546 Reset.n42 SARlogic_0.dffrs_9.nand3_8.B 5.09593
R6547 Reset.n48 SARlogic_0.dffrs_3.nand3_8.B 5.09593
R6548 Reset.n28 SARlogic_0.dffrs_10.nand3_8.B 5.09593
R6549 Reset.n34 SARlogic_0.dffrs_4.nand3_8.B 5.09593
R6550 Reset.n14 SARlogic_0.dffrs_11.nand3_8.B 5.09593
R6551 Reset.n20 SARlogic_0.dffrs_5.nand3_8.B 5.09593
R6552 Reset.n8 SARlogic_0.dffrs_12.nand3_8.B 5.09593
R6553 Reset.n23 Reset.n22 4.5005
R6554 Reset.n37 Reset.n36 4.5005
R6555 Reset.n51 Reset.n50 4.5005
R6556 Reset.n65 Reset.n64 4.5005
R6557 Reset.n79 Reset.n78 4.5005
R6558 Reset.n93 Reset.n92 4.5005
R6559 Reset.n37 Reset.n23 3.6383
R6560 Reset.n51 Reset.n37 3.6383
R6561 Reset.n65 Reset.n51 3.6383
R6562 Reset.n79 Reset.n65 3.6383
R6563 Reset.n93 Reset.n79 3.6113
R6564 SARlogic_0.dffrs_13.setb SARlogic_0.dffrs_13.nand3_0.C 0.783821
R6565 SARlogic_0.reset Reset 0.18425
R6566 SARlogic_0.reset Reset.n94 0.13775
R6567 SARlogic_0.dffrs_14.resetb Reset.n85 0.136036
R6568 SARlogic_0.dffrs_0.resetb Reset.n91 0.136036
R6569 SARlogic_0.dffrs_7.resetb Reset.n71 0.136036
R6570 SARlogic_0.dffrs_1.resetb Reset.n77 0.136036
R6571 SARlogic_0.dffrs_8.resetb Reset.n57 0.136036
R6572 SARlogic_0.dffrs_2.resetb Reset.n63 0.136036
R6573 SARlogic_0.dffrs_9.resetb Reset.n43 0.136036
R6574 SARlogic_0.dffrs_3.resetb Reset.n49 0.136036
R6575 SARlogic_0.dffrs_10.resetb Reset.n29 0.136036
R6576 SARlogic_0.dffrs_4.resetb Reset.n35 0.136036
R6577 SARlogic_0.dffrs_11.resetb Reset.n15 0.136036
R6578 SARlogic_0.dffrs_5.resetb Reset.n21 0.136036
R6579 SARlogic_0.dffrs_12.resetb Reset.n9 0.136036
R6580 Reset.n1 SARlogic_0.dffrs_13.nand3_2.C 0.0455
R6581 Reset.n81 SARlogic_0.dffrs_14.nand3_7.A 0.0455
R6582 Reset.n87 SARlogic_0.dffrs_0.nand3_7.A 0.0455
R6583 Reset.n67 SARlogic_0.dffrs_7.nand3_7.A 0.0455
R6584 Reset.n73 SARlogic_0.dffrs_1.nand3_7.A 0.0455
R6585 Reset.n53 SARlogic_0.dffrs_8.nand3_7.A 0.0455
R6586 Reset.n59 SARlogic_0.dffrs_2.nand3_7.A 0.0455
R6587 Reset.n39 SARlogic_0.dffrs_9.nand3_7.A 0.0455
R6588 Reset.n45 SARlogic_0.dffrs_3.nand3_7.A 0.0455
R6589 Reset.n25 SARlogic_0.dffrs_10.nand3_7.A 0.0455
R6590 Reset.n31 SARlogic_0.dffrs_4.nand3_7.A 0.0455
R6591 Reset.n11 SARlogic_0.dffrs_11.nand3_7.A 0.0455
R6592 Reset.n17 SARlogic_0.dffrs_5.nand3_7.A 0.0455
R6593 Reset.n5 SARlogic_0.dffrs_12.nand3_7.A 0.0455
R6594 SARlogic_0.dffrs_13.nand3_0.C Reset.n3 0.0374643
R6595 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t5 41.0041
R6596 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t4 40.8177
R6597 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t9 40.6313
R6598 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t8 27.3166
R6599 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t6 27.1302
R6600 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t7 26.9438
R6601 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.t0 10.0473
R6602 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n4 9.90747
R6603 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n2 9.90116
R6604 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.t2 6.51042
R6605 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.n7 6.04952
R6606 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_6.C.n1 5.7305
R6607 SARlogic_0.dffrs_14.nand3_2.B SARlogic_0.dffrs_14.nand3_6.C.n0 5.47979
R6608 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C.n3 5.13907
R6609 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n9 4.72925
R6610 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_6.C.n5 4.5005
R6611 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.n8 0.732092
R6612 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t3 0.7285
R6613 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t1 0.7285
R6614 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n6 0.449758
R6615 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_2.B 0.166901
R6616 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_0.A 0.0455
R6617 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C 0.0455
R6618 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t8 41.0041
R6619 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t7 40.8177
R6620 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t6 40.6313
R6621 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t5 27.3166
R6622 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t9 27.1302
R6623 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t4 26.9438
R6624 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.t1 10.0473
R6625 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n4 9.90747
R6626 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n2 9.90116
R6627 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.t0 6.51042
R6628 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.n7 6.04952
R6629 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_6.C.n1 5.7305
R6630 SARlogic_0.dffrs_2.nand3_2.B SARlogic_0.dffrs_2.nand3_6.C.n0 5.47979
R6631 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C.n3 5.13907
R6632 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n9 4.72925
R6633 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_6.C.n5 4.5005
R6634 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.n8 0.732092
R6635 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t2 0.7285
R6636 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t3 0.7285
R6637 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n6 0.449758
R6638 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_2.B 0.166901
R6639 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_0.A 0.0455
R6640 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C 0.0455
R6641 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t4 40.6313
R6642 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t5 27.3166
R6643 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n1 14.2854
R6644 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.t0 10.0473
R6645 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.t1 6.51042
R6646 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.n2 6.04952
R6647 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C.n0 5.13907
R6648 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n4 4.72925
R6649 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.n3 0.732092
R6650 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t3 0.7285
R6651 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t2 0.7285
R6652 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C 0.0455
R6653 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t8 41.0041
R6654 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t5 40.6313
R6655 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t4 40.6313
R6656 SARlogic_0.dffrs_1.Qb SARlogic_0.dffrs_8.setb 28.021
R6657 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t7 27.3166
R6658 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t6 27.3166
R6659 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t9 26.9438
R6660 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.t3 10.0473
R6661 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb.n1 9.84255
R6662 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n3 9.22229
R6663 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.t2 6.51042
R6664 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.n7 6.04952
R6665 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.Qb.n0 5.7305
R6666 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n4 5.14711
R6667 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_1.Qb.n2 5.13907
R6668 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n6 4.94976
R6669 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n9 4.72925
R6670 SARlogic_0.dffrs_8.setb SARlogic_0.dffrs_8.nand3_0.C 0.784786
R6671 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.n8 0.732092
R6672 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t0 0.7285
R6673 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t1 0.7285
R6674 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb 0.175225
R6675 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.nand3_2.A 0.0455
R6676 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_8.nand3_2.C 0.0455
R6677 SARlogic_0.dffrs_8.nand3_0.C SARlogic_0.dffrs_1.Qb.n5 0.0374643
R6678 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t6 41.0041
R6679 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t5 40.8177
R6680 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t7 27.1302
R6681 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t4 26.9438
R6682 SARlogic_0.dffrs_4.nand3_6.A SARlogic_0.dffrs_4.nand3_0.B 17.0041
R6683 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n2 14.8493
R6684 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.t0 10.0473
R6685 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.t1 6.51042
R6686 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.n3 6.04952
R6687 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_8.Z.n0 5.7305
R6688 SARlogic_0.dffrs_4.nand3_0.B SARlogic_0.dffrs_4.nand3_8.Z.n1 5.47979
R6689 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n5 4.72925
R6690 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.n4 0.732092
R6691 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t3 0.7285
R6692 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t2 0.7285
R6693 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_6.A 0.0455
R6694 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t7 40.8177
R6695 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t5 40.6313
R6696 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t6 27.3166
R6697 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t4 27.1302
R6698 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_8.C.n2 14.119
R6699 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.t0 10.0473
R6700 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.t1 6.51042
R6701 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.n4 6.04952
R6702 SARlogic_0.dffrs_4.nand3_7.B SARlogic_0.dffrs_4.nand3_8.C.n0 5.47979
R6703 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C.n1 5.13907
R6704 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n6 4.72925
R6705 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.n5 0.732092
R6706 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t3 0.7285
R6707 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t2 0.7285
R6708 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_7.B 0.438233
R6709 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n3 0.166901
R6710 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C 0.0455
R6711 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t4 40.8177
R6712 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t6 40.6313
R6713 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t7 27.3166
R6714 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t5 27.1302
R6715 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_8.C.n2 14.119
R6716 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.t1 10.0473
R6717 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.t0 6.51042
R6718 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.n4 6.04952
R6719 SARlogic_0.dffrs_1.nand3_7.B SARlogic_0.dffrs_1.nand3_8.C.n0 5.47979
R6720 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C.n1 5.13907
R6721 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n6 4.72925
R6722 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.n5 0.732092
R6723 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t2 0.7285
R6724 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t3 0.7285
R6725 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_7.B 0.438233
R6726 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n3 0.166901
R6727 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C 0.0455
R6728 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t6 40.8177
R6729 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t7 40.6313
R6730 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t4 27.3166
R6731 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t5 27.1302
R6732 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_8.C.n2 14.119
R6733 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.t0 10.0473
R6734 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.t1 6.51042
R6735 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.n4 6.04952
R6736 SARlogic_0.dffrs_5.nand3_7.B SARlogic_0.dffrs_5.nand3_8.C.n0 5.47979
R6737 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C.n1 5.13907
R6738 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n6 4.72925
R6739 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.n5 0.732092
R6740 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t3 0.7285
R6741 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t2 0.7285
R6742 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_7.B 0.438233
R6743 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n3 0.166901
R6744 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C 0.0455
R6745 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t4 41.0041
R6746 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t7 40.8177
R6747 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t6 27.1302
R6748 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t5 26.9438
R6749 SARlogic_0.dffrs_3.nand3_6.A SARlogic_0.dffrs_3.nand3_0.B 17.0041
R6750 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n2 14.8493
R6751 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.t3 10.0473
R6752 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.t1 6.51042
R6753 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.n3 6.04952
R6754 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_8.Z.n0 5.7305
R6755 SARlogic_0.dffrs_3.nand3_0.B SARlogic_0.dffrs_3.nand3_8.Z.n1 5.47979
R6756 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n5 4.72925
R6757 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.n4 0.732092
R6758 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t2 0.7285
R6759 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t0 0.7285
R6760 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_6.A 0.0455
R6761 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t7 40.8177
R6762 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t5 40.6313
R6763 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t6 27.3166
R6764 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t4 27.1302
R6765 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_8.C.n2 14.119
R6766 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.t0 10.0473
R6767 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.t1 6.51042
R6768 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.n4 6.04952
R6769 SARlogic_0.dffrs_3.nand3_7.B SARlogic_0.dffrs_3.nand3_8.C.n0 5.47979
R6770 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C.n1 5.13907
R6771 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n6 4.72925
R6772 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.n5 0.732092
R6773 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t2 0.7285
R6774 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t3 0.7285
R6775 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_7.B 0.438233
R6776 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n3 0.166901
R6777 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C 0.0455
R6778 a_33257_31423.n1 a_33257_31423.t5 41.0041
R6779 a_33257_31423.n0 a_33257_31423.t6 40.8177
R6780 a_33257_31423.n2 a_33257_31423.t9 40.6313
R6781 a_33257_31423.n2 a_33257_31423.t4 27.3166
R6782 a_33257_31423.n0 a_33257_31423.t8 27.1302
R6783 a_33257_31423.n1 a_33257_31423.t7 26.9438
R6784 a_33257_31423.n3 a_33257_31423.n1 15.6312
R6785 a_33257_31423.n3 a_33257_31423.n2 15.046
R6786 a_33257_31423.n5 a_33257_31423.t1 10.0473
R6787 a_33257_31423.n6 a_33257_31423.t3 6.51042
R6788 a_33257_31423.n7 a_33257_31423.n6 6.04952
R6789 a_33257_31423.n4 a_33257_31423.n0 5.64619
R6790 a_33257_31423.n5 a_33257_31423.n4 5.17851
R6791 a_33257_31423.n4 a_33257_31423.n3 4.5005
R6792 a_33257_31423.n6 a_33257_31423.n5 0.732092
R6793 a_33257_31423.n7 a_33257_31423.t2 0.7285
R6794 a_33257_31423.t0 a_33257_31423.n7 0.7285
R6795 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t8 41.0041
R6796 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t7 40.8177
R6797 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t4 40.6313
R6798 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t5 27.3166
R6799 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t9 27.1302
R6800 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t6 26.9438
R6801 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.t2 10.0473
R6802 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n4 9.90747
R6803 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n2 9.90116
R6804 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.t1 6.51042
R6805 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.n7 6.04952
R6806 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_6.C.n1 5.7305
R6807 SARlogic_0.dffrs_5.nand3_2.B SARlogic_0.dffrs_5.nand3_6.C.n0 5.47979
R6808 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C.n3 5.13907
R6809 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n9 4.72925
R6810 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_6.C.n5 4.5005
R6811 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.n8 0.732092
R6812 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t3 0.7285
R6813 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t0 0.7285
R6814 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n6 0.449758
R6815 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_2.B 0.166901
R6816 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_0.A 0.0455
R6817 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C 0.0455
R6818 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t6 40.8177
R6819 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t5 40.6313
R6820 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t7 27.3166
R6821 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t4 27.1302
R6822 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_8.C.n2 14.119
R6823 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.t0 10.0473
R6824 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.t1 6.51042
R6825 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.n4 6.04952
R6826 SARlogic_0.dffrs_12.nand3_7.B SARlogic_0.dffrs_12.nand3_8.C.n0 5.47979
R6827 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C.n1 5.13907
R6828 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n6 4.72925
R6829 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.n5 0.732092
R6830 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t2 0.7285
R6831 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t3 0.7285
R6832 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_7.B 0.438233
R6833 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n3 0.166901
R6834 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C 0.0455
R6835 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t16 49.7997
R6836 comparator_no_offsetcal_0.x3.in comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t11 31.5367
R6837 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t9 19.735
R6838 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 18.0852
R6839 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t8 16.9998
R6840 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t15 14.5537
R6841 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 14.2885
R6842 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t17 13.6729
R6843 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t12 13.3844
R6844 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t14 13.3445
R6845 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 11.24
R6846 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 7.16477
R6847 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 6.95627
R6848 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 6.75194
R6849 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 6.32624
R6850 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t10 5.04666
R6851 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t13 4.84137
R6852 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 2.836
R6853 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 2.75432
R6854 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t2 1.8205
R6855 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t4 1.8205
R6856 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t6 1.8205
R6857 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t0 1.8205
R6858 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t5 0.8195
R6859 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t3 0.8195
R6860 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t7 0.8195
R6861 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t1 0.8195
R6862 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 0.733357
R6863 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 0.440894
R6864 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 0.426875
R6865 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 0.289009
R6866 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 0.0607115
R6867 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 comparator_no_offsetcal_0.x3.in 0.014
R6868 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t16 49.7997
R6869 comparator_no_offsetcal_0.x5.in comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t12 31.5367
R6870 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t10 19.735
R6871 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t9 18.9075
R6872 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t8 16.9998
R6873 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t14 13.6729
R6874 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t11 13.3844
R6875 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t17 13.3445
R6876 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 12.247
R6877 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 11.2403
R6878 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 9.4181
R6879 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 7.4449
R6880 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 6.95074
R6881 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 6.75194
R6882 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 6.32761
R6883 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t15 5.04666
R6884 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 4.94262
R6885 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t13 4.84137
R6886 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 2.836
R6887 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 2.75432
R6888 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t6 1.8205
R6889 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t5 1.8205
R6890 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t7 1.8205
R6891 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t4 1.8205
R6892 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t1 0.8195
R6893 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t2 0.8195
R6894 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t3 0.8195
R6895 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t0 0.8195
R6896 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 0.733357
R6897 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 0.5315
R6898 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 0.289009
R6899 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 0.184462
R6900 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 comparator_no_offsetcal_0.x5.in 0.014
R6901 Clk.n0 Clk.t23 41.0041
R6902 Clk.n22 Clk.t5 41.0041
R6903 Clk.n18 Clk.t24 41.0041
R6904 Clk.n14 Clk.t14 41.0041
R6905 Clk.n10 Clk.t1 41.0041
R6906 Clk.n6 Clk.t10 41.0041
R6907 Clk.n3 Clk.t28 41.0041
R6908 Clk.n1 Clk.t25 40.8177
R6909 Clk.n23 Clk.t8 40.8177
R6910 Clk.n19 Clk.t20 40.8177
R6911 Clk.n15 Clk.t17 40.8177
R6912 Clk.n11 Clk.t29 40.8177
R6913 Clk.n7 Clk.t6 40.8177
R6914 Clk.n4 Clk.t2 40.8177
R6915 Clk.n1 Clk.t19 27.1302
R6916 Clk.n23 Clk.t26 27.1302
R6917 Clk.n19 Clk.t4 27.1302
R6918 Clk.n15 Clk.t15 27.1302
R6919 Clk.n11 Clk.t32 27.1302
R6920 Clk.n7 Clk.t30 27.1302
R6921 Clk.n4 Clk.t13 27.1302
R6922 Clk.n0 Clk.t31 26.9438
R6923 Clk.n22 Clk.t16 26.9438
R6924 Clk.n18 Clk.t0 26.9438
R6925 Clk.n14 Clk.t21 26.9438
R6926 Clk.n10 Clk.t7 26.9438
R6927 Clk.n6 Clk.t18 26.9438
R6928 Clk.n3 Clk.t3 26.9438
R6929 Clk.n31 Clk.t12 21.1483
R6930 Clk.n30 Clk.t11 21.1483
R6931 Clk.n29 Clk.t22 21.1483
R6932 Clk.n28 Clk.t9 21.1483
R6933 Clk.n27 Clk.t27 20.5929
R6934 Clk.n9 SARlogic_0.dffrs_5.clk 20.5278
R6935 Clk.n28 Clk.n27 19.1491
R6936 Clk.n21 SARlogic_0.dffrs_1.clk 16.89
R6937 Clk.n17 SARlogic_0.dffrs_2.clk 16.89
R6938 Clk.n13 SARlogic_0.dffrs_3.clk 16.89
R6939 Clk.n9 SARlogic_0.dffrs_4.clk 16.89
R6940 Clk.n25 SARlogic_0.dffrs_0.clk 16.8417
R6941 Clk.n32 Clk.n31 15.5861
R6942 Clk.n26 SARlogic_0.dffrs_13.clk 12.2453
R6943 SARlogic_0.clk Clk.n33 11.0885
R6944 Clk.n26 Clk.n25 8.1113
R6945 SARlogic_0.dffrs_13.nand3_1.A Clk.n0 5.7755
R6946 SARlogic_0.dffrs_0.nand3_1.A Clk.n22 5.7755
R6947 SARlogic_0.dffrs_1.nand3_1.A Clk.n18 5.7755
R6948 SARlogic_0.dffrs_2.nand3_1.A Clk.n14 5.7755
R6949 SARlogic_0.dffrs_3.nand3_1.A Clk.n10 5.7755
R6950 SARlogic_0.dffrs_4.nand3_1.A Clk.n6 5.7755
R6951 SARlogic_0.dffrs_5.nand3_1.A Clk.n3 5.7755
R6952 SARlogic_0.dffrs_13.nand3_6.B Clk.n1 5.47979
R6953 SARlogic_0.dffrs_0.nand3_6.B Clk.n23 5.47979
R6954 SARlogic_0.dffrs_1.nand3_6.B Clk.n19 5.47979
R6955 SARlogic_0.dffrs_2.nand3_6.B Clk.n15 5.47979
R6956 SARlogic_0.dffrs_3.nand3_6.B Clk.n11 5.47979
R6957 SARlogic_0.dffrs_4.nand3_6.B Clk.n7 5.47979
R6958 SARlogic_0.dffrs_5.nand3_6.B Clk.n4 5.47979
R6959 Clk.n33 comparator_no_offsetcal_0.CLK 5.39581
R6960 Clk.n30 Clk.n29 4.47208
R6961 Clk.n13 Clk.n9 3.6383
R6962 Clk.n17 Clk.n13 3.6383
R6963 Clk.n21 Clk.n17 3.6383
R6964 Clk.n25 Clk.n21 3.6113
R6965 Clk.n32 Clk.n27 3.56405
R6966 Clk.n2 SARlogic_0.dffrs_13.nand3_6.B 2.17818
R6967 Clk.n24 SARlogic_0.dffrs_0.nand3_6.B 2.17818
R6968 Clk.n20 SARlogic_0.dffrs_1.nand3_6.B 2.17818
R6969 Clk.n16 SARlogic_0.dffrs_2.nand3_6.B 2.17818
R6970 Clk.n12 SARlogic_0.dffrs_3.nand3_6.B 2.17818
R6971 Clk.n8 SARlogic_0.dffrs_4.nand3_6.B 2.17818
R6972 Clk.n5 SARlogic_0.dffrs_5.nand3_6.B 2.17818
R6973 Clk.n2 SARlogic_0.dffrs_13.nand3_1.A 1.34729
R6974 Clk.n24 SARlogic_0.dffrs_0.nand3_1.A 1.34729
R6975 Clk.n20 SARlogic_0.dffrs_1.nand3_1.A 1.34729
R6976 Clk.n16 SARlogic_0.dffrs_2.nand3_1.A 1.34729
R6977 Clk.n12 SARlogic_0.dffrs_3.nand3_1.A 1.34729
R6978 Clk.n8 SARlogic_0.dffrs_4.nand3_1.A 1.34729
R6979 Clk.n5 SARlogic_0.dffrs_5.nand3_1.A 1.34729
R6980 comparator_no_offsetcal_0.CLK Clk.n32 1.32418
R6981 Clk.n29 Clk.n28 1.01892
R6982 Clk.n31 Clk.n30 1.01892
R6983 SARlogic_0.dffrs_13.clk Clk.n2 0.611214
R6984 SARlogic_0.dffrs_0.clk Clk.n24 0.611214
R6985 SARlogic_0.dffrs_1.clk Clk.n20 0.611214
R6986 SARlogic_0.dffrs_2.clk Clk.n16 0.611214
R6987 SARlogic_0.dffrs_3.clk Clk.n12 0.611214
R6988 SARlogic_0.dffrs_4.clk Clk.n8 0.611214
R6989 SARlogic_0.dffrs_5.clk Clk.n5 0.611214
R6990 Clk.n33 Clk 0.514034
R6991 SARlogic_0.clk Clk.n26 0.13775
R6992 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t8 41.0041
R6993 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t6 40.8177
R6994 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t7 40.6313
R6995 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t4 27.3166
R6996 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t9 27.1302
R6997 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t5 26.9438
R6998 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.t1 10.0473
R6999 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n4 9.90747
R7000 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n2 9.90116
R7001 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.t2 6.51042
R7002 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.n7 6.04952
R7003 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_6.C.n1 5.7305
R7004 SARlogic_0.dffrs_1.nand3_2.B SARlogic_0.dffrs_1.nand3_6.C.n0 5.47979
R7005 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C.n3 5.13907
R7006 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n9 4.72925
R7007 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_6.C.n5 4.5005
R7008 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.n8 0.732092
R7009 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t3 0.7285
R7010 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t0 0.7285
R7011 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n6 0.449758
R7012 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_2.B 0.166901
R7013 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_0.A 0.0455
R7014 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C 0.0455
R7015 adc_PISO_0.B3.n3 adc_PISO_0.B3.t5 41.0041
R7016 adc_PISO_0.B3.n4 adc_PISO_0.B3.t11 40.8177
R7017 adc_PISO_0.B3.n7 adc_PISO_0.B3.t4 40.6313
R7018 adc_PISO_0.B3.n1 adc_PISO_0.B3.t6 34.2529
R7019 adc_PISO_0.B3.n6 SARlogic_0.dffrs_8.clk 34.1594
R7020 adc_PISO_0.B3.n7 adc_PISO_0.B3.t10 27.3166
R7021 adc_PISO_0.B3.n4 adc_PISO_0.B3.t9 27.1302
R7022 adc_PISO_0.B3.n3 adc_PISO_0.B3.t7 26.9438
R7023 adc_PISO_0.B3.n0 adc_PISO_0.B3.t8 19.673
R7024 adc_PISO_0.B3.n0 adc_PISO_0.B3.t12 19.4007
R7025 SARlogic_0.d2 adc_PISO_0.B3 17.5376
R7026 adc_PISO_0.B3.n9 adc_PISO_0.B3.n8 14.0582
R7027 adc_PISO_0.B3.n9 adc_PISO_0.B3.n6 12.0118
R7028 adc_PISO_0.B3.n12 adc_PISO_0.B3.t0 10.0473
R7029 adc_PISO_0.B3.n2 adc_PISO_0.B3.n1 8.05164
R7030 adc_PISO_0.B3.n11 adc_PISO_0.B3.t1 6.51042
R7031 adc_PISO_0.B3.n11 adc_PISO_0.B3.n10 6.04952
R7032 SARlogic_0.dffrs_8.nand3_1.A adc_PISO_0.B3.n3 5.7755
R7033 SARlogic_0.dffrs_8.nand3_6.B adc_PISO_0.B3.n4 5.47979
R7034 adc_PISO_0.B3.n8 adc_PISO_0.B3.n7 5.13907
R7035 SARlogic_0.dffrs_9.nand3_2.Z adc_PISO_0.B3.n12 4.72925
R7036 adc_PISO_0.B3.n5 SARlogic_0.dffrs_8.nand3_6.B 2.17818
R7037 adc_PISO_0.B3 adc_PISO_0.B3.n2 1.87121
R7038 adc_PISO_0.B3.n5 SARlogic_0.dffrs_8.nand3_1.A 1.34729
R7039 adc_PISO_0.B3.n12 adc_PISO_0.B3.n11 0.732092
R7040 adc_PISO_0.B3.n10 adc_PISO_0.B3.t3 0.7285
R7041 adc_PISO_0.B3.n10 adc_PISO_0.B3.t2 0.7285
R7042 adc_PISO_0.B3.n6 SARlogic_0.d2 0.698
R7043 SARlogic_0.dffrs_8.clk adc_PISO_0.B3.n5 0.610571
R7044 SARlogic_0.dffrs_9.nand3_2.Z adc_PISO_0.B3.n9 0.166901
R7045 adc_PISO_0.B3.n1 adc_PISO_0.B3.n0 0.106438
R7046 adc_PISO_0.B3.n8 SARlogic_0.dffrs_9.nand3_7.C 0.0455
R7047 adc_PISO_0.B3.n2 adc_PISO_0.2inmux_4.In 0.0455
R7048 a_4841_31422.n1 a_4841_31422.t4 41.0041
R7049 a_4841_31422.n0 a_4841_31422.t6 40.8177
R7050 a_4841_31422.n2 a_4841_31422.t7 40.6313
R7051 a_4841_31422.n2 a_4841_31422.t9 27.3166
R7052 a_4841_31422.n0 a_4841_31422.t8 27.1302
R7053 a_4841_31422.n1 a_4841_31422.t5 26.9438
R7054 a_4841_31422.n3 a_4841_31422.n1 15.6312
R7055 a_4841_31422.n3 a_4841_31422.n2 15.046
R7056 a_4841_31422.n5 a_4841_31422.t2 10.0473
R7057 a_4841_31422.t0 a_4841_31422.n7 6.51042
R7058 a_4841_31422.n7 a_4841_31422.n6 6.04952
R7059 a_4841_31422.n4 a_4841_31422.n0 5.64619
R7060 a_4841_31422.n5 a_4841_31422.n4 5.17851
R7061 a_4841_31422.n4 a_4841_31422.n3 4.5005
R7062 a_4841_31422.n7 a_4841_31422.n5 0.732092
R7063 a_4841_31422.n6 a_4841_31422.t1 0.7285
R7064 a_4841_31422.n6 a_4841_31422.t3 0.7285
R7065 a_4841_33627.n0 a_4841_33627.t4 40.6313
R7066 a_4841_33627.n0 a_4841_33627.t5 27.3166
R7067 a_4841_33627.n1 a_4841_33627.n0 24.1527
R7068 a_4841_33627.n1 a_4841_33627.t1 10.0473
R7069 a_4841_33627.t0 a_4841_33627.n3 6.51042
R7070 a_4841_33627.n3 a_4841_33627.n2 6.04952
R7071 a_4841_33627.n3 a_4841_33627.n1 0.732092
R7072 a_4841_33627.n2 a_4841_33627.t3 0.7285
R7073 a_4841_33627.n2 a_4841_33627.t2 0.7285
R7074 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t6 40.6313
R7075 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.t4 34.1066
R7076 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t7 27.3166
R7077 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t5 19.673
R7078 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t8 19.4007
R7079 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n3 14.6967
R7080 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.t3 10.0473
R7081 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n6 9.39565
R7082 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit.n1 6.70486
R7083 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.t2 6.51042
R7084 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.n4 6.04952
R7085 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n2 5.81514
R7086 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.n5 0.732092
R7087 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t0 0.7285
R7088 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t1 0.7285
R7089 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n7 0.458082
R7090 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.n0 0.252687
R7091 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit 0.0519286
R7092 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t4 40.6313
R7093 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t5 27.3166
R7094 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n1 14.2854
R7095 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.t1 10.0473
R7096 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.t2 6.51042
R7097 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.n2 6.04952
R7098 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C.n0 5.13907
R7099 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n4 4.72925
R7100 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.n3 0.732092
R7101 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t0 0.7285
R7102 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t3 0.7285
R7103 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C 0.0455
R7104 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t5 41.0041
R7105 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t6 40.8177
R7106 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t4 40.6313
R7107 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t9 27.3166
R7108 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t7 27.1302
R7109 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t8 26.9438
R7110 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.t1 10.0473
R7111 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n4 9.90747
R7112 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n2 9.90116
R7113 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.t2 6.51042
R7114 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.n7 6.04952
R7115 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_6.C.n1 5.7305
R7116 SARlogic_0.dffrs_3.nand3_2.B SARlogic_0.dffrs_3.nand3_6.C.n0 5.47979
R7117 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C.n3 5.13907
R7118 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n9 4.72925
R7119 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_6.C.n5 4.5005
R7120 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.n8 0.732092
R7121 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t3 0.7285
R7122 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t0 0.7285
R7123 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n6 0.449758
R7124 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_2.B 0.166901
R7125 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_0.A 0.0455
R7126 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C 0.0455
R7127 a_33337_30170.n0 a_33337_30170.t7 41.0041
R7128 a_33337_30170.n1 a_33337_30170.t4 40.8177
R7129 a_33337_30170.n1 a_33337_30170.t6 27.1302
R7130 a_33337_30170.n0 a_33337_30170.t5 26.9438
R7131 a_33337_30170.n2 a_33337_30170.n1 22.5284
R7132 a_33337_30170.n3 a_33337_30170.n2 19.5781
R7133 a_33337_30170.n3 a_33337_30170.t3 10.0473
R7134 a_33337_30170.t0 a_33337_30170.n5 6.51042
R7135 a_33337_30170.n5 a_33337_30170.n4 6.04952
R7136 a_33337_30170.n2 a_33337_30170.n0 5.7305
R7137 a_33337_30170.n5 a_33337_30170.n3 0.732092
R7138 a_33337_30170.n4 a_33337_30170.t2 0.7285
R7139 a_33337_30170.n4 a_33337_30170.t1 0.7285
R7140 a_33257_33628.n0 a_33257_33628.t4 40.6313
R7141 a_33257_33628.n0 a_33257_33628.t5 27.3166
R7142 a_33257_33628.n1 a_33257_33628.n0 24.1527
R7143 a_33257_33628.n1 a_33257_33628.t2 10.0473
R7144 a_33257_33628.n2 a_33257_33628.t1 6.51042
R7145 a_33257_33628.n3 a_33257_33628.n2 6.04952
R7146 a_33257_33628.n2 a_33257_33628.n1 0.732092
R7147 a_33257_33628.t0 a_33257_33628.n3 0.7285
R7148 a_33257_33628.n3 a_33257_33628.t3 0.7285
R7149 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t5 41.0041
R7150 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t4 40.6313
R7151 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t6 27.3166
R7152 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t7 26.9438
R7153 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d 17.5022
R7154 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d.n2 14.0582
R7155 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.t1 10.0473
R7156 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.t0 6.51042
R7157 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.n4 6.04952
R7158 SARlogic_0.dffrs_0.nand3_8.A SARlogic_0.dffrs_0.d.n0 5.7755
R7159 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_0.d.n1 5.13907
R7160 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n6 4.72925
R7161 SARlogic_0.dffrs_0.d SARlogic_0.dffrs_0.nand3_8.A 0.783821
R7162 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.n5 0.732092
R7163 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t2 0.7285
R7164 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t3 0.7285
R7165 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n3 0.166901
R7166 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_13.nand3_7.C 0.0455
R7167 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t7 41.0041
R7168 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t4 40.6313
R7169 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t8 40.6313
R7170 SARlogic_0.dffrs_13.Qb SARlogic_0.dffrs_14.setb 27.9776
R7171 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t6 27.3166
R7172 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t5 27.3166
R7173 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t9 26.9438
R7174 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.t1 10.0473
R7175 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb.n1 9.84255
R7176 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n3 9.22229
R7177 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.t2 6.51042
R7178 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.n7 6.04952
R7179 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.Qb.n0 5.7305
R7180 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n4 5.14711
R7181 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_13.Qb.n2 5.13907
R7182 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n6 4.94976
R7183 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n9 4.72925
R7184 SARlogic_0.dffrs_14.setb SARlogic_0.dffrs_14.nand3_0.C 0.784786
R7185 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.n8 0.732092
R7186 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t3 0.7285
R7187 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t0 0.7285
R7188 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb 0.175225
R7189 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.nand3_2.A 0.0455
R7190 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_14.nand3_2.C 0.0455
R7191 SARlogic_0.dffrs_14.nand3_0.C SARlogic_0.dffrs_13.Qb.n5 0.0374643
R7192 Comp_out.n9 Comp_out 11.2807
R7193 Comp_out.n5 Comp_out.n4 6.5435
R7194 Comp_out.n2 Comp_out.n1 6.5435
R7195 comparator_no_offsetcal_0.x4.Y Comp_out.n8 4.5005
R7196 Comp_out.n9 comparator_no_offsetcal_0.x4.Y 2.3842
R7197 Comp_out.n6 Comp_out.n3 2.17483
R7198 Comp_out.n4 Comp_out.t1 2.03874
R7199 Comp_out.n4 Comp_out.t2 2.03874
R7200 Comp_out.n1 Comp_out.t0 2.03874
R7201 Comp_out.n1 Comp_out.t3 2.03874
R7202 Comp_out.n8 Comp_out.n0 2.00383
R7203 Comp_out.n0 Comp_out.t7 1.13285
R7204 Comp_out.n0 Comp_out.t6 1.13285
R7205 Comp_out.n3 Comp_out.t4 1.13285
R7206 Comp_out.n3 Comp_out.t5 1.13285
R7207 Comp_out.n5 Comp_out.n2 0.5105
R7208 Comp_out.n7 Comp_out.n6 0.5105
R7209 Comp_out.n7 Comp_out.n2 0.2165
R7210 Comp_out.n6 Comp_out.n5 0.2165
R7211 Comp_out.n8 Comp_out.n7 0.1175
R7212 comparator_no_offsetcal_0.Vout Comp_out.n9 0.0311818
R7213 a_9083_28820.n0 a_9083_28820.t4 34.1797
R7214 a_9083_28820.n0 a_9083_28820.t5 19.5798
R7215 a_9083_28820.t1 a_9083_28820.n3 18.7717
R7216 a_9083_28820.n3 a_9083_28820.t0 9.2885
R7217 a_9083_28820.n2 a_9083_28820.n0 4.93379
R7218 a_9083_28820.n1 a_9083_28820.t3 4.23346
R7219 a_9083_28820.n1 a_9083_28820.t2 3.85546
R7220 a_9083_28820.n3 a_9083_28820.n2 0.4055
R7221 a_9083_28820.n2 a_9083_28820.n1 0.352625
R7222 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t7 41.0041
R7223 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t8 40.8177
R7224 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t6 40.6313
R7225 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t5 27.3166
R7226 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t4 27.1302
R7227 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t9 26.9438
R7228 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.t1 10.0473
R7229 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n4 9.90747
R7230 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n2 9.90116
R7231 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.t2 6.51042
R7232 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.n7 6.04952
R7233 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_6.C.n1 5.7305
R7234 SARlogic_0.dffrs_9.nand3_2.B SARlogic_0.dffrs_9.nand3_6.C.n0 5.47979
R7235 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C.n3 5.13907
R7236 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n9 4.72925
R7237 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_6.C.n5 4.5005
R7238 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.n8 0.732092
R7239 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t3 0.7285
R7240 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t0 0.7285
R7241 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n6 0.449758
R7242 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_2.B 0.166901
R7243 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_0.A 0.0455
R7244 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C 0.0455
R7245 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t6 40.8177
R7246 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t7 40.6313
R7247 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t4 27.3166
R7248 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t5 27.1302
R7249 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_8.C.n2 14.119
R7250 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.t2 10.0473
R7251 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.t1 6.51042
R7252 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.n4 6.04952
R7253 SARlogic_0.dffrs_2.nand3_7.B SARlogic_0.dffrs_2.nand3_8.C.n0 5.47979
R7254 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C.n1 5.13907
R7255 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n6 4.72925
R7256 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.n5 0.732092
R7257 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t3 0.7285
R7258 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t0 0.7285
R7259 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_7.B 0.438233
R7260 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n3 0.166901
R7261 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C 0.0455
R7262 a_30255_29264.n0 a_30255_29264.t5 34.1797
R7263 a_30255_29264.n0 a_30255_29264.t4 19.5798
R7264 a_30255_29264.n1 a_30255_29264.t3 10.3401
R7265 a_30255_29264.n1 a_30255_29264.t2 9.2885
R7266 a_30255_29264.n2 a_30255_29264.n0 4.93379
R7267 a_30255_29264.n3 a_30255_29264.t0 4.09202
R7268 a_30255_29264.t1 a_30255_29264.n3 3.95079
R7269 a_30255_29264.n2 a_30255_29264.n1 0.599711
R7270 a_30255_29264.n3 a_30255_29264.n2 0.296375
R7271 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t3 41.0041
R7272 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t2 26.9438
R7273 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t0 9.6935
R7274 adc_PISO_0.dffrs_4.d adc_PISO_0.2inmux_5.OUT.n0 6.55979
R7275 adc_PISO_0.2inmux_5.OUT adc_PISO_0.dffrs_4.d 4.883
R7276 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t1 4.35383
R7277 adc_PISO_0.2inmux_5.OUT adc_PISO_0.2inmux_5.OUT.n1 0.350857
R7278 adc_PISO_0.B1.n3 adc_PISO_0.B1.t4 41.0041
R7279 adc_PISO_0.B1.n4 adc_PISO_0.B1.t10 40.8177
R7280 adc_PISO_0.B1.n7 adc_PISO_0.B1.t5 40.6313
R7281 adc_PISO_0.B1.n6 adc_PISO_0.B1 36.2544
R7282 adc_PISO_0.B1.n1 adc_PISO_0.B1.t9 34.2529
R7283 adc_PISO_0.B1.n6 SARlogic_0.dffrs_10.clk 33.5936
R7284 adc_PISO_0.B1.n7 adc_PISO_0.B1.t12 27.3166
R7285 adc_PISO_0.B1.n4 adc_PISO_0.B1.t7 27.1302
R7286 adc_PISO_0.B1.n3 adc_PISO_0.B1.t6 26.9438
R7287 adc_PISO_0.B1.n0 adc_PISO_0.B1.t11 19.673
R7288 adc_PISO_0.B1.n0 adc_PISO_0.B1.t8 19.4007
R7289 adc_PISO_0.B1.n9 adc_PISO_0.B1.n8 14.0582
R7290 adc_PISO_0.B1.n9 adc_PISO_0.B1.n6 11.4461
R7291 adc_PISO_0.B1.n12 adc_PISO_0.B1.t0 10.0473
R7292 adc_PISO_0.B1.n2 adc_PISO_0.B1.n1 8.05164
R7293 adc_PISO_0.B1.n11 adc_PISO_0.B1.t1 6.51042
R7294 adc_PISO_0.B1.n11 adc_PISO_0.B1.n10 6.04952
R7295 SARlogic_0.dffrs_10.nand3_1.A adc_PISO_0.B1.n3 5.7755
R7296 SARlogic_0.dffrs_10.nand3_6.B adc_PISO_0.B1.n4 5.47979
R7297 adc_PISO_0.B1.n8 adc_PISO_0.B1.n7 5.13907
R7298 SARlogic_0.dffrs_11.nand3_2.Z adc_PISO_0.B1.n12 4.72925
R7299 adc_PISO_0.B1.n5 SARlogic_0.dffrs_10.nand3_6.B 2.17818
R7300 adc_PISO_0.B1 adc_PISO_0.B1.n2 1.87121
R7301 adc_PISO_0.B1.n5 SARlogic_0.dffrs_10.nand3_1.A 1.34729
R7302 adc_PISO_0.B1.n12 adc_PISO_0.B1.n11 0.732092
R7303 adc_PISO_0.B1.n10 adc_PISO_0.B1.t3 0.7285
R7304 adc_PISO_0.B1.n10 adc_PISO_0.B1.t2 0.7285
R7305 SARlogic_0.dffrs_10.clk adc_PISO_0.B1.n5 0.610571
R7306 SARlogic_0.dffrs_11.nand3_2.Z adc_PISO_0.B1.n9 0.166901
R7307 adc_PISO_0.B1.n1 adc_PISO_0.B1.n0 0.106438
R7308 adc_PISO_0.B1.n8 SARlogic_0.dffrs_11.nand3_7.C 0.0455
R7309 adc_PISO_0.B1.n2 adc_PISO_0.2inmux_1.In 0.0455
R7310 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t4 41.0041
R7311 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t5 40.8177
R7312 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t9 40.6313
R7313 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t8 27.3166
R7314 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t7 27.1302
R7315 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t6 26.9438
R7316 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.t1 10.0473
R7317 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n4 9.90747
R7318 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n2 9.90116
R7319 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.t2 6.51042
R7320 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.n7 6.04952
R7321 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_6.C.n1 5.7305
R7322 SARlogic_0.dffrs_10.nand3_2.B SARlogic_0.dffrs_10.nand3_6.C.n0 5.47979
R7323 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C.n3 5.13907
R7324 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n9 4.72925
R7325 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_6.C.n5 4.5005
R7326 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.n8 0.732092
R7327 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t3 0.7285
R7328 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t0 0.7285
R7329 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n6 0.449758
R7330 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_2.B 0.166901
R7331 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_0.A 0.0455
R7332 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C 0.0455
R7333 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t8 41.0041
R7334 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t5 40.6313
R7335 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t4 40.6313
R7336 SARlogic_0.dffrs_3.Qb SARlogic_0.dffrs_10.setb 28.021
R7337 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t7 27.3166
R7338 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t6 27.3166
R7339 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t9 26.9438
R7340 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.t2 10.0473
R7341 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb.n1 9.84255
R7342 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n3 9.22229
R7343 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.t3 6.51042
R7344 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.n7 6.04952
R7345 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.Qb.n0 5.7305
R7346 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n4 5.14711
R7347 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_3.Qb.n2 5.13907
R7348 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n6 4.94976
R7349 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n9 4.72925
R7350 SARlogic_0.dffrs_10.setb SARlogic_0.dffrs_10.nand3_0.C 0.784786
R7351 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.n8 0.732092
R7352 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t1 0.7285
R7353 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t0 0.7285
R7354 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb 0.175225
R7355 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.nand3_2.A 0.0455
R7356 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_10.nand3_2.C 0.0455
R7357 SARlogic_0.dffrs_10.nand3_0.C SARlogic_0.dffrs_3.Qb.n5 0.0374643
R7358 a_14313_33628.n0 a_14313_33628.t5 40.6313
R7359 a_14313_33628.n0 a_14313_33628.t4 27.3166
R7360 a_14313_33628.n1 a_14313_33628.n0 24.1527
R7361 a_14313_33628.n1 a_14313_33628.t2 10.0473
R7362 a_14313_33628.n2 a_14313_33628.t3 6.51042
R7363 a_14313_33628.n3 a_14313_33628.n2 6.04952
R7364 a_14313_33628.n2 a_14313_33628.n1 0.732092
R7365 a_14313_33628.t0 a_14313_33628.n3 0.7285
R7366 a_14313_33628.n3 a_14313_33628.t1 0.7285
R7367 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t8 41.0041
R7368 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t4 40.6313
R7369 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t5 40.6313
R7370 SARlogic_0.dffrs_5.Qb SARlogic_0.dffrs_12.setb 28.013
R7371 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t6 27.3166
R7372 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t7 27.3166
R7373 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t9 26.9438
R7374 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.t2 10.0473
R7375 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb.n1 9.84255
R7376 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n3 9.22229
R7377 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.t3 6.51042
R7378 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.n7 6.04952
R7379 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.Qb.n0 5.7305
R7380 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n4 5.14711
R7381 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_5.Qb.n2 5.13907
R7382 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n6 4.94976
R7383 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n9 4.72925
R7384 SARlogic_0.dffrs_12.setb SARlogic_0.dffrs_12.nand3_0.C 0.784786
R7385 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.n8 0.732092
R7386 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t1 0.7285
R7387 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t0 0.7285
R7388 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb 0.175225
R7389 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.nand3_2.A 0.0455
R7390 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_12.nand3_2.C 0.0455
R7391 SARlogic_0.dffrs_12.nand3_0.C SARlogic_0.dffrs_5.Qb.n5 0.0374643
R7392 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t4 40.6313
R7393 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.t8 34.1066
R7394 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t5 27.3166
R7395 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t6 19.673
R7396 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t7 19.4007
R7397 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n3 14.6967
R7398 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.t1 10.0473
R7399 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n6 9.39565
R7400 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.dffrs_1.Q.n1 6.70486
R7401 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.t0 6.51042
R7402 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.n4 6.04952
R7403 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n2 5.81354
R7404 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.n5 0.732092
R7405 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t2 0.7285
R7406 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t3 0.7285
R7407 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n7 0.458082
R7408 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.n0 0.252687
R7409 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.2inmux_3.Bit 0.0519286
R7410 adc_PISO_0.B6.n3 adc_PISO_0.B6.t4 40.6313
R7411 adc_PISO_0.B6.n1 adc_PISO_0.B6.t6 34.2529
R7412 adc_PISO_0.B6.n3 adc_PISO_0.B6.t8 27.3166
R7413 adc_PISO_0.B6.n5 adc_PISO_0.B6 23.5656
R7414 adc_PISO_0.B6.n0 adc_PISO_0.B6.t7 19.673
R7415 adc_PISO_0.B6.n0 adc_PISO_0.B6.t5 19.4007
R7416 adc_PISO_0.B6.n5 adc_PISO_0.B6.n4 14.0582
R7417 adc_PISO_0.B6.n8 adc_PISO_0.B6.t3 10.0473
R7418 adc_PISO_0.B6.n2 adc_PISO_0.B6.n1 8.05164
R7419 adc_PISO_0.B6.n7 adc_PISO_0.B6.t2 6.51042
R7420 adc_PISO_0.B6.n7 adc_PISO_0.B6.n6 6.04952
R7421 adc_PISO_0.B6.n4 adc_PISO_0.B6.n3 5.13907
R7422 SARlogic_0.dffrs_14.nand3_2.Z adc_PISO_0.B6.n8 4.72925
R7423 adc_PISO_0.B6 adc_PISO_0.B6.n2 1.87121
R7424 adc_PISO_0.B6.n8 adc_PISO_0.B6.n7 0.732092
R7425 adc_PISO_0.B6.n6 adc_PISO_0.B6.t0 0.7285
R7426 adc_PISO_0.B6.n6 adc_PISO_0.B6.t1 0.7285
R7427 SARlogic_0.dffrs_14.nand3_2.Z adc_PISO_0.B6.n5 0.166901
R7428 adc_PISO_0.B6.n1 adc_PISO_0.B6.n0 0.106438
R7429 adc_PISO_0.B6.n4 SARlogic_0.dffrs_14.nand3_7.C 0.0455
R7430 adc_PISO_0.B6.n2 adc_PISO_0.2inmux_0.In 0.0455
R7431 a_33257_29218.n2 a_33257_29218.t4 40.8177
R7432 a_33257_29218.n3 a_33257_29218.t7 40.6313
R7433 a_33257_29218.n3 a_33257_29218.t6 27.3166
R7434 a_33257_29218.n2 a_33257_29218.t5 27.1302
R7435 a_33257_29218.n4 a_33257_29218.n3 19.2576
R7436 a_33257_29218.t0 a_33257_29218.n5 10.0473
R7437 a_33257_29218.n1 a_33257_29218.t1 6.51042
R7438 a_33257_29218.n1 a_33257_29218.n0 6.04952
R7439 a_33257_29218.n4 a_33257_29218.n2 5.91752
R7440 a_33257_29218.n5 a_33257_29218.n4 4.89565
R7441 a_33257_29218.n5 a_33257_29218.n1 0.732092
R7442 a_33257_29218.n0 a_33257_29218.t3 0.7285
R7443 a_33257_29218.n0 a_33257_29218.t2 0.7285
R7444 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t5 41.0041
R7445 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t6 40.6313
R7446 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t4 40.6313
R7447 SARlogic_0.dffrs_0.Qb SARlogic_0.dffrs_7.setb 28.021
R7448 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t9 27.3166
R7449 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t7 27.3166
R7450 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t8 26.9438
R7451 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.t3 10.0473
R7452 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb.n1 9.84255
R7453 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n3 9.22229
R7454 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.t2 6.51042
R7455 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.n7 6.04952
R7456 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.Qb.n0 5.7305
R7457 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n4 5.14711
R7458 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_0.Qb.n2 5.13907
R7459 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n6 4.94976
R7460 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n9 4.72925
R7461 SARlogic_0.dffrs_7.setb SARlogic_0.dffrs_7.nand3_0.C 0.784786
R7462 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.n8 0.732092
R7463 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t0 0.7285
R7464 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t1 0.7285
R7465 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb 0.175225
R7466 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.nand3_2.A 0.0455
R7467 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_7.nand3_2.C 0.0455
R7468 SARlogic_0.dffrs_7.nand3_0.C SARlogic_0.dffrs_0.Qb.n5 0.0374643
R7469 a_9083_31160.n0 a_9083_31160.t5 34.1797
R7470 a_9083_31160.n0 a_9083_31160.t4 19.5798
R7471 a_9083_31160.n1 a_9083_31160.t1 18.7717
R7472 a_9083_31160.n1 a_9083_31160.t2 9.2885
R7473 a_9083_31160.n2 a_9083_31160.n0 4.93379
R7474 a_9083_31160.t0 a_9083_31160.n3 4.23346
R7475 a_9083_31160.n3 a_9083_31160.t3 3.85546
R7476 a_9083_31160.n2 a_9083_31160.n1 0.4055
R7477 a_9083_31160.n3 a_9083_31160.n2 0.352625
R7478 a_23785_29218.n0 a_23785_29218.t5 40.8177
R7479 a_23785_29218.n1 a_23785_29218.t4 40.6313
R7480 a_23785_29218.n1 a_23785_29218.t7 27.3166
R7481 a_23785_29218.n0 a_23785_29218.t6 27.1302
R7482 a_23785_29218.n2 a_23785_29218.n1 19.2576
R7483 a_23785_29218.n3 a_23785_29218.t3 10.0473
R7484 a_23785_29218.t0 a_23785_29218.n5 6.51042
R7485 a_23785_29218.n5 a_23785_29218.n4 6.04952
R7486 a_23785_29218.n2 a_23785_29218.n0 5.91752
R7487 a_23785_29218.n3 a_23785_29218.n2 4.89565
R7488 a_23785_29218.n5 a_23785_29218.n3 0.732092
R7489 a_23785_29218.n4 a_23785_29218.t1 0.7285
R7490 a_23785_29218.n4 a_23785_29218.t2 0.7285
R7491 a_23865_30170.n0 a_23865_30170.t7 41.0041
R7492 a_23865_30170.n1 a_23865_30170.t5 40.8177
R7493 a_23865_30170.n1 a_23865_30170.t6 27.1302
R7494 a_23865_30170.n0 a_23865_30170.t4 26.9438
R7495 a_23865_30170.n2 a_23865_30170.n1 22.5284
R7496 a_23865_30170.n3 a_23865_30170.n2 19.5781
R7497 a_23865_30170.n3 a_23865_30170.t1 10.0473
R7498 a_23865_30170.n4 a_23865_30170.t2 6.51042
R7499 a_23865_30170.n5 a_23865_30170.n4 6.04952
R7500 a_23865_30170.n2 a_23865_30170.n0 5.7305
R7501 a_23865_30170.n4 a_23865_30170.n3 0.732092
R7502 a_23865_30170.n5 a_23865_30170.t3 0.7285
R7503 a_23865_30170.t0 a_23865_30170.n5 0.7285
R7504 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t4 40.6313
R7505 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t5 27.3166
R7506 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n1 14.2854
R7507 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.t1 10.0473
R7508 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.t2 6.51042
R7509 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.n2 6.04952
R7510 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C.n0 5.13907
R7511 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n4 4.72925
R7512 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.n3 0.732092
R7513 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t0 0.7285
R7514 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t3 0.7285
R7515 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C 0.0455
R7516 a_42729_33628.n0 a_42729_33628.t4 40.6313
R7517 a_42729_33628.n0 a_42729_33628.t5 27.3166
R7518 a_42729_33628.n1 a_42729_33628.n0 24.1527
R7519 a_42729_33628.n1 a_42729_33628.t1 10.0473
R7520 a_42729_33628.t0 a_42729_33628.n3 6.51042
R7521 a_42729_33628.n3 a_42729_33628.n2 6.04952
R7522 a_42729_33628.n3 a_42729_33628.n1 0.732092
R7523 a_42729_33628.n2 a_42729_33628.t3 0.7285
R7524 a_42729_33628.n2 a_42729_33628.t2 0.7285
R7525 a_42729_31423.n3 a_42729_31423.t4 41.0041
R7526 a_42729_31423.n2 a_42729_31423.t5 40.8177
R7527 a_42729_31423.n4 a_42729_31423.t6 40.6313
R7528 a_42729_31423.n4 a_42729_31423.t9 27.3166
R7529 a_42729_31423.n2 a_42729_31423.t8 27.1302
R7530 a_42729_31423.n3 a_42729_31423.t7 26.9438
R7531 a_42729_31423.n5 a_42729_31423.n3 15.6312
R7532 a_42729_31423.n5 a_42729_31423.n4 15.046
R7533 a_42729_31423.t0 a_42729_31423.n7 10.0473
R7534 a_42729_31423.n1 a_42729_31423.t3 6.51042
R7535 a_42729_31423.n1 a_42729_31423.n0 6.04952
R7536 a_42729_31423.n6 a_42729_31423.n2 5.64619
R7537 a_42729_31423.n7 a_42729_31423.n6 5.17851
R7538 a_42729_31423.n6 a_42729_31423.n5 4.5005
R7539 a_42729_31423.n7 a_42729_31423.n1 0.732092
R7540 a_42729_31423.n0 a_42729_31423.t2 0.7285
R7541 a_42729_31423.n0 a_42729_31423.t1 0.7285
R7542 a_28027_31160.n0 a_28027_31160.t4 34.1797
R7543 a_28027_31160.n0 a_28027_31160.t5 19.5798
R7544 a_28027_31160.n1 a_28027_31160.t1 18.7717
R7545 a_28027_31160.n1 a_28027_31160.t2 9.2885
R7546 a_28027_31160.n2 a_28027_31160.n0 4.93379
R7547 a_28027_31160.t0 a_28027_31160.n3 4.23346
R7548 a_28027_31160.n3 a_28027_31160.t3 3.85546
R7549 a_28027_31160.n2 a_28027_31160.n1 0.4055
R7550 a_28027_31160.n3 a_28027_31160.n2 0.352625
R7551 a_23785_31423.n1 a_23785_31423.t5 41.0041
R7552 a_23785_31423.n0 a_23785_31423.t7 40.8177
R7553 a_23785_31423.n2 a_23785_31423.t4 40.6313
R7554 a_23785_31423.n2 a_23785_31423.t6 27.3166
R7555 a_23785_31423.n0 a_23785_31423.t9 27.1302
R7556 a_23785_31423.n1 a_23785_31423.t8 26.9438
R7557 a_23785_31423.n3 a_23785_31423.n1 15.6312
R7558 a_23785_31423.n3 a_23785_31423.n2 15.046
R7559 a_23785_31423.n5 a_23785_31423.t1 10.0473
R7560 a_23785_31423.t0 a_23785_31423.n7 6.51042
R7561 a_23785_31423.n7 a_23785_31423.n6 6.04952
R7562 a_23785_31423.n4 a_23785_31423.n0 5.64619
R7563 a_23785_31423.n5 a_23785_31423.n4 5.17851
R7564 a_23785_31423.n4 a_23785_31423.n3 4.5005
R7565 a_23785_31423.n7 a_23785_31423.n5 0.732092
R7566 a_23785_31423.n6 a_23785_31423.t2 0.7285
R7567 a_23785_31423.n6 a_23785_31423.t3 0.7285
R7568 Vin1.n7 Vin1.n6 23.1032
R7569 Vin1.n3 Vin1.n2 23.1032
R7570 Vin1.n0 Vin1.t8 22.5295
R7571 Vin1.n2 Vin1.t2 16.3641
R7572 Vin1.n6 Vin1.t6 16.3626
R7573 Vin1.n2 Vin1.t7 16.0225
R7574 Vin1.n6 Vin1.t1 16.021
R7575 Vin1.n8 Vin1.t4 11.5195
R7576 Vin1.n5 Vin1.t3 11.5195
R7577 Vin1.n4 Vin1.t9 11.5195
R7578 Vin1.n1 Vin1.t5 11.5195
R7579 Vin1.n0 Vin1.t0 11.5195
R7580 comparator_no_offsetcal_0.Vin1 Vin1 6.1115
R7581 Vin1.n1 Vin1.n0 4.00673
R7582 comparator_no_offsetcal_0.Vin1 Vin1.n8 3.5169
R7583 Vin1.n7 Vin1.n5 3.16619
R7584 Vin1.n3 Vin1.n1 0.650658
R7585 Vin1.n8 Vin1.n7 0.280193
R7586 Vin1.n4 Vin1.n3 0.279681
R7587 Vin1.n5 Vin1.n4 0.231705
R7588 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t14 19.5626
R7589 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 11.9065
R7590 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 11.2495
R7591 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 11.243
R7592 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 8.80104
R7593 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 6.60725
R7594 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 6.52262
R7595 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 6.386
R7596 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 5.44213
R7597 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 4.36738
R7598 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 4.36738
R7599 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 4.3505
R7600 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 2.2505
R7601 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 2.14009
R7602 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 1.50001
R7603 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 1.49326
R7604 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t8 1.0925
R7605 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t16 1.0925
R7606 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t6 1.0925
R7607 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t11 1.0925
R7608 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t13 1.0925
R7609 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t4 1.0925
R7610 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t10 1.0925
R7611 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t5 1.0925
R7612 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t12 1.0925
R7613 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t7 1.0925
R7614 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t3 1.0925
R7615 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t9 1.0925
R7616 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t1 0.8195
R7617 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t15 0.8195
R7618 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 0.8195
R7619 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t0 0.8195
R7620 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 0.314375
R7621 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 0.16025
R7622 a_n4631_31422.n3 a_n4631_31422.t9 41.0041
R7623 a_n4631_31422.n2 a_n4631_31422.t6 40.8177
R7624 a_n4631_31422.n4 a_n4631_31422.t5 40.6313
R7625 a_n4631_31422.n4 a_n4631_31422.t7 27.3166
R7626 a_n4631_31422.n2 a_n4631_31422.t8 27.1302
R7627 a_n4631_31422.n3 a_n4631_31422.t4 26.9438
R7628 a_n4631_31422.n5 a_n4631_31422.n3 15.6312
R7629 a_n4631_31422.n5 a_n4631_31422.n4 15.046
R7630 a_n4631_31422.t0 a_n4631_31422.n7 10.0473
R7631 a_n4631_31422.n1 a_n4631_31422.t3 6.51042
R7632 a_n4631_31422.n1 a_n4631_31422.n0 6.04952
R7633 a_n4631_31422.n6 a_n4631_31422.n2 5.64619
R7634 a_n4631_31422.n7 a_n4631_31422.n6 5.17851
R7635 a_n4631_31422.n6 a_n4631_31422.n5 4.5005
R7636 a_n4631_31422.n7 a_n4631_31422.n1 0.732092
R7637 a_n4631_31422.n0 a_n4631_31422.t2 0.7285
R7638 a_n4631_31422.n0 a_n4631_31422.t1 0.7285
R7639 a_n4631_33627.n0 a_n4631_33627.t4 40.6313
R7640 a_n4631_33627.n0 a_n4631_33627.t5 27.3166
R7641 a_n4631_33627.n1 a_n4631_33627.n0 24.1527
R7642 a_n4631_33627.n1 a_n4631_33627.t1 10.0473
R7643 a_n4631_33627.t0 a_n4631_33627.n3 6.51042
R7644 a_n4631_33627.n3 a_n4631_33627.n2 6.04952
R7645 a_n4631_33627.n3 a_n4631_33627.n1 0.732092
R7646 a_n4631_33627.n2 a_n4631_33627.t3 0.7285
R7647 a_n4631_33627.n2 a_n4631_33627.t2 0.7285
R7648 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t6 40.8177
R7649 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t7 40.6313
R7650 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t4 27.3166
R7651 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t5 27.1302
R7652 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_8.C.n2 14.119
R7653 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.t0 10.0473
R7654 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.t1 6.51042
R7655 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.n4 6.04952
R7656 SARlogic_0.dffrs_11.nand3_7.B SARlogic_0.dffrs_11.nand3_8.C.n0 5.47979
R7657 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C.n1 5.13907
R7658 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n6 4.72925
R7659 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.n5 0.732092
R7660 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t3 0.7285
R7661 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t2 0.7285
R7662 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_7.B 0.438233
R7663 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n3 0.166901
R7664 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C 0.0455
R7665 SAR_in.n9 SAR_in.t11 41.0041
R7666 SAR_in.n7 SAR_in.t6 41.0041
R7667 SAR_in.n5 SAR_in.t2 41.0041
R7668 SAR_in.n3 SAR_in.t8 41.0041
R7669 SAR_in.n1 SAR_in.t1 41.0041
R7670 SAR_in.n0 SAR_in.t7 41.0041
R7671 SAR_in.n9 SAR_in.t3 26.9438
R7672 SAR_in.n7 SAR_in.t9 26.9438
R7673 SAR_in.n5 SAR_in.t5 26.9438
R7674 SAR_in.n3 SAR_in.t0 26.9438
R7675 SAR_in.n1 SAR_in.t4 26.9438
R7676 SAR_in.n0 SAR_in.t10 26.9438
R7677 SAR_in.n2 SARlogic_0.dffrs_11.d 15.3544
R7678 SAR_in.n8 SARlogic_0.dffrs_7.d 11.7166
R7679 SAR_in.n6 SARlogic_0.dffrs_8.d 11.7166
R7680 SAR_in.n4 SARlogic_0.dffrs_9.d 11.7166
R7681 SAR_in.n2 SARlogic_0.dffrs_10.d 11.7166
R7682 SAR_in.n10 SARlogic_0.dffrs_14.d 11.6732
R7683 SARlogic_0.comp_in SAR_in.n10 7.63655
R7684 SARlogic_0.dffrs_14.nand3_8.A SAR_in.n9 5.7755
R7685 SARlogic_0.dffrs_7.nand3_8.A SAR_in.n7 5.7755
R7686 SARlogic_0.dffrs_8.nand3_8.A SAR_in.n5 5.7755
R7687 SARlogic_0.dffrs_9.nand3_8.A SAR_in.n3 5.7755
R7688 SARlogic_0.dffrs_10.nand3_8.A SAR_in.n1 5.7755
R7689 SARlogic_0.dffrs_11.nand3_8.A SAR_in.n0 5.7755
R7690 SAR_in.n4 SAR_in.n2 3.6383
R7691 SAR_in.n6 SAR_in.n4 3.6383
R7692 SAR_in.n8 SAR_in.n6 3.6383
R7693 SAR_in.n10 SAR_in.n8 3.6113
R7694 SARlogic_0.dffrs_14.d SARlogic_0.dffrs_14.nand3_8.A 0.784786
R7695 SARlogic_0.dffrs_7.d SARlogic_0.dffrs_7.nand3_8.A 0.784786
R7696 SARlogic_0.dffrs_8.d SARlogic_0.dffrs_8.nand3_8.A 0.784786
R7697 SARlogic_0.dffrs_9.d SARlogic_0.dffrs_9.nand3_8.A 0.784786
R7698 SARlogic_0.dffrs_10.d SARlogic_0.dffrs_10.nand3_8.A 0.784786
R7699 SARlogic_0.dffrs_11.d SARlogic_0.dffrs_11.nand3_8.A 0.784786
R7700 SARlogic_0.comp_in SAR_in 0.1775
R7701 a_n9861_31159.n0 a_n9861_31159.t4 34.1797
R7702 a_n9861_31159.n0 a_n9861_31159.t5 19.5798
R7703 a_n9861_31159.n1 a_n9861_31159.t1 18.7717
R7704 a_n9861_31159.n1 a_n9861_31159.t2 9.2885
R7705 a_n9861_31159.n2 a_n9861_31159.n0 4.93379
R7706 a_n9861_31159.t0 a_n9861_31159.n3 4.23346
R7707 a_n9861_31159.n3 a_n9861_31159.t3 3.85546
R7708 a_n9861_31159.n2 a_n9861_31159.n1 0.4055
R7709 a_n9861_31159.n3 a_n9861_31159.n2 0.352625
R7710 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t6 40.8177
R7711 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t7 40.6313
R7712 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t5 27.3166
R7713 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t4 27.1302
R7714 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_8.C.n2 14.119
R7715 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.t3 10.0473
R7716 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.t2 6.51042
R7717 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.n4 6.04952
R7718 SARlogic_0.dffrs_14.nand3_7.B SARlogic_0.dffrs_14.nand3_8.C.n0 5.47979
R7719 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C.n1 5.13907
R7720 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n6 4.72925
R7721 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.n5 0.732092
R7722 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t0 0.7285
R7723 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t1 0.7285
R7724 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_7.B 0.438233
R7725 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n3 0.166901
R7726 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C 0.0455
R7727 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t6 41.0041
R7728 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t7 40.8177
R7729 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t4 27.1302
R7730 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t5 26.9438
R7731 SARlogic_0.dffrs_13.nand3_6.A SARlogic_0.dffrs_13.nand3_0.B 17.0041
R7732 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n2 14.8493
R7733 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.t0 10.0473
R7734 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.t1 6.51042
R7735 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.n3 6.04952
R7736 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_8.Z.n0 5.7305
R7737 SARlogic_0.dffrs_13.nand3_0.B SARlogic_0.dffrs_13.nand3_8.Z.n1 5.47979
R7738 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n5 4.72925
R7739 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.n4 0.732092
R7740 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t3 0.7285
R7741 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t2 0.7285
R7742 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_6.A 0.0455
R7743 a_n389_31159.n0 a_n389_31159.t4 34.1797
R7744 a_n389_31159.n0 a_n389_31159.t5 19.5798
R7745 a_n389_31159.n1 a_n389_31159.t2 18.7717
R7746 a_n389_31159.n1 a_n389_31159.t1 9.2885
R7747 a_n389_31159.n2 a_n389_31159.n0 4.93379
R7748 a_n389_31159.t0 a_n389_31159.n3 4.23346
R7749 a_n389_31159.n3 a_n389_31159.t3 3.85546
R7750 a_n389_31159.n2 a_n389_31159.n1 0.4055
R7751 a_n389_31159.n3 a_n389_31159.n2 0.352625
R7752 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t5 40.8177
R7753 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t7 40.6313
R7754 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t4 27.3166
R7755 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t6 27.1302
R7756 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_8.C.n2 14.119
R7757 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.t2 10.0473
R7758 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.t3 6.51042
R7759 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.n4 6.04952
R7760 SARlogic_0.dffrs_9.nand3_7.B SARlogic_0.dffrs_9.nand3_8.C.n0 5.47979
R7761 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C.n1 5.13907
R7762 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n6 4.72925
R7763 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.n5 0.732092
R7764 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t1 0.7285
R7765 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t0 0.7285
R7766 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_7.B 0.438233
R7767 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n3 0.166901
R7768 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C 0.0455
R7769 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t6 41.0041
R7770 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t7 40.8177
R7771 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t4 40.6313
R7772 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t5 27.3166
R7773 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t8 27.1302
R7774 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t9 26.9438
R7775 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.t2 10.0473
R7776 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n4 9.90747
R7777 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n2 9.90116
R7778 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.t1 6.51042
R7779 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.n7 6.04952
R7780 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_6.C.n1 5.7305
R7781 SARlogic_0.dffrs_0.nand3_2.B SARlogic_0.dffrs_0.nand3_6.C.n0 5.47979
R7782 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C.n3 5.13907
R7783 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n9 4.72925
R7784 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_6.C.n5 4.5005
R7785 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.n8 0.732092
R7786 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t3 0.7285
R7787 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t0 0.7285
R7788 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n6 0.449758
R7789 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_2.B 0.166901
R7790 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_0.A 0.0455
R7791 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C 0.0455
R7792 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t6 40.8177
R7793 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t5 40.6313
R7794 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t7 27.3166
R7795 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t4 27.1302
R7796 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_8.C.n2 14.119
R7797 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.t1 10.0473
R7798 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.t3 6.51042
R7799 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.n4 6.04952
R7800 SARlogic_0.dffrs_0.nand3_7.B SARlogic_0.dffrs_0.nand3_8.C.n0 5.47979
R7801 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C.n1 5.13907
R7802 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n6 4.72925
R7803 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.n5 0.732092
R7804 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t2 0.7285
R7805 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t0 0.7285
R7806 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_7.B 0.438233
R7807 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n3 0.166901
R7808 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C 0.0455
R7809 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t7 41.0041
R7810 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t6 40.8177
R7811 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t5 40.6313
R7812 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t4 27.3166
R7813 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t8 27.1302
R7814 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t9 26.9438
R7815 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.t1 10.0473
R7816 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n4 9.90747
R7817 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n2 9.90116
R7818 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.t3 6.51042
R7819 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.n7 6.04952
R7820 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_6.C.n1 5.7305
R7821 SARlogic_0.dffrs_11.nand3_2.B SARlogic_0.dffrs_11.nand3_6.C.n0 5.47979
R7822 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C.n3 5.13907
R7823 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n9 4.72925
R7824 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_6.C.n5 4.5005
R7825 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.n8 0.732092
R7826 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t2 0.7285
R7827 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t0 0.7285
R7828 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n6 0.449758
R7829 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_2.B 0.166901
R7830 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_0.A 0.0455
R7831 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C 0.0455
R7832 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t4 41.0041
R7833 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t5 40.8177
R7834 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t9 40.6313
R7835 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t8 27.3166
R7836 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t7 27.1302
R7837 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t6 26.9438
R7838 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.t3 10.0473
R7839 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n4 9.90747
R7840 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n2 9.90116
R7841 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.t2 6.51042
R7842 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.n7 6.04952
R7843 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_6.C.n1 5.7305
R7844 SARlogic_0.dffrs_8.nand3_2.B SARlogic_0.dffrs_8.nand3_6.C.n0 5.47979
R7845 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C.n3 5.13907
R7846 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n9 4.72925
R7847 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_6.C.n5 4.5005
R7848 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.n8 0.732092
R7849 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t1 0.7285
R7850 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t0 0.7285
R7851 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n6 0.449758
R7852 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_2.B 0.166901
R7853 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_0.A 0.0455
R7854 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C 0.0455
R7855 a_n389_28819.n0 a_n389_28819.t5 34.1797
R7856 a_n389_28819.n0 a_n389_28819.t4 19.5798
R7857 a_n389_28819.n1 a_n389_28819.t1 18.7717
R7858 a_n389_28819.n1 a_n389_28819.t2 9.2885
R7859 a_n389_28819.n2 a_n389_28819.n0 4.93379
R7860 a_n389_28819.t0 a_n389_28819.n3 4.23346
R7861 a_n389_28819.n3 a_n389_28819.t3 3.85546
R7862 a_n389_28819.n2 a_n389_28819.n1 0.4055
R7863 a_n389_28819.n3 a_n389_28819.n2 0.352625
R7864 a_1839_29263.n0 a_1839_29263.t5 34.1797
R7865 a_1839_29263.n0 a_1839_29263.t4 19.5798
R7866 a_1839_29263.n1 a_1839_29263.t3 10.3401
R7867 a_1839_29263.n1 a_1839_29263.t2 9.2885
R7868 a_1839_29263.n2 a_1839_29263.n0 4.93379
R7869 a_1839_29263.n3 a_1839_29263.t0 4.09202
R7870 a_1839_29263.t1 a_1839_29263.n3 3.95079
R7871 a_1839_29263.n2 a_1839_29263.n1 0.599711
R7872 a_1839_29263.n3 a_1839_29263.n2 0.296375
R7873 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t4 40.6313
R7874 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t5 27.3166
R7875 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n1 14.2854
R7876 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.t1 10.0473
R7877 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.t0 6.51042
R7878 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.n2 6.04952
R7879 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C.n0 5.13907
R7880 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n4 4.72925
R7881 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.n3 0.732092
R7882 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t3 0.7285
R7883 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t2 0.7285
R7884 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C 0.0455
R7885 a_20783_29264.n0 a_20783_29264.t5 34.1797
R7886 a_20783_29264.n0 a_20783_29264.t4 19.5798
R7887 a_20783_29264.t0 a_20783_29264.n3 10.3401
R7888 a_20783_29264.n3 a_20783_29264.t3 9.2885
R7889 a_20783_29264.n2 a_20783_29264.n0 4.93379
R7890 a_20783_29264.n1 a_20783_29264.t2 4.09202
R7891 a_20783_29264.n1 a_20783_29264.t1 3.95079
R7892 a_20783_29264.n3 a_20783_29264.n2 0.599711
R7893 a_20783_29264.n2 a_20783_29264.n1 0.296375
R7894 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t8 40.6313
R7895 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.t6 34.1066
R7896 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t4 27.3166
R7897 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t7 19.673
R7898 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t5 19.4007
R7899 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n3 14.6967
R7900 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.t1 10.0473
R7901 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n6 9.39565
R7902 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit.n1 6.70486
R7903 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.t2 6.51042
R7904 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.n4 6.04952
R7905 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n2 5.81514
R7906 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.n5 0.732092
R7907 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t0 0.7285
R7908 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t3 0.7285
R7909 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n7 0.458082
R7910 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.n0 0.252687
R7911 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit 0.0519286
R7912 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_11.clk 44.4671
R7913 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t7 41.0041
R7914 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t6 40.8177
R7915 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t8 40.6313
R7916 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t5 27.3166
R7917 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t4 27.1302
R7918 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t9 26.9438
R7919 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_12.Q.n4 14.0582
R7920 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.t1 10.0473
R7921 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.t2 6.51042
R7922 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.n6 6.04952
R7923 SARlogic_0.dffrs_11.nand3_1.A SARlogic_0.dffrs_12.Q.n0 5.7755
R7924 SARlogic_0.dffrs_11.nand3_6.B SARlogic_0.dffrs_12.Q.n1 5.47979
R7925 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.Q.n3 5.13907
R7926 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n8 4.72925
R7927 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_6.B 2.17818
R7928 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_1.A 1.34729
R7929 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.n7 0.732092
R7930 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t3 0.7285
R7931 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t0 0.7285
R7932 SARlogic_0.dffrs_11.clk SARlogic_0.dffrs_12.Q.n2 0.610571
R7933 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n5 0.166901
R7934 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.nand3_7.C 0.0455
R7935 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t3 41.0041
R7936 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t2 26.9438
R7937 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t0 9.6935
R7938 adc_PISO_0.dffrs_1.d adc_PISO_0.2inmux_2.OUT.n0 6.55979
R7939 adc_PISO_0.2inmux_2.OUT adc_PISO_0.dffrs_1.d 4.883
R7940 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t1 4.35383
R7941 adc_PISO_0.2inmux_2.OUT adc_PISO_0.2inmux_2.OUT.n1 0.350857
R7942 a_4921_30169.n0 a_4921_30169.t5 41.0041
R7943 a_4921_30169.n1 a_4921_30169.t6 40.8177
R7944 a_4921_30169.n1 a_4921_30169.t4 27.1302
R7945 a_4921_30169.n0 a_4921_30169.t7 26.9438
R7946 a_4921_30169.n2 a_4921_30169.n1 22.5284
R7947 a_4921_30169.n3 a_4921_30169.n2 19.5781
R7948 a_4921_30169.n3 a_4921_30169.t1 10.0473
R7949 a_4921_30169.t0 a_4921_30169.n5 6.51042
R7950 a_4921_30169.n5 a_4921_30169.n4 6.04952
R7951 a_4921_30169.n2 a_4921_30169.n0 5.7305
R7952 a_4921_30169.n5 a_4921_30169.n3 0.732092
R7953 a_4921_30169.n4 a_4921_30169.t3 0.7285
R7954 a_4921_30169.n4 a_4921_30169.t2 0.7285
R7955 a_n4631_29217.n0 a_n4631_29217.t6 40.8177
R7956 a_n4631_29217.n1 a_n4631_29217.t5 40.6313
R7957 a_n4631_29217.n1 a_n4631_29217.t7 27.3166
R7958 a_n4631_29217.n0 a_n4631_29217.t4 27.1302
R7959 a_n4631_29217.n2 a_n4631_29217.n1 19.2576
R7960 a_n4631_29217.n3 a_n4631_29217.t3 10.0473
R7961 a_n4631_29217.n4 a_n4631_29217.t2 6.51042
R7962 a_n4631_29217.n5 a_n4631_29217.n4 6.04952
R7963 a_n4631_29217.n2 a_n4631_29217.n0 5.91752
R7964 a_n4631_29217.n3 a_n4631_29217.n2 4.89565
R7965 a_n4631_29217.n4 a_n4631_29217.n3 0.732092
R7966 a_n4631_29217.n5 a_n4631_29217.t1 0.7285
R7967 a_n4631_29217.t0 a_n4631_29217.n5 0.7285
R7968 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t6 41.0041
R7969 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t5 40.8177
R7970 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t4 40.6313
R7971 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t9 27.3166
R7972 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t7 27.1302
R7973 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t8 26.9438
R7974 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.t1 10.0473
R7975 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n4 9.90747
R7976 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n2 9.90116
R7977 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.t0 6.51042
R7978 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.n7 6.04952
R7979 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_6.C.n1 5.7305
R7980 SARlogic_0.dffrs_7.nand3_2.B SARlogic_0.dffrs_7.nand3_6.C.n0 5.47979
R7981 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C.n3 5.13907
R7982 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n9 4.72925
R7983 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_6.C.n5 4.5005
R7984 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.n8 0.732092
R7985 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t3 0.7285
R7986 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t2 0.7285
R7987 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n6 0.449758
R7988 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_2.B 0.166901
R7989 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_0.A 0.0455
R7990 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C 0.0455
R7991 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t2 41.0041
R7992 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t3 26.9438
R7993 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t0 9.6935
R7994 adc_PISO_0.dffrs_2.d adc_PISO_0.2inmux_3.OUT.n0 6.55979
R7995 adc_PISO_0.2inmux_3.OUT adc_PISO_0.dffrs_2.d 4.883
R7996 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t1 4.35383
R7997 adc_PISO_0.2inmux_3.OUT adc_PISO_0.2inmux_3.OUT.n1 0.350857
R7998 a_14393_30170.n0 a_14393_30170.t4 41.0041
R7999 a_14393_30170.n1 a_14393_30170.t6 40.8177
R8000 a_14393_30170.n1 a_14393_30170.t7 27.1302
R8001 a_14393_30170.n0 a_14393_30170.t5 26.9438
R8002 a_14393_30170.n2 a_14393_30170.n1 22.5284
R8003 a_14393_30170.n3 a_14393_30170.n2 19.5781
R8004 a_14393_30170.n3 a_14393_30170.t1 10.0473
R8005 a_14393_30170.t0 a_14393_30170.n5 6.51042
R8006 a_14393_30170.n5 a_14393_30170.n4 6.04952
R8007 a_14393_30170.n2 a_14393_30170.n0 5.7305
R8008 a_14393_30170.n5 a_14393_30170.n3 0.732092
R8009 a_14393_30170.n4 a_14393_30170.t2 0.7285
R8010 a_14393_30170.n4 a_14393_30170.t3 0.7285
R8011 Vin2.n7 Vin2.n6 23.1032
R8012 Vin2.n3 Vin2.n2 23.1032
R8013 Vin2.n0 Vin2.t6 22.8502
R8014 Vin2.n2 Vin2.t5 16.3656
R8015 Vin2.n6 Vin2.t1 16.3641
R8016 Vin2.n2 Vin2.t2 16.021
R8017 Vin2.n6 Vin2.t4 16.0195
R8018 Vin2.n8 Vin2.t8 11.5195
R8019 Vin2.n5 Vin2.t7 11.5195
R8020 Vin2.n4 Vin2.t0 11.5195
R8021 Vin2.n1 Vin2.t9 11.5195
R8022 Vin2.n0 Vin2.t3 11.5195
R8023 comparator_no_offsetcal_0.Vin2 Vin2 6.1091
R8024 comparator_no_offsetcal_0.Vin2 Vin2.n8 3.51835
R8025 Vin2.n7 Vin2.n5 2.53166
R8026 Vin2.n1 Vin2.n0 2.48408
R8027 Vin2.n3 Vin2.n1 1.40666
R8028 Vin2.n8 Vin2.n7 0.647658
R8029 Vin2.n4 Vin2.n3 0.647132
R8030 Vin2.n5 Vin2.n4 0.234605
R8031 Clk_piso.n19 Clk_piso.t9 41.0041
R8032 Clk_piso.n15 Clk_piso.t16 41.0041
R8033 Clk_piso.n11 Clk_piso.t6 41.0041
R8034 Clk_piso.n7 Clk_piso.t2 41.0041
R8035 Clk_piso.n3 Clk_piso.t0 41.0041
R8036 Clk_piso.n0 Clk_piso.t10 41.0041
R8037 Clk_piso.n20 Clk_piso.t13 40.8177
R8038 Clk_piso.n16 Clk_piso.t11 40.8177
R8039 Clk_piso.n12 Clk_piso.t3 40.8177
R8040 Clk_piso.n8 Clk_piso.t1 40.8177
R8041 Clk_piso.n4 Clk_piso.t15 40.8177
R8042 Clk_piso.n1 Clk_piso.t12 40.8177
R8043 Clk_piso.n20 Clk_piso.t21 27.1302
R8044 Clk_piso.n16 Clk_piso.t19 27.1302
R8045 Clk_piso.n12 Clk_piso.t8 27.1302
R8046 Clk_piso.n8 Clk_piso.t5 27.1302
R8047 Clk_piso.n4 Clk_piso.t22 27.1302
R8048 Clk_piso.n1 Clk_piso.t20 27.1302
R8049 Clk_piso.n19 Clk_piso.t17 26.9438
R8050 Clk_piso.n15 Clk_piso.t23 26.9438
R8051 Clk_piso.n11 Clk_piso.t14 26.9438
R8052 Clk_piso.n7 Clk_piso.t7 26.9438
R8053 Clk_piso.n3 Clk_piso.t4 26.9438
R8054 Clk_piso.n0 Clk_piso.t18 26.9438
R8055 Clk_piso.n6 adc_PISO_0.dffrs_5.clk 23.2034
R8056 Clk_piso.n22 Clk_piso.n18 13.9468
R8057 Clk_piso.n18 Clk_piso.n14 13.9463
R8058 Clk_piso.n10 Clk_piso.n6 13.9457
R8059 Clk_piso.n14 Clk_piso.n10 13.9457
R8060 Clk_piso.n23 Clk_piso 13.1341
R8061 Clk_piso.n22 adc_PISO_0.dffrs_0.clk 9.25764
R8062 Clk_piso.n18 adc_PISO_0.dffrs_1.clk 9.25764
R8063 Clk_piso.n14 adc_PISO_0.dffrs_2.clk 9.25764
R8064 Clk_piso.n10 adc_PISO_0.dffrs_3.clk 9.25764
R8065 Clk_piso.n6 adc_PISO_0.dffrs_4.clk 9.25764
R8066 Clk_piso.n21 Clk_piso.n20 7.65746
R8067 Clk_piso.n17 Clk_piso.n16 7.65746
R8068 Clk_piso.n13 Clk_piso.n12 7.65746
R8069 Clk_piso.n9 Clk_piso.n8 7.65746
R8070 Clk_piso.n5 Clk_piso.n4 7.65746
R8071 Clk_piso.n2 Clk_piso.n1 7.65746
R8072 Clk_piso.n21 Clk_piso.n19 7.12229
R8073 Clk_piso.n17 Clk_piso.n15 7.12229
R8074 Clk_piso.n13 Clk_piso.n11 7.12229
R8075 Clk_piso.n9 Clk_piso.n7 7.12229
R8076 Clk_piso.n5 Clk_piso.n3 7.12229
R8077 Clk_piso.n2 Clk_piso.n0 7.12229
R8078 Clk_piso.n23 Clk_piso.n22 3.49505
R8079 adc_PISO_0.dffrs_0.clk Clk_piso.n21 0.611214
R8080 adc_PISO_0.dffrs_1.clk Clk_piso.n17 0.611214
R8081 adc_PISO_0.dffrs_2.clk Clk_piso.n13 0.611214
R8082 adc_PISO_0.dffrs_3.clk Clk_piso.n9 0.611214
R8083 adc_PISO_0.dffrs_4.clk Clk_piso.n5 0.611214
R8084 adc_PISO_0.dffrs_5.clk Clk_piso.n2 0.611214
R8085 adc_PISO_0.clk Clk_piso.n23 0.0336579
R8086 a_14313_29218.n0 a_14313_29218.t6 40.8177
R8087 a_14313_29218.n1 a_14313_29218.t5 40.6313
R8088 a_14313_29218.n1 a_14313_29218.t4 27.3166
R8089 a_14313_29218.n0 a_14313_29218.t7 27.1302
R8090 a_14313_29218.n2 a_14313_29218.n1 19.2576
R8091 a_14313_29218.n3 a_14313_29218.t1 10.0473
R8092 a_14313_29218.n4 a_14313_29218.t2 6.51042
R8093 a_14313_29218.n5 a_14313_29218.n4 6.04952
R8094 a_14313_29218.n2 a_14313_29218.n0 5.91752
R8095 a_14313_29218.n3 a_14313_29218.n2 4.89565
R8096 a_14313_29218.n4 a_14313_29218.n3 0.732092
R8097 a_14313_29218.t0 a_14313_29218.n5 0.7285
R8098 a_14313_29218.n5 a_14313_29218.t3 0.7285
R8099 a_4841_29217.n0 a_4841_29217.t6 40.8177
R8100 a_4841_29217.n1 a_4841_29217.t5 40.6313
R8101 a_4841_29217.n1 a_4841_29217.t7 27.3166
R8102 a_4841_29217.n0 a_4841_29217.t4 27.1302
R8103 a_4841_29217.n2 a_4841_29217.n1 19.2576
R8104 a_4841_29217.n3 a_4841_29217.t3 10.0473
R8105 a_4841_29217.n4 a_4841_29217.t2 6.51042
R8106 a_4841_29217.n5 a_4841_29217.n4 6.04952
R8107 a_4841_29217.n2 a_4841_29217.n0 5.91752
R8108 a_4841_29217.n3 a_4841_29217.n2 4.89565
R8109 a_4841_29217.n4 a_4841_29217.n3 0.732092
R8110 a_4841_29217.t0 a_4841_29217.n5 0.7285
R8111 a_4841_29217.n5 a_4841_29217.t1 0.7285
R8112 adc_PISO_0.B5.n3 adc_PISO_0.B5.t11 41.0041
R8113 adc_PISO_0.B5.n4 adc_PISO_0.B5.t12 40.8177
R8114 adc_PISO_0.B5.n7 adc_PISO_0.B5.t7 40.6313
R8115 adc_PISO_0.B5.n1 adc_PISO_0.B5.t10 34.2529
R8116 adc_PISO_0.B5.n6 SARlogic_0.dffrs_14.clk 33.675
R8117 adc_PISO_0.B5.n7 adc_PISO_0.B5.t5 27.3166
R8118 adc_PISO_0.B5.n4 adc_PISO_0.B5.t8 27.1302
R8119 adc_PISO_0.B5.n3 adc_PISO_0.B5.t4 26.9438
R8120 adc_PISO_0.B5.n0 adc_PISO_0.B5.t6 19.673
R8121 adc_PISO_0.B5.n0 adc_PISO_0.B5.t9 19.4007
R8122 adc_PISO_0.B5.n9 adc_PISO_0.B5.n8 14.0582
R8123 adc_PISO_0.B5.n9 adc_PISO_0.B5.n6 11.3593
R8124 adc_PISO_0.B5.n12 adc_PISO_0.B5.t3 10.0473
R8125 adc_PISO_0.B5.n2 adc_PISO_0.B5.n1 8.05164
R8126 adc_PISO_0.B5.n11 adc_PISO_0.B5.t2 6.51042
R8127 adc_PISO_0.B5.n11 adc_PISO_0.B5.n10 6.04952
R8128 SARlogic_0.dffrs_14.nand3_1.A adc_PISO_0.B5.n3 5.7755
R8129 SARlogic_0.dffrs_14.nand3_6.B adc_PISO_0.B5.n4 5.47979
R8130 adc_PISO_0.B5.n8 adc_PISO_0.B5.n7 5.13907
R8131 SARlogic_0.dffrs_7.nand3_2.Z adc_PISO_0.B5.n12 4.72925
R8132 adc_PISO_0.B5.n6 adc_PISO_0.B5 3.49604
R8133 adc_PISO_0.B5.n5 SARlogic_0.dffrs_14.nand3_6.B 2.17818
R8134 adc_PISO_0.B5 adc_PISO_0.B5.n2 1.87121
R8135 adc_PISO_0.B5.n5 SARlogic_0.dffrs_14.nand3_1.A 1.34729
R8136 adc_PISO_0.B5.n12 adc_PISO_0.B5.n11 0.732092
R8137 adc_PISO_0.B5.n10 adc_PISO_0.B5.t1 0.7285
R8138 adc_PISO_0.B5.n10 adc_PISO_0.B5.t0 0.7285
R8139 SARlogic_0.dffrs_14.clk adc_PISO_0.B5.n5 0.611214
R8140 SARlogic_0.dffrs_7.nand3_2.Z adc_PISO_0.B5.n9 0.166901
R8141 adc_PISO_0.B5.n1 adc_PISO_0.B5.n0 0.106438
R8142 adc_PISO_0.B5.n8 SARlogic_0.dffrs_7.nand3_7.C 0.0455
R8143 adc_PISO_0.B5.n2 adc_PISO_0.2inmux_2.In 0.0455
R8144 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t5 41.0041
R8145 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t7 40.6313
R8146 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t8 40.6313
R8147 SARlogic_0.dffrs_4.Qb SARlogic_0.dffrs_11.setb 28.021
R8148 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t9 27.3166
R8149 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t4 27.3166
R8150 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t6 26.9438
R8151 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.t3 10.0473
R8152 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb.n1 9.84255
R8153 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n3 9.22229
R8154 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.t2 6.51042
R8155 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.n7 6.04952
R8156 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.Qb.n0 5.7305
R8157 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n4 5.14711
R8158 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_4.Qb.n2 5.13907
R8159 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n6 4.94976
R8160 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n9 4.72925
R8161 SARlogic_0.dffrs_11.setb SARlogic_0.dffrs_11.nand3_0.C 0.784786
R8162 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.n8 0.732092
R8163 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t0 0.7285
R8164 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t1 0.7285
R8165 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb 0.175225
R8166 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.nand3_2.A 0.0455
R8167 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_11.nand3_2.C 0.0455
R8168 SARlogic_0.dffrs_11.nand3_0.C SARlogic_0.dffrs_4.Qb.n5 0.0374643
R8169 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t6 40.8177
R8170 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t5 40.6313
R8171 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t7 27.3166
R8172 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t4 27.1302
R8173 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_8.C.n2 14.119
R8174 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.t0 10.0473
R8175 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.t1 6.51042
R8176 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.n4 6.04952
R8177 SARlogic_0.dffrs_8.nand3_7.B SARlogic_0.dffrs_8.nand3_8.C.n0 5.47979
R8178 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C.n1 5.13907
R8179 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n6 4.72925
R8180 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.n5 0.732092
R8181 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t3 0.7285
R8182 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t2 0.7285
R8183 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_7.B 0.438233
R8184 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n3 0.166901
R8185 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C 0.0455
R8186 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t5 41.0041
R8187 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t6 40.8177
R8188 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t4 27.1302
R8189 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t7 26.9438
R8190 SARlogic_0.dffrs_2.nand3_6.A SARlogic_0.dffrs_2.nand3_0.B 17.0041
R8191 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n2 14.8493
R8192 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.t2 10.0473
R8193 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.t1 6.51042
R8194 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.n3 6.04952
R8195 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_8.Z.n0 5.7305
R8196 SARlogic_0.dffrs_2.nand3_0.B SARlogic_0.dffrs_2.nand3_8.Z.n1 5.47979
R8197 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n5 4.72925
R8198 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.n4 0.732092
R8199 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t3 0.7285
R8200 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t0 0.7285
R8201 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_6.A 0.0455
R8202 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t5 40.6313
R8203 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.t6 34.1066
R8204 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t7 27.3166
R8205 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t8 19.673
R8206 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t4 19.4007
R8207 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n3 14.6967
R8208 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.t1 10.0473
R8209 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n6 9.39565
R8210 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.dffrs_3.Q.n1 6.70486
R8211 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.t2 6.51042
R8212 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.n4 6.04952
R8213 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n2 5.81514
R8214 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.n5 0.732092
R8215 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t0 0.7285
R8216 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t3 0.7285
R8217 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n7 0.458082
R8218 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.n0 0.252687
R8219 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.2inmux_5.Bit 0.0519286
R8220 a_39727_29264.n0 a_39727_29264.t5 34.1797
R8221 a_39727_29264.n0 a_39727_29264.t4 19.5798
R8222 a_39727_29264.n3 a_39727_29264.t3 10.3401
R8223 a_39727_29264.t0 a_39727_29264.n3 9.2885
R8224 a_39727_29264.n2 a_39727_29264.n0 4.93379
R8225 a_39727_29264.n1 a_39727_29264.t1 4.09202
R8226 a_39727_29264.n1 a_39727_29264.t2 3.95079
R8227 a_39727_29264.n3 a_39727_29264.n2 0.599711
R8228 a_39727_29264.n2 a_39727_29264.n1 0.296375
R8229 a_42809_30170.n0 a_42809_30170.t5 41.0041
R8230 a_42809_30170.n1 a_42809_30170.t7 40.8177
R8231 a_42809_30170.n1 a_42809_30170.t4 27.1302
R8232 a_42809_30170.n0 a_42809_30170.t6 26.9438
R8233 a_42809_30170.n2 a_42809_30170.n1 22.5284
R8234 a_42809_30170.n3 a_42809_30170.n2 19.5781
R8235 a_42809_30170.n3 a_42809_30170.t2 10.0473
R8236 a_42809_30170.n4 a_42809_30170.t1 6.51042
R8237 a_42809_30170.n5 a_42809_30170.n4 6.04952
R8238 a_42809_30170.n2 a_42809_30170.n0 5.7305
R8239 a_42809_30170.n4 a_42809_30170.n3 0.732092
R8240 a_42809_30170.n5 a_42809_30170.t3 0.7285
R8241 a_42809_30170.t0 a_42809_30170.n5 0.7285
R8242 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t7 40.8177
R8243 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t5 40.6313
R8244 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t6 27.3166
R8245 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t4 27.1302
R8246 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_8.C.n2 14.119
R8247 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.t1 10.0473
R8248 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.t2 6.51042
R8249 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.n4 6.04952
R8250 SARlogic_0.dffrs_10.nand3_7.B SARlogic_0.dffrs_10.nand3_8.C.n0 5.47979
R8251 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C.n1 5.13907
R8252 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n6 4.72925
R8253 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.n5 0.732092
R8254 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t3 0.7285
R8255 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t0 0.7285
R8256 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_7.B 0.438233
R8257 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n3 0.166901
R8258 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C 0.0455
R8259 adc_PISO_0.serial_out Piso_out 68.5339
R8260 Piso_out.n0 Piso_out.t5 40.6313
R8261 Piso_out.n0 Piso_out.t4 27.3166
R8262 Piso_out.n4 Piso_out.n0 14.6967
R8263 Piso_out.n3 Piso_out.t1 10.0473
R8264 Piso_out.n4 Piso_out.n3 9.39565
R8265 Piso_out.n2 Piso_out.t0 6.51042
R8266 Piso_out.n2 Piso_out.n1 6.04952
R8267 adc_PISO_0.serial_out adc_PISO_0.dffrs_5.Q 5.90514
R8268 Piso_out.n3 Piso_out.n2 0.732092
R8269 Piso_out.n1 Piso_out.t3 0.7285
R8270 Piso_out.n1 Piso_out.t2 0.7285
R8271 adc_PISO_0.dffrs_5.Q Piso_out.n4 0.458082
R8272 a_n4551_30169.n0 a_n4551_30169.t5 41.0041
R8273 a_n4551_30169.n1 a_n4551_30169.t7 40.8177
R8274 a_n4551_30169.n1 a_n4551_30169.t4 27.1302
R8275 a_n4551_30169.n0 a_n4551_30169.t6 26.9438
R8276 a_n4551_30169.n2 a_n4551_30169.n1 22.5284
R8277 a_n4551_30169.n3 a_n4551_30169.n2 19.5781
R8278 a_n4551_30169.n3 a_n4551_30169.t1 10.0473
R8279 a_n4551_30169.n4 a_n4551_30169.t3 6.51042
R8280 a_n4551_30169.n5 a_n4551_30169.n4 6.04952
R8281 a_n4551_30169.n2 a_n4551_30169.n0 5.7305
R8282 a_n4551_30169.n4 a_n4551_30169.n3 0.732092
R8283 a_n4551_30169.n5 a_n4551_30169.t2 0.7285
R8284 a_n4551_30169.t0 a_n4551_30169.n5 0.7285
R8285 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t4 41.0041
R8286 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t5 40.8177
R8287 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t7 27.1302
R8288 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t6 26.9438
R8289 SARlogic_0.dffrs_0.nand3_6.A SARlogic_0.dffrs_0.nand3_0.B 17.0041
R8290 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n2 14.8493
R8291 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.t0 10.0473
R8292 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.t1 6.51042
R8293 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.n3 6.04952
R8294 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_8.Z.n0 5.7305
R8295 SARlogic_0.dffrs_0.nand3_0.B SARlogic_0.dffrs_0.nand3_8.Z.n1 5.47979
R8296 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n5 4.72925
R8297 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.n4 0.732092
R8298 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t3 0.7285
R8299 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t2 0.7285
R8300 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_6.A 0.0455
R8301 a_11311_29264.n0 a_11311_29264.t5 34.1797
R8302 a_11311_29264.n0 a_11311_29264.t4 19.5798
R8303 a_11311_29264.n1 a_11311_29264.t3 10.3401
R8304 a_11311_29264.n1 a_11311_29264.t2 9.2885
R8305 a_11311_29264.n2 a_11311_29264.n0 4.93379
R8306 a_11311_29264.t1 a_11311_29264.n3 4.09202
R8307 a_11311_29264.n3 a_11311_29264.t0 3.95079
R8308 a_11311_29264.n2 a_11311_29264.n1 0.599711
R8309 a_11311_29264.n3 a_11311_29264.n2 0.296375
R8310 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t7 41.0041
R8311 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t4 40.8177
R8312 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t5 27.1302
R8313 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t6 26.9438
R8314 SARlogic_0.dffrs_5.nand3_6.A SARlogic_0.dffrs_5.nand3_0.B 17.0041
R8315 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n2 14.8493
R8316 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.t2 10.0473
R8317 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.t1 6.51042
R8318 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.n3 6.04952
R8319 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_8.Z.n0 5.7305
R8320 SARlogic_0.dffrs_5.nand3_0.B SARlogic_0.dffrs_5.nand3_8.Z.n1 5.47979
R8321 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n5 4.72925
R8322 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.n4 0.732092
R8323 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t3 0.7285
R8324 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t0 0.7285
R8325 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_6.A 0.0455
R8326 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t7 40.8177
R8327 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t5 40.6313
R8328 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t6 27.3166
R8329 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t4 27.1302
R8330 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_8.C.n2 14.119
R8331 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.t0 10.0473
R8332 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.t1 6.51042
R8333 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.n4 6.04952
R8334 SARlogic_0.dffrs_13.nand3_7.B SARlogic_0.dffrs_13.nand3_8.C.n0 5.47979
R8335 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C.n1 5.13907
R8336 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n6 4.72925
R8337 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.n5 0.732092
R8338 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t3 0.7285
R8339 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t2 0.7285
R8340 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_7.B 0.438233
R8341 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n3 0.166901
R8342 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C 0.0455
R8343 a_n7633_29263.n0 a_n7633_29263.t4 34.1797
R8344 a_n7633_29263.n0 a_n7633_29263.t5 19.5798
R8345 a_n7633_29263.t0 a_n7633_29263.n3 10.3401
R8346 a_n7633_29263.n3 a_n7633_29263.t3 9.2885
R8347 a_n7633_29263.n2 a_n7633_29263.n0 4.93379
R8348 a_n7633_29263.n1 a_n7633_29263.t1 4.09202
R8349 a_n7633_29263.n1 a_n7633_29263.t2 3.95079
R8350 a_n7633_29263.n3 a_n7633_29263.n2 0.599711
R8351 a_n7633_29263.n2 a_n7633_29263.n1 0.296375
R8352 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t2 41.0041
R8353 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t3 26.9438
R8354 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t0 9.6935
R8355 adc_PISO_0.dffrs_0.d adc_PISO_0.2inmux_0.OUT.n0 6.55979
R8356 adc_PISO_0.2inmux_0.OUT adc_PISO_0.dffrs_0.d 4.883
R8357 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t1 4.35383
R8358 adc_PISO_0.2inmux_0.OUT adc_PISO_0.2inmux_0.OUT.n1 0.350857
R8359 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t4 41.0041
R8360 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t6 40.6313
R8361 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t7 27.3166
R8362 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t5 26.9438
R8363 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_5.d 17.5382
R8364 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_4.Q.n2 14.0582
R8365 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.t2 10.0473
R8366 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.t3 6.51042
R8367 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.n4 6.04952
R8368 SARlogic_0.dffrs_5.nand3_8.A SARlogic_0.dffrs_4.Q.n0 5.7755
R8369 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.Q.n1 5.13907
R8370 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n6 4.72925
R8371 SARlogic_0.dffrs_5.d SARlogic_0.dffrs_5.nand3_8.A 0.784786
R8372 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.n5 0.732092
R8373 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t1 0.7285
R8374 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t0 0.7285
R8375 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n3 0.166901
R8376 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.nand3_7.C 0.0455
R8377 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t4 41.0041
R8378 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t7 40.6313
R8379 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t6 27.3166
R8380 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t5 26.9438
R8381 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_1.d 17.5382
R8382 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_0.Q.n2 14.0582
R8383 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.t1 10.0473
R8384 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.t0 6.51042
R8385 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.n4 6.04952
R8386 SARlogic_0.dffrs_1.nand3_8.A SARlogic_0.dffrs_0.Q.n0 5.7755
R8387 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.Q.n1 5.13907
R8388 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n6 4.72925
R8389 SARlogic_0.dffrs_1.d SARlogic_0.dffrs_1.nand3_8.A 0.784786
R8390 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.n5 0.732092
R8391 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t2 0.7285
R8392 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t3 0.7285
R8393 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n3 0.166901
R8394 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.nand3_7.C 0.0455
R8395 a_18555_28820.n0 a_18555_28820.t5 34.1797
R8396 a_18555_28820.n0 a_18555_28820.t4 19.5798
R8397 a_18555_28820.n1 a_18555_28820.t2 18.7717
R8398 a_18555_28820.n1 a_18555_28820.t1 9.2885
R8399 a_18555_28820.n2 a_18555_28820.n0 4.93379
R8400 a_18555_28820.t0 a_18555_28820.n3 4.23346
R8401 a_18555_28820.n3 a_18555_28820.t3 3.85546
R8402 a_18555_28820.n2 a_18555_28820.n1 0.4055
R8403 a_18555_28820.n3 a_18555_28820.n2 0.352625
R8404 a_23785_33628.n0 a_23785_33628.t4 40.6313
R8405 a_23785_33628.n0 a_23785_33628.t5 27.3166
R8406 a_23785_33628.n1 a_23785_33628.n0 24.1527
R8407 a_23785_33628.n1 a_23785_33628.t1 10.0473
R8408 a_23785_33628.n2 a_23785_33628.t2 6.51042
R8409 a_23785_33628.n3 a_23785_33628.n2 6.04952
R8410 a_23785_33628.n2 a_23785_33628.n1 0.732092
R8411 a_23785_33628.t0 a_23785_33628.n3 0.7285
R8412 a_23785_33628.n3 a_23785_33628.t3 0.7285
R8413 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t6 41.0041
R8414 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t5 40.8177
R8415 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t4 27.1302
R8416 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t7 26.9438
R8417 SARlogic_0.dffrs_1.nand3_6.A SARlogic_0.dffrs_1.nand3_0.B 17.0041
R8418 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n2 14.8493
R8419 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.t2 10.0473
R8420 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.t1 6.51042
R8421 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.n3 6.04952
R8422 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_8.Z.n0 5.7305
R8423 SARlogic_0.dffrs_1.nand3_0.B SARlogic_0.dffrs_1.nand3_8.Z.n1 5.47979
R8424 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n5 4.72925
R8425 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.n4 0.732092
R8426 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t3 0.7285
R8427 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t0 0.7285
R8428 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_6.A 0.0455
R8429 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t4 41.0041
R8430 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t7 40.6313
R8431 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t6 27.3166
R8432 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t5 26.9438
R8433 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d 17.5382
R8434 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d.n2 14.0582
R8435 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.t2 10.0473
R8436 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.t1 6.51042
R8437 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.n4 6.04952
R8438 SARlogic_0.dffrs_2.nand3_8.A SARlogic_0.dffrs_2.d.n0 5.7755
R8439 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_2.d.n1 5.13907
R8440 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n6 4.72925
R8441 SARlogic_0.dffrs_2.d SARlogic_0.dffrs_2.nand3_8.A 0.784786
R8442 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.n5 0.732092
R8443 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t0 0.7285
R8444 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t3 0.7285
R8445 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n3 0.166901
R8446 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_1.nand3_7.C 0.0455
R8447 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t5 40.6313
R8448 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t4 27.3166
R8449 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n1 14.2246
R8450 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.t1 10.0473
R8451 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.t0 6.51042
R8452 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.n2 6.04952
R8453 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.Q.n0 5.13907
R8454 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n4 4.72925
R8455 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.n3 0.732092
R8456 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t2 0.7285
R8457 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t3 0.7285
R8458 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.nand3_7.C 0.0455
R8459 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t5 41.0041
R8460 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t6 40.8177
R8461 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t4 40.6313
R8462 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t7 27.3166
R8463 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t8 27.1302
R8464 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t9 26.9438
R8465 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.t0 10.0473
R8466 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n4 9.90747
R8467 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n2 9.90116
R8468 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.t1 6.51042
R8469 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.n7 6.04952
R8470 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_6.C.n1 5.7305
R8471 SARlogic_0.dffrs_4.nand3_2.B SARlogic_0.dffrs_4.nand3_6.C.n0 5.47979
R8472 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C.n3 5.13907
R8473 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n9 4.72925
R8474 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_6.C.n5 4.5005
R8475 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.n8 0.732092
R8476 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t2 0.7285
R8477 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t3 0.7285
R8478 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n6 0.449758
R8479 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_2.B 0.166901
R8480 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_0.A 0.0455
R8481 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C 0.0455
R8482 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t2 41.0041
R8483 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t3 26.9438
R8484 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t0 9.6935
R8485 adc_PISO_0.dffrs_5.d adc_PISO_0.2inmux_1.OUT.n0 6.55979
R8486 adc_PISO_0.2inmux_1.OUT adc_PISO_0.dffrs_5.d 4.883
R8487 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t1 4.35383
R8488 adc_PISO_0.2inmux_1.OUT adc_PISO_0.2inmux_1.OUT.n1 0.350857
R8489 Load.n0 Load.t1 34.1797
R8490 Load.n0 Load.t0 19.5798
R8491 inv2_0.in Load.n0 4.87271
R8492 inv2_0.in Load 0.868357
R8493 a_42729_29218.n0 a_42729_29218.t5 40.8177
R8494 a_42729_29218.n1 a_42729_29218.t6 40.6313
R8495 a_42729_29218.n1 a_42729_29218.t4 27.3166
R8496 a_42729_29218.n0 a_42729_29218.t7 27.1302
R8497 a_42729_29218.n2 a_42729_29218.n1 19.2576
R8498 a_42729_29218.n3 a_42729_29218.t1 10.0473
R8499 a_42729_29218.n4 a_42729_29218.t2 6.51042
R8500 a_42729_29218.n5 a_42729_29218.n4 6.04952
R8501 a_42729_29218.n2 a_42729_29218.n0 5.91752
R8502 a_42729_29218.n3 a_42729_29218.n2 4.89565
R8503 a_42729_29218.n4 a_42729_29218.n3 0.732092
R8504 a_42729_29218.t0 a_42729_29218.n5 0.7285
R8505 a_42729_29218.n5 a_42729_29218.t3 0.7285
R8506 a_18555_31160.n0 a_18555_31160.t5 34.1797
R8507 a_18555_31160.n0 a_18555_31160.t4 19.5798
R8508 a_18555_31160.n1 a_18555_31160.t1 18.7717
R8509 a_18555_31160.n1 a_18555_31160.t2 9.2885
R8510 a_18555_31160.n2 a_18555_31160.n0 4.93379
R8511 a_18555_31160.t0 a_18555_31160.n3 4.23346
R8512 a_18555_31160.n3 a_18555_31160.t3 3.85546
R8513 a_18555_31160.n2 a_18555_31160.n1 0.4055
R8514 a_18555_31160.n3 a_18555_31160.n2 0.352625
R8515 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t7 41.0041
R8516 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t5 40.8177
R8517 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t6 40.6313
R8518 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t9 27.3166
R8519 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t8 27.1302
R8520 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t4 26.9438
R8521 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.t2 10.0473
R8522 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n4 9.90747
R8523 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n2 9.90116
R8524 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.t3 6.51042
R8525 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.n7 6.04952
R8526 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_6.C.n1 5.7305
R8527 SARlogic_0.dffrs_13.nand3_2.B SARlogic_0.dffrs_13.nand3_6.C.n0 5.47979
R8528 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C.n3 5.13907
R8529 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n9 4.72925
R8530 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_6.C.n5 4.5005
R8531 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.n8 0.732092
R8532 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t0 0.7285
R8533 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t1 0.7285
R8534 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n6 0.449758
R8535 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_2.B 0.166901
R8536 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_0.A 0.0455
R8537 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C 0.0455
R8538 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t4 40.6313
R8539 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t5 27.3166
R8540 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n1 14.2854
R8541 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.t0 10.0473
R8542 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.t1 6.51042
R8543 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.n2 6.04952
R8544 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C.n0 5.13907
R8545 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n4 4.72925
R8546 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.n3 0.732092
R8547 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t2 0.7285
R8548 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t3 0.7285
R8549 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C 0.0455
R8550 a_n9861_28819.n0 a_n9861_28819.t5 34.1797
R8551 a_n9861_28819.n0 a_n9861_28819.t4 19.5798
R8552 a_n9861_28819.n1 a_n9861_28819.t2 18.7717
R8553 a_n9861_28819.n1 a_n9861_28819.t3 9.2885
R8554 a_n9861_28819.n2 a_n9861_28819.n0 4.93379
R8555 a_n9861_28819.t0 a_n9861_28819.n3 4.23346
R8556 a_n9861_28819.n3 a_n9861_28819.t1 3.85546
R8557 a_n9861_28819.n2 a_n9861_28819.n1 0.4055
R8558 a_n9861_28819.n3 a_n9861_28819.n2 0.352625
R8559 a_37499_28820.n0 a_37499_28820.t5 34.1797
R8560 a_37499_28820.n0 a_37499_28820.t4 19.5798
R8561 a_37499_28820.n1 a_37499_28820.t1 18.7717
R8562 a_37499_28820.n1 a_37499_28820.t2 9.2885
R8563 a_37499_28820.n2 a_37499_28820.n0 4.93379
R8564 a_37499_28820.t0 a_37499_28820.n3 4.23346
R8565 a_37499_28820.n3 a_37499_28820.t3 3.85546
R8566 a_37499_28820.n2 a_37499_28820.n1 0.4055
R8567 a_37499_28820.n3 a_37499_28820.n2 0.352625
R8568 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t4 40.6313
R8569 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t5 27.3166
R8570 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n1 14.2854
R8571 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.t2 10.0473
R8572 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.t3 6.51042
R8573 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.n2 6.04952
R8574 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C.n0 5.13907
R8575 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n4 4.72925
R8576 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.n3 0.732092
R8577 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t0 0.7285
R8578 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t1 0.7285
R8579 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C 0.0455
R8580 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t5 41.0041
R8581 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t6 40.6313
R8582 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t4 27.3166
R8583 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t7 26.9438
R8584 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_3.d 17.5382
R8585 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_2.Q.n2 14.0582
R8586 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.t3 10.0473
R8587 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.t2 6.51042
R8588 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.n4 6.04952
R8589 SARlogic_0.dffrs_3.nand3_8.A SARlogic_0.dffrs_2.Q.n0 5.7755
R8590 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.Q.n1 5.13907
R8591 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n6 4.72925
R8592 SARlogic_0.dffrs_3.d SARlogic_0.dffrs_3.nand3_8.A 0.784786
R8593 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.n5 0.732092
R8594 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t0 0.7285
R8595 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t1 0.7285
R8596 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n3 0.166901
R8597 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.nand3_7.C 0.0455
R8598 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t6 40.6313
R8599 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.t5 34.1066
R8600 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t7 27.3166
R8601 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t8 19.673
R8602 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t4 19.4007
R8603 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n3 14.6967
R8604 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.t1 10.0473
R8605 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n6 9.39565
R8606 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.dffrs_2.Q.n1 6.70486
R8607 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.t0 6.51042
R8608 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.n4 6.04952
R8609 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n2 5.81514
R8610 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.n5 0.732092
R8611 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t3 0.7285
R8612 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t2 0.7285
R8613 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n7 0.458082
R8614 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.n0 0.252687
R8615 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.2inmux_4.Bit 0.0519286
R8616 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t4 40.6313
R8617 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t5 27.3166
R8618 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n1 14.2854
R8619 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.t1 10.0473
R8620 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.t2 6.51042
R8621 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.n2 6.04952
R8622 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C.n0 5.13907
R8623 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n4 4.72925
R8624 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.n3 0.732092
R8625 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t0 0.7285
R8626 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t3 0.7285
R8627 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C 0.0455
R8628 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t3 41.0041
R8629 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t2 26.9438
R8630 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t0 9.6935
R8631 adc_PISO_0.dffrs_3.d adc_PISO_0.2inmux_4.OUT.n0 6.55979
R8632 adc_PISO_0.2inmux_4.OUT adc_PISO_0.dffrs_3.d 4.883
R8633 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t1 4.35383
R8634 adc_PISO_0.2inmux_4.OUT adc_PISO_0.2inmux_4.OUT.n1 0.350857
R8635 a_14313_31423.n3 a_14313_31423.t4 41.0041
R8636 a_14313_31423.n2 a_14313_31423.t6 40.8177
R8637 a_14313_31423.n4 a_14313_31423.t5 40.6313
R8638 a_14313_31423.n4 a_14313_31423.t8 27.3166
R8639 a_14313_31423.n2 a_14313_31423.t9 27.1302
R8640 a_14313_31423.n3 a_14313_31423.t7 26.9438
R8641 a_14313_31423.n5 a_14313_31423.n3 15.6312
R8642 a_14313_31423.n5 a_14313_31423.n4 15.046
R8643 a_14313_31423.t0 a_14313_31423.n7 10.0473
R8644 a_14313_31423.n1 a_14313_31423.t1 6.51042
R8645 a_14313_31423.n1 a_14313_31423.n0 6.04952
R8646 a_14313_31423.n6 a_14313_31423.n2 5.64619
R8647 a_14313_31423.n7 a_14313_31423.n6 5.17851
R8648 a_14313_31423.n6 a_14313_31423.n5 4.5005
R8649 a_14313_31423.n7 a_14313_31423.n1 0.732092
R8650 a_14313_31423.n0 a_14313_31423.t3 0.7285
R8651 a_14313_31423.n0 a_14313_31423.t2 0.7285
R8652 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t4 41.0041
R8653 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t7 40.6313
R8654 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t6 40.6313
R8655 SARlogic_0.dffrs_2.Qb SARlogic_0.dffrs_9.setb 28.021
R8656 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t9 27.3166
R8657 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t8 27.3166
R8658 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t5 26.9438
R8659 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.t2 10.0473
R8660 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb.n1 9.84255
R8661 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n3 9.22229
R8662 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.t3 6.51042
R8663 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.n7 6.04952
R8664 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.Qb.n0 5.7305
R8665 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n4 5.14711
R8666 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_2.Qb.n2 5.13907
R8667 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n6 4.94976
R8668 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n9 4.72925
R8669 SARlogic_0.dffrs_9.setb SARlogic_0.dffrs_9.nand3_0.C 0.784786
R8670 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.n8 0.732092
R8671 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t0 0.7285
R8672 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t1 0.7285
R8673 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb 0.175225
R8674 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.nand3_2.A 0.0455
R8675 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_9.nand3_2.C 0.0455
R8676 SARlogic_0.dffrs_9.nand3_0.C SARlogic_0.dffrs_2.Qb.n5 0.0374643
.ends

