magic
tech gf180mcuD
magscale 1 10
timestamp 1755268346
<< error_p >>
rect -34 113 -23 159
rect 23 113 34 124
rect -80 -78 -57 -67
rect 57 -78 80 -67
rect -34 -159 -23 -113
<< nwell >>
rect -278 -290 278 290
<< pmos >>
rect -28 -80 28 80
<< pdiff >>
rect -116 67 -28 80
rect -116 -67 -103 67
rect -57 -67 -28 67
rect -116 -80 -28 -67
rect 28 67 116 80
rect 28 -67 57 67
rect 103 -67 116 67
rect 28 -80 116 -67
<< pdiffc >>
rect -103 -67 -57 67
rect 57 -67 103 67
<< nsubdiff >>
rect -254 194 254 266
rect -254 150 -182 194
rect -254 -150 -241 150
rect -195 -150 -182 150
rect 182 150 254 194
rect -254 -194 -182 -150
rect 182 -150 195 150
rect 241 -150 254 150
rect 182 -194 254 -150
rect -254 -266 254 -194
<< nsubdiffcont >>
rect -241 -150 -195 150
rect 195 -150 241 150
<< polysilicon >>
rect -36 159 36 172
rect -36 113 -23 159
rect 23 113 36 159
rect -36 100 36 113
rect -28 80 28 100
rect -28 -100 28 -80
rect -36 -113 36 -100
rect -36 -159 -23 -113
rect 23 -159 36 -113
rect -36 -172 36 -159
<< polycontact >>
rect -23 113 23 159
rect -23 -159 23 -113
<< metal1 >>
rect -241 207 241 253
rect -241 150 -195 207
rect -34 113 -23 159
rect 23 113 34 159
rect 195 150 241 207
rect -103 67 -57 78
rect -103 -78 -57 -67
rect 57 67 103 78
rect 57 -78 103 -67
rect -241 -207 -195 -150
rect -34 -159 -23 -113
rect 23 -159 34 -113
rect 195 -207 241 -150
rect -241 -253 241 -207
<< properties >>
string FIXED_BBOX -218 -230 218 230
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.8 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
