magic
tech gf180mcuD
magscale 1 10
timestamp 1757551291
<< error_s >>
rect 635 -937 667 -891
rect 154 -1000 192 -971
rect 376 -1017 387 -971
rect 633 -1040 667 -992
rect 681 -1040 713 -937
rect 1339 -960 1371 -951
rect 1339 -997 1408 -960
rect 376 -1929 387 -1883
rect 681 -1920 715 -1040
rect 896 -1077 907 -1031
rect 1080 -1077 1091 -1031
rect 1348 -1052 1417 -997
rect 1337 -1100 1417 -1052
rect 2043 -1057 2075 -1011
rect 681 -2023 713 -1920
rect 896 -1989 907 -1943
rect 1080 -1989 1091 -1943
rect 1348 -1980 1419 -1100
rect 1600 -1137 1611 -1091
rect 1784 -1137 1795 -1091
rect 2041 -1160 2075 -1112
rect 2089 -1160 2121 -1057
rect 1348 -2083 1417 -1980
rect 1600 -2049 1611 -2003
rect 1784 -2049 1795 -2003
rect 2089 -2040 2123 -1160
rect 2304 -1197 2315 -1151
rect 2488 -1197 2499 -1151
rect 2840 -1435 2848 -988
rect 2784 -1492 2792 -1436
rect 1348 -2120 1408 -2083
rect 2089 -2143 2121 -2040
rect 2304 -2109 2315 -2063
rect 2488 -2109 2499 -2063
rect 2840 -2216 2848 -1492
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use CDAC_INV_V0  x1v
timestamp 1757551132
transform 1 0 1853 0 1 -920
box 963 -1320 1714 633
use nfet_03v3_W5K4UP  XM1
timestamp 0
transform 1 0 322 0 1 -1450
box -382 -610 382 610
use pfet_03v3_LS6D84  XM2
timestamp 0
transform 1 0 2434 0 1 -1630
box -382 -610 382 610
use nfet_03v3_W5K4UP  XM3
timestamp 0
transform 1 0 1026 0 1 -1510
box -382 -610 382 610
use pfet_03v3_LS6D84  XM4
timestamp 0
transform 1 0 1730 0 1 -1570
box -382 -610 382 610
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 sw_vout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 sw_bit
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 avss
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 avdd
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 sw_Vref
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 1280 0 0 0 vreflow
port 5 nsew
<< end >>
