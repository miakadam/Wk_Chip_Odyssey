magic
tech gf180mcuD
magscale 1 10
timestamp 1757675171
<< nwell >>
rect 2060 -1120 3100 -500
<< pwell >>
rect 2060 -1940 3100 -1320
<< nmos >>
rect 2310 -1730 2390 -1530
rect 2770 -1730 2850 -1530
<< pmos >>
rect 2310 -910 2390 -710
rect 2770 -910 2850 -710
<< ndiff >>
rect 2222 -1543 2310 -1530
rect 2222 -1717 2235 -1543
rect 2281 -1717 2310 -1543
rect 2222 -1730 2310 -1717
rect 2390 -1543 2478 -1530
rect 2390 -1717 2419 -1543
rect 2465 -1717 2478 -1543
rect 2390 -1730 2478 -1717
rect 2682 -1543 2770 -1530
rect 2682 -1717 2695 -1543
rect 2741 -1717 2770 -1543
rect 2682 -1730 2770 -1717
rect 2850 -1543 2938 -1530
rect 2850 -1717 2879 -1543
rect 2925 -1717 2938 -1543
rect 2850 -1730 2938 -1717
<< pdiff >>
rect 2222 -723 2310 -710
rect 2222 -897 2235 -723
rect 2281 -897 2310 -723
rect 2222 -910 2310 -897
rect 2390 -723 2478 -710
rect 2390 -897 2419 -723
rect 2465 -897 2478 -723
rect 2390 -910 2478 -897
rect 2682 -723 2770 -710
rect 2682 -897 2695 -723
rect 2741 -897 2770 -723
rect 2682 -910 2770 -897
rect 2850 -723 2938 -710
rect 2850 -897 2879 -723
rect 2925 -897 2938 -723
rect 2850 -910 2938 -897
<< ndiffc >>
rect 2235 -1717 2281 -1543
rect 2419 -1717 2465 -1543
rect 2695 -1717 2741 -1543
rect 2879 -1717 2925 -1543
<< pdiffc >>
rect 2235 -897 2281 -723
rect 2419 -897 2465 -723
rect 2695 -897 2741 -723
rect 2879 -897 2925 -723
<< psubdiff >>
rect 2084 -1416 3076 -1344
rect 2084 -1460 2156 -1416
rect 2084 -1800 2097 -1460
rect 2143 -1800 2156 -1460
rect 2544 -1460 2616 -1416
rect 2084 -1844 2156 -1800
rect 2544 -1800 2557 -1460
rect 2603 -1800 2616 -1460
rect 3004 -1460 3076 -1416
rect 2544 -1844 2616 -1800
rect 3004 -1800 3017 -1460
rect 3063 -1800 3076 -1460
rect 3004 -1844 3076 -1800
rect 2084 -1916 3076 -1844
<< nsubdiff >>
rect 2084 -596 3076 -524
rect 2084 -640 2156 -596
rect 2084 -980 2097 -640
rect 2143 -980 2156 -640
rect 2544 -640 2616 -596
rect 2084 -1024 2156 -980
rect 2544 -980 2557 -640
rect 2603 -980 2616 -640
rect 3004 -640 3076 -596
rect 2544 -1024 2616 -980
rect 3004 -980 3017 -640
rect 3063 -980 3076 -640
rect 3004 -1024 3076 -980
rect 2084 -1096 3076 -1024
<< psubdiffcont >>
rect 2097 -1800 2143 -1460
rect 2557 -1800 2603 -1460
rect 3017 -1800 3063 -1460
<< nsubdiffcont >>
rect 2097 -980 2143 -640
rect 2557 -980 2603 -640
rect 3017 -980 3063 -640
<< polysilicon >>
rect 2310 -631 2390 -618
rect 2310 -677 2323 -631
rect 2377 -677 2390 -631
rect 2310 -710 2390 -677
rect 2310 -943 2390 -910
rect 2310 -989 2323 -943
rect 2377 -989 2390 -943
rect 2310 -1002 2390 -989
rect 2770 -631 2850 -618
rect 2770 -677 2783 -631
rect 2837 -677 2850 -631
rect 2770 -710 2850 -677
rect 2770 -943 2850 -910
rect 2770 -989 2783 -943
rect 2837 -989 2850 -943
rect 2770 -1002 2850 -989
rect 2310 -1451 2390 -1438
rect 2310 -1497 2323 -1451
rect 2377 -1497 2390 -1451
rect 2310 -1530 2390 -1497
rect 2310 -1763 2390 -1730
rect 2310 -1809 2323 -1763
rect 2377 -1809 2390 -1763
rect 2310 -1822 2390 -1809
rect 2770 -1451 2850 -1438
rect 2770 -1497 2783 -1451
rect 2837 -1497 2850 -1451
rect 2770 -1530 2850 -1497
rect 2770 -1763 2850 -1730
rect 2770 -1809 2783 -1763
rect 2837 -1809 2850 -1763
rect 2770 -1822 2850 -1809
<< polycontact >>
rect 2323 -677 2377 -631
rect 2323 -989 2377 -943
rect 2783 -677 2837 -631
rect 2783 -989 2837 -943
rect 2323 -1497 2377 -1451
rect 2323 -1809 2377 -1763
rect 2783 -1497 2837 -1451
rect 2783 -1809 2837 -1763
<< metal1 >>
rect 2097 -500 3063 -420
rect 2097 -640 2143 -500
rect 2312 -631 2388 -598
rect 2312 -677 2323 -631
rect 2377 -677 2388 -631
rect 2557 -640 2603 -629
rect 2235 -723 2281 -712
rect 2143 -897 2235 -723
rect 2419 -723 2465 -712
rect 2402 -782 2419 -772
rect 2465 -782 2482 -772
rect 2402 -838 2414 -782
rect 2470 -838 2482 -782
rect 2402 -848 2419 -838
rect 2235 -908 2281 -897
rect 2465 -848 2482 -838
rect 2419 -908 2465 -897
rect 2097 -991 2143 -980
rect 2312 -989 2323 -943
rect 2377 -989 2388 -943
rect 2772 -631 2848 -598
rect 2772 -677 2783 -631
rect 2837 -677 2848 -631
rect 3017 -640 3063 -500
rect 2695 -723 2741 -712
rect 2678 -782 2695 -772
rect 2879 -723 2925 -712
rect 2741 -782 2758 -772
rect 2678 -838 2690 -782
rect 2746 -838 2758 -782
rect 2678 -848 2695 -838
rect 2741 -848 2758 -838
rect 2695 -908 2741 -897
rect 2925 -897 3017 -723
rect 2879 -908 2925 -897
rect 2322 -1176 2378 -989
rect 2557 -991 2603 -980
rect 2772 -989 2783 -943
rect 2837 -989 2848 -943
rect 2540 -1040 2610 -1038
rect 2782 -1040 2838 -989
rect 3017 -991 3063 -980
rect 2540 -1096 2552 -1040
rect 2608 -1096 2838 -1040
rect 2540 -1098 2610 -1096
rect 2322 -1178 2620 -1176
rect 2322 -1234 2552 -1178
rect 2608 -1234 2620 -1178
rect 2322 -1236 2620 -1234
rect 2097 -1460 2143 -1449
rect 2312 -1451 2388 -1418
rect 2312 -1497 2323 -1451
rect 2377 -1497 2388 -1451
rect 2557 -1460 2603 -1449
rect 2235 -1543 2281 -1532
rect 2143 -1717 2235 -1543
rect 2419 -1543 2465 -1532
rect 2402 -1602 2419 -1592
rect 2465 -1602 2482 -1592
rect 2402 -1658 2414 -1602
rect 2470 -1658 2482 -1602
rect 2402 -1668 2419 -1658
rect 2235 -1728 2281 -1717
rect 2465 -1668 2482 -1658
rect 2419 -1728 2465 -1717
rect 2312 -1768 2323 -1763
rect 2097 -1940 2143 -1800
rect 2310 -1778 2323 -1768
rect 2377 -1768 2388 -1763
rect 2377 -1778 2390 -1768
rect 2310 -1834 2322 -1778
rect 2378 -1834 2390 -1778
rect 2772 -1451 2848 -1418
rect 2772 -1497 2783 -1451
rect 2837 -1497 2848 -1451
rect 3017 -1460 3063 -1449
rect 2695 -1543 2741 -1532
rect 2678 -1602 2695 -1592
rect 2879 -1543 2925 -1532
rect 2741 -1602 2758 -1592
rect 2678 -1658 2690 -1602
rect 2746 -1658 2758 -1602
rect 2678 -1668 2695 -1658
rect 2741 -1668 2758 -1658
rect 2695 -1728 2741 -1717
rect 2925 -1717 3017 -1543
rect 2879 -1728 2925 -1717
rect 2772 -1768 2783 -1763
rect 2557 -1811 2603 -1800
rect 2770 -1778 2783 -1768
rect 2837 -1768 2848 -1763
rect 2837 -1778 2850 -1768
rect 2310 -1844 2390 -1834
rect 2770 -1834 2782 -1778
rect 2838 -1834 2850 -1778
rect 2770 -1844 2850 -1834
rect 3017 -1940 3063 -1800
rect 2097 -2020 3063 -1940
<< via1 >>
rect 2414 -838 2419 -782
rect 2419 -838 2465 -782
rect 2465 -838 2470 -782
rect 2690 -838 2695 -782
rect 2695 -838 2741 -782
rect 2741 -838 2746 -782
rect 2552 -1096 2608 -1040
rect 2552 -1234 2608 -1178
rect 2414 -1658 2419 -1602
rect 2419 -1658 2465 -1602
rect 2465 -1658 2470 -1602
rect 2322 -1809 2323 -1778
rect 2323 -1809 2377 -1778
rect 2377 -1809 2378 -1778
rect 2322 -1834 2378 -1809
rect 2690 -1658 2695 -1602
rect 2695 -1658 2741 -1602
rect 2741 -1658 2746 -1602
rect 2782 -1809 2783 -1778
rect 2783 -1809 2837 -1778
rect 2837 -1809 2838 -1778
rect 2782 -1834 2838 -1809
<< metal2 >>
rect 2402 -782 2482 -772
rect 2402 -838 2414 -782
rect 2470 -838 2482 -782
rect 2402 -848 2482 -838
rect 2678 -782 2758 -772
rect 2678 -838 2690 -782
rect 2746 -838 2758 -782
rect 2678 -848 2758 -838
rect 2414 -1040 2470 -848
rect 2539 -1040 2619 -1028
rect 2414 -1096 2552 -1040
rect 2608 -1096 2619 -1040
rect 2414 -1288 2470 -1096
rect 2539 -1108 2619 -1096
rect 2540 -1178 2620 -1168
rect 2690 -1178 2746 -848
rect 2540 -1234 2552 -1178
rect 2608 -1234 2746 -1178
rect 2540 -1244 2620 -1234
rect 1870 -1344 2470 -1288
rect 2414 -1592 2470 -1344
rect 2690 -1288 2746 -1234
rect 2690 -1344 3290 -1288
rect 2690 -1592 2746 -1344
rect 2402 -1602 2482 -1592
rect 2402 -1658 2414 -1602
rect 2470 -1658 2482 -1602
rect 2402 -1668 2482 -1658
rect 2678 -1602 2758 -1592
rect 2678 -1658 2690 -1602
rect 2746 -1658 2758 -1602
rect 2678 -1668 2758 -1658
rect 2310 -1778 2390 -1768
rect 2310 -1834 2322 -1778
rect 2378 -1834 2390 -1778
rect 2310 -1844 2390 -1834
rect 2770 -1778 2850 -1768
rect 2770 -1834 2782 -1778
rect 2838 -1834 2850 -1778
rect 2770 -1844 2850 -1834
rect 2322 -2178 2378 -1844
rect 2782 -2178 2838 -1844
<< labels >>
rlabel metal1 2578 -420 2578 -420 1 VDD
port 0 n
rlabel metal2 1870 -1318 1870 -1318 7 Vout1
port 1 w
rlabel metal2 3290 -1318 3290 -1318 3 Vout2
port 2 e
rlabel metal2 2350 -2178 2350 -2178 5 Vin1
port 3 s
rlabel metal2 2811 -2178 2811 -2178 5 Vin2
port 4 s
rlabel metal1 2583 -2020 2583 -2020 5 VSS
port 5 s
<< end >>
