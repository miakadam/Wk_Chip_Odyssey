magic
tech gf180mcuD
magscale 1 5
timestamp 1757048890
use nfet_03v3_3TMVZR  XM9
timestamp 1757048890
transform 1 0 1374 0 1 560
box -479 -180 479 180
use nfet_03v3_3TMVZR  XM10
timestamp 1757048890
transform 1 0 1377 0 1 120
box -479 -180 479 180
use nfet_03v3_3TMVZR  XM20
timestamp 1757048890
transform 1 0 2454 0 1 130
box -479 -180 479 180
use nfet_03v3_3TMVZR  XM21
timestamp 1757048890
transform 1 0 2469 0 1 575
box -479 -180 479 180
<< end >>
