magic
tech gf180mcuD
magscale 1 10
timestamp 1757846348
<< nwell >>
rect 4648 17287 5596 18207
rect 8690 17284 9638 18204
rect 12732 17284 13680 18204
rect 16774 17284 17722 18204
rect 20816 17284 21764 18204
rect 24858 17284 25806 18204
rect 28900 17284 29848 18204
rect 4648 15082 5596 16002
rect 6134 15082 7082 16002
rect 8690 15079 9638 15999
rect 10176 15079 11124 15999
rect 12732 15079 13680 15999
rect 14218 15079 15166 15999
rect 16774 15079 17722 15999
rect 18260 15079 19208 15999
rect 20816 15079 21764 15999
rect 22302 15079 23250 15999
rect 24858 15079 25806 15999
rect 26344 15079 27292 15999
rect 28900 15079 29848 15999
rect 30386 15079 31334 15999
rect 4648 12877 5596 13797
rect 6134 12878 7082 13798
rect 8690 12874 9638 13794
rect 10176 12875 11124 13795
rect 12732 12874 13680 13794
rect 14218 12875 15166 13795
rect 16774 12874 17722 13794
rect 18260 12875 19208 13795
rect 20816 12874 21764 13794
rect 22302 12875 23250 13795
rect 24858 12874 25806 13794
rect 26344 12875 27292 13795
rect 28900 12874 29848 13794
rect 30386 12875 31334 13795
rect 4648 10672 5596 11592
rect 8690 10669 9638 11589
rect 12732 10669 13680 11589
rect 16774 10669 17722 11589
rect 20816 10669 21764 11589
rect 24858 10669 25806 11589
rect 28900 10669 29848 11589
rect 636 7708 1584 8628
rect 4648 7708 5596 8628
rect 8690 7708 9638 8628
rect 12732 7708 13680 8628
rect 16774 7708 17722 8628
rect 20816 7708 21764 8628
rect 24858 7708 25806 8628
rect 636 5503 1584 6423
rect 2122 5503 3070 6423
rect 4648 5503 5596 6423
rect 6134 5503 7082 6423
rect 8690 5503 9638 6423
rect 10176 5503 11124 6423
rect 12732 5503 13680 6423
rect 14218 5503 15166 6423
rect 16774 5503 17722 6423
rect 18260 5503 19208 6423
rect 20816 5503 21764 6423
rect 22302 5503 23250 6423
rect 24858 5503 25806 6423
rect 26344 5503 27292 6423
rect 636 3298 1584 4218
rect 2122 3299 3070 4219
rect 4648 3298 5596 4218
rect 6134 3299 7082 4219
rect 8690 3298 9638 4218
rect 10176 3299 11124 4219
rect 12732 3298 13680 4218
rect 14218 3299 15166 4219
rect 16774 3298 17722 4218
rect 18260 3299 19208 4219
rect 20816 3298 21764 4218
rect 22302 3299 23250 4219
rect 24858 3298 25806 4218
rect 26344 3299 27292 4219
rect 636 1093 1584 2013
rect 4648 1093 5596 2013
rect 8690 1093 9638 2013
rect 12732 1093 13680 2013
rect 16774 1093 17722 2013
rect 20816 1093 21764 2013
rect 24858 1093 25806 2013
<< pwell >>
rect 5411 17047 5479 17287
rect 4648 16427 5596 17047
rect 9453 17044 9521 17284
rect 13495 17044 13563 17284
rect 17537 17044 17605 17284
rect 21579 17044 21647 17284
rect 25621 17044 25689 17284
rect 29663 17044 29731 17284
rect 8690 16424 9638 17044
rect 12732 16424 13680 17044
rect 16774 16424 17722 17044
rect 20816 16424 21764 17044
rect 24858 16424 25806 17044
rect 28900 16424 29848 17044
rect 5411 14842 5479 15082
rect 6897 14842 6965 15082
rect 4648 14222 5596 14842
rect 6134 14222 7082 14842
rect 9453 14839 9521 15079
rect 10939 14839 11007 15079
rect 13495 14839 13563 15079
rect 14981 14839 15049 15079
rect 17537 14839 17605 15079
rect 19023 14839 19091 15079
rect 21579 14839 21647 15079
rect 23065 14839 23133 15079
rect 25621 14839 25689 15079
rect 27107 14839 27175 15079
rect 29663 14839 29731 15079
rect 31149 14839 31217 15079
rect 8690 14219 9638 14839
rect 10176 14219 11124 14839
rect 12732 14219 13680 14839
rect 14218 14219 15166 14839
rect 16774 14219 17722 14839
rect 18260 14219 19208 14839
rect 20816 14219 21764 14839
rect 22302 14219 23250 14839
rect 24858 14219 25806 14839
rect 26344 14219 27292 14839
rect 28900 14219 29848 14839
rect 30386 14219 31334 14839
rect 5411 12637 5479 12877
rect 6897 12638 6965 12878
rect 4648 12017 5596 12637
rect 6134 12018 7082 12638
rect 9453 12634 9521 12874
rect 10939 12635 11007 12875
rect 8690 12014 9638 12634
rect 10176 12015 11124 12635
rect 13495 12634 13563 12874
rect 14981 12635 15049 12875
rect 12732 12014 13680 12634
rect 14218 12015 15166 12635
rect 17537 12634 17605 12874
rect 19023 12635 19091 12875
rect 16774 12014 17722 12634
rect 18260 12015 19208 12635
rect 21579 12634 21647 12874
rect 23065 12635 23133 12875
rect 20816 12014 21764 12634
rect 22302 12015 23250 12635
rect 25621 12634 25689 12874
rect 27107 12635 27175 12875
rect 24858 12014 25806 12634
rect 26344 12015 27292 12635
rect 29663 12634 29731 12874
rect 31149 12635 31217 12875
rect 28900 12014 29848 12634
rect 30386 12015 31334 12635
rect 5411 10432 5479 10672
rect 4648 9812 5596 10432
rect 9453 10429 9521 10669
rect 13495 10429 13563 10669
rect 17537 10429 17605 10669
rect 21579 10429 21647 10669
rect 25621 10429 25689 10669
rect 29663 10429 29731 10669
rect 8690 9809 9638 10429
rect 12732 9809 13680 10429
rect 16774 9809 17722 10429
rect 20816 9809 21764 10429
rect 24858 9809 25806 10429
rect 28900 9809 29848 10429
rect 1399 7468 1467 7708
rect 5411 7468 5479 7708
rect 9453 7468 9521 7708
rect 13495 7468 13563 7708
rect 17537 7468 17605 7708
rect 21579 7468 21647 7708
rect 25621 7468 25689 7708
rect 636 6848 1584 7468
rect 4648 6848 5596 7468
rect 8690 6848 9638 7468
rect 12732 6848 13680 7468
rect 16774 6848 17722 7468
rect 20816 6848 21764 7468
rect 24858 6848 25806 7468
rect 1399 5263 1467 5503
rect 2885 5263 2953 5503
rect 5411 5263 5479 5503
rect 6897 5263 6965 5503
rect 9453 5263 9521 5503
rect 10939 5263 11007 5503
rect 13495 5263 13563 5503
rect 14981 5263 15049 5503
rect 17537 5263 17605 5503
rect 19023 5263 19091 5503
rect 21579 5263 21647 5503
rect 23065 5263 23133 5503
rect 25621 5263 25689 5503
rect 27107 5263 27175 5503
rect 636 4643 1584 5263
rect 2122 4643 3070 5263
rect 4648 4643 5596 5263
rect 6134 4643 7082 5263
rect 8690 4643 9638 5263
rect 10176 4643 11124 5263
rect 12732 4643 13680 5263
rect 14218 4643 15166 5263
rect 16774 4643 17722 5263
rect 18260 4643 19208 5263
rect 20816 4643 21764 5263
rect 22302 4643 23250 5263
rect 24858 4643 25806 5263
rect 26344 4643 27292 5263
rect 1399 3058 1467 3298
rect 2885 3059 2953 3299
rect 636 2438 1584 3058
rect 2122 2439 3070 3059
rect 5411 3058 5479 3298
rect 6897 3059 6965 3299
rect 4648 2438 5596 3058
rect 6134 2439 7082 3059
rect 9453 3058 9521 3298
rect 10939 3059 11007 3299
rect 8690 2438 9638 3058
rect 10176 2439 11124 3059
rect 13495 3058 13563 3298
rect 14981 3059 15049 3299
rect 12732 2438 13680 3058
rect 14218 2439 15166 3059
rect 17537 3058 17605 3298
rect 19023 3059 19091 3299
rect 16774 2438 17722 3058
rect 18260 2439 19208 3059
rect 21579 3058 21647 3298
rect 23065 3059 23133 3299
rect 20816 2438 21764 3058
rect 22302 2439 23250 3059
rect 25621 3058 25689 3298
rect 27107 3059 27175 3299
rect 24858 2438 25806 3058
rect 26344 2439 27292 3059
rect 1399 853 1467 1093
rect 5411 853 5479 1093
rect 9453 853 9521 1093
rect 13495 853 13563 1093
rect 17537 853 17605 1093
rect 21579 853 21647 1093
rect 25621 853 25689 1093
rect 636 233 1584 853
rect 4648 233 5596 853
rect 8690 233 9638 853
rect 12732 233 13680 853
rect 16774 233 17722 853
rect 20816 233 21764 853
rect 24858 233 25806 853
<< nmos >>
rect 4898 16637 4978 16837
rect 5082 16637 5162 16837
rect 5266 16637 5346 16837
rect 8940 16634 9020 16834
rect 9124 16634 9204 16834
rect 9308 16634 9388 16834
rect 12982 16634 13062 16834
rect 13166 16634 13246 16834
rect 13350 16634 13430 16834
rect 17024 16634 17104 16834
rect 17208 16634 17288 16834
rect 17392 16634 17472 16834
rect 21066 16634 21146 16834
rect 21250 16634 21330 16834
rect 21434 16634 21514 16834
rect 25108 16634 25188 16834
rect 25292 16634 25372 16834
rect 25476 16634 25556 16834
rect 29150 16634 29230 16834
rect 29334 16634 29414 16834
rect 29518 16634 29598 16834
rect 4898 14432 4978 14632
rect 5082 14432 5162 14632
rect 5266 14432 5346 14632
rect 6384 14432 6464 14632
rect 6568 14432 6648 14632
rect 6752 14432 6832 14632
rect 8940 14429 9020 14629
rect 9124 14429 9204 14629
rect 9308 14429 9388 14629
rect 10426 14429 10506 14629
rect 10610 14429 10690 14629
rect 10794 14429 10874 14629
rect 12982 14429 13062 14629
rect 13166 14429 13246 14629
rect 13350 14429 13430 14629
rect 14468 14429 14548 14629
rect 14652 14429 14732 14629
rect 14836 14429 14916 14629
rect 17024 14429 17104 14629
rect 17208 14429 17288 14629
rect 17392 14429 17472 14629
rect 18510 14429 18590 14629
rect 18694 14429 18774 14629
rect 18878 14429 18958 14629
rect 21066 14429 21146 14629
rect 21250 14429 21330 14629
rect 21434 14429 21514 14629
rect 22552 14429 22632 14629
rect 22736 14429 22816 14629
rect 22920 14429 23000 14629
rect 25108 14429 25188 14629
rect 25292 14429 25372 14629
rect 25476 14429 25556 14629
rect 26594 14429 26674 14629
rect 26778 14429 26858 14629
rect 26962 14429 27042 14629
rect 29150 14429 29230 14629
rect 29334 14429 29414 14629
rect 29518 14429 29598 14629
rect 30636 14429 30716 14629
rect 30820 14429 30900 14629
rect 31004 14429 31084 14629
rect 4898 12227 4978 12427
rect 5082 12227 5162 12427
rect 5266 12227 5346 12427
rect 6384 12228 6464 12428
rect 6568 12228 6648 12428
rect 6752 12228 6832 12428
rect 8940 12224 9020 12424
rect 9124 12224 9204 12424
rect 9308 12224 9388 12424
rect 10426 12225 10506 12425
rect 10610 12225 10690 12425
rect 10794 12225 10874 12425
rect 12982 12224 13062 12424
rect 13166 12224 13246 12424
rect 13350 12224 13430 12424
rect 14468 12225 14548 12425
rect 14652 12225 14732 12425
rect 14836 12225 14916 12425
rect 17024 12224 17104 12424
rect 17208 12224 17288 12424
rect 17392 12224 17472 12424
rect 18510 12225 18590 12425
rect 18694 12225 18774 12425
rect 18878 12225 18958 12425
rect 21066 12224 21146 12424
rect 21250 12224 21330 12424
rect 21434 12224 21514 12424
rect 22552 12225 22632 12425
rect 22736 12225 22816 12425
rect 22920 12225 23000 12425
rect 25108 12224 25188 12424
rect 25292 12224 25372 12424
rect 25476 12224 25556 12424
rect 26594 12225 26674 12425
rect 26778 12225 26858 12425
rect 26962 12225 27042 12425
rect 29150 12224 29230 12424
rect 29334 12224 29414 12424
rect 29518 12224 29598 12424
rect 30636 12225 30716 12425
rect 30820 12225 30900 12425
rect 31004 12225 31084 12425
rect 4898 10022 4978 10222
rect 5082 10022 5162 10222
rect 5266 10022 5346 10222
rect 8940 10019 9020 10219
rect 9124 10019 9204 10219
rect 9308 10019 9388 10219
rect 12982 10019 13062 10219
rect 13166 10019 13246 10219
rect 13350 10019 13430 10219
rect 17024 10019 17104 10219
rect 17208 10019 17288 10219
rect 17392 10019 17472 10219
rect 21066 10019 21146 10219
rect 21250 10019 21330 10219
rect 21434 10019 21514 10219
rect 25108 10019 25188 10219
rect 25292 10019 25372 10219
rect 25476 10019 25556 10219
rect 29150 10019 29230 10219
rect 29334 10019 29414 10219
rect 29518 10019 29598 10219
rect 886 7058 966 7258
rect 1070 7058 1150 7258
rect 1254 7058 1334 7258
rect 4898 7058 4978 7258
rect 5082 7058 5162 7258
rect 5266 7058 5346 7258
rect 8940 7058 9020 7258
rect 9124 7058 9204 7258
rect 9308 7058 9388 7258
rect 12982 7058 13062 7258
rect 13166 7058 13246 7258
rect 13350 7058 13430 7258
rect 17024 7058 17104 7258
rect 17208 7058 17288 7258
rect 17392 7058 17472 7258
rect 21066 7058 21146 7258
rect 21250 7058 21330 7258
rect 21434 7058 21514 7258
rect 25108 7058 25188 7258
rect 25292 7058 25372 7258
rect 25476 7058 25556 7258
rect 886 4853 966 5053
rect 1070 4853 1150 5053
rect 1254 4853 1334 5053
rect 2372 4853 2452 5053
rect 2556 4853 2636 5053
rect 2740 4853 2820 5053
rect 4898 4853 4978 5053
rect 5082 4853 5162 5053
rect 5266 4853 5346 5053
rect 6384 4853 6464 5053
rect 6568 4853 6648 5053
rect 6752 4853 6832 5053
rect 8940 4853 9020 5053
rect 9124 4853 9204 5053
rect 9308 4853 9388 5053
rect 10426 4853 10506 5053
rect 10610 4853 10690 5053
rect 10794 4853 10874 5053
rect 12982 4853 13062 5053
rect 13166 4853 13246 5053
rect 13350 4853 13430 5053
rect 14468 4853 14548 5053
rect 14652 4853 14732 5053
rect 14836 4853 14916 5053
rect 17024 4853 17104 5053
rect 17208 4853 17288 5053
rect 17392 4853 17472 5053
rect 18510 4853 18590 5053
rect 18694 4853 18774 5053
rect 18878 4853 18958 5053
rect 21066 4853 21146 5053
rect 21250 4853 21330 5053
rect 21434 4853 21514 5053
rect 22552 4853 22632 5053
rect 22736 4853 22816 5053
rect 22920 4853 23000 5053
rect 25108 4853 25188 5053
rect 25292 4853 25372 5053
rect 25476 4853 25556 5053
rect 26594 4853 26674 5053
rect 26778 4853 26858 5053
rect 26962 4853 27042 5053
rect 886 2648 966 2848
rect 1070 2648 1150 2848
rect 1254 2648 1334 2848
rect 2372 2649 2452 2849
rect 2556 2649 2636 2849
rect 2740 2649 2820 2849
rect 4898 2648 4978 2848
rect 5082 2648 5162 2848
rect 5266 2648 5346 2848
rect 6384 2649 6464 2849
rect 6568 2649 6648 2849
rect 6752 2649 6832 2849
rect 8940 2648 9020 2848
rect 9124 2648 9204 2848
rect 9308 2648 9388 2848
rect 10426 2649 10506 2849
rect 10610 2649 10690 2849
rect 10794 2649 10874 2849
rect 12982 2648 13062 2848
rect 13166 2648 13246 2848
rect 13350 2648 13430 2848
rect 14468 2649 14548 2849
rect 14652 2649 14732 2849
rect 14836 2649 14916 2849
rect 17024 2648 17104 2848
rect 17208 2648 17288 2848
rect 17392 2648 17472 2848
rect 18510 2649 18590 2849
rect 18694 2649 18774 2849
rect 18878 2649 18958 2849
rect 21066 2648 21146 2848
rect 21250 2648 21330 2848
rect 21434 2648 21514 2848
rect 22552 2649 22632 2849
rect 22736 2649 22816 2849
rect 22920 2649 23000 2849
rect 25108 2648 25188 2848
rect 25292 2648 25372 2848
rect 25476 2648 25556 2848
rect 26594 2649 26674 2849
rect 26778 2649 26858 2849
rect 26962 2649 27042 2849
rect 886 443 966 643
rect 1070 443 1150 643
rect 1254 443 1334 643
rect 4898 443 4978 643
rect 5082 443 5162 643
rect 5266 443 5346 643
rect 8940 443 9020 643
rect 9124 443 9204 643
rect 9308 443 9388 643
rect 12982 443 13062 643
rect 13166 443 13246 643
rect 13350 443 13430 643
rect 17024 443 17104 643
rect 17208 443 17288 643
rect 17392 443 17472 643
rect 21066 443 21146 643
rect 21250 443 21330 643
rect 21434 443 21514 643
rect 25108 443 25188 643
rect 25292 443 25372 643
rect 25476 443 25556 643
<< pmos >>
rect 4898 17497 4978 17997
rect 5082 17497 5162 17997
rect 5266 17497 5346 17997
rect 8940 17494 9020 17994
rect 9124 17494 9204 17994
rect 9308 17494 9388 17994
rect 12982 17494 13062 17994
rect 13166 17494 13246 17994
rect 13350 17494 13430 17994
rect 17024 17494 17104 17994
rect 17208 17494 17288 17994
rect 17392 17494 17472 17994
rect 21066 17494 21146 17994
rect 21250 17494 21330 17994
rect 21434 17494 21514 17994
rect 25108 17494 25188 17994
rect 25292 17494 25372 17994
rect 25476 17494 25556 17994
rect 29150 17494 29230 17994
rect 29334 17494 29414 17994
rect 29518 17494 29598 17994
rect 4898 15292 4978 15792
rect 5082 15292 5162 15792
rect 5266 15292 5346 15792
rect 6384 15292 6464 15792
rect 6568 15292 6648 15792
rect 6752 15292 6832 15792
rect 8940 15289 9020 15789
rect 9124 15289 9204 15789
rect 9308 15289 9388 15789
rect 10426 15289 10506 15789
rect 10610 15289 10690 15789
rect 10794 15289 10874 15789
rect 12982 15289 13062 15789
rect 13166 15289 13246 15789
rect 13350 15289 13430 15789
rect 14468 15289 14548 15789
rect 14652 15289 14732 15789
rect 14836 15289 14916 15789
rect 17024 15289 17104 15789
rect 17208 15289 17288 15789
rect 17392 15289 17472 15789
rect 18510 15289 18590 15789
rect 18694 15289 18774 15789
rect 18878 15289 18958 15789
rect 21066 15289 21146 15789
rect 21250 15289 21330 15789
rect 21434 15289 21514 15789
rect 22552 15289 22632 15789
rect 22736 15289 22816 15789
rect 22920 15289 23000 15789
rect 25108 15289 25188 15789
rect 25292 15289 25372 15789
rect 25476 15289 25556 15789
rect 26594 15289 26674 15789
rect 26778 15289 26858 15789
rect 26962 15289 27042 15789
rect 29150 15289 29230 15789
rect 29334 15289 29414 15789
rect 29518 15289 29598 15789
rect 30636 15289 30716 15789
rect 30820 15289 30900 15789
rect 31004 15289 31084 15789
rect 4898 13087 4978 13587
rect 5082 13087 5162 13587
rect 5266 13087 5346 13587
rect 6384 13088 6464 13588
rect 6568 13088 6648 13588
rect 6752 13088 6832 13588
rect 8940 13084 9020 13584
rect 9124 13084 9204 13584
rect 9308 13084 9388 13584
rect 10426 13085 10506 13585
rect 10610 13085 10690 13585
rect 10794 13085 10874 13585
rect 12982 13084 13062 13584
rect 13166 13084 13246 13584
rect 13350 13084 13430 13584
rect 14468 13085 14548 13585
rect 14652 13085 14732 13585
rect 14836 13085 14916 13585
rect 17024 13084 17104 13584
rect 17208 13084 17288 13584
rect 17392 13084 17472 13584
rect 18510 13085 18590 13585
rect 18694 13085 18774 13585
rect 18878 13085 18958 13585
rect 21066 13084 21146 13584
rect 21250 13084 21330 13584
rect 21434 13084 21514 13584
rect 22552 13085 22632 13585
rect 22736 13085 22816 13585
rect 22920 13085 23000 13585
rect 25108 13084 25188 13584
rect 25292 13084 25372 13584
rect 25476 13084 25556 13584
rect 26594 13085 26674 13585
rect 26778 13085 26858 13585
rect 26962 13085 27042 13585
rect 29150 13084 29230 13584
rect 29334 13084 29414 13584
rect 29518 13084 29598 13584
rect 30636 13085 30716 13585
rect 30820 13085 30900 13585
rect 31004 13085 31084 13585
rect 4898 10882 4978 11382
rect 5082 10882 5162 11382
rect 5266 10882 5346 11382
rect 8940 10879 9020 11379
rect 9124 10879 9204 11379
rect 9308 10879 9388 11379
rect 12982 10879 13062 11379
rect 13166 10879 13246 11379
rect 13350 10879 13430 11379
rect 17024 10879 17104 11379
rect 17208 10879 17288 11379
rect 17392 10879 17472 11379
rect 21066 10879 21146 11379
rect 21250 10879 21330 11379
rect 21434 10879 21514 11379
rect 25108 10879 25188 11379
rect 25292 10879 25372 11379
rect 25476 10879 25556 11379
rect 29150 10879 29230 11379
rect 29334 10879 29414 11379
rect 29518 10879 29598 11379
rect 886 7918 966 8418
rect 1070 7918 1150 8418
rect 1254 7918 1334 8418
rect 4898 7918 4978 8418
rect 5082 7918 5162 8418
rect 5266 7918 5346 8418
rect 8940 7918 9020 8418
rect 9124 7918 9204 8418
rect 9308 7918 9388 8418
rect 12982 7918 13062 8418
rect 13166 7918 13246 8418
rect 13350 7918 13430 8418
rect 17024 7918 17104 8418
rect 17208 7918 17288 8418
rect 17392 7918 17472 8418
rect 21066 7918 21146 8418
rect 21250 7918 21330 8418
rect 21434 7918 21514 8418
rect 25108 7918 25188 8418
rect 25292 7918 25372 8418
rect 25476 7918 25556 8418
rect 886 5713 966 6213
rect 1070 5713 1150 6213
rect 1254 5713 1334 6213
rect 2372 5713 2452 6213
rect 2556 5713 2636 6213
rect 2740 5713 2820 6213
rect 4898 5713 4978 6213
rect 5082 5713 5162 6213
rect 5266 5713 5346 6213
rect 6384 5713 6464 6213
rect 6568 5713 6648 6213
rect 6752 5713 6832 6213
rect 8940 5713 9020 6213
rect 9124 5713 9204 6213
rect 9308 5713 9388 6213
rect 10426 5713 10506 6213
rect 10610 5713 10690 6213
rect 10794 5713 10874 6213
rect 12982 5713 13062 6213
rect 13166 5713 13246 6213
rect 13350 5713 13430 6213
rect 14468 5713 14548 6213
rect 14652 5713 14732 6213
rect 14836 5713 14916 6213
rect 17024 5713 17104 6213
rect 17208 5713 17288 6213
rect 17392 5713 17472 6213
rect 18510 5713 18590 6213
rect 18694 5713 18774 6213
rect 18878 5713 18958 6213
rect 21066 5713 21146 6213
rect 21250 5713 21330 6213
rect 21434 5713 21514 6213
rect 22552 5713 22632 6213
rect 22736 5713 22816 6213
rect 22920 5713 23000 6213
rect 25108 5713 25188 6213
rect 25292 5713 25372 6213
rect 25476 5713 25556 6213
rect 26594 5713 26674 6213
rect 26778 5713 26858 6213
rect 26962 5713 27042 6213
rect 886 3508 966 4008
rect 1070 3508 1150 4008
rect 1254 3508 1334 4008
rect 2372 3509 2452 4009
rect 2556 3509 2636 4009
rect 2740 3509 2820 4009
rect 4898 3508 4978 4008
rect 5082 3508 5162 4008
rect 5266 3508 5346 4008
rect 6384 3509 6464 4009
rect 6568 3509 6648 4009
rect 6752 3509 6832 4009
rect 8940 3508 9020 4008
rect 9124 3508 9204 4008
rect 9308 3508 9388 4008
rect 10426 3509 10506 4009
rect 10610 3509 10690 4009
rect 10794 3509 10874 4009
rect 12982 3508 13062 4008
rect 13166 3508 13246 4008
rect 13350 3508 13430 4008
rect 14468 3509 14548 4009
rect 14652 3509 14732 4009
rect 14836 3509 14916 4009
rect 17024 3508 17104 4008
rect 17208 3508 17288 4008
rect 17392 3508 17472 4008
rect 18510 3509 18590 4009
rect 18694 3509 18774 4009
rect 18878 3509 18958 4009
rect 21066 3508 21146 4008
rect 21250 3508 21330 4008
rect 21434 3508 21514 4008
rect 22552 3509 22632 4009
rect 22736 3509 22816 4009
rect 22920 3509 23000 4009
rect 25108 3508 25188 4008
rect 25292 3508 25372 4008
rect 25476 3508 25556 4008
rect 26594 3509 26674 4009
rect 26778 3509 26858 4009
rect 26962 3509 27042 4009
rect 886 1303 966 1803
rect 1070 1303 1150 1803
rect 1254 1303 1334 1803
rect 4898 1303 4978 1803
rect 5082 1303 5162 1803
rect 5266 1303 5346 1803
rect 8940 1303 9020 1803
rect 9124 1303 9204 1803
rect 9308 1303 9388 1803
rect 12982 1303 13062 1803
rect 13166 1303 13246 1803
rect 13350 1303 13430 1803
rect 17024 1303 17104 1803
rect 17208 1303 17288 1803
rect 17392 1303 17472 1803
rect 21066 1303 21146 1803
rect 21250 1303 21330 1803
rect 21434 1303 21514 1803
rect 25108 1303 25188 1803
rect 25292 1303 25372 1803
rect 25476 1303 25556 1803
<< ndiff >>
rect 4810 16824 4898 16837
rect 4810 16650 4823 16824
rect 4869 16650 4898 16824
rect 4810 16637 4898 16650
rect 4978 16824 5082 16837
rect 4978 16650 5007 16824
rect 5053 16650 5082 16824
rect 4978 16637 5082 16650
rect 5162 16824 5266 16837
rect 5162 16650 5191 16824
rect 5237 16650 5266 16824
rect 5162 16637 5266 16650
rect 5346 16824 5434 16837
rect 5346 16650 5375 16824
rect 5421 16650 5434 16824
rect 5346 16637 5434 16650
rect 8852 16821 8940 16834
rect 8852 16647 8865 16821
rect 8911 16647 8940 16821
rect 8852 16634 8940 16647
rect 9020 16821 9124 16834
rect 9020 16647 9049 16821
rect 9095 16647 9124 16821
rect 9020 16634 9124 16647
rect 9204 16821 9308 16834
rect 9204 16647 9233 16821
rect 9279 16647 9308 16821
rect 9204 16634 9308 16647
rect 9388 16821 9476 16834
rect 9388 16647 9417 16821
rect 9463 16647 9476 16821
rect 9388 16634 9476 16647
rect 12894 16821 12982 16834
rect 12894 16647 12907 16821
rect 12953 16647 12982 16821
rect 12894 16634 12982 16647
rect 13062 16821 13166 16834
rect 13062 16647 13091 16821
rect 13137 16647 13166 16821
rect 13062 16634 13166 16647
rect 13246 16821 13350 16834
rect 13246 16647 13275 16821
rect 13321 16647 13350 16821
rect 13246 16634 13350 16647
rect 13430 16821 13518 16834
rect 13430 16647 13459 16821
rect 13505 16647 13518 16821
rect 13430 16634 13518 16647
rect 16936 16821 17024 16834
rect 16936 16647 16949 16821
rect 16995 16647 17024 16821
rect 16936 16634 17024 16647
rect 17104 16821 17208 16834
rect 17104 16647 17133 16821
rect 17179 16647 17208 16821
rect 17104 16634 17208 16647
rect 17288 16821 17392 16834
rect 17288 16647 17317 16821
rect 17363 16647 17392 16821
rect 17288 16634 17392 16647
rect 17472 16821 17560 16834
rect 17472 16647 17501 16821
rect 17547 16647 17560 16821
rect 17472 16634 17560 16647
rect 20978 16821 21066 16834
rect 20978 16647 20991 16821
rect 21037 16647 21066 16821
rect 20978 16634 21066 16647
rect 21146 16821 21250 16834
rect 21146 16647 21175 16821
rect 21221 16647 21250 16821
rect 21146 16634 21250 16647
rect 21330 16821 21434 16834
rect 21330 16647 21359 16821
rect 21405 16647 21434 16821
rect 21330 16634 21434 16647
rect 21514 16821 21602 16834
rect 21514 16647 21543 16821
rect 21589 16647 21602 16821
rect 21514 16634 21602 16647
rect 25020 16821 25108 16834
rect 25020 16647 25033 16821
rect 25079 16647 25108 16821
rect 25020 16634 25108 16647
rect 25188 16821 25292 16834
rect 25188 16647 25217 16821
rect 25263 16647 25292 16821
rect 25188 16634 25292 16647
rect 25372 16821 25476 16834
rect 25372 16647 25401 16821
rect 25447 16647 25476 16821
rect 25372 16634 25476 16647
rect 25556 16821 25644 16834
rect 25556 16647 25585 16821
rect 25631 16647 25644 16821
rect 25556 16634 25644 16647
rect 29062 16821 29150 16834
rect 29062 16647 29075 16821
rect 29121 16647 29150 16821
rect 29062 16634 29150 16647
rect 29230 16821 29334 16834
rect 29230 16647 29259 16821
rect 29305 16647 29334 16821
rect 29230 16634 29334 16647
rect 29414 16821 29518 16834
rect 29414 16647 29443 16821
rect 29489 16647 29518 16821
rect 29414 16634 29518 16647
rect 29598 16821 29686 16834
rect 29598 16647 29627 16821
rect 29673 16647 29686 16821
rect 29598 16634 29686 16647
rect 4810 14619 4898 14632
rect 4810 14445 4823 14619
rect 4869 14445 4898 14619
rect 4810 14432 4898 14445
rect 4978 14619 5082 14632
rect 4978 14445 5007 14619
rect 5053 14445 5082 14619
rect 4978 14432 5082 14445
rect 5162 14619 5266 14632
rect 5162 14445 5191 14619
rect 5237 14445 5266 14619
rect 5162 14432 5266 14445
rect 5346 14619 5434 14632
rect 5346 14445 5375 14619
rect 5421 14445 5434 14619
rect 5346 14432 5434 14445
rect 6296 14619 6384 14632
rect 6296 14445 6309 14619
rect 6355 14445 6384 14619
rect 6296 14432 6384 14445
rect 6464 14619 6568 14632
rect 6464 14445 6493 14619
rect 6539 14445 6568 14619
rect 6464 14432 6568 14445
rect 6648 14619 6752 14632
rect 6648 14445 6677 14619
rect 6723 14445 6752 14619
rect 6648 14432 6752 14445
rect 6832 14619 6920 14632
rect 6832 14445 6861 14619
rect 6907 14445 6920 14619
rect 6832 14432 6920 14445
rect 8852 14616 8940 14629
rect 8852 14442 8865 14616
rect 8911 14442 8940 14616
rect 8852 14429 8940 14442
rect 9020 14616 9124 14629
rect 9020 14442 9049 14616
rect 9095 14442 9124 14616
rect 9020 14429 9124 14442
rect 9204 14616 9308 14629
rect 9204 14442 9233 14616
rect 9279 14442 9308 14616
rect 9204 14429 9308 14442
rect 9388 14616 9476 14629
rect 9388 14442 9417 14616
rect 9463 14442 9476 14616
rect 9388 14429 9476 14442
rect 10338 14616 10426 14629
rect 10338 14442 10351 14616
rect 10397 14442 10426 14616
rect 10338 14429 10426 14442
rect 10506 14616 10610 14629
rect 10506 14442 10535 14616
rect 10581 14442 10610 14616
rect 10506 14429 10610 14442
rect 10690 14616 10794 14629
rect 10690 14442 10719 14616
rect 10765 14442 10794 14616
rect 10690 14429 10794 14442
rect 10874 14616 10962 14629
rect 10874 14442 10903 14616
rect 10949 14442 10962 14616
rect 10874 14429 10962 14442
rect 12894 14616 12982 14629
rect 12894 14442 12907 14616
rect 12953 14442 12982 14616
rect 12894 14429 12982 14442
rect 13062 14616 13166 14629
rect 13062 14442 13091 14616
rect 13137 14442 13166 14616
rect 13062 14429 13166 14442
rect 13246 14616 13350 14629
rect 13246 14442 13275 14616
rect 13321 14442 13350 14616
rect 13246 14429 13350 14442
rect 13430 14616 13518 14629
rect 13430 14442 13459 14616
rect 13505 14442 13518 14616
rect 13430 14429 13518 14442
rect 14380 14616 14468 14629
rect 14380 14442 14393 14616
rect 14439 14442 14468 14616
rect 14380 14429 14468 14442
rect 14548 14616 14652 14629
rect 14548 14442 14577 14616
rect 14623 14442 14652 14616
rect 14548 14429 14652 14442
rect 14732 14616 14836 14629
rect 14732 14442 14761 14616
rect 14807 14442 14836 14616
rect 14732 14429 14836 14442
rect 14916 14616 15004 14629
rect 14916 14442 14945 14616
rect 14991 14442 15004 14616
rect 14916 14429 15004 14442
rect 16936 14616 17024 14629
rect 16936 14442 16949 14616
rect 16995 14442 17024 14616
rect 16936 14429 17024 14442
rect 17104 14616 17208 14629
rect 17104 14442 17133 14616
rect 17179 14442 17208 14616
rect 17104 14429 17208 14442
rect 17288 14616 17392 14629
rect 17288 14442 17317 14616
rect 17363 14442 17392 14616
rect 17288 14429 17392 14442
rect 17472 14616 17560 14629
rect 17472 14442 17501 14616
rect 17547 14442 17560 14616
rect 17472 14429 17560 14442
rect 18422 14616 18510 14629
rect 18422 14442 18435 14616
rect 18481 14442 18510 14616
rect 18422 14429 18510 14442
rect 18590 14616 18694 14629
rect 18590 14442 18619 14616
rect 18665 14442 18694 14616
rect 18590 14429 18694 14442
rect 18774 14616 18878 14629
rect 18774 14442 18803 14616
rect 18849 14442 18878 14616
rect 18774 14429 18878 14442
rect 18958 14616 19046 14629
rect 18958 14442 18987 14616
rect 19033 14442 19046 14616
rect 18958 14429 19046 14442
rect 20978 14616 21066 14629
rect 20978 14442 20991 14616
rect 21037 14442 21066 14616
rect 20978 14429 21066 14442
rect 21146 14616 21250 14629
rect 21146 14442 21175 14616
rect 21221 14442 21250 14616
rect 21146 14429 21250 14442
rect 21330 14616 21434 14629
rect 21330 14442 21359 14616
rect 21405 14442 21434 14616
rect 21330 14429 21434 14442
rect 21514 14616 21602 14629
rect 21514 14442 21543 14616
rect 21589 14442 21602 14616
rect 21514 14429 21602 14442
rect 22464 14616 22552 14629
rect 22464 14442 22477 14616
rect 22523 14442 22552 14616
rect 22464 14429 22552 14442
rect 22632 14616 22736 14629
rect 22632 14442 22661 14616
rect 22707 14442 22736 14616
rect 22632 14429 22736 14442
rect 22816 14616 22920 14629
rect 22816 14442 22845 14616
rect 22891 14442 22920 14616
rect 22816 14429 22920 14442
rect 23000 14616 23088 14629
rect 23000 14442 23029 14616
rect 23075 14442 23088 14616
rect 23000 14429 23088 14442
rect 25020 14616 25108 14629
rect 25020 14442 25033 14616
rect 25079 14442 25108 14616
rect 25020 14429 25108 14442
rect 25188 14616 25292 14629
rect 25188 14442 25217 14616
rect 25263 14442 25292 14616
rect 25188 14429 25292 14442
rect 25372 14616 25476 14629
rect 25372 14442 25401 14616
rect 25447 14442 25476 14616
rect 25372 14429 25476 14442
rect 25556 14616 25644 14629
rect 25556 14442 25585 14616
rect 25631 14442 25644 14616
rect 25556 14429 25644 14442
rect 26506 14616 26594 14629
rect 26506 14442 26519 14616
rect 26565 14442 26594 14616
rect 26506 14429 26594 14442
rect 26674 14616 26778 14629
rect 26674 14442 26703 14616
rect 26749 14442 26778 14616
rect 26674 14429 26778 14442
rect 26858 14616 26962 14629
rect 26858 14442 26887 14616
rect 26933 14442 26962 14616
rect 26858 14429 26962 14442
rect 27042 14616 27130 14629
rect 27042 14442 27071 14616
rect 27117 14442 27130 14616
rect 27042 14429 27130 14442
rect 29062 14616 29150 14629
rect 29062 14442 29075 14616
rect 29121 14442 29150 14616
rect 29062 14429 29150 14442
rect 29230 14616 29334 14629
rect 29230 14442 29259 14616
rect 29305 14442 29334 14616
rect 29230 14429 29334 14442
rect 29414 14616 29518 14629
rect 29414 14442 29443 14616
rect 29489 14442 29518 14616
rect 29414 14429 29518 14442
rect 29598 14616 29686 14629
rect 29598 14442 29627 14616
rect 29673 14442 29686 14616
rect 29598 14429 29686 14442
rect 30548 14616 30636 14629
rect 30548 14442 30561 14616
rect 30607 14442 30636 14616
rect 30548 14429 30636 14442
rect 30716 14616 30820 14629
rect 30716 14442 30745 14616
rect 30791 14442 30820 14616
rect 30716 14429 30820 14442
rect 30900 14616 31004 14629
rect 30900 14442 30929 14616
rect 30975 14442 31004 14616
rect 30900 14429 31004 14442
rect 31084 14616 31172 14629
rect 31084 14442 31113 14616
rect 31159 14442 31172 14616
rect 31084 14429 31172 14442
rect 4810 12414 4898 12427
rect 4810 12240 4823 12414
rect 4869 12240 4898 12414
rect 4810 12227 4898 12240
rect 4978 12414 5082 12427
rect 4978 12240 5007 12414
rect 5053 12240 5082 12414
rect 4978 12227 5082 12240
rect 5162 12414 5266 12427
rect 5162 12240 5191 12414
rect 5237 12240 5266 12414
rect 5162 12227 5266 12240
rect 5346 12414 5434 12427
rect 5346 12240 5375 12414
rect 5421 12240 5434 12414
rect 5346 12227 5434 12240
rect 6296 12415 6384 12428
rect 6296 12241 6309 12415
rect 6355 12241 6384 12415
rect 6296 12228 6384 12241
rect 6464 12415 6568 12428
rect 6464 12241 6493 12415
rect 6539 12241 6568 12415
rect 6464 12228 6568 12241
rect 6648 12415 6752 12428
rect 6648 12241 6677 12415
rect 6723 12241 6752 12415
rect 6648 12228 6752 12241
rect 6832 12415 6920 12428
rect 6832 12241 6861 12415
rect 6907 12241 6920 12415
rect 6832 12228 6920 12241
rect 8852 12411 8940 12424
rect 8852 12237 8865 12411
rect 8911 12237 8940 12411
rect 8852 12224 8940 12237
rect 9020 12411 9124 12424
rect 9020 12237 9049 12411
rect 9095 12237 9124 12411
rect 9020 12224 9124 12237
rect 9204 12411 9308 12424
rect 9204 12237 9233 12411
rect 9279 12237 9308 12411
rect 9204 12224 9308 12237
rect 9388 12411 9476 12424
rect 9388 12237 9417 12411
rect 9463 12237 9476 12411
rect 9388 12224 9476 12237
rect 10338 12412 10426 12425
rect 10338 12238 10351 12412
rect 10397 12238 10426 12412
rect 10338 12225 10426 12238
rect 10506 12412 10610 12425
rect 10506 12238 10535 12412
rect 10581 12238 10610 12412
rect 10506 12225 10610 12238
rect 10690 12412 10794 12425
rect 10690 12238 10719 12412
rect 10765 12238 10794 12412
rect 10690 12225 10794 12238
rect 10874 12412 10962 12425
rect 10874 12238 10903 12412
rect 10949 12238 10962 12412
rect 10874 12225 10962 12238
rect 12894 12411 12982 12424
rect 12894 12237 12907 12411
rect 12953 12237 12982 12411
rect 12894 12224 12982 12237
rect 13062 12411 13166 12424
rect 13062 12237 13091 12411
rect 13137 12237 13166 12411
rect 13062 12224 13166 12237
rect 13246 12411 13350 12424
rect 13246 12237 13275 12411
rect 13321 12237 13350 12411
rect 13246 12224 13350 12237
rect 13430 12411 13518 12424
rect 13430 12237 13459 12411
rect 13505 12237 13518 12411
rect 13430 12224 13518 12237
rect 14380 12412 14468 12425
rect 14380 12238 14393 12412
rect 14439 12238 14468 12412
rect 14380 12225 14468 12238
rect 14548 12412 14652 12425
rect 14548 12238 14577 12412
rect 14623 12238 14652 12412
rect 14548 12225 14652 12238
rect 14732 12412 14836 12425
rect 14732 12238 14761 12412
rect 14807 12238 14836 12412
rect 14732 12225 14836 12238
rect 14916 12412 15004 12425
rect 14916 12238 14945 12412
rect 14991 12238 15004 12412
rect 14916 12225 15004 12238
rect 16936 12411 17024 12424
rect 16936 12237 16949 12411
rect 16995 12237 17024 12411
rect 16936 12224 17024 12237
rect 17104 12411 17208 12424
rect 17104 12237 17133 12411
rect 17179 12237 17208 12411
rect 17104 12224 17208 12237
rect 17288 12411 17392 12424
rect 17288 12237 17317 12411
rect 17363 12237 17392 12411
rect 17288 12224 17392 12237
rect 17472 12411 17560 12424
rect 17472 12237 17501 12411
rect 17547 12237 17560 12411
rect 17472 12224 17560 12237
rect 18422 12412 18510 12425
rect 18422 12238 18435 12412
rect 18481 12238 18510 12412
rect 18422 12225 18510 12238
rect 18590 12412 18694 12425
rect 18590 12238 18619 12412
rect 18665 12238 18694 12412
rect 18590 12225 18694 12238
rect 18774 12412 18878 12425
rect 18774 12238 18803 12412
rect 18849 12238 18878 12412
rect 18774 12225 18878 12238
rect 18958 12412 19046 12425
rect 18958 12238 18987 12412
rect 19033 12238 19046 12412
rect 18958 12225 19046 12238
rect 20978 12411 21066 12424
rect 20978 12237 20991 12411
rect 21037 12237 21066 12411
rect 20978 12224 21066 12237
rect 21146 12411 21250 12424
rect 21146 12237 21175 12411
rect 21221 12237 21250 12411
rect 21146 12224 21250 12237
rect 21330 12411 21434 12424
rect 21330 12237 21359 12411
rect 21405 12237 21434 12411
rect 21330 12224 21434 12237
rect 21514 12411 21602 12424
rect 21514 12237 21543 12411
rect 21589 12237 21602 12411
rect 21514 12224 21602 12237
rect 22464 12412 22552 12425
rect 22464 12238 22477 12412
rect 22523 12238 22552 12412
rect 22464 12225 22552 12238
rect 22632 12412 22736 12425
rect 22632 12238 22661 12412
rect 22707 12238 22736 12412
rect 22632 12225 22736 12238
rect 22816 12412 22920 12425
rect 22816 12238 22845 12412
rect 22891 12238 22920 12412
rect 22816 12225 22920 12238
rect 23000 12412 23088 12425
rect 23000 12238 23029 12412
rect 23075 12238 23088 12412
rect 23000 12225 23088 12238
rect 25020 12411 25108 12424
rect 25020 12237 25033 12411
rect 25079 12237 25108 12411
rect 25020 12224 25108 12237
rect 25188 12411 25292 12424
rect 25188 12237 25217 12411
rect 25263 12237 25292 12411
rect 25188 12224 25292 12237
rect 25372 12411 25476 12424
rect 25372 12237 25401 12411
rect 25447 12237 25476 12411
rect 25372 12224 25476 12237
rect 25556 12411 25644 12424
rect 25556 12237 25585 12411
rect 25631 12237 25644 12411
rect 25556 12224 25644 12237
rect 26506 12412 26594 12425
rect 26506 12238 26519 12412
rect 26565 12238 26594 12412
rect 26506 12225 26594 12238
rect 26674 12412 26778 12425
rect 26674 12238 26703 12412
rect 26749 12238 26778 12412
rect 26674 12225 26778 12238
rect 26858 12412 26962 12425
rect 26858 12238 26887 12412
rect 26933 12238 26962 12412
rect 26858 12225 26962 12238
rect 27042 12412 27130 12425
rect 27042 12238 27071 12412
rect 27117 12238 27130 12412
rect 27042 12225 27130 12238
rect 29062 12411 29150 12424
rect 29062 12237 29075 12411
rect 29121 12237 29150 12411
rect 29062 12224 29150 12237
rect 29230 12411 29334 12424
rect 29230 12237 29259 12411
rect 29305 12237 29334 12411
rect 29230 12224 29334 12237
rect 29414 12411 29518 12424
rect 29414 12237 29443 12411
rect 29489 12237 29518 12411
rect 29414 12224 29518 12237
rect 29598 12411 29686 12424
rect 29598 12237 29627 12411
rect 29673 12237 29686 12411
rect 29598 12224 29686 12237
rect 30548 12412 30636 12425
rect 30548 12238 30561 12412
rect 30607 12238 30636 12412
rect 30548 12225 30636 12238
rect 30716 12412 30820 12425
rect 30716 12238 30745 12412
rect 30791 12238 30820 12412
rect 30716 12225 30820 12238
rect 30900 12412 31004 12425
rect 30900 12238 30929 12412
rect 30975 12238 31004 12412
rect 30900 12225 31004 12238
rect 31084 12412 31172 12425
rect 31084 12238 31113 12412
rect 31159 12238 31172 12412
rect 31084 12225 31172 12238
rect 4810 10209 4898 10222
rect 4810 10035 4823 10209
rect 4869 10035 4898 10209
rect 4810 10022 4898 10035
rect 4978 10209 5082 10222
rect 4978 10035 5007 10209
rect 5053 10035 5082 10209
rect 4978 10022 5082 10035
rect 5162 10209 5266 10222
rect 5162 10035 5191 10209
rect 5237 10035 5266 10209
rect 5162 10022 5266 10035
rect 5346 10209 5434 10222
rect 5346 10035 5375 10209
rect 5421 10035 5434 10209
rect 5346 10022 5434 10035
rect 8852 10206 8940 10219
rect 8852 10032 8865 10206
rect 8911 10032 8940 10206
rect 8852 10019 8940 10032
rect 9020 10206 9124 10219
rect 9020 10032 9049 10206
rect 9095 10032 9124 10206
rect 9020 10019 9124 10032
rect 9204 10206 9308 10219
rect 9204 10032 9233 10206
rect 9279 10032 9308 10206
rect 9204 10019 9308 10032
rect 9388 10206 9476 10219
rect 9388 10032 9417 10206
rect 9463 10032 9476 10206
rect 9388 10019 9476 10032
rect 12894 10206 12982 10219
rect 12894 10032 12907 10206
rect 12953 10032 12982 10206
rect 12894 10019 12982 10032
rect 13062 10206 13166 10219
rect 13062 10032 13091 10206
rect 13137 10032 13166 10206
rect 13062 10019 13166 10032
rect 13246 10206 13350 10219
rect 13246 10032 13275 10206
rect 13321 10032 13350 10206
rect 13246 10019 13350 10032
rect 13430 10206 13518 10219
rect 13430 10032 13459 10206
rect 13505 10032 13518 10206
rect 13430 10019 13518 10032
rect 16936 10206 17024 10219
rect 16936 10032 16949 10206
rect 16995 10032 17024 10206
rect 16936 10019 17024 10032
rect 17104 10206 17208 10219
rect 17104 10032 17133 10206
rect 17179 10032 17208 10206
rect 17104 10019 17208 10032
rect 17288 10206 17392 10219
rect 17288 10032 17317 10206
rect 17363 10032 17392 10206
rect 17288 10019 17392 10032
rect 17472 10206 17560 10219
rect 17472 10032 17501 10206
rect 17547 10032 17560 10206
rect 17472 10019 17560 10032
rect 20978 10206 21066 10219
rect 20978 10032 20991 10206
rect 21037 10032 21066 10206
rect 20978 10019 21066 10032
rect 21146 10206 21250 10219
rect 21146 10032 21175 10206
rect 21221 10032 21250 10206
rect 21146 10019 21250 10032
rect 21330 10206 21434 10219
rect 21330 10032 21359 10206
rect 21405 10032 21434 10206
rect 21330 10019 21434 10032
rect 21514 10206 21602 10219
rect 21514 10032 21543 10206
rect 21589 10032 21602 10206
rect 21514 10019 21602 10032
rect 25020 10206 25108 10219
rect 25020 10032 25033 10206
rect 25079 10032 25108 10206
rect 25020 10019 25108 10032
rect 25188 10206 25292 10219
rect 25188 10032 25217 10206
rect 25263 10032 25292 10206
rect 25188 10019 25292 10032
rect 25372 10206 25476 10219
rect 25372 10032 25401 10206
rect 25447 10032 25476 10206
rect 25372 10019 25476 10032
rect 25556 10206 25644 10219
rect 25556 10032 25585 10206
rect 25631 10032 25644 10206
rect 25556 10019 25644 10032
rect 29062 10206 29150 10219
rect 29062 10032 29075 10206
rect 29121 10032 29150 10206
rect 29062 10019 29150 10032
rect 29230 10206 29334 10219
rect 29230 10032 29259 10206
rect 29305 10032 29334 10206
rect 29230 10019 29334 10032
rect 29414 10206 29518 10219
rect 29414 10032 29443 10206
rect 29489 10032 29518 10206
rect 29414 10019 29518 10032
rect 29598 10206 29686 10219
rect 29598 10032 29627 10206
rect 29673 10032 29686 10206
rect 29598 10019 29686 10032
rect 798 7245 886 7258
rect 798 7071 811 7245
rect 857 7071 886 7245
rect 798 7058 886 7071
rect 966 7245 1070 7258
rect 966 7071 995 7245
rect 1041 7071 1070 7245
rect 966 7058 1070 7071
rect 1150 7245 1254 7258
rect 1150 7071 1179 7245
rect 1225 7071 1254 7245
rect 1150 7058 1254 7071
rect 1334 7245 1422 7258
rect 1334 7071 1363 7245
rect 1409 7071 1422 7245
rect 1334 7058 1422 7071
rect 4810 7245 4898 7258
rect 4810 7071 4823 7245
rect 4869 7071 4898 7245
rect 4810 7058 4898 7071
rect 4978 7245 5082 7258
rect 4978 7071 5007 7245
rect 5053 7071 5082 7245
rect 4978 7058 5082 7071
rect 5162 7245 5266 7258
rect 5162 7071 5191 7245
rect 5237 7071 5266 7245
rect 5162 7058 5266 7071
rect 5346 7245 5434 7258
rect 5346 7071 5375 7245
rect 5421 7071 5434 7245
rect 5346 7058 5434 7071
rect 8852 7245 8940 7258
rect 8852 7071 8865 7245
rect 8911 7071 8940 7245
rect 8852 7058 8940 7071
rect 9020 7245 9124 7258
rect 9020 7071 9049 7245
rect 9095 7071 9124 7245
rect 9020 7058 9124 7071
rect 9204 7245 9308 7258
rect 9204 7071 9233 7245
rect 9279 7071 9308 7245
rect 9204 7058 9308 7071
rect 9388 7245 9476 7258
rect 9388 7071 9417 7245
rect 9463 7071 9476 7245
rect 9388 7058 9476 7071
rect 12894 7245 12982 7258
rect 12894 7071 12907 7245
rect 12953 7071 12982 7245
rect 12894 7058 12982 7071
rect 13062 7245 13166 7258
rect 13062 7071 13091 7245
rect 13137 7071 13166 7245
rect 13062 7058 13166 7071
rect 13246 7245 13350 7258
rect 13246 7071 13275 7245
rect 13321 7071 13350 7245
rect 13246 7058 13350 7071
rect 13430 7245 13518 7258
rect 13430 7071 13459 7245
rect 13505 7071 13518 7245
rect 13430 7058 13518 7071
rect 16936 7245 17024 7258
rect 16936 7071 16949 7245
rect 16995 7071 17024 7245
rect 16936 7058 17024 7071
rect 17104 7245 17208 7258
rect 17104 7071 17133 7245
rect 17179 7071 17208 7245
rect 17104 7058 17208 7071
rect 17288 7245 17392 7258
rect 17288 7071 17317 7245
rect 17363 7071 17392 7245
rect 17288 7058 17392 7071
rect 17472 7245 17560 7258
rect 17472 7071 17501 7245
rect 17547 7071 17560 7245
rect 17472 7058 17560 7071
rect 20978 7245 21066 7258
rect 20978 7071 20991 7245
rect 21037 7071 21066 7245
rect 20978 7058 21066 7071
rect 21146 7245 21250 7258
rect 21146 7071 21175 7245
rect 21221 7071 21250 7245
rect 21146 7058 21250 7071
rect 21330 7245 21434 7258
rect 21330 7071 21359 7245
rect 21405 7071 21434 7245
rect 21330 7058 21434 7071
rect 21514 7245 21602 7258
rect 21514 7071 21543 7245
rect 21589 7071 21602 7245
rect 21514 7058 21602 7071
rect 25020 7245 25108 7258
rect 25020 7071 25033 7245
rect 25079 7071 25108 7245
rect 25020 7058 25108 7071
rect 25188 7245 25292 7258
rect 25188 7071 25217 7245
rect 25263 7071 25292 7245
rect 25188 7058 25292 7071
rect 25372 7245 25476 7258
rect 25372 7071 25401 7245
rect 25447 7071 25476 7245
rect 25372 7058 25476 7071
rect 25556 7245 25644 7258
rect 25556 7071 25585 7245
rect 25631 7071 25644 7245
rect 25556 7058 25644 7071
rect 798 5040 886 5053
rect 798 4866 811 5040
rect 857 4866 886 5040
rect 798 4853 886 4866
rect 966 5040 1070 5053
rect 966 4866 995 5040
rect 1041 4866 1070 5040
rect 966 4853 1070 4866
rect 1150 5040 1254 5053
rect 1150 4866 1179 5040
rect 1225 4866 1254 5040
rect 1150 4853 1254 4866
rect 1334 5040 1422 5053
rect 1334 4866 1363 5040
rect 1409 4866 1422 5040
rect 1334 4853 1422 4866
rect 2284 5040 2372 5053
rect 2284 4866 2297 5040
rect 2343 4866 2372 5040
rect 2284 4853 2372 4866
rect 2452 5040 2556 5053
rect 2452 4866 2481 5040
rect 2527 4866 2556 5040
rect 2452 4853 2556 4866
rect 2636 5040 2740 5053
rect 2636 4866 2665 5040
rect 2711 4866 2740 5040
rect 2636 4853 2740 4866
rect 2820 5040 2908 5053
rect 2820 4866 2849 5040
rect 2895 4866 2908 5040
rect 2820 4853 2908 4866
rect 4810 5040 4898 5053
rect 4810 4866 4823 5040
rect 4869 4866 4898 5040
rect 4810 4853 4898 4866
rect 4978 5040 5082 5053
rect 4978 4866 5007 5040
rect 5053 4866 5082 5040
rect 4978 4853 5082 4866
rect 5162 5040 5266 5053
rect 5162 4866 5191 5040
rect 5237 4866 5266 5040
rect 5162 4853 5266 4866
rect 5346 5040 5434 5053
rect 5346 4866 5375 5040
rect 5421 4866 5434 5040
rect 5346 4853 5434 4866
rect 6296 5040 6384 5053
rect 6296 4866 6309 5040
rect 6355 4866 6384 5040
rect 6296 4853 6384 4866
rect 6464 5040 6568 5053
rect 6464 4866 6493 5040
rect 6539 4866 6568 5040
rect 6464 4853 6568 4866
rect 6648 5040 6752 5053
rect 6648 4866 6677 5040
rect 6723 4866 6752 5040
rect 6648 4853 6752 4866
rect 6832 5040 6920 5053
rect 6832 4866 6861 5040
rect 6907 4866 6920 5040
rect 6832 4853 6920 4866
rect 8852 5040 8940 5053
rect 8852 4866 8865 5040
rect 8911 4866 8940 5040
rect 8852 4853 8940 4866
rect 9020 5040 9124 5053
rect 9020 4866 9049 5040
rect 9095 4866 9124 5040
rect 9020 4853 9124 4866
rect 9204 5040 9308 5053
rect 9204 4866 9233 5040
rect 9279 4866 9308 5040
rect 9204 4853 9308 4866
rect 9388 5040 9476 5053
rect 9388 4866 9417 5040
rect 9463 4866 9476 5040
rect 9388 4853 9476 4866
rect 10338 5040 10426 5053
rect 10338 4866 10351 5040
rect 10397 4866 10426 5040
rect 10338 4853 10426 4866
rect 10506 5040 10610 5053
rect 10506 4866 10535 5040
rect 10581 4866 10610 5040
rect 10506 4853 10610 4866
rect 10690 5040 10794 5053
rect 10690 4866 10719 5040
rect 10765 4866 10794 5040
rect 10690 4853 10794 4866
rect 10874 5040 10962 5053
rect 10874 4866 10903 5040
rect 10949 4866 10962 5040
rect 10874 4853 10962 4866
rect 12894 5040 12982 5053
rect 12894 4866 12907 5040
rect 12953 4866 12982 5040
rect 12894 4853 12982 4866
rect 13062 5040 13166 5053
rect 13062 4866 13091 5040
rect 13137 4866 13166 5040
rect 13062 4853 13166 4866
rect 13246 5040 13350 5053
rect 13246 4866 13275 5040
rect 13321 4866 13350 5040
rect 13246 4853 13350 4866
rect 13430 5040 13518 5053
rect 13430 4866 13459 5040
rect 13505 4866 13518 5040
rect 13430 4853 13518 4866
rect 14380 5040 14468 5053
rect 14380 4866 14393 5040
rect 14439 4866 14468 5040
rect 14380 4853 14468 4866
rect 14548 5040 14652 5053
rect 14548 4866 14577 5040
rect 14623 4866 14652 5040
rect 14548 4853 14652 4866
rect 14732 5040 14836 5053
rect 14732 4866 14761 5040
rect 14807 4866 14836 5040
rect 14732 4853 14836 4866
rect 14916 5040 15004 5053
rect 14916 4866 14945 5040
rect 14991 4866 15004 5040
rect 14916 4853 15004 4866
rect 16936 5040 17024 5053
rect 16936 4866 16949 5040
rect 16995 4866 17024 5040
rect 16936 4853 17024 4866
rect 17104 5040 17208 5053
rect 17104 4866 17133 5040
rect 17179 4866 17208 5040
rect 17104 4853 17208 4866
rect 17288 5040 17392 5053
rect 17288 4866 17317 5040
rect 17363 4866 17392 5040
rect 17288 4853 17392 4866
rect 17472 5040 17560 5053
rect 17472 4866 17501 5040
rect 17547 4866 17560 5040
rect 17472 4853 17560 4866
rect 18422 5040 18510 5053
rect 18422 4866 18435 5040
rect 18481 4866 18510 5040
rect 18422 4853 18510 4866
rect 18590 5040 18694 5053
rect 18590 4866 18619 5040
rect 18665 4866 18694 5040
rect 18590 4853 18694 4866
rect 18774 5040 18878 5053
rect 18774 4866 18803 5040
rect 18849 4866 18878 5040
rect 18774 4853 18878 4866
rect 18958 5040 19046 5053
rect 18958 4866 18987 5040
rect 19033 4866 19046 5040
rect 18958 4853 19046 4866
rect 20978 5040 21066 5053
rect 20978 4866 20991 5040
rect 21037 4866 21066 5040
rect 20978 4853 21066 4866
rect 21146 5040 21250 5053
rect 21146 4866 21175 5040
rect 21221 4866 21250 5040
rect 21146 4853 21250 4866
rect 21330 5040 21434 5053
rect 21330 4866 21359 5040
rect 21405 4866 21434 5040
rect 21330 4853 21434 4866
rect 21514 5040 21602 5053
rect 21514 4866 21543 5040
rect 21589 4866 21602 5040
rect 21514 4853 21602 4866
rect 22464 5040 22552 5053
rect 22464 4866 22477 5040
rect 22523 4866 22552 5040
rect 22464 4853 22552 4866
rect 22632 5040 22736 5053
rect 22632 4866 22661 5040
rect 22707 4866 22736 5040
rect 22632 4853 22736 4866
rect 22816 5040 22920 5053
rect 22816 4866 22845 5040
rect 22891 4866 22920 5040
rect 22816 4853 22920 4866
rect 23000 5040 23088 5053
rect 23000 4866 23029 5040
rect 23075 4866 23088 5040
rect 23000 4853 23088 4866
rect 25020 5040 25108 5053
rect 25020 4866 25033 5040
rect 25079 4866 25108 5040
rect 25020 4853 25108 4866
rect 25188 5040 25292 5053
rect 25188 4866 25217 5040
rect 25263 4866 25292 5040
rect 25188 4853 25292 4866
rect 25372 5040 25476 5053
rect 25372 4866 25401 5040
rect 25447 4866 25476 5040
rect 25372 4853 25476 4866
rect 25556 5040 25644 5053
rect 25556 4866 25585 5040
rect 25631 4866 25644 5040
rect 25556 4853 25644 4866
rect 26506 5040 26594 5053
rect 26506 4866 26519 5040
rect 26565 4866 26594 5040
rect 26506 4853 26594 4866
rect 26674 5040 26778 5053
rect 26674 4866 26703 5040
rect 26749 4866 26778 5040
rect 26674 4853 26778 4866
rect 26858 5040 26962 5053
rect 26858 4866 26887 5040
rect 26933 4866 26962 5040
rect 26858 4853 26962 4866
rect 27042 5040 27130 5053
rect 27042 4866 27071 5040
rect 27117 4866 27130 5040
rect 27042 4853 27130 4866
rect 798 2835 886 2848
rect 798 2661 811 2835
rect 857 2661 886 2835
rect 798 2648 886 2661
rect 966 2835 1070 2848
rect 966 2661 995 2835
rect 1041 2661 1070 2835
rect 966 2648 1070 2661
rect 1150 2835 1254 2848
rect 1150 2661 1179 2835
rect 1225 2661 1254 2835
rect 1150 2648 1254 2661
rect 1334 2835 1422 2848
rect 1334 2661 1363 2835
rect 1409 2661 1422 2835
rect 1334 2648 1422 2661
rect 2284 2836 2372 2849
rect 2284 2662 2297 2836
rect 2343 2662 2372 2836
rect 2284 2649 2372 2662
rect 2452 2836 2556 2849
rect 2452 2662 2481 2836
rect 2527 2662 2556 2836
rect 2452 2649 2556 2662
rect 2636 2836 2740 2849
rect 2636 2662 2665 2836
rect 2711 2662 2740 2836
rect 2636 2649 2740 2662
rect 2820 2836 2908 2849
rect 2820 2662 2849 2836
rect 2895 2662 2908 2836
rect 2820 2649 2908 2662
rect 4810 2835 4898 2848
rect 4810 2661 4823 2835
rect 4869 2661 4898 2835
rect 4810 2648 4898 2661
rect 4978 2835 5082 2848
rect 4978 2661 5007 2835
rect 5053 2661 5082 2835
rect 4978 2648 5082 2661
rect 5162 2835 5266 2848
rect 5162 2661 5191 2835
rect 5237 2661 5266 2835
rect 5162 2648 5266 2661
rect 5346 2835 5434 2848
rect 5346 2661 5375 2835
rect 5421 2661 5434 2835
rect 5346 2648 5434 2661
rect 6296 2836 6384 2849
rect 6296 2662 6309 2836
rect 6355 2662 6384 2836
rect 6296 2649 6384 2662
rect 6464 2836 6568 2849
rect 6464 2662 6493 2836
rect 6539 2662 6568 2836
rect 6464 2649 6568 2662
rect 6648 2836 6752 2849
rect 6648 2662 6677 2836
rect 6723 2662 6752 2836
rect 6648 2649 6752 2662
rect 6832 2836 6920 2849
rect 6832 2662 6861 2836
rect 6907 2662 6920 2836
rect 6832 2649 6920 2662
rect 8852 2835 8940 2848
rect 8852 2661 8865 2835
rect 8911 2661 8940 2835
rect 8852 2648 8940 2661
rect 9020 2835 9124 2848
rect 9020 2661 9049 2835
rect 9095 2661 9124 2835
rect 9020 2648 9124 2661
rect 9204 2835 9308 2848
rect 9204 2661 9233 2835
rect 9279 2661 9308 2835
rect 9204 2648 9308 2661
rect 9388 2835 9476 2848
rect 9388 2661 9417 2835
rect 9463 2661 9476 2835
rect 9388 2648 9476 2661
rect 10338 2836 10426 2849
rect 10338 2662 10351 2836
rect 10397 2662 10426 2836
rect 10338 2649 10426 2662
rect 10506 2836 10610 2849
rect 10506 2662 10535 2836
rect 10581 2662 10610 2836
rect 10506 2649 10610 2662
rect 10690 2836 10794 2849
rect 10690 2662 10719 2836
rect 10765 2662 10794 2836
rect 10690 2649 10794 2662
rect 10874 2836 10962 2849
rect 10874 2662 10903 2836
rect 10949 2662 10962 2836
rect 10874 2649 10962 2662
rect 12894 2835 12982 2848
rect 12894 2661 12907 2835
rect 12953 2661 12982 2835
rect 12894 2648 12982 2661
rect 13062 2835 13166 2848
rect 13062 2661 13091 2835
rect 13137 2661 13166 2835
rect 13062 2648 13166 2661
rect 13246 2835 13350 2848
rect 13246 2661 13275 2835
rect 13321 2661 13350 2835
rect 13246 2648 13350 2661
rect 13430 2835 13518 2848
rect 13430 2661 13459 2835
rect 13505 2661 13518 2835
rect 13430 2648 13518 2661
rect 14380 2836 14468 2849
rect 14380 2662 14393 2836
rect 14439 2662 14468 2836
rect 14380 2649 14468 2662
rect 14548 2836 14652 2849
rect 14548 2662 14577 2836
rect 14623 2662 14652 2836
rect 14548 2649 14652 2662
rect 14732 2836 14836 2849
rect 14732 2662 14761 2836
rect 14807 2662 14836 2836
rect 14732 2649 14836 2662
rect 14916 2836 15004 2849
rect 14916 2662 14945 2836
rect 14991 2662 15004 2836
rect 14916 2649 15004 2662
rect 16936 2835 17024 2848
rect 16936 2661 16949 2835
rect 16995 2661 17024 2835
rect 16936 2648 17024 2661
rect 17104 2835 17208 2848
rect 17104 2661 17133 2835
rect 17179 2661 17208 2835
rect 17104 2648 17208 2661
rect 17288 2835 17392 2848
rect 17288 2661 17317 2835
rect 17363 2661 17392 2835
rect 17288 2648 17392 2661
rect 17472 2835 17560 2848
rect 17472 2661 17501 2835
rect 17547 2661 17560 2835
rect 17472 2648 17560 2661
rect 18422 2836 18510 2849
rect 18422 2662 18435 2836
rect 18481 2662 18510 2836
rect 18422 2649 18510 2662
rect 18590 2836 18694 2849
rect 18590 2662 18619 2836
rect 18665 2662 18694 2836
rect 18590 2649 18694 2662
rect 18774 2836 18878 2849
rect 18774 2662 18803 2836
rect 18849 2662 18878 2836
rect 18774 2649 18878 2662
rect 18958 2836 19046 2849
rect 18958 2662 18987 2836
rect 19033 2662 19046 2836
rect 18958 2649 19046 2662
rect 20978 2835 21066 2848
rect 20978 2661 20991 2835
rect 21037 2661 21066 2835
rect 20978 2648 21066 2661
rect 21146 2835 21250 2848
rect 21146 2661 21175 2835
rect 21221 2661 21250 2835
rect 21146 2648 21250 2661
rect 21330 2835 21434 2848
rect 21330 2661 21359 2835
rect 21405 2661 21434 2835
rect 21330 2648 21434 2661
rect 21514 2835 21602 2848
rect 21514 2661 21543 2835
rect 21589 2661 21602 2835
rect 21514 2648 21602 2661
rect 22464 2836 22552 2849
rect 22464 2662 22477 2836
rect 22523 2662 22552 2836
rect 22464 2649 22552 2662
rect 22632 2836 22736 2849
rect 22632 2662 22661 2836
rect 22707 2662 22736 2836
rect 22632 2649 22736 2662
rect 22816 2836 22920 2849
rect 22816 2662 22845 2836
rect 22891 2662 22920 2836
rect 22816 2649 22920 2662
rect 23000 2836 23088 2849
rect 23000 2662 23029 2836
rect 23075 2662 23088 2836
rect 23000 2649 23088 2662
rect 25020 2835 25108 2848
rect 25020 2661 25033 2835
rect 25079 2661 25108 2835
rect 25020 2648 25108 2661
rect 25188 2835 25292 2848
rect 25188 2661 25217 2835
rect 25263 2661 25292 2835
rect 25188 2648 25292 2661
rect 25372 2835 25476 2848
rect 25372 2661 25401 2835
rect 25447 2661 25476 2835
rect 25372 2648 25476 2661
rect 25556 2835 25644 2848
rect 25556 2661 25585 2835
rect 25631 2661 25644 2835
rect 25556 2648 25644 2661
rect 26506 2836 26594 2849
rect 26506 2662 26519 2836
rect 26565 2662 26594 2836
rect 26506 2649 26594 2662
rect 26674 2836 26778 2849
rect 26674 2662 26703 2836
rect 26749 2662 26778 2836
rect 26674 2649 26778 2662
rect 26858 2836 26962 2849
rect 26858 2662 26887 2836
rect 26933 2662 26962 2836
rect 26858 2649 26962 2662
rect 27042 2836 27130 2849
rect 27042 2662 27071 2836
rect 27117 2662 27130 2836
rect 27042 2649 27130 2662
rect 798 630 886 643
rect 798 456 811 630
rect 857 456 886 630
rect 798 443 886 456
rect 966 630 1070 643
rect 966 456 995 630
rect 1041 456 1070 630
rect 966 443 1070 456
rect 1150 630 1254 643
rect 1150 456 1179 630
rect 1225 456 1254 630
rect 1150 443 1254 456
rect 1334 630 1422 643
rect 1334 456 1363 630
rect 1409 456 1422 630
rect 1334 443 1422 456
rect 4810 630 4898 643
rect 4810 456 4823 630
rect 4869 456 4898 630
rect 4810 443 4898 456
rect 4978 630 5082 643
rect 4978 456 5007 630
rect 5053 456 5082 630
rect 4978 443 5082 456
rect 5162 630 5266 643
rect 5162 456 5191 630
rect 5237 456 5266 630
rect 5162 443 5266 456
rect 5346 630 5434 643
rect 5346 456 5375 630
rect 5421 456 5434 630
rect 5346 443 5434 456
rect 8852 630 8940 643
rect 8852 456 8865 630
rect 8911 456 8940 630
rect 8852 443 8940 456
rect 9020 630 9124 643
rect 9020 456 9049 630
rect 9095 456 9124 630
rect 9020 443 9124 456
rect 9204 630 9308 643
rect 9204 456 9233 630
rect 9279 456 9308 630
rect 9204 443 9308 456
rect 9388 630 9476 643
rect 9388 456 9417 630
rect 9463 456 9476 630
rect 9388 443 9476 456
rect 12894 630 12982 643
rect 12894 456 12907 630
rect 12953 456 12982 630
rect 12894 443 12982 456
rect 13062 630 13166 643
rect 13062 456 13091 630
rect 13137 456 13166 630
rect 13062 443 13166 456
rect 13246 630 13350 643
rect 13246 456 13275 630
rect 13321 456 13350 630
rect 13246 443 13350 456
rect 13430 630 13518 643
rect 13430 456 13459 630
rect 13505 456 13518 630
rect 13430 443 13518 456
rect 16936 630 17024 643
rect 16936 456 16949 630
rect 16995 456 17024 630
rect 16936 443 17024 456
rect 17104 630 17208 643
rect 17104 456 17133 630
rect 17179 456 17208 630
rect 17104 443 17208 456
rect 17288 630 17392 643
rect 17288 456 17317 630
rect 17363 456 17392 630
rect 17288 443 17392 456
rect 17472 630 17560 643
rect 17472 456 17501 630
rect 17547 456 17560 630
rect 17472 443 17560 456
rect 20978 630 21066 643
rect 20978 456 20991 630
rect 21037 456 21066 630
rect 20978 443 21066 456
rect 21146 630 21250 643
rect 21146 456 21175 630
rect 21221 456 21250 630
rect 21146 443 21250 456
rect 21330 630 21434 643
rect 21330 456 21359 630
rect 21405 456 21434 630
rect 21330 443 21434 456
rect 21514 630 21602 643
rect 21514 456 21543 630
rect 21589 456 21602 630
rect 21514 443 21602 456
rect 25020 630 25108 643
rect 25020 456 25033 630
rect 25079 456 25108 630
rect 25020 443 25108 456
rect 25188 630 25292 643
rect 25188 456 25217 630
rect 25263 456 25292 630
rect 25188 443 25292 456
rect 25372 630 25476 643
rect 25372 456 25401 630
rect 25447 456 25476 630
rect 25372 443 25476 456
rect 25556 630 25644 643
rect 25556 456 25585 630
rect 25631 456 25644 630
rect 25556 443 25644 456
<< pdiff >>
rect 4810 17984 4898 17997
rect 4810 17510 4823 17984
rect 4869 17510 4898 17984
rect 4810 17497 4898 17510
rect 4978 17984 5082 17997
rect 4978 17510 5007 17984
rect 5053 17510 5082 17984
rect 4978 17497 5082 17510
rect 5162 17984 5266 17997
rect 5162 17510 5191 17984
rect 5237 17510 5266 17984
rect 5162 17497 5266 17510
rect 5346 17984 5434 17997
rect 5346 17510 5375 17984
rect 5421 17510 5434 17984
rect 5346 17497 5434 17510
rect 8852 17981 8940 17994
rect 8852 17507 8865 17981
rect 8911 17507 8940 17981
rect 8852 17494 8940 17507
rect 9020 17981 9124 17994
rect 9020 17507 9049 17981
rect 9095 17507 9124 17981
rect 9020 17494 9124 17507
rect 9204 17981 9308 17994
rect 9204 17507 9233 17981
rect 9279 17507 9308 17981
rect 9204 17494 9308 17507
rect 9388 17981 9476 17994
rect 9388 17507 9417 17981
rect 9463 17507 9476 17981
rect 9388 17494 9476 17507
rect 12894 17981 12982 17994
rect 12894 17507 12907 17981
rect 12953 17507 12982 17981
rect 12894 17494 12982 17507
rect 13062 17981 13166 17994
rect 13062 17507 13091 17981
rect 13137 17507 13166 17981
rect 13062 17494 13166 17507
rect 13246 17981 13350 17994
rect 13246 17507 13275 17981
rect 13321 17507 13350 17981
rect 13246 17494 13350 17507
rect 13430 17981 13518 17994
rect 13430 17507 13459 17981
rect 13505 17507 13518 17981
rect 13430 17494 13518 17507
rect 16936 17981 17024 17994
rect 16936 17507 16949 17981
rect 16995 17507 17024 17981
rect 16936 17494 17024 17507
rect 17104 17981 17208 17994
rect 17104 17507 17133 17981
rect 17179 17507 17208 17981
rect 17104 17494 17208 17507
rect 17288 17981 17392 17994
rect 17288 17507 17317 17981
rect 17363 17507 17392 17981
rect 17288 17494 17392 17507
rect 17472 17981 17560 17994
rect 17472 17507 17501 17981
rect 17547 17507 17560 17981
rect 17472 17494 17560 17507
rect 20978 17981 21066 17994
rect 20978 17507 20991 17981
rect 21037 17507 21066 17981
rect 20978 17494 21066 17507
rect 21146 17981 21250 17994
rect 21146 17507 21175 17981
rect 21221 17507 21250 17981
rect 21146 17494 21250 17507
rect 21330 17981 21434 17994
rect 21330 17507 21359 17981
rect 21405 17507 21434 17981
rect 21330 17494 21434 17507
rect 21514 17981 21602 17994
rect 21514 17507 21543 17981
rect 21589 17507 21602 17981
rect 21514 17494 21602 17507
rect 25020 17981 25108 17994
rect 25020 17507 25033 17981
rect 25079 17507 25108 17981
rect 25020 17494 25108 17507
rect 25188 17981 25292 17994
rect 25188 17507 25217 17981
rect 25263 17507 25292 17981
rect 25188 17494 25292 17507
rect 25372 17981 25476 17994
rect 25372 17507 25401 17981
rect 25447 17507 25476 17981
rect 25372 17494 25476 17507
rect 25556 17981 25644 17994
rect 25556 17507 25585 17981
rect 25631 17507 25644 17981
rect 25556 17494 25644 17507
rect 29062 17981 29150 17994
rect 29062 17507 29075 17981
rect 29121 17507 29150 17981
rect 29062 17494 29150 17507
rect 29230 17981 29334 17994
rect 29230 17507 29259 17981
rect 29305 17507 29334 17981
rect 29230 17494 29334 17507
rect 29414 17981 29518 17994
rect 29414 17507 29443 17981
rect 29489 17507 29518 17981
rect 29414 17494 29518 17507
rect 29598 17981 29686 17994
rect 29598 17507 29627 17981
rect 29673 17507 29686 17981
rect 29598 17494 29686 17507
rect 4810 15779 4898 15792
rect 4810 15305 4823 15779
rect 4869 15305 4898 15779
rect 4810 15292 4898 15305
rect 4978 15779 5082 15792
rect 4978 15305 5007 15779
rect 5053 15305 5082 15779
rect 4978 15292 5082 15305
rect 5162 15779 5266 15792
rect 5162 15305 5191 15779
rect 5237 15305 5266 15779
rect 5162 15292 5266 15305
rect 5346 15779 5434 15792
rect 5346 15305 5375 15779
rect 5421 15305 5434 15779
rect 5346 15292 5434 15305
rect 6296 15779 6384 15792
rect 6296 15305 6309 15779
rect 6355 15305 6384 15779
rect 6296 15292 6384 15305
rect 6464 15779 6568 15792
rect 6464 15305 6493 15779
rect 6539 15305 6568 15779
rect 6464 15292 6568 15305
rect 6648 15779 6752 15792
rect 6648 15305 6677 15779
rect 6723 15305 6752 15779
rect 6648 15292 6752 15305
rect 6832 15779 6920 15792
rect 6832 15305 6861 15779
rect 6907 15305 6920 15779
rect 6832 15292 6920 15305
rect 8852 15776 8940 15789
rect 8852 15302 8865 15776
rect 8911 15302 8940 15776
rect 8852 15289 8940 15302
rect 9020 15776 9124 15789
rect 9020 15302 9049 15776
rect 9095 15302 9124 15776
rect 9020 15289 9124 15302
rect 9204 15776 9308 15789
rect 9204 15302 9233 15776
rect 9279 15302 9308 15776
rect 9204 15289 9308 15302
rect 9388 15776 9476 15789
rect 9388 15302 9417 15776
rect 9463 15302 9476 15776
rect 9388 15289 9476 15302
rect 10338 15776 10426 15789
rect 10338 15302 10351 15776
rect 10397 15302 10426 15776
rect 10338 15289 10426 15302
rect 10506 15776 10610 15789
rect 10506 15302 10535 15776
rect 10581 15302 10610 15776
rect 10506 15289 10610 15302
rect 10690 15776 10794 15789
rect 10690 15302 10719 15776
rect 10765 15302 10794 15776
rect 10690 15289 10794 15302
rect 10874 15776 10962 15789
rect 10874 15302 10903 15776
rect 10949 15302 10962 15776
rect 10874 15289 10962 15302
rect 12894 15776 12982 15789
rect 12894 15302 12907 15776
rect 12953 15302 12982 15776
rect 12894 15289 12982 15302
rect 13062 15776 13166 15789
rect 13062 15302 13091 15776
rect 13137 15302 13166 15776
rect 13062 15289 13166 15302
rect 13246 15776 13350 15789
rect 13246 15302 13275 15776
rect 13321 15302 13350 15776
rect 13246 15289 13350 15302
rect 13430 15776 13518 15789
rect 13430 15302 13459 15776
rect 13505 15302 13518 15776
rect 13430 15289 13518 15302
rect 14380 15776 14468 15789
rect 14380 15302 14393 15776
rect 14439 15302 14468 15776
rect 14380 15289 14468 15302
rect 14548 15776 14652 15789
rect 14548 15302 14577 15776
rect 14623 15302 14652 15776
rect 14548 15289 14652 15302
rect 14732 15776 14836 15789
rect 14732 15302 14761 15776
rect 14807 15302 14836 15776
rect 14732 15289 14836 15302
rect 14916 15776 15004 15789
rect 14916 15302 14945 15776
rect 14991 15302 15004 15776
rect 14916 15289 15004 15302
rect 16936 15776 17024 15789
rect 16936 15302 16949 15776
rect 16995 15302 17024 15776
rect 16936 15289 17024 15302
rect 17104 15776 17208 15789
rect 17104 15302 17133 15776
rect 17179 15302 17208 15776
rect 17104 15289 17208 15302
rect 17288 15776 17392 15789
rect 17288 15302 17317 15776
rect 17363 15302 17392 15776
rect 17288 15289 17392 15302
rect 17472 15776 17560 15789
rect 17472 15302 17501 15776
rect 17547 15302 17560 15776
rect 17472 15289 17560 15302
rect 18422 15776 18510 15789
rect 18422 15302 18435 15776
rect 18481 15302 18510 15776
rect 18422 15289 18510 15302
rect 18590 15776 18694 15789
rect 18590 15302 18619 15776
rect 18665 15302 18694 15776
rect 18590 15289 18694 15302
rect 18774 15776 18878 15789
rect 18774 15302 18803 15776
rect 18849 15302 18878 15776
rect 18774 15289 18878 15302
rect 18958 15776 19046 15789
rect 18958 15302 18987 15776
rect 19033 15302 19046 15776
rect 18958 15289 19046 15302
rect 20978 15776 21066 15789
rect 20978 15302 20991 15776
rect 21037 15302 21066 15776
rect 20978 15289 21066 15302
rect 21146 15776 21250 15789
rect 21146 15302 21175 15776
rect 21221 15302 21250 15776
rect 21146 15289 21250 15302
rect 21330 15776 21434 15789
rect 21330 15302 21359 15776
rect 21405 15302 21434 15776
rect 21330 15289 21434 15302
rect 21514 15776 21602 15789
rect 21514 15302 21543 15776
rect 21589 15302 21602 15776
rect 21514 15289 21602 15302
rect 22464 15776 22552 15789
rect 22464 15302 22477 15776
rect 22523 15302 22552 15776
rect 22464 15289 22552 15302
rect 22632 15776 22736 15789
rect 22632 15302 22661 15776
rect 22707 15302 22736 15776
rect 22632 15289 22736 15302
rect 22816 15776 22920 15789
rect 22816 15302 22845 15776
rect 22891 15302 22920 15776
rect 22816 15289 22920 15302
rect 23000 15776 23088 15789
rect 23000 15302 23029 15776
rect 23075 15302 23088 15776
rect 23000 15289 23088 15302
rect 25020 15776 25108 15789
rect 25020 15302 25033 15776
rect 25079 15302 25108 15776
rect 25020 15289 25108 15302
rect 25188 15776 25292 15789
rect 25188 15302 25217 15776
rect 25263 15302 25292 15776
rect 25188 15289 25292 15302
rect 25372 15776 25476 15789
rect 25372 15302 25401 15776
rect 25447 15302 25476 15776
rect 25372 15289 25476 15302
rect 25556 15776 25644 15789
rect 25556 15302 25585 15776
rect 25631 15302 25644 15776
rect 25556 15289 25644 15302
rect 26506 15776 26594 15789
rect 26506 15302 26519 15776
rect 26565 15302 26594 15776
rect 26506 15289 26594 15302
rect 26674 15776 26778 15789
rect 26674 15302 26703 15776
rect 26749 15302 26778 15776
rect 26674 15289 26778 15302
rect 26858 15776 26962 15789
rect 26858 15302 26887 15776
rect 26933 15302 26962 15776
rect 26858 15289 26962 15302
rect 27042 15776 27130 15789
rect 27042 15302 27071 15776
rect 27117 15302 27130 15776
rect 27042 15289 27130 15302
rect 29062 15776 29150 15789
rect 29062 15302 29075 15776
rect 29121 15302 29150 15776
rect 29062 15289 29150 15302
rect 29230 15776 29334 15789
rect 29230 15302 29259 15776
rect 29305 15302 29334 15776
rect 29230 15289 29334 15302
rect 29414 15776 29518 15789
rect 29414 15302 29443 15776
rect 29489 15302 29518 15776
rect 29414 15289 29518 15302
rect 29598 15776 29686 15789
rect 29598 15302 29627 15776
rect 29673 15302 29686 15776
rect 29598 15289 29686 15302
rect 30548 15776 30636 15789
rect 30548 15302 30561 15776
rect 30607 15302 30636 15776
rect 30548 15289 30636 15302
rect 30716 15776 30820 15789
rect 30716 15302 30745 15776
rect 30791 15302 30820 15776
rect 30716 15289 30820 15302
rect 30900 15776 31004 15789
rect 30900 15302 30929 15776
rect 30975 15302 31004 15776
rect 30900 15289 31004 15302
rect 31084 15776 31172 15789
rect 31084 15302 31113 15776
rect 31159 15302 31172 15776
rect 31084 15289 31172 15302
rect 4810 13574 4898 13587
rect 4810 13100 4823 13574
rect 4869 13100 4898 13574
rect 4810 13087 4898 13100
rect 4978 13574 5082 13587
rect 4978 13100 5007 13574
rect 5053 13100 5082 13574
rect 4978 13087 5082 13100
rect 5162 13574 5266 13587
rect 5162 13100 5191 13574
rect 5237 13100 5266 13574
rect 5162 13087 5266 13100
rect 5346 13574 5434 13587
rect 5346 13100 5375 13574
rect 5421 13100 5434 13574
rect 5346 13087 5434 13100
rect 6296 13575 6384 13588
rect 6296 13101 6309 13575
rect 6355 13101 6384 13575
rect 6296 13088 6384 13101
rect 6464 13575 6568 13588
rect 6464 13101 6493 13575
rect 6539 13101 6568 13575
rect 6464 13088 6568 13101
rect 6648 13575 6752 13588
rect 6648 13101 6677 13575
rect 6723 13101 6752 13575
rect 6648 13088 6752 13101
rect 6832 13575 6920 13588
rect 6832 13101 6861 13575
rect 6907 13101 6920 13575
rect 6832 13088 6920 13101
rect 8852 13571 8940 13584
rect 8852 13097 8865 13571
rect 8911 13097 8940 13571
rect 8852 13084 8940 13097
rect 9020 13571 9124 13584
rect 9020 13097 9049 13571
rect 9095 13097 9124 13571
rect 9020 13084 9124 13097
rect 9204 13571 9308 13584
rect 9204 13097 9233 13571
rect 9279 13097 9308 13571
rect 9204 13084 9308 13097
rect 9388 13571 9476 13584
rect 9388 13097 9417 13571
rect 9463 13097 9476 13571
rect 9388 13084 9476 13097
rect 10338 13572 10426 13585
rect 10338 13098 10351 13572
rect 10397 13098 10426 13572
rect 10338 13085 10426 13098
rect 10506 13572 10610 13585
rect 10506 13098 10535 13572
rect 10581 13098 10610 13572
rect 10506 13085 10610 13098
rect 10690 13572 10794 13585
rect 10690 13098 10719 13572
rect 10765 13098 10794 13572
rect 10690 13085 10794 13098
rect 10874 13572 10962 13585
rect 10874 13098 10903 13572
rect 10949 13098 10962 13572
rect 10874 13085 10962 13098
rect 12894 13571 12982 13584
rect 12894 13097 12907 13571
rect 12953 13097 12982 13571
rect 12894 13084 12982 13097
rect 13062 13571 13166 13584
rect 13062 13097 13091 13571
rect 13137 13097 13166 13571
rect 13062 13084 13166 13097
rect 13246 13571 13350 13584
rect 13246 13097 13275 13571
rect 13321 13097 13350 13571
rect 13246 13084 13350 13097
rect 13430 13571 13518 13584
rect 13430 13097 13459 13571
rect 13505 13097 13518 13571
rect 13430 13084 13518 13097
rect 14380 13572 14468 13585
rect 14380 13098 14393 13572
rect 14439 13098 14468 13572
rect 14380 13085 14468 13098
rect 14548 13572 14652 13585
rect 14548 13098 14577 13572
rect 14623 13098 14652 13572
rect 14548 13085 14652 13098
rect 14732 13572 14836 13585
rect 14732 13098 14761 13572
rect 14807 13098 14836 13572
rect 14732 13085 14836 13098
rect 14916 13572 15004 13585
rect 14916 13098 14945 13572
rect 14991 13098 15004 13572
rect 14916 13085 15004 13098
rect 16936 13571 17024 13584
rect 16936 13097 16949 13571
rect 16995 13097 17024 13571
rect 16936 13084 17024 13097
rect 17104 13571 17208 13584
rect 17104 13097 17133 13571
rect 17179 13097 17208 13571
rect 17104 13084 17208 13097
rect 17288 13571 17392 13584
rect 17288 13097 17317 13571
rect 17363 13097 17392 13571
rect 17288 13084 17392 13097
rect 17472 13571 17560 13584
rect 17472 13097 17501 13571
rect 17547 13097 17560 13571
rect 17472 13084 17560 13097
rect 18422 13572 18510 13585
rect 18422 13098 18435 13572
rect 18481 13098 18510 13572
rect 18422 13085 18510 13098
rect 18590 13572 18694 13585
rect 18590 13098 18619 13572
rect 18665 13098 18694 13572
rect 18590 13085 18694 13098
rect 18774 13572 18878 13585
rect 18774 13098 18803 13572
rect 18849 13098 18878 13572
rect 18774 13085 18878 13098
rect 18958 13572 19046 13585
rect 18958 13098 18987 13572
rect 19033 13098 19046 13572
rect 18958 13085 19046 13098
rect 20978 13571 21066 13584
rect 20978 13097 20991 13571
rect 21037 13097 21066 13571
rect 20978 13084 21066 13097
rect 21146 13571 21250 13584
rect 21146 13097 21175 13571
rect 21221 13097 21250 13571
rect 21146 13084 21250 13097
rect 21330 13571 21434 13584
rect 21330 13097 21359 13571
rect 21405 13097 21434 13571
rect 21330 13084 21434 13097
rect 21514 13571 21602 13584
rect 21514 13097 21543 13571
rect 21589 13097 21602 13571
rect 21514 13084 21602 13097
rect 22464 13572 22552 13585
rect 22464 13098 22477 13572
rect 22523 13098 22552 13572
rect 22464 13085 22552 13098
rect 22632 13572 22736 13585
rect 22632 13098 22661 13572
rect 22707 13098 22736 13572
rect 22632 13085 22736 13098
rect 22816 13572 22920 13585
rect 22816 13098 22845 13572
rect 22891 13098 22920 13572
rect 22816 13085 22920 13098
rect 23000 13572 23088 13585
rect 23000 13098 23029 13572
rect 23075 13098 23088 13572
rect 23000 13085 23088 13098
rect 25020 13571 25108 13584
rect 25020 13097 25033 13571
rect 25079 13097 25108 13571
rect 25020 13084 25108 13097
rect 25188 13571 25292 13584
rect 25188 13097 25217 13571
rect 25263 13097 25292 13571
rect 25188 13084 25292 13097
rect 25372 13571 25476 13584
rect 25372 13097 25401 13571
rect 25447 13097 25476 13571
rect 25372 13084 25476 13097
rect 25556 13571 25644 13584
rect 25556 13097 25585 13571
rect 25631 13097 25644 13571
rect 25556 13084 25644 13097
rect 26506 13572 26594 13585
rect 26506 13098 26519 13572
rect 26565 13098 26594 13572
rect 26506 13085 26594 13098
rect 26674 13572 26778 13585
rect 26674 13098 26703 13572
rect 26749 13098 26778 13572
rect 26674 13085 26778 13098
rect 26858 13572 26962 13585
rect 26858 13098 26887 13572
rect 26933 13098 26962 13572
rect 26858 13085 26962 13098
rect 27042 13572 27130 13585
rect 27042 13098 27071 13572
rect 27117 13098 27130 13572
rect 27042 13085 27130 13098
rect 29062 13571 29150 13584
rect 29062 13097 29075 13571
rect 29121 13097 29150 13571
rect 29062 13084 29150 13097
rect 29230 13571 29334 13584
rect 29230 13097 29259 13571
rect 29305 13097 29334 13571
rect 29230 13084 29334 13097
rect 29414 13571 29518 13584
rect 29414 13097 29443 13571
rect 29489 13097 29518 13571
rect 29414 13084 29518 13097
rect 29598 13571 29686 13584
rect 29598 13097 29627 13571
rect 29673 13097 29686 13571
rect 29598 13084 29686 13097
rect 30548 13572 30636 13585
rect 30548 13098 30561 13572
rect 30607 13098 30636 13572
rect 30548 13085 30636 13098
rect 30716 13572 30820 13585
rect 30716 13098 30745 13572
rect 30791 13098 30820 13572
rect 30716 13085 30820 13098
rect 30900 13572 31004 13585
rect 30900 13098 30929 13572
rect 30975 13098 31004 13572
rect 30900 13085 31004 13098
rect 31084 13572 31172 13585
rect 31084 13098 31113 13572
rect 31159 13098 31172 13572
rect 31084 13085 31172 13098
rect 4810 11369 4898 11382
rect 4810 10895 4823 11369
rect 4869 10895 4898 11369
rect 4810 10882 4898 10895
rect 4978 11369 5082 11382
rect 4978 10895 5007 11369
rect 5053 10895 5082 11369
rect 4978 10882 5082 10895
rect 5162 11369 5266 11382
rect 5162 10895 5191 11369
rect 5237 10895 5266 11369
rect 5162 10882 5266 10895
rect 5346 11369 5434 11382
rect 5346 10895 5375 11369
rect 5421 10895 5434 11369
rect 5346 10882 5434 10895
rect 8852 11366 8940 11379
rect 8852 10892 8865 11366
rect 8911 10892 8940 11366
rect 8852 10879 8940 10892
rect 9020 11366 9124 11379
rect 9020 10892 9049 11366
rect 9095 10892 9124 11366
rect 9020 10879 9124 10892
rect 9204 11366 9308 11379
rect 9204 10892 9233 11366
rect 9279 10892 9308 11366
rect 9204 10879 9308 10892
rect 9388 11366 9476 11379
rect 9388 10892 9417 11366
rect 9463 10892 9476 11366
rect 9388 10879 9476 10892
rect 12894 11366 12982 11379
rect 12894 10892 12907 11366
rect 12953 10892 12982 11366
rect 12894 10879 12982 10892
rect 13062 11366 13166 11379
rect 13062 10892 13091 11366
rect 13137 10892 13166 11366
rect 13062 10879 13166 10892
rect 13246 11366 13350 11379
rect 13246 10892 13275 11366
rect 13321 10892 13350 11366
rect 13246 10879 13350 10892
rect 13430 11366 13518 11379
rect 13430 10892 13459 11366
rect 13505 10892 13518 11366
rect 13430 10879 13518 10892
rect 16936 11366 17024 11379
rect 16936 10892 16949 11366
rect 16995 10892 17024 11366
rect 16936 10879 17024 10892
rect 17104 11366 17208 11379
rect 17104 10892 17133 11366
rect 17179 10892 17208 11366
rect 17104 10879 17208 10892
rect 17288 11366 17392 11379
rect 17288 10892 17317 11366
rect 17363 10892 17392 11366
rect 17288 10879 17392 10892
rect 17472 11366 17560 11379
rect 17472 10892 17501 11366
rect 17547 10892 17560 11366
rect 17472 10879 17560 10892
rect 20978 11366 21066 11379
rect 20978 10892 20991 11366
rect 21037 10892 21066 11366
rect 20978 10879 21066 10892
rect 21146 11366 21250 11379
rect 21146 10892 21175 11366
rect 21221 10892 21250 11366
rect 21146 10879 21250 10892
rect 21330 11366 21434 11379
rect 21330 10892 21359 11366
rect 21405 10892 21434 11366
rect 21330 10879 21434 10892
rect 21514 11366 21602 11379
rect 21514 10892 21543 11366
rect 21589 10892 21602 11366
rect 21514 10879 21602 10892
rect 25020 11366 25108 11379
rect 25020 10892 25033 11366
rect 25079 10892 25108 11366
rect 25020 10879 25108 10892
rect 25188 11366 25292 11379
rect 25188 10892 25217 11366
rect 25263 10892 25292 11366
rect 25188 10879 25292 10892
rect 25372 11366 25476 11379
rect 25372 10892 25401 11366
rect 25447 10892 25476 11366
rect 25372 10879 25476 10892
rect 25556 11366 25644 11379
rect 25556 10892 25585 11366
rect 25631 10892 25644 11366
rect 25556 10879 25644 10892
rect 29062 11366 29150 11379
rect 29062 10892 29075 11366
rect 29121 10892 29150 11366
rect 29062 10879 29150 10892
rect 29230 11366 29334 11379
rect 29230 10892 29259 11366
rect 29305 10892 29334 11366
rect 29230 10879 29334 10892
rect 29414 11366 29518 11379
rect 29414 10892 29443 11366
rect 29489 10892 29518 11366
rect 29414 10879 29518 10892
rect 29598 11366 29686 11379
rect 29598 10892 29627 11366
rect 29673 10892 29686 11366
rect 29598 10879 29686 10892
rect 798 8405 886 8418
rect 798 7931 811 8405
rect 857 7931 886 8405
rect 798 7918 886 7931
rect 966 8405 1070 8418
rect 966 7931 995 8405
rect 1041 7931 1070 8405
rect 966 7918 1070 7931
rect 1150 8405 1254 8418
rect 1150 7931 1179 8405
rect 1225 7931 1254 8405
rect 1150 7918 1254 7931
rect 1334 8405 1422 8418
rect 1334 7931 1363 8405
rect 1409 7931 1422 8405
rect 1334 7918 1422 7931
rect 4810 8405 4898 8418
rect 4810 7931 4823 8405
rect 4869 7931 4898 8405
rect 4810 7918 4898 7931
rect 4978 8405 5082 8418
rect 4978 7931 5007 8405
rect 5053 7931 5082 8405
rect 4978 7918 5082 7931
rect 5162 8405 5266 8418
rect 5162 7931 5191 8405
rect 5237 7931 5266 8405
rect 5162 7918 5266 7931
rect 5346 8405 5434 8418
rect 5346 7931 5375 8405
rect 5421 7931 5434 8405
rect 5346 7918 5434 7931
rect 8852 8405 8940 8418
rect 8852 7931 8865 8405
rect 8911 7931 8940 8405
rect 8852 7918 8940 7931
rect 9020 8405 9124 8418
rect 9020 7931 9049 8405
rect 9095 7931 9124 8405
rect 9020 7918 9124 7931
rect 9204 8405 9308 8418
rect 9204 7931 9233 8405
rect 9279 7931 9308 8405
rect 9204 7918 9308 7931
rect 9388 8405 9476 8418
rect 9388 7931 9417 8405
rect 9463 7931 9476 8405
rect 9388 7918 9476 7931
rect 12894 8405 12982 8418
rect 12894 7931 12907 8405
rect 12953 7931 12982 8405
rect 12894 7918 12982 7931
rect 13062 8405 13166 8418
rect 13062 7931 13091 8405
rect 13137 7931 13166 8405
rect 13062 7918 13166 7931
rect 13246 8405 13350 8418
rect 13246 7931 13275 8405
rect 13321 7931 13350 8405
rect 13246 7918 13350 7931
rect 13430 8405 13518 8418
rect 13430 7931 13459 8405
rect 13505 7931 13518 8405
rect 13430 7918 13518 7931
rect 16936 8405 17024 8418
rect 16936 7931 16949 8405
rect 16995 7931 17024 8405
rect 16936 7918 17024 7931
rect 17104 8405 17208 8418
rect 17104 7931 17133 8405
rect 17179 7931 17208 8405
rect 17104 7918 17208 7931
rect 17288 8405 17392 8418
rect 17288 7931 17317 8405
rect 17363 7931 17392 8405
rect 17288 7918 17392 7931
rect 17472 8405 17560 8418
rect 17472 7931 17501 8405
rect 17547 7931 17560 8405
rect 17472 7918 17560 7931
rect 20978 8405 21066 8418
rect 20978 7931 20991 8405
rect 21037 7931 21066 8405
rect 20978 7918 21066 7931
rect 21146 8405 21250 8418
rect 21146 7931 21175 8405
rect 21221 7931 21250 8405
rect 21146 7918 21250 7931
rect 21330 8405 21434 8418
rect 21330 7931 21359 8405
rect 21405 7931 21434 8405
rect 21330 7918 21434 7931
rect 21514 8405 21602 8418
rect 21514 7931 21543 8405
rect 21589 7931 21602 8405
rect 21514 7918 21602 7931
rect 25020 8405 25108 8418
rect 25020 7931 25033 8405
rect 25079 7931 25108 8405
rect 25020 7918 25108 7931
rect 25188 8405 25292 8418
rect 25188 7931 25217 8405
rect 25263 7931 25292 8405
rect 25188 7918 25292 7931
rect 25372 8405 25476 8418
rect 25372 7931 25401 8405
rect 25447 7931 25476 8405
rect 25372 7918 25476 7931
rect 25556 8405 25644 8418
rect 25556 7931 25585 8405
rect 25631 7931 25644 8405
rect 25556 7918 25644 7931
rect 798 6200 886 6213
rect 798 5726 811 6200
rect 857 5726 886 6200
rect 798 5713 886 5726
rect 966 6200 1070 6213
rect 966 5726 995 6200
rect 1041 5726 1070 6200
rect 966 5713 1070 5726
rect 1150 6200 1254 6213
rect 1150 5726 1179 6200
rect 1225 5726 1254 6200
rect 1150 5713 1254 5726
rect 1334 6200 1422 6213
rect 1334 5726 1363 6200
rect 1409 5726 1422 6200
rect 1334 5713 1422 5726
rect 2284 6200 2372 6213
rect 2284 5726 2297 6200
rect 2343 5726 2372 6200
rect 2284 5713 2372 5726
rect 2452 6200 2556 6213
rect 2452 5726 2481 6200
rect 2527 5726 2556 6200
rect 2452 5713 2556 5726
rect 2636 6200 2740 6213
rect 2636 5726 2665 6200
rect 2711 5726 2740 6200
rect 2636 5713 2740 5726
rect 2820 6200 2908 6213
rect 2820 5726 2849 6200
rect 2895 5726 2908 6200
rect 2820 5713 2908 5726
rect 4810 6200 4898 6213
rect 4810 5726 4823 6200
rect 4869 5726 4898 6200
rect 4810 5713 4898 5726
rect 4978 6200 5082 6213
rect 4978 5726 5007 6200
rect 5053 5726 5082 6200
rect 4978 5713 5082 5726
rect 5162 6200 5266 6213
rect 5162 5726 5191 6200
rect 5237 5726 5266 6200
rect 5162 5713 5266 5726
rect 5346 6200 5434 6213
rect 5346 5726 5375 6200
rect 5421 5726 5434 6200
rect 5346 5713 5434 5726
rect 6296 6200 6384 6213
rect 6296 5726 6309 6200
rect 6355 5726 6384 6200
rect 6296 5713 6384 5726
rect 6464 6200 6568 6213
rect 6464 5726 6493 6200
rect 6539 5726 6568 6200
rect 6464 5713 6568 5726
rect 6648 6200 6752 6213
rect 6648 5726 6677 6200
rect 6723 5726 6752 6200
rect 6648 5713 6752 5726
rect 6832 6200 6920 6213
rect 6832 5726 6861 6200
rect 6907 5726 6920 6200
rect 6832 5713 6920 5726
rect 8852 6200 8940 6213
rect 8852 5726 8865 6200
rect 8911 5726 8940 6200
rect 8852 5713 8940 5726
rect 9020 6200 9124 6213
rect 9020 5726 9049 6200
rect 9095 5726 9124 6200
rect 9020 5713 9124 5726
rect 9204 6200 9308 6213
rect 9204 5726 9233 6200
rect 9279 5726 9308 6200
rect 9204 5713 9308 5726
rect 9388 6200 9476 6213
rect 9388 5726 9417 6200
rect 9463 5726 9476 6200
rect 9388 5713 9476 5726
rect 10338 6200 10426 6213
rect 10338 5726 10351 6200
rect 10397 5726 10426 6200
rect 10338 5713 10426 5726
rect 10506 6200 10610 6213
rect 10506 5726 10535 6200
rect 10581 5726 10610 6200
rect 10506 5713 10610 5726
rect 10690 6200 10794 6213
rect 10690 5726 10719 6200
rect 10765 5726 10794 6200
rect 10690 5713 10794 5726
rect 10874 6200 10962 6213
rect 10874 5726 10903 6200
rect 10949 5726 10962 6200
rect 10874 5713 10962 5726
rect 12894 6200 12982 6213
rect 12894 5726 12907 6200
rect 12953 5726 12982 6200
rect 12894 5713 12982 5726
rect 13062 6200 13166 6213
rect 13062 5726 13091 6200
rect 13137 5726 13166 6200
rect 13062 5713 13166 5726
rect 13246 6200 13350 6213
rect 13246 5726 13275 6200
rect 13321 5726 13350 6200
rect 13246 5713 13350 5726
rect 13430 6200 13518 6213
rect 13430 5726 13459 6200
rect 13505 5726 13518 6200
rect 13430 5713 13518 5726
rect 14380 6200 14468 6213
rect 14380 5726 14393 6200
rect 14439 5726 14468 6200
rect 14380 5713 14468 5726
rect 14548 6200 14652 6213
rect 14548 5726 14577 6200
rect 14623 5726 14652 6200
rect 14548 5713 14652 5726
rect 14732 6200 14836 6213
rect 14732 5726 14761 6200
rect 14807 5726 14836 6200
rect 14732 5713 14836 5726
rect 14916 6200 15004 6213
rect 14916 5726 14945 6200
rect 14991 5726 15004 6200
rect 14916 5713 15004 5726
rect 16936 6200 17024 6213
rect 16936 5726 16949 6200
rect 16995 5726 17024 6200
rect 16936 5713 17024 5726
rect 17104 6200 17208 6213
rect 17104 5726 17133 6200
rect 17179 5726 17208 6200
rect 17104 5713 17208 5726
rect 17288 6200 17392 6213
rect 17288 5726 17317 6200
rect 17363 5726 17392 6200
rect 17288 5713 17392 5726
rect 17472 6200 17560 6213
rect 17472 5726 17501 6200
rect 17547 5726 17560 6200
rect 17472 5713 17560 5726
rect 18422 6200 18510 6213
rect 18422 5726 18435 6200
rect 18481 5726 18510 6200
rect 18422 5713 18510 5726
rect 18590 6200 18694 6213
rect 18590 5726 18619 6200
rect 18665 5726 18694 6200
rect 18590 5713 18694 5726
rect 18774 6200 18878 6213
rect 18774 5726 18803 6200
rect 18849 5726 18878 6200
rect 18774 5713 18878 5726
rect 18958 6200 19046 6213
rect 18958 5726 18987 6200
rect 19033 5726 19046 6200
rect 18958 5713 19046 5726
rect 20978 6200 21066 6213
rect 20978 5726 20991 6200
rect 21037 5726 21066 6200
rect 20978 5713 21066 5726
rect 21146 6200 21250 6213
rect 21146 5726 21175 6200
rect 21221 5726 21250 6200
rect 21146 5713 21250 5726
rect 21330 6200 21434 6213
rect 21330 5726 21359 6200
rect 21405 5726 21434 6200
rect 21330 5713 21434 5726
rect 21514 6200 21602 6213
rect 21514 5726 21543 6200
rect 21589 5726 21602 6200
rect 21514 5713 21602 5726
rect 22464 6200 22552 6213
rect 22464 5726 22477 6200
rect 22523 5726 22552 6200
rect 22464 5713 22552 5726
rect 22632 6200 22736 6213
rect 22632 5726 22661 6200
rect 22707 5726 22736 6200
rect 22632 5713 22736 5726
rect 22816 6200 22920 6213
rect 22816 5726 22845 6200
rect 22891 5726 22920 6200
rect 22816 5713 22920 5726
rect 23000 6200 23088 6213
rect 23000 5726 23029 6200
rect 23075 5726 23088 6200
rect 23000 5713 23088 5726
rect 25020 6200 25108 6213
rect 25020 5726 25033 6200
rect 25079 5726 25108 6200
rect 25020 5713 25108 5726
rect 25188 6200 25292 6213
rect 25188 5726 25217 6200
rect 25263 5726 25292 6200
rect 25188 5713 25292 5726
rect 25372 6200 25476 6213
rect 25372 5726 25401 6200
rect 25447 5726 25476 6200
rect 25372 5713 25476 5726
rect 25556 6200 25644 6213
rect 25556 5726 25585 6200
rect 25631 5726 25644 6200
rect 25556 5713 25644 5726
rect 26506 6200 26594 6213
rect 26506 5726 26519 6200
rect 26565 5726 26594 6200
rect 26506 5713 26594 5726
rect 26674 6200 26778 6213
rect 26674 5726 26703 6200
rect 26749 5726 26778 6200
rect 26674 5713 26778 5726
rect 26858 6200 26962 6213
rect 26858 5726 26887 6200
rect 26933 5726 26962 6200
rect 26858 5713 26962 5726
rect 27042 6200 27130 6213
rect 27042 5726 27071 6200
rect 27117 5726 27130 6200
rect 27042 5713 27130 5726
rect 798 3995 886 4008
rect 798 3521 811 3995
rect 857 3521 886 3995
rect 798 3508 886 3521
rect 966 3995 1070 4008
rect 966 3521 995 3995
rect 1041 3521 1070 3995
rect 966 3508 1070 3521
rect 1150 3995 1254 4008
rect 1150 3521 1179 3995
rect 1225 3521 1254 3995
rect 1150 3508 1254 3521
rect 1334 3995 1422 4008
rect 1334 3521 1363 3995
rect 1409 3521 1422 3995
rect 1334 3508 1422 3521
rect 2284 3996 2372 4009
rect 2284 3522 2297 3996
rect 2343 3522 2372 3996
rect 2284 3509 2372 3522
rect 2452 3996 2556 4009
rect 2452 3522 2481 3996
rect 2527 3522 2556 3996
rect 2452 3509 2556 3522
rect 2636 3996 2740 4009
rect 2636 3522 2665 3996
rect 2711 3522 2740 3996
rect 2636 3509 2740 3522
rect 2820 3996 2908 4009
rect 2820 3522 2849 3996
rect 2895 3522 2908 3996
rect 2820 3509 2908 3522
rect 4810 3995 4898 4008
rect 4810 3521 4823 3995
rect 4869 3521 4898 3995
rect 4810 3508 4898 3521
rect 4978 3995 5082 4008
rect 4978 3521 5007 3995
rect 5053 3521 5082 3995
rect 4978 3508 5082 3521
rect 5162 3995 5266 4008
rect 5162 3521 5191 3995
rect 5237 3521 5266 3995
rect 5162 3508 5266 3521
rect 5346 3995 5434 4008
rect 5346 3521 5375 3995
rect 5421 3521 5434 3995
rect 5346 3508 5434 3521
rect 6296 3996 6384 4009
rect 6296 3522 6309 3996
rect 6355 3522 6384 3996
rect 6296 3509 6384 3522
rect 6464 3996 6568 4009
rect 6464 3522 6493 3996
rect 6539 3522 6568 3996
rect 6464 3509 6568 3522
rect 6648 3996 6752 4009
rect 6648 3522 6677 3996
rect 6723 3522 6752 3996
rect 6648 3509 6752 3522
rect 6832 3996 6920 4009
rect 6832 3522 6861 3996
rect 6907 3522 6920 3996
rect 6832 3509 6920 3522
rect 8852 3995 8940 4008
rect 8852 3521 8865 3995
rect 8911 3521 8940 3995
rect 8852 3508 8940 3521
rect 9020 3995 9124 4008
rect 9020 3521 9049 3995
rect 9095 3521 9124 3995
rect 9020 3508 9124 3521
rect 9204 3995 9308 4008
rect 9204 3521 9233 3995
rect 9279 3521 9308 3995
rect 9204 3508 9308 3521
rect 9388 3995 9476 4008
rect 9388 3521 9417 3995
rect 9463 3521 9476 3995
rect 9388 3508 9476 3521
rect 10338 3996 10426 4009
rect 10338 3522 10351 3996
rect 10397 3522 10426 3996
rect 10338 3509 10426 3522
rect 10506 3996 10610 4009
rect 10506 3522 10535 3996
rect 10581 3522 10610 3996
rect 10506 3509 10610 3522
rect 10690 3996 10794 4009
rect 10690 3522 10719 3996
rect 10765 3522 10794 3996
rect 10690 3509 10794 3522
rect 10874 3996 10962 4009
rect 10874 3522 10903 3996
rect 10949 3522 10962 3996
rect 10874 3509 10962 3522
rect 12894 3995 12982 4008
rect 12894 3521 12907 3995
rect 12953 3521 12982 3995
rect 12894 3508 12982 3521
rect 13062 3995 13166 4008
rect 13062 3521 13091 3995
rect 13137 3521 13166 3995
rect 13062 3508 13166 3521
rect 13246 3995 13350 4008
rect 13246 3521 13275 3995
rect 13321 3521 13350 3995
rect 13246 3508 13350 3521
rect 13430 3995 13518 4008
rect 13430 3521 13459 3995
rect 13505 3521 13518 3995
rect 13430 3508 13518 3521
rect 14380 3996 14468 4009
rect 14380 3522 14393 3996
rect 14439 3522 14468 3996
rect 14380 3509 14468 3522
rect 14548 3996 14652 4009
rect 14548 3522 14577 3996
rect 14623 3522 14652 3996
rect 14548 3509 14652 3522
rect 14732 3996 14836 4009
rect 14732 3522 14761 3996
rect 14807 3522 14836 3996
rect 14732 3509 14836 3522
rect 14916 3996 15004 4009
rect 14916 3522 14945 3996
rect 14991 3522 15004 3996
rect 14916 3509 15004 3522
rect 16936 3995 17024 4008
rect 16936 3521 16949 3995
rect 16995 3521 17024 3995
rect 16936 3508 17024 3521
rect 17104 3995 17208 4008
rect 17104 3521 17133 3995
rect 17179 3521 17208 3995
rect 17104 3508 17208 3521
rect 17288 3995 17392 4008
rect 17288 3521 17317 3995
rect 17363 3521 17392 3995
rect 17288 3508 17392 3521
rect 17472 3995 17560 4008
rect 17472 3521 17501 3995
rect 17547 3521 17560 3995
rect 17472 3508 17560 3521
rect 18422 3996 18510 4009
rect 18422 3522 18435 3996
rect 18481 3522 18510 3996
rect 18422 3509 18510 3522
rect 18590 3996 18694 4009
rect 18590 3522 18619 3996
rect 18665 3522 18694 3996
rect 18590 3509 18694 3522
rect 18774 3996 18878 4009
rect 18774 3522 18803 3996
rect 18849 3522 18878 3996
rect 18774 3509 18878 3522
rect 18958 3996 19046 4009
rect 18958 3522 18987 3996
rect 19033 3522 19046 3996
rect 18958 3509 19046 3522
rect 20978 3995 21066 4008
rect 20978 3521 20991 3995
rect 21037 3521 21066 3995
rect 20978 3508 21066 3521
rect 21146 3995 21250 4008
rect 21146 3521 21175 3995
rect 21221 3521 21250 3995
rect 21146 3508 21250 3521
rect 21330 3995 21434 4008
rect 21330 3521 21359 3995
rect 21405 3521 21434 3995
rect 21330 3508 21434 3521
rect 21514 3995 21602 4008
rect 21514 3521 21543 3995
rect 21589 3521 21602 3995
rect 21514 3508 21602 3521
rect 22464 3996 22552 4009
rect 22464 3522 22477 3996
rect 22523 3522 22552 3996
rect 22464 3509 22552 3522
rect 22632 3996 22736 4009
rect 22632 3522 22661 3996
rect 22707 3522 22736 3996
rect 22632 3509 22736 3522
rect 22816 3996 22920 4009
rect 22816 3522 22845 3996
rect 22891 3522 22920 3996
rect 22816 3509 22920 3522
rect 23000 3996 23088 4009
rect 23000 3522 23029 3996
rect 23075 3522 23088 3996
rect 23000 3509 23088 3522
rect 25020 3995 25108 4008
rect 25020 3521 25033 3995
rect 25079 3521 25108 3995
rect 25020 3508 25108 3521
rect 25188 3995 25292 4008
rect 25188 3521 25217 3995
rect 25263 3521 25292 3995
rect 25188 3508 25292 3521
rect 25372 3995 25476 4008
rect 25372 3521 25401 3995
rect 25447 3521 25476 3995
rect 25372 3508 25476 3521
rect 25556 3995 25644 4008
rect 25556 3521 25585 3995
rect 25631 3521 25644 3995
rect 25556 3508 25644 3521
rect 26506 3996 26594 4009
rect 26506 3522 26519 3996
rect 26565 3522 26594 3996
rect 26506 3509 26594 3522
rect 26674 3996 26778 4009
rect 26674 3522 26703 3996
rect 26749 3522 26778 3996
rect 26674 3509 26778 3522
rect 26858 3996 26962 4009
rect 26858 3522 26887 3996
rect 26933 3522 26962 3996
rect 26858 3509 26962 3522
rect 27042 3996 27130 4009
rect 27042 3522 27071 3996
rect 27117 3522 27130 3996
rect 27042 3509 27130 3522
rect 798 1790 886 1803
rect 798 1316 811 1790
rect 857 1316 886 1790
rect 798 1303 886 1316
rect 966 1790 1070 1803
rect 966 1316 995 1790
rect 1041 1316 1070 1790
rect 966 1303 1070 1316
rect 1150 1790 1254 1803
rect 1150 1316 1179 1790
rect 1225 1316 1254 1790
rect 1150 1303 1254 1316
rect 1334 1790 1422 1803
rect 1334 1316 1363 1790
rect 1409 1316 1422 1790
rect 1334 1303 1422 1316
rect 4810 1790 4898 1803
rect 4810 1316 4823 1790
rect 4869 1316 4898 1790
rect 4810 1303 4898 1316
rect 4978 1790 5082 1803
rect 4978 1316 5007 1790
rect 5053 1316 5082 1790
rect 4978 1303 5082 1316
rect 5162 1790 5266 1803
rect 5162 1316 5191 1790
rect 5237 1316 5266 1790
rect 5162 1303 5266 1316
rect 5346 1790 5434 1803
rect 5346 1316 5375 1790
rect 5421 1316 5434 1790
rect 5346 1303 5434 1316
rect 8852 1790 8940 1803
rect 8852 1316 8865 1790
rect 8911 1316 8940 1790
rect 8852 1303 8940 1316
rect 9020 1790 9124 1803
rect 9020 1316 9049 1790
rect 9095 1316 9124 1790
rect 9020 1303 9124 1316
rect 9204 1790 9308 1803
rect 9204 1316 9233 1790
rect 9279 1316 9308 1790
rect 9204 1303 9308 1316
rect 9388 1790 9476 1803
rect 9388 1316 9417 1790
rect 9463 1316 9476 1790
rect 9388 1303 9476 1316
rect 12894 1790 12982 1803
rect 12894 1316 12907 1790
rect 12953 1316 12982 1790
rect 12894 1303 12982 1316
rect 13062 1790 13166 1803
rect 13062 1316 13091 1790
rect 13137 1316 13166 1790
rect 13062 1303 13166 1316
rect 13246 1790 13350 1803
rect 13246 1316 13275 1790
rect 13321 1316 13350 1790
rect 13246 1303 13350 1316
rect 13430 1790 13518 1803
rect 13430 1316 13459 1790
rect 13505 1316 13518 1790
rect 13430 1303 13518 1316
rect 16936 1790 17024 1803
rect 16936 1316 16949 1790
rect 16995 1316 17024 1790
rect 16936 1303 17024 1316
rect 17104 1790 17208 1803
rect 17104 1316 17133 1790
rect 17179 1316 17208 1790
rect 17104 1303 17208 1316
rect 17288 1790 17392 1803
rect 17288 1316 17317 1790
rect 17363 1316 17392 1790
rect 17288 1303 17392 1316
rect 17472 1790 17560 1803
rect 17472 1316 17501 1790
rect 17547 1316 17560 1790
rect 17472 1303 17560 1316
rect 20978 1790 21066 1803
rect 20978 1316 20991 1790
rect 21037 1316 21066 1790
rect 20978 1303 21066 1316
rect 21146 1790 21250 1803
rect 21146 1316 21175 1790
rect 21221 1316 21250 1790
rect 21146 1303 21250 1316
rect 21330 1790 21434 1803
rect 21330 1316 21359 1790
rect 21405 1316 21434 1790
rect 21330 1303 21434 1316
rect 21514 1790 21602 1803
rect 21514 1316 21543 1790
rect 21589 1316 21602 1790
rect 21514 1303 21602 1316
rect 25020 1790 25108 1803
rect 25020 1316 25033 1790
rect 25079 1316 25108 1790
rect 25020 1303 25108 1316
rect 25188 1790 25292 1803
rect 25188 1316 25217 1790
rect 25263 1316 25292 1790
rect 25188 1303 25292 1316
rect 25372 1790 25476 1803
rect 25372 1316 25401 1790
rect 25447 1316 25476 1790
rect 25372 1303 25476 1316
rect 25556 1790 25644 1803
rect 25556 1316 25585 1790
rect 25631 1316 25644 1790
rect 25556 1303 25644 1316
<< ndiffc >>
rect 4823 16650 4869 16824
rect 5007 16650 5053 16824
rect 5191 16650 5237 16824
rect 5375 16650 5421 16824
rect 8865 16647 8911 16821
rect 9049 16647 9095 16821
rect 9233 16647 9279 16821
rect 9417 16647 9463 16821
rect 12907 16647 12953 16821
rect 13091 16647 13137 16821
rect 13275 16647 13321 16821
rect 13459 16647 13505 16821
rect 16949 16647 16995 16821
rect 17133 16647 17179 16821
rect 17317 16647 17363 16821
rect 17501 16647 17547 16821
rect 20991 16647 21037 16821
rect 21175 16647 21221 16821
rect 21359 16647 21405 16821
rect 21543 16647 21589 16821
rect 25033 16647 25079 16821
rect 25217 16647 25263 16821
rect 25401 16647 25447 16821
rect 25585 16647 25631 16821
rect 29075 16647 29121 16821
rect 29259 16647 29305 16821
rect 29443 16647 29489 16821
rect 29627 16647 29673 16821
rect 4823 14445 4869 14619
rect 5007 14445 5053 14619
rect 5191 14445 5237 14619
rect 5375 14445 5421 14619
rect 6309 14445 6355 14619
rect 6493 14445 6539 14619
rect 6677 14445 6723 14619
rect 6861 14445 6907 14619
rect 8865 14442 8911 14616
rect 9049 14442 9095 14616
rect 9233 14442 9279 14616
rect 9417 14442 9463 14616
rect 10351 14442 10397 14616
rect 10535 14442 10581 14616
rect 10719 14442 10765 14616
rect 10903 14442 10949 14616
rect 12907 14442 12953 14616
rect 13091 14442 13137 14616
rect 13275 14442 13321 14616
rect 13459 14442 13505 14616
rect 14393 14442 14439 14616
rect 14577 14442 14623 14616
rect 14761 14442 14807 14616
rect 14945 14442 14991 14616
rect 16949 14442 16995 14616
rect 17133 14442 17179 14616
rect 17317 14442 17363 14616
rect 17501 14442 17547 14616
rect 18435 14442 18481 14616
rect 18619 14442 18665 14616
rect 18803 14442 18849 14616
rect 18987 14442 19033 14616
rect 20991 14442 21037 14616
rect 21175 14442 21221 14616
rect 21359 14442 21405 14616
rect 21543 14442 21589 14616
rect 22477 14442 22523 14616
rect 22661 14442 22707 14616
rect 22845 14442 22891 14616
rect 23029 14442 23075 14616
rect 25033 14442 25079 14616
rect 25217 14442 25263 14616
rect 25401 14442 25447 14616
rect 25585 14442 25631 14616
rect 26519 14442 26565 14616
rect 26703 14442 26749 14616
rect 26887 14442 26933 14616
rect 27071 14442 27117 14616
rect 29075 14442 29121 14616
rect 29259 14442 29305 14616
rect 29443 14442 29489 14616
rect 29627 14442 29673 14616
rect 30561 14442 30607 14616
rect 30745 14442 30791 14616
rect 30929 14442 30975 14616
rect 31113 14442 31159 14616
rect 4823 12240 4869 12414
rect 5007 12240 5053 12414
rect 5191 12240 5237 12414
rect 5375 12240 5421 12414
rect 6309 12241 6355 12415
rect 6493 12241 6539 12415
rect 6677 12241 6723 12415
rect 6861 12241 6907 12415
rect 8865 12237 8911 12411
rect 9049 12237 9095 12411
rect 9233 12237 9279 12411
rect 9417 12237 9463 12411
rect 10351 12238 10397 12412
rect 10535 12238 10581 12412
rect 10719 12238 10765 12412
rect 10903 12238 10949 12412
rect 12907 12237 12953 12411
rect 13091 12237 13137 12411
rect 13275 12237 13321 12411
rect 13459 12237 13505 12411
rect 14393 12238 14439 12412
rect 14577 12238 14623 12412
rect 14761 12238 14807 12412
rect 14945 12238 14991 12412
rect 16949 12237 16995 12411
rect 17133 12237 17179 12411
rect 17317 12237 17363 12411
rect 17501 12237 17547 12411
rect 18435 12238 18481 12412
rect 18619 12238 18665 12412
rect 18803 12238 18849 12412
rect 18987 12238 19033 12412
rect 20991 12237 21037 12411
rect 21175 12237 21221 12411
rect 21359 12237 21405 12411
rect 21543 12237 21589 12411
rect 22477 12238 22523 12412
rect 22661 12238 22707 12412
rect 22845 12238 22891 12412
rect 23029 12238 23075 12412
rect 25033 12237 25079 12411
rect 25217 12237 25263 12411
rect 25401 12237 25447 12411
rect 25585 12237 25631 12411
rect 26519 12238 26565 12412
rect 26703 12238 26749 12412
rect 26887 12238 26933 12412
rect 27071 12238 27117 12412
rect 29075 12237 29121 12411
rect 29259 12237 29305 12411
rect 29443 12237 29489 12411
rect 29627 12237 29673 12411
rect 30561 12238 30607 12412
rect 30745 12238 30791 12412
rect 30929 12238 30975 12412
rect 31113 12238 31159 12412
rect 4823 10035 4869 10209
rect 5007 10035 5053 10209
rect 5191 10035 5237 10209
rect 5375 10035 5421 10209
rect 8865 10032 8911 10206
rect 9049 10032 9095 10206
rect 9233 10032 9279 10206
rect 9417 10032 9463 10206
rect 12907 10032 12953 10206
rect 13091 10032 13137 10206
rect 13275 10032 13321 10206
rect 13459 10032 13505 10206
rect 16949 10032 16995 10206
rect 17133 10032 17179 10206
rect 17317 10032 17363 10206
rect 17501 10032 17547 10206
rect 20991 10032 21037 10206
rect 21175 10032 21221 10206
rect 21359 10032 21405 10206
rect 21543 10032 21589 10206
rect 25033 10032 25079 10206
rect 25217 10032 25263 10206
rect 25401 10032 25447 10206
rect 25585 10032 25631 10206
rect 29075 10032 29121 10206
rect 29259 10032 29305 10206
rect 29443 10032 29489 10206
rect 29627 10032 29673 10206
rect 811 7071 857 7245
rect 995 7071 1041 7245
rect 1179 7071 1225 7245
rect 1363 7071 1409 7245
rect 4823 7071 4869 7245
rect 5007 7071 5053 7245
rect 5191 7071 5237 7245
rect 5375 7071 5421 7245
rect 8865 7071 8911 7245
rect 9049 7071 9095 7245
rect 9233 7071 9279 7245
rect 9417 7071 9463 7245
rect 12907 7071 12953 7245
rect 13091 7071 13137 7245
rect 13275 7071 13321 7245
rect 13459 7071 13505 7245
rect 16949 7071 16995 7245
rect 17133 7071 17179 7245
rect 17317 7071 17363 7245
rect 17501 7071 17547 7245
rect 20991 7071 21037 7245
rect 21175 7071 21221 7245
rect 21359 7071 21405 7245
rect 21543 7071 21589 7245
rect 25033 7071 25079 7245
rect 25217 7071 25263 7245
rect 25401 7071 25447 7245
rect 25585 7071 25631 7245
rect 811 4866 857 5040
rect 995 4866 1041 5040
rect 1179 4866 1225 5040
rect 1363 4866 1409 5040
rect 2297 4866 2343 5040
rect 2481 4866 2527 5040
rect 2665 4866 2711 5040
rect 2849 4866 2895 5040
rect 4823 4866 4869 5040
rect 5007 4866 5053 5040
rect 5191 4866 5237 5040
rect 5375 4866 5421 5040
rect 6309 4866 6355 5040
rect 6493 4866 6539 5040
rect 6677 4866 6723 5040
rect 6861 4866 6907 5040
rect 8865 4866 8911 5040
rect 9049 4866 9095 5040
rect 9233 4866 9279 5040
rect 9417 4866 9463 5040
rect 10351 4866 10397 5040
rect 10535 4866 10581 5040
rect 10719 4866 10765 5040
rect 10903 4866 10949 5040
rect 12907 4866 12953 5040
rect 13091 4866 13137 5040
rect 13275 4866 13321 5040
rect 13459 4866 13505 5040
rect 14393 4866 14439 5040
rect 14577 4866 14623 5040
rect 14761 4866 14807 5040
rect 14945 4866 14991 5040
rect 16949 4866 16995 5040
rect 17133 4866 17179 5040
rect 17317 4866 17363 5040
rect 17501 4866 17547 5040
rect 18435 4866 18481 5040
rect 18619 4866 18665 5040
rect 18803 4866 18849 5040
rect 18987 4866 19033 5040
rect 20991 4866 21037 5040
rect 21175 4866 21221 5040
rect 21359 4866 21405 5040
rect 21543 4866 21589 5040
rect 22477 4866 22523 5040
rect 22661 4866 22707 5040
rect 22845 4866 22891 5040
rect 23029 4866 23075 5040
rect 25033 4866 25079 5040
rect 25217 4866 25263 5040
rect 25401 4866 25447 5040
rect 25585 4866 25631 5040
rect 26519 4866 26565 5040
rect 26703 4866 26749 5040
rect 26887 4866 26933 5040
rect 27071 4866 27117 5040
rect 811 2661 857 2835
rect 995 2661 1041 2835
rect 1179 2661 1225 2835
rect 1363 2661 1409 2835
rect 2297 2662 2343 2836
rect 2481 2662 2527 2836
rect 2665 2662 2711 2836
rect 2849 2662 2895 2836
rect 4823 2661 4869 2835
rect 5007 2661 5053 2835
rect 5191 2661 5237 2835
rect 5375 2661 5421 2835
rect 6309 2662 6355 2836
rect 6493 2662 6539 2836
rect 6677 2662 6723 2836
rect 6861 2662 6907 2836
rect 8865 2661 8911 2835
rect 9049 2661 9095 2835
rect 9233 2661 9279 2835
rect 9417 2661 9463 2835
rect 10351 2662 10397 2836
rect 10535 2662 10581 2836
rect 10719 2662 10765 2836
rect 10903 2662 10949 2836
rect 12907 2661 12953 2835
rect 13091 2661 13137 2835
rect 13275 2661 13321 2835
rect 13459 2661 13505 2835
rect 14393 2662 14439 2836
rect 14577 2662 14623 2836
rect 14761 2662 14807 2836
rect 14945 2662 14991 2836
rect 16949 2661 16995 2835
rect 17133 2661 17179 2835
rect 17317 2661 17363 2835
rect 17501 2661 17547 2835
rect 18435 2662 18481 2836
rect 18619 2662 18665 2836
rect 18803 2662 18849 2836
rect 18987 2662 19033 2836
rect 20991 2661 21037 2835
rect 21175 2661 21221 2835
rect 21359 2661 21405 2835
rect 21543 2661 21589 2835
rect 22477 2662 22523 2836
rect 22661 2662 22707 2836
rect 22845 2662 22891 2836
rect 23029 2662 23075 2836
rect 25033 2661 25079 2835
rect 25217 2661 25263 2835
rect 25401 2661 25447 2835
rect 25585 2661 25631 2835
rect 26519 2662 26565 2836
rect 26703 2662 26749 2836
rect 26887 2662 26933 2836
rect 27071 2662 27117 2836
rect 811 456 857 630
rect 995 456 1041 630
rect 1179 456 1225 630
rect 1363 456 1409 630
rect 4823 456 4869 630
rect 5007 456 5053 630
rect 5191 456 5237 630
rect 5375 456 5421 630
rect 8865 456 8911 630
rect 9049 456 9095 630
rect 9233 456 9279 630
rect 9417 456 9463 630
rect 12907 456 12953 630
rect 13091 456 13137 630
rect 13275 456 13321 630
rect 13459 456 13505 630
rect 16949 456 16995 630
rect 17133 456 17179 630
rect 17317 456 17363 630
rect 17501 456 17547 630
rect 20991 456 21037 630
rect 21175 456 21221 630
rect 21359 456 21405 630
rect 21543 456 21589 630
rect 25033 456 25079 630
rect 25217 456 25263 630
rect 25401 456 25447 630
rect 25585 456 25631 630
<< pdiffc >>
rect 4823 17510 4869 17984
rect 5007 17510 5053 17984
rect 5191 17510 5237 17984
rect 5375 17510 5421 17984
rect 8865 17507 8911 17981
rect 9049 17507 9095 17981
rect 9233 17507 9279 17981
rect 9417 17507 9463 17981
rect 12907 17507 12953 17981
rect 13091 17507 13137 17981
rect 13275 17507 13321 17981
rect 13459 17507 13505 17981
rect 16949 17507 16995 17981
rect 17133 17507 17179 17981
rect 17317 17507 17363 17981
rect 17501 17507 17547 17981
rect 20991 17507 21037 17981
rect 21175 17507 21221 17981
rect 21359 17507 21405 17981
rect 21543 17507 21589 17981
rect 25033 17507 25079 17981
rect 25217 17507 25263 17981
rect 25401 17507 25447 17981
rect 25585 17507 25631 17981
rect 29075 17507 29121 17981
rect 29259 17507 29305 17981
rect 29443 17507 29489 17981
rect 29627 17507 29673 17981
rect 4823 15305 4869 15779
rect 5007 15305 5053 15779
rect 5191 15305 5237 15779
rect 5375 15305 5421 15779
rect 6309 15305 6355 15779
rect 6493 15305 6539 15779
rect 6677 15305 6723 15779
rect 6861 15305 6907 15779
rect 8865 15302 8911 15776
rect 9049 15302 9095 15776
rect 9233 15302 9279 15776
rect 9417 15302 9463 15776
rect 10351 15302 10397 15776
rect 10535 15302 10581 15776
rect 10719 15302 10765 15776
rect 10903 15302 10949 15776
rect 12907 15302 12953 15776
rect 13091 15302 13137 15776
rect 13275 15302 13321 15776
rect 13459 15302 13505 15776
rect 14393 15302 14439 15776
rect 14577 15302 14623 15776
rect 14761 15302 14807 15776
rect 14945 15302 14991 15776
rect 16949 15302 16995 15776
rect 17133 15302 17179 15776
rect 17317 15302 17363 15776
rect 17501 15302 17547 15776
rect 18435 15302 18481 15776
rect 18619 15302 18665 15776
rect 18803 15302 18849 15776
rect 18987 15302 19033 15776
rect 20991 15302 21037 15776
rect 21175 15302 21221 15776
rect 21359 15302 21405 15776
rect 21543 15302 21589 15776
rect 22477 15302 22523 15776
rect 22661 15302 22707 15776
rect 22845 15302 22891 15776
rect 23029 15302 23075 15776
rect 25033 15302 25079 15776
rect 25217 15302 25263 15776
rect 25401 15302 25447 15776
rect 25585 15302 25631 15776
rect 26519 15302 26565 15776
rect 26703 15302 26749 15776
rect 26887 15302 26933 15776
rect 27071 15302 27117 15776
rect 29075 15302 29121 15776
rect 29259 15302 29305 15776
rect 29443 15302 29489 15776
rect 29627 15302 29673 15776
rect 30561 15302 30607 15776
rect 30745 15302 30791 15776
rect 30929 15302 30975 15776
rect 31113 15302 31159 15776
rect 4823 13100 4869 13574
rect 5007 13100 5053 13574
rect 5191 13100 5237 13574
rect 5375 13100 5421 13574
rect 6309 13101 6355 13575
rect 6493 13101 6539 13575
rect 6677 13101 6723 13575
rect 6861 13101 6907 13575
rect 8865 13097 8911 13571
rect 9049 13097 9095 13571
rect 9233 13097 9279 13571
rect 9417 13097 9463 13571
rect 10351 13098 10397 13572
rect 10535 13098 10581 13572
rect 10719 13098 10765 13572
rect 10903 13098 10949 13572
rect 12907 13097 12953 13571
rect 13091 13097 13137 13571
rect 13275 13097 13321 13571
rect 13459 13097 13505 13571
rect 14393 13098 14439 13572
rect 14577 13098 14623 13572
rect 14761 13098 14807 13572
rect 14945 13098 14991 13572
rect 16949 13097 16995 13571
rect 17133 13097 17179 13571
rect 17317 13097 17363 13571
rect 17501 13097 17547 13571
rect 18435 13098 18481 13572
rect 18619 13098 18665 13572
rect 18803 13098 18849 13572
rect 18987 13098 19033 13572
rect 20991 13097 21037 13571
rect 21175 13097 21221 13571
rect 21359 13097 21405 13571
rect 21543 13097 21589 13571
rect 22477 13098 22523 13572
rect 22661 13098 22707 13572
rect 22845 13098 22891 13572
rect 23029 13098 23075 13572
rect 25033 13097 25079 13571
rect 25217 13097 25263 13571
rect 25401 13097 25447 13571
rect 25585 13097 25631 13571
rect 26519 13098 26565 13572
rect 26703 13098 26749 13572
rect 26887 13098 26933 13572
rect 27071 13098 27117 13572
rect 29075 13097 29121 13571
rect 29259 13097 29305 13571
rect 29443 13097 29489 13571
rect 29627 13097 29673 13571
rect 30561 13098 30607 13572
rect 30745 13098 30791 13572
rect 30929 13098 30975 13572
rect 31113 13098 31159 13572
rect 4823 10895 4869 11369
rect 5007 10895 5053 11369
rect 5191 10895 5237 11369
rect 5375 10895 5421 11369
rect 8865 10892 8911 11366
rect 9049 10892 9095 11366
rect 9233 10892 9279 11366
rect 9417 10892 9463 11366
rect 12907 10892 12953 11366
rect 13091 10892 13137 11366
rect 13275 10892 13321 11366
rect 13459 10892 13505 11366
rect 16949 10892 16995 11366
rect 17133 10892 17179 11366
rect 17317 10892 17363 11366
rect 17501 10892 17547 11366
rect 20991 10892 21037 11366
rect 21175 10892 21221 11366
rect 21359 10892 21405 11366
rect 21543 10892 21589 11366
rect 25033 10892 25079 11366
rect 25217 10892 25263 11366
rect 25401 10892 25447 11366
rect 25585 10892 25631 11366
rect 29075 10892 29121 11366
rect 29259 10892 29305 11366
rect 29443 10892 29489 11366
rect 29627 10892 29673 11366
rect 811 7931 857 8405
rect 995 7931 1041 8405
rect 1179 7931 1225 8405
rect 1363 7931 1409 8405
rect 4823 7931 4869 8405
rect 5007 7931 5053 8405
rect 5191 7931 5237 8405
rect 5375 7931 5421 8405
rect 8865 7931 8911 8405
rect 9049 7931 9095 8405
rect 9233 7931 9279 8405
rect 9417 7931 9463 8405
rect 12907 7931 12953 8405
rect 13091 7931 13137 8405
rect 13275 7931 13321 8405
rect 13459 7931 13505 8405
rect 16949 7931 16995 8405
rect 17133 7931 17179 8405
rect 17317 7931 17363 8405
rect 17501 7931 17547 8405
rect 20991 7931 21037 8405
rect 21175 7931 21221 8405
rect 21359 7931 21405 8405
rect 21543 7931 21589 8405
rect 25033 7931 25079 8405
rect 25217 7931 25263 8405
rect 25401 7931 25447 8405
rect 25585 7931 25631 8405
rect 811 5726 857 6200
rect 995 5726 1041 6200
rect 1179 5726 1225 6200
rect 1363 5726 1409 6200
rect 2297 5726 2343 6200
rect 2481 5726 2527 6200
rect 2665 5726 2711 6200
rect 2849 5726 2895 6200
rect 4823 5726 4869 6200
rect 5007 5726 5053 6200
rect 5191 5726 5237 6200
rect 5375 5726 5421 6200
rect 6309 5726 6355 6200
rect 6493 5726 6539 6200
rect 6677 5726 6723 6200
rect 6861 5726 6907 6200
rect 8865 5726 8911 6200
rect 9049 5726 9095 6200
rect 9233 5726 9279 6200
rect 9417 5726 9463 6200
rect 10351 5726 10397 6200
rect 10535 5726 10581 6200
rect 10719 5726 10765 6200
rect 10903 5726 10949 6200
rect 12907 5726 12953 6200
rect 13091 5726 13137 6200
rect 13275 5726 13321 6200
rect 13459 5726 13505 6200
rect 14393 5726 14439 6200
rect 14577 5726 14623 6200
rect 14761 5726 14807 6200
rect 14945 5726 14991 6200
rect 16949 5726 16995 6200
rect 17133 5726 17179 6200
rect 17317 5726 17363 6200
rect 17501 5726 17547 6200
rect 18435 5726 18481 6200
rect 18619 5726 18665 6200
rect 18803 5726 18849 6200
rect 18987 5726 19033 6200
rect 20991 5726 21037 6200
rect 21175 5726 21221 6200
rect 21359 5726 21405 6200
rect 21543 5726 21589 6200
rect 22477 5726 22523 6200
rect 22661 5726 22707 6200
rect 22845 5726 22891 6200
rect 23029 5726 23075 6200
rect 25033 5726 25079 6200
rect 25217 5726 25263 6200
rect 25401 5726 25447 6200
rect 25585 5726 25631 6200
rect 26519 5726 26565 6200
rect 26703 5726 26749 6200
rect 26887 5726 26933 6200
rect 27071 5726 27117 6200
rect 811 3521 857 3995
rect 995 3521 1041 3995
rect 1179 3521 1225 3995
rect 1363 3521 1409 3995
rect 2297 3522 2343 3996
rect 2481 3522 2527 3996
rect 2665 3522 2711 3996
rect 2849 3522 2895 3996
rect 4823 3521 4869 3995
rect 5007 3521 5053 3995
rect 5191 3521 5237 3995
rect 5375 3521 5421 3995
rect 6309 3522 6355 3996
rect 6493 3522 6539 3996
rect 6677 3522 6723 3996
rect 6861 3522 6907 3996
rect 8865 3521 8911 3995
rect 9049 3521 9095 3995
rect 9233 3521 9279 3995
rect 9417 3521 9463 3995
rect 10351 3522 10397 3996
rect 10535 3522 10581 3996
rect 10719 3522 10765 3996
rect 10903 3522 10949 3996
rect 12907 3521 12953 3995
rect 13091 3521 13137 3995
rect 13275 3521 13321 3995
rect 13459 3521 13505 3995
rect 14393 3522 14439 3996
rect 14577 3522 14623 3996
rect 14761 3522 14807 3996
rect 14945 3522 14991 3996
rect 16949 3521 16995 3995
rect 17133 3521 17179 3995
rect 17317 3521 17363 3995
rect 17501 3521 17547 3995
rect 18435 3522 18481 3996
rect 18619 3522 18665 3996
rect 18803 3522 18849 3996
rect 18987 3522 19033 3996
rect 20991 3521 21037 3995
rect 21175 3521 21221 3995
rect 21359 3521 21405 3995
rect 21543 3521 21589 3995
rect 22477 3522 22523 3996
rect 22661 3522 22707 3996
rect 22845 3522 22891 3996
rect 23029 3522 23075 3996
rect 25033 3521 25079 3995
rect 25217 3521 25263 3995
rect 25401 3521 25447 3995
rect 25585 3521 25631 3995
rect 26519 3522 26565 3996
rect 26703 3522 26749 3996
rect 26887 3522 26933 3996
rect 27071 3522 27117 3996
rect 811 1316 857 1790
rect 995 1316 1041 1790
rect 1179 1316 1225 1790
rect 1363 1316 1409 1790
rect 4823 1316 4869 1790
rect 5007 1316 5053 1790
rect 5191 1316 5237 1790
rect 5375 1316 5421 1790
rect 8865 1316 8911 1790
rect 9049 1316 9095 1790
rect 9233 1316 9279 1790
rect 9417 1316 9463 1790
rect 12907 1316 12953 1790
rect 13091 1316 13137 1790
rect 13275 1316 13321 1790
rect 13459 1316 13505 1790
rect 16949 1316 16995 1790
rect 17133 1316 17179 1790
rect 17317 1316 17363 1790
rect 17501 1316 17547 1790
rect 20991 1316 21037 1790
rect 21175 1316 21221 1790
rect 21359 1316 21405 1790
rect 21543 1316 21589 1790
rect 25033 1316 25079 1790
rect 25217 1316 25263 1790
rect 25401 1316 25447 1790
rect 25585 1316 25631 1790
<< psubdiff >>
rect 4672 16951 5572 17023
rect 4672 16907 4744 16951
rect 4672 16567 4685 16907
rect 4731 16567 4744 16907
rect 5500 16907 5572 16951
rect 4672 16523 4744 16567
rect 5500 16567 5513 16907
rect 5559 16567 5572 16907
rect 5500 16523 5572 16567
rect 4672 16451 5572 16523
rect 8714 16948 9614 17020
rect 8714 16904 8786 16948
rect 8714 16564 8727 16904
rect 8773 16564 8786 16904
rect 9542 16904 9614 16948
rect 8714 16520 8786 16564
rect 9542 16564 9555 16904
rect 9601 16564 9614 16904
rect 9542 16520 9614 16564
rect 8714 16448 9614 16520
rect 12756 16948 13656 17020
rect 12756 16904 12828 16948
rect 12756 16564 12769 16904
rect 12815 16564 12828 16904
rect 13584 16904 13656 16948
rect 12756 16520 12828 16564
rect 13584 16564 13597 16904
rect 13643 16564 13656 16904
rect 13584 16520 13656 16564
rect 12756 16448 13656 16520
rect 16798 16948 17698 17020
rect 16798 16904 16870 16948
rect 16798 16564 16811 16904
rect 16857 16564 16870 16904
rect 17626 16904 17698 16948
rect 16798 16520 16870 16564
rect 17626 16564 17639 16904
rect 17685 16564 17698 16904
rect 17626 16520 17698 16564
rect 16798 16448 17698 16520
rect 20840 16948 21740 17020
rect 20840 16904 20912 16948
rect 20840 16564 20853 16904
rect 20899 16564 20912 16904
rect 21668 16904 21740 16948
rect 20840 16520 20912 16564
rect 21668 16564 21681 16904
rect 21727 16564 21740 16904
rect 21668 16520 21740 16564
rect 20840 16448 21740 16520
rect 24882 16948 25782 17020
rect 24882 16904 24954 16948
rect 24882 16564 24895 16904
rect 24941 16564 24954 16904
rect 25710 16904 25782 16948
rect 24882 16520 24954 16564
rect 25710 16564 25723 16904
rect 25769 16564 25782 16904
rect 25710 16520 25782 16564
rect 24882 16448 25782 16520
rect 28924 16948 29824 17020
rect 28924 16904 28996 16948
rect 28924 16564 28937 16904
rect 28983 16564 28996 16904
rect 29752 16904 29824 16948
rect 28924 16520 28996 16564
rect 29752 16564 29765 16904
rect 29811 16564 29824 16904
rect 29752 16520 29824 16564
rect 28924 16448 29824 16520
rect 4672 14746 5572 14818
rect 4672 14702 4744 14746
rect 4672 14362 4685 14702
rect 4731 14362 4744 14702
rect 5500 14702 5572 14746
rect 4672 14318 4744 14362
rect 5500 14362 5513 14702
rect 5559 14362 5572 14702
rect 5500 14318 5572 14362
rect 4672 14246 5572 14318
rect 6158 14746 7058 14818
rect 6158 14702 6230 14746
rect 6158 14362 6171 14702
rect 6217 14362 6230 14702
rect 6986 14702 7058 14746
rect 6158 14318 6230 14362
rect 6986 14362 6999 14702
rect 7045 14362 7058 14702
rect 6986 14318 7058 14362
rect 6158 14246 7058 14318
rect 8714 14743 9614 14815
rect 8714 14699 8786 14743
rect 8714 14359 8727 14699
rect 8773 14359 8786 14699
rect 9542 14699 9614 14743
rect 8714 14315 8786 14359
rect 9542 14359 9555 14699
rect 9601 14359 9614 14699
rect 9542 14315 9614 14359
rect 8714 14243 9614 14315
rect 10200 14743 11100 14815
rect 10200 14699 10272 14743
rect 10200 14359 10213 14699
rect 10259 14359 10272 14699
rect 11028 14699 11100 14743
rect 10200 14315 10272 14359
rect 11028 14359 11041 14699
rect 11087 14359 11100 14699
rect 11028 14315 11100 14359
rect 10200 14243 11100 14315
rect 12756 14743 13656 14815
rect 12756 14699 12828 14743
rect 12756 14359 12769 14699
rect 12815 14359 12828 14699
rect 13584 14699 13656 14743
rect 12756 14315 12828 14359
rect 13584 14359 13597 14699
rect 13643 14359 13656 14699
rect 13584 14315 13656 14359
rect 12756 14243 13656 14315
rect 14242 14743 15142 14815
rect 14242 14699 14314 14743
rect 14242 14359 14255 14699
rect 14301 14359 14314 14699
rect 15070 14699 15142 14743
rect 14242 14315 14314 14359
rect 15070 14359 15083 14699
rect 15129 14359 15142 14699
rect 15070 14315 15142 14359
rect 14242 14243 15142 14315
rect 16798 14743 17698 14815
rect 16798 14699 16870 14743
rect 16798 14359 16811 14699
rect 16857 14359 16870 14699
rect 17626 14699 17698 14743
rect 16798 14315 16870 14359
rect 17626 14359 17639 14699
rect 17685 14359 17698 14699
rect 17626 14315 17698 14359
rect 16798 14243 17698 14315
rect 18284 14743 19184 14815
rect 18284 14699 18356 14743
rect 18284 14359 18297 14699
rect 18343 14359 18356 14699
rect 19112 14699 19184 14743
rect 18284 14315 18356 14359
rect 19112 14359 19125 14699
rect 19171 14359 19184 14699
rect 19112 14315 19184 14359
rect 18284 14243 19184 14315
rect 20840 14743 21740 14815
rect 20840 14699 20912 14743
rect 20840 14359 20853 14699
rect 20899 14359 20912 14699
rect 21668 14699 21740 14743
rect 20840 14315 20912 14359
rect 21668 14359 21681 14699
rect 21727 14359 21740 14699
rect 21668 14315 21740 14359
rect 20840 14243 21740 14315
rect 22326 14743 23226 14815
rect 22326 14699 22398 14743
rect 22326 14359 22339 14699
rect 22385 14359 22398 14699
rect 23154 14699 23226 14743
rect 22326 14315 22398 14359
rect 23154 14359 23167 14699
rect 23213 14359 23226 14699
rect 23154 14315 23226 14359
rect 22326 14243 23226 14315
rect 24882 14743 25782 14815
rect 24882 14699 24954 14743
rect 24882 14359 24895 14699
rect 24941 14359 24954 14699
rect 25710 14699 25782 14743
rect 24882 14315 24954 14359
rect 25710 14359 25723 14699
rect 25769 14359 25782 14699
rect 25710 14315 25782 14359
rect 24882 14243 25782 14315
rect 26368 14743 27268 14815
rect 26368 14699 26440 14743
rect 26368 14359 26381 14699
rect 26427 14359 26440 14699
rect 27196 14699 27268 14743
rect 26368 14315 26440 14359
rect 27196 14359 27209 14699
rect 27255 14359 27268 14699
rect 27196 14315 27268 14359
rect 26368 14243 27268 14315
rect 28924 14743 29824 14815
rect 28924 14699 28996 14743
rect 28924 14359 28937 14699
rect 28983 14359 28996 14699
rect 29752 14699 29824 14743
rect 28924 14315 28996 14359
rect 29752 14359 29765 14699
rect 29811 14359 29824 14699
rect 29752 14315 29824 14359
rect 28924 14243 29824 14315
rect 30410 14743 31310 14815
rect 30410 14699 30482 14743
rect 30410 14359 30423 14699
rect 30469 14359 30482 14699
rect 31238 14699 31310 14743
rect 30410 14315 30482 14359
rect 31238 14359 31251 14699
rect 31297 14359 31310 14699
rect 31238 14315 31310 14359
rect 30410 14243 31310 14315
rect 4672 12541 5572 12613
rect 4672 12497 4744 12541
rect 4672 12157 4685 12497
rect 4731 12157 4744 12497
rect 5500 12497 5572 12541
rect 4672 12113 4744 12157
rect 5500 12157 5513 12497
rect 5559 12157 5572 12497
rect 5500 12113 5572 12157
rect 4672 12041 5572 12113
rect 6158 12542 7058 12614
rect 6158 12498 6230 12542
rect 6158 12158 6171 12498
rect 6217 12158 6230 12498
rect 6986 12498 7058 12542
rect 6158 12114 6230 12158
rect 6986 12158 6999 12498
rect 7045 12158 7058 12498
rect 6986 12114 7058 12158
rect 6158 12042 7058 12114
rect 8714 12538 9614 12610
rect 8714 12494 8786 12538
rect 8714 12154 8727 12494
rect 8773 12154 8786 12494
rect 9542 12494 9614 12538
rect 8714 12110 8786 12154
rect 9542 12154 9555 12494
rect 9601 12154 9614 12494
rect 9542 12110 9614 12154
rect 8714 12038 9614 12110
rect 10200 12539 11100 12611
rect 10200 12495 10272 12539
rect 10200 12155 10213 12495
rect 10259 12155 10272 12495
rect 11028 12495 11100 12539
rect 10200 12111 10272 12155
rect 11028 12155 11041 12495
rect 11087 12155 11100 12495
rect 11028 12111 11100 12155
rect 10200 12039 11100 12111
rect 12756 12538 13656 12610
rect 12756 12494 12828 12538
rect 12756 12154 12769 12494
rect 12815 12154 12828 12494
rect 13584 12494 13656 12538
rect 12756 12110 12828 12154
rect 13584 12154 13597 12494
rect 13643 12154 13656 12494
rect 13584 12110 13656 12154
rect 12756 12038 13656 12110
rect 14242 12539 15142 12611
rect 14242 12495 14314 12539
rect 14242 12155 14255 12495
rect 14301 12155 14314 12495
rect 15070 12495 15142 12539
rect 14242 12111 14314 12155
rect 15070 12155 15083 12495
rect 15129 12155 15142 12495
rect 15070 12111 15142 12155
rect 14242 12039 15142 12111
rect 16798 12538 17698 12610
rect 16798 12494 16870 12538
rect 16798 12154 16811 12494
rect 16857 12154 16870 12494
rect 17626 12494 17698 12538
rect 16798 12110 16870 12154
rect 17626 12154 17639 12494
rect 17685 12154 17698 12494
rect 17626 12110 17698 12154
rect 16798 12038 17698 12110
rect 18284 12539 19184 12611
rect 18284 12495 18356 12539
rect 18284 12155 18297 12495
rect 18343 12155 18356 12495
rect 19112 12495 19184 12539
rect 18284 12111 18356 12155
rect 19112 12155 19125 12495
rect 19171 12155 19184 12495
rect 19112 12111 19184 12155
rect 18284 12039 19184 12111
rect 20840 12538 21740 12610
rect 20840 12494 20912 12538
rect 20840 12154 20853 12494
rect 20899 12154 20912 12494
rect 21668 12494 21740 12538
rect 20840 12110 20912 12154
rect 21668 12154 21681 12494
rect 21727 12154 21740 12494
rect 21668 12110 21740 12154
rect 20840 12038 21740 12110
rect 22326 12539 23226 12611
rect 22326 12495 22398 12539
rect 22326 12155 22339 12495
rect 22385 12155 22398 12495
rect 23154 12495 23226 12539
rect 22326 12111 22398 12155
rect 23154 12155 23167 12495
rect 23213 12155 23226 12495
rect 23154 12111 23226 12155
rect 22326 12039 23226 12111
rect 24882 12538 25782 12610
rect 24882 12494 24954 12538
rect 24882 12154 24895 12494
rect 24941 12154 24954 12494
rect 25710 12494 25782 12538
rect 24882 12110 24954 12154
rect 25710 12154 25723 12494
rect 25769 12154 25782 12494
rect 25710 12110 25782 12154
rect 24882 12038 25782 12110
rect 26368 12539 27268 12611
rect 26368 12495 26440 12539
rect 26368 12155 26381 12495
rect 26427 12155 26440 12495
rect 27196 12495 27268 12539
rect 26368 12111 26440 12155
rect 27196 12155 27209 12495
rect 27255 12155 27268 12495
rect 27196 12111 27268 12155
rect 26368 12039 27268 12111
rect 28924 12538 29824 12610
rect 28924 12494 28996 12538
rect 28924 12154 28937 12494
rect 28983 12154 28996 12494
rect 29752 12494 29824 12538
rect 28924 12110 28996 12154
rect 29752 12154 29765 12494
rect 29811 12154 29824 12494
rect 29752 12110 29824 12154
rect 28924 12038 29824 12110
rect 30410 12539 31310 12611
rect 30410 12495 30482 12539
rect 30410 12155 30423 12495
rect 30469 12155 30482 12495
rect 31238 12495 31310 12539
rect 30410 12111 30482 12155
rect 31238 12155 31251 12495
rect 31297 12155 31310 12495
rect 31238 12111 31310 12155
rect 30410 12039 31310 12111
rect 4672 10336 5572 10408
rect 4672 10292 4744 10336
rect 4672 9952 4685 10292
rect 4731 9952 4744 10292
rect 5500 10292 5572 10336
rect 4672 9908 4744 9952
rect 5500 9952 5513 10292
rect 5559 9952 5572 10292
rect 5500 9908 5572 9952
rect 4672 9836 5572 9908
rect 8714 10333 9614 10405
rect 8714 10289 8786 10333
rect 8714 9949 8727 10289
rect 8773 9949 8786 10289
rect 9542 10289 9614 10333
rect 8714 9905 8786 9949
rect 9542 9949 9555 10289
rect 9601 9949 9614 10289
rect 9542 9905 9614 9949
rect 8714 9833 9614 9905
rect 12756 10333 13656 10405
rect 12756 10289 12828 10333
rect 12756 9949 12769 10289
rect 12815 9949 12828 10289
rect 13584 10289 13656 10333
rect 12756 9905 12828 9949
rect 13584 9949 13597 10289
rect 13643 9949 13656 10289
rect 13584 9905 13656 9949
rect 12756 9833 13656 9905
rect 16798 10333 17698 10405
rect 16798 10289 16870 10333
rect 16798 9949 16811 10289
rect 16857 9949 16870 10289
rect 17626 10289 17698 10333
rect 16798 9905 16870 9949
rect 17626 9949 17639 10289
rect 17685 9949 17698 10289
rect 17626 9905 17698 9949
rect 16798 9833 17698 9905
rect 20840 10333 21740 10405
rect 20840 10289 20912 10333
rect 20840 9949 20853 10289
rect 20899 9949 20912 10289
rect 21668 10289 21740 10333
rect 20840 9905 20912 9949
rect 21668 9949 21681 10289
rect 21727 9949 21740 10289
rect 21668 9905 21740 9949
rect 20840 9833 21740 9905
rect 24882 10333 25782 10405
rect 24882 10289 24954 10333
rect 24882 9949 24895 10289
rect 24941 9949 24954 10289
rect 25710 10289 25782 10333
rect 24882 9905 24954 9949
rect 25710 9949 25723 10289
rect 25769 9949 25782 10289
rect 25710 9905 25782 9949
rect 24882 9833 25782 9905
rect 28924 10333 29824 10405
rect 28924 10289 28996 10333
rect 28924 9949 28937 10289
rect 28983 9949 28996 10289
rect 29752 10289 29824 10333
rect 28924 9905 28996 9949
rect 29752 9949 29765 10289
rect 29811 9949 29824 10289
rect 29752 9905 29824 9949
rect 28924 9833 29824 9905
rect 660 7372 1560 7444
rect 660 7328 732 7372
rect 660 6988 673 7328
rect 719 6988 732 7328
rect 1488 7328 1560 7372
rect 660 6944 732 6988
rect 1488 6988 1501 7328
rect 1547 6988 1560 7328
rect 1488 6944 1560 6988
rect 660 6872 1560 6944
rect 4672 7372 5572 7444
rect 4672 7328 4744 7372
rect 4672 6988 4685 7328
rect 4731 6988 4744 7328
rect 5500 7328 5572 7372
rect 4672 6944 4744 6988
rect 5500 6988 5513 7328
rect 5559 6988 5572 7328
rect 5500 6944 5572 6988
rect 4672 6872 5572 6944
rect 8714 7372 9614 7444
rect 8714 7328 8786 7372
rect 8714 6988 8727 7328
rect 8773 6988 8786 7328
rect 9542 7328 9614 7372
rect 8714 6944 8786 6988
rect 9542 6988 9555 7328
rect 9601 6988 9614 7328
rect 9542 6944 9614 6988
rect 8714 6872 9614 6944
rect 12756 7372 13656 7444
rect 12756 7328 12828 7372
rect 12756 6988 12769 7328
rect 12815 6988 12828 7328
rect 13584 7328 13656 7372
rect 12756 6944 12828 6988
rect 13584 6988 13597 7328
rect 13643 6988 13656 7328
rect 13584 6944 13656 6988
rect 12756 6872 13656 6944
rect 16798 7372 17698 7444
rect 16798 7328 16870 7372
rect 16798 6988 16811 7328
rect 16857 6988 16870 7328
rect 17626 7328 17698 7372
rect 16798 6944 16870 6988
rect 17626 6988 17639 7328
rect 17685 6988 17698 7328
rect 17626 6944 17698 6988
rect 16798 6872 17698 6944
rect 20840 7372 21740 7444
rect 20840 7328 20912 7372
rect 20840 6988 20853 7328
rect 20899 6988 20912 7328
rect 21668 7328 21740 7372
rect 20840 6944 20912 6988
rect 21668 6988 21681 7328
rect 21727 6988 21740 7328
rect 21668 6944 21740 6988
rect 20840 6872 21740 6944
rect 24882 7372 25782 7444
rect 24882 7328 24954 7372
rect 24882 6988 24895 7328
rect 24941 6988 24954 7328
rect 25710 7328 25782 7372
rect 24882 6944 24954 6988
rect 25710 6988 25723 7328
rect 25769 6988 25782 7328
rect 25710 6944 25782 6988
rect 24882 6872 25782 6944
rect 660 5167 1560 5239
rect 660 5123 732 5167
rect 660 4783 673 5123
rect 719 4783 732 5123
rect 1488 5123 1560 5167
rect 660 4739 732 4783
rect 1488 4783 1501 5123
rect 1547 4783 1560 5123
rect 1488 4739 1560 4783
rect 660 4667 1560 4739
rect 2146 5167 3046 5239
rect 2146 5123 2218 5167
rect 2146 4783 2159 5123
rect 2205 4783 2218 5123
rect 2974 5123 3046 5167
rect 2146 4739 2218 4783
rect 2974 4783 2987 5123
rect 3033 4783 3046 5123
rect 2974 4739 3046 4783
rect 2146 4667 3046 4739
rect 4672 5167 5572 5239
rect 4672 5123 4744 5167
rect 4672 4783 4685 5123
rect 4731 4783 4744 5123
rect 5500 5123 5572 5167
rect 4672 4739 4744 4783
rect 5500 4783 5513 5123
rect 5559 4783 5572 5123
rect 5500 4739 5572 4783
rect 4672 4667 5572 4739
rect 6158 5167 7058 5239
rect 6158 5123 6230 5167
rect 6158 4783 6171 5123
rect 6217 4783 6230 5123
rect 6986 5123 7058 5167
rect 6158 4739 6230 4783
rect 6986 4783 6999 5123
rect 7045 4783 7058 5123
rect 6986 4739 7058 4783
rect 6158 4667 7058 4739
rect 8714 5167 9614 5239
rect 8714 5123 8786 5167
rect 8714 4783 8727 5123
rect 8773 4783 8786 5123
rect 9542 5123 9614 5167
rect 8714 4739 8786 4783
rect 9542 4783 9555 5123
rect 9601 4783 9614 5123
rect 9542 4739 9614 4783
rect 8714 4667 9614 4739
rect 10200 5167 11100 5239
rect 10200 5123 10272 5167
rect 10200 4783 10213 5123
rect 10259 4783 10272 5123
rect 11028 5123 11100 5167
rect 10200 4739 10272 4783
rect 11028 4783 11041 5123
rect 11087 4783 11100 5123
rect 11028 4739 11100 4783
rect 10200 4667 11100 4739
rect 12756 5167 13656 5239
rect 12756 5123 12828 5167
rect 12756 4783 12769 5123
rect 12815 4783 12828 5123
rect 13584 5123 13656 5167
rect 12756 4739 12828 4783
rect 13584 4783 13597 5123
rect 13643 4783 13656 5123
rect 13584 4739 13656 4783
rect 12756 4667 13656 4739
rect 14242 5167 15142 5239
rect 14242 5123 14314 5167
rect 14242 4783 14255 5123
rect 14301 4783 14314 5123
rect 15070 5123 15142 5167
rect 14242 4739 14314 4783
rect 15070 4783 15083 5123
rect 15129 4783 15142 5123
rect 15070 4739 15142 4783
rect 14242 4667 15142 4739
rect 16798 5167 17698 5239
rect 16798 5123 16870 5167
rect 16798 4783 16811 5123
rect 16857 4783 16870 5123
rect 17626 5123 17698 5167
rect 16798 4739 16870 4783
rect 17626 4783 17639 5123
rect 17685 4783 17698 5123
rect 17626 4739 17698 4783
rect 16798 4667 17698 4739
rect 18284 5167 19184 5239
rect 18284 5123 18356 5167
rect 18284 4783 18297 5123
rect 18343 4783 18356 5123
rect 19112 5123 19184 5167
rect 18284 4739 18356 4783
rect 19112 4783 19125 5123
rect 19171 4783 19184 5123
rect 19112 4739 19184 4783
rect 18284 4667 19184 4739
rect 20840 5167 21740 5239
rect 20840 5123 20912 5167
rect 20840 4783 20853 5123
rect 20899 4783 20912 5123
rect 21668 5123 21740 5167
rect 20840 4739 20912 4783
rect 21668 4783 21681 5123
rect 21727 4783 21740 5123
rect 21668 4739 21740 4783
rect 20840 4667 21740 4739
rect 22326 5167 23226 5239
rect 22326 5123 22398 5167
rect 22326 4783 22339 5123
rect 22385 4783 22398 5123
rect 23154 5123 23226 5167
rect 22326 4739 22398 4783
rect 23154 4783 23167 5123
rect 23213 4783 23226 5123
rect 23154 4739 23226 4783
rect 22326 4667 23226 4739
rect 24882 5167 25782 5239
rect 24882 5123 24954 5167
rect 24882 4783 24895 5123
rect 24941 4783 24954 5123
rect 25710 5123 25782 5167
rect 24882 4739 24954 4783
rect 25710 4783 25723 5123
rect 25769 4783 25782 5123
rect 25710 4739 25782 4783
rect 24882 4667 25782 4739
rect 26368 5167 27268 5239
rect 26368 5123 26440 5167
rect 26368 4783 26381 5123
rect 26427 4783 26440 5123
rect 27196 5123 27268 5167
rect 26368 4739 26440 4783
rect 27196 4783 27209 5123
rect 27255 4783 27268 5123
rect 27196 4739 27268 4783
rect 26368 4667 27268 4739
rect 660 2962 1560 3034
rect 660 2918 732 2962
rect 660 2578 673 2918
rect 719 2578 732 2918
rect 1488 2918 1560 2962
rect 660 2534 732 2578
rect 1488 2578 1501 2918
rect 1547 2578 1560 2918
rect 1488 2534 1560 2578
rect 660 2462 1560 2534
rect 2146 2963 3046 3035
rect 2146 2919 2218 2963
rect 2146 2579 2159 2919
rect 2205 2579 2218 2919
rect 2974 2919 3046 2963
rect 2146 2535 2218 2579
rect 2974 2579 2987 2919
rect 3033 2579 3046 2919
rect 2974 2535 3046 2579
rect 2146 2463 3046 2535
rect 4672 2962 5572 3034
rect 4672 2918 4744 2962
rect 4672 2578 4685 2918
rect 4731 2578 4744 2918
rect 5500 2918 5572 2962
rect 4672 2534 4744 2578
rect 5500 2578 5513 2918
rect 5559 2578 5572 2918
rect 5500 2534 5572 2578
rect 4672 2462 5572 2534
rect 6158 2963 7058 3035
rect 6158 2919 6230 2963
rect 6158 2579 6171 2919
rect 6217 2579 6230 2919
rect 6986 2919 7058 2963
rect 6158 2535 6230 2579
rect 6986 2579 6999 2919
rect 7045 2579 7058 2919
rect 6986 2535 7058 2579
rect 6158 2463 7058 2535
rect 8714 2962 9614 3034
rect 8714 2918 8786 2962
rect 8714 2578 8727 2918
rect 8773 2578 8786 2918
rect 9542 2918 9614 2962
rect 8714 2534 8786 2578
rect 9542 2578 9555 2918
rect 9601 2578 9614 2918
rect 9542 2534 9614 2578
rect 8714 2462 9614 2534
rect 10200 2963 11100 3035
rect 10200 2919 10272 2963
rect 10200 2579 10213 2919
rect 10259 2579 10272 2919
rect 11028 2919 11100 2963
rect 10200 2535 10272 2579
rect 11028 2579 11041 2919
rect 11087 2579 11100 2919
rect 11028 2535 11100 2579
rect 10200 2463 11100 2535
rect 12756 2962 13656 3034
rect 12756 2918 12828 2962
rect 12756 2578 12769 2918
rect 12815 2578 12828 2918
rect 13584 2918 13656 2962
rect 12756 2534 12828 2578
rect 13584 2578 13597 2918
rect 13643 2578 13656 2918
rect 13584 2534 13656 2578
rect 12756 2462 13656 2534
rect 14242 2963 15142 3035
rect 14242 2919 14314 2963
rect 14242 2579 14255 2919
rect 14301 2579 14314 2919
rect 15070 2919 15142 2963
rect 14242 2535 14314 2579
rect 15070 2579 15083 2919
rect 15129 2579 15142 2919
rect 15070 2535 15142 2579
rect 14242 2463 15142 2535
rect 16798 2962 17698 3034
rect 16798 2918 16870 2962
rect 16798 2578 16811 2918
rect 16857 2578 16870 2918
rect 17626 2918 17698 2962
rect 16798 2534 16870 2578
rect 17626 2578 17639 2918
rect 17685 2578 17698 2918
rect 17626 2534 17698 2578
rect 16798 2462 17698 2534
rect 18284 2963 19184 3035
rect 18284 2919 18356 2963
rect 18284 2579 18297 2919
rect 18343 2579 18356 2919
rect 19112 2919 19184 2963
rect 18284 2535 18356 2579
rect 19112 2579 19125 2919
rect 19171 2579 19184 2919
rect 19112 2535 19184 2579
rect 18284 2463 19184 2535
rect 20840 2962 21740 3034
rect 20840 2918 20912 2962
rect 20840 2578 20853 2918
rect 20899 2578 20912 2918
rect 21668 2918 21740 2962
rect 20840 2534 20912 2578
rect 21668 2578 21681 2918
rect 21727 2578 21740 2918
rect 21668 2534 21740 2578
rect 20840 2462 21740 2534
rect 22326 2963 23226 3035
rect 22326 2919 22398 2963
rect 22326 2579 22339 2919
rect 22385 2579 22398 2919
rect 23154 2919 23226 2963
rect 22326 2535 22398 2579
rect 23154 2579 23167 2919
rect 23213 2579 23226 2919
rect 23154 2535 23226 2579
rect 22326 2463 23226 2535
rect 24882 2962 25782 3034
rect 24882 2918 24954 2962
rect 24882 2578 24895 2918
rect 24941 2578 24954 2918
rect 25710 2918 25782 2962
rect 24882 2534 24954 2578
rect 25710 2578 25723 2918
rect 25769 2578 25782 2918
rect 25710 2534 25782 2578
rect 24882 2462 25782 2534
rect 26368 2963 27268 3035
rect 26368 2919 26440 2963
rect 26368 2579 26381 2919
rect 26427 2579 26440 2919
rect 27196 2919 27268 2963
rect 26368 2535 26440 2579
rect 27196 2579 27209 2919
rect 27255 2579 27268 2919
rect 27196 2535 27268 2579
rect 26368 2463 27268 2535
rect 660 757 1560 829
rect 660 713 732 757
rect 660 373 673 713
rect 719 373 732 713
rect 1488 713 1560 757
rect 660 329 732 373
rect 1488 373 1501 713
rect 1547 373 1560 713
rect 1488 329 1560 373
rect 660 257 1560 329
rect 4672 757 5572 829
rect 4672 713 4744 757
rect 4672 373 4685 713
rect 4731 373 4744 713
rect 5500 713 5572 757
rect 4672 329 4744 373
rect 5500 373 5513 713
rect 5559 373 5572 713
rect 5500 329 5572 373
rect 4672 257 5572 329
rect 8714 757 9614 829
rect 8714 713 8786 757
rect 8714 373 8727 713
rect 8773 373 8786 713
rect 9542 713 9614 757
rect 8714 329 8786 373
rect 9542 373 9555 713
rect 9601 373 9614 713
rect 9542 329 9614 373
rect 8714 257 9614 329
rect 12756 757 13656 829
rect 12756 713 12828 757
rect 12756 373 12769 713
rect 12815 373 12828 713
rect 13584 713 13656 757
rect 12756 329 12828 373
rect 13584 373 13597 713
rect 13643 373 13656 713
rect 13584 329 13656 373
rect 12756 257 13656 329
rect 16798 757 17698 829
rect 16798 713 16870 757
rect 16798 373 16811 713
rect 16857 373 16870 713
rect 17626 713 17698 757
rect 16798 329 16870 373
rect 17626 373 17639 713
rect 17685 373 17698 713
rect 17626 329 17698 373
rect 16798 257 17698 329
rect 20840 757 21740 829
rect 20840 713 20912 757
rect 20840 373 20853 713
rect 20899 373 20912 713
rect 21668 713 21740 757
rect 20840 329 20912 373
rect 21668 373 21681 713
rect 21727 373 21740 713
rect 21668 329 21740 373
rect 20840 257 21740 329
rect 24882 757 25782 829
rect 24882 713 24954 757
rect 24882 373 24895 713
rect 24941 373 24954 713
rect 25710 713 25782 757
rect 24882 329 24954 373
rect 25710 373 25723 713
rect 25769 373 25782 713
rect 25710 329 25782 373
rect 24882 257 25782 329
<< nsubdiff >>
rect 4672 18111 5572 18183
rect 4672 18067 4744 18111
rect 4672 17427 4685 18067
rect 4731 17427 4744 18067
rect 5500 18067 5572 18111
rect 4672 17383 4744 17427
rect 5500 17427 5513 18067
rect 5559 17427 5572 18067
rect 5500 17383 5572 17427
rect 4672 17311 5572 17383
rect 8714 18108 9614 18180
rect 8714 18064 8786 18108
rect 8714 17424 8727 18064
rect 8773 17424 8786 18064
rect 9542 18064 9614 18108
rect 8714 17380 8786 17424
rect 9542 17424 9555 18064
rect 9601 17424 9614 18064
rect 9542 17380 9614 17424
rect 8714 17308 9614 17380
rect 12756 18108 13656 18180
rect 12756 18064 12828 18108
rect 12756 17424 12769 18064
rect 12815 17424 12828 18064
rect 13584 18064 13656 18108
rect 12756 17380 12828 17424
rect 13584 17424 13597 18064
rect 13643 17424 13656 18064
rect 13584 17380 13656 17424
rect 12756 17308 13656 17380
rect 16798 18108 17698 18180
rect 16798 18064 16870 18108
rect 16798 17424 16811 18064
rect 16857 17424 16870 18064
rect 17626 18064 17698 18108
rect 16798 17380 16870 17424
rect 17626 17424 17639 18064
rect 17685 17424 17698 18064
rect 17626 17380 17698 17424
rect 16798 17308 17698 17380
rect 20840 18108 21740 18180
rect 20840 18064 20912 18108
rect 20840 17424 20853 18064
rect 20899 17424 20912 18064
rect 21668 18064 21740 18108
rect 20840 17380 20912 17424
rect 21668 17424 21681 18064
rect 21727 17424 21740 18064
rect 21668 17380 21740 17424
rect 20840 17308 21740 17380
rect 24882 18108 25782 18180
rect 24882 18064 24954 18108
rect 24882 17424 24895 18064
rect 24941 17424 24954 18064
rect 25710 18064 25782 18108
rect 24882 17380 24954 17424
rect 25710 17424 25723 18064
rect 25769 17424 25782 18064
rect 25710 17380 25782 17424
rect 24882 17308 25782 17380
rect 28924 18108 29824 18180
rect 28924 18064 28996 18108
rect 28924 17424 28937 18064
rect 28983 17424 28996 18064
rect 29752 18064 29824 18108
rect 28924 17380 28996 17424
rect 29752 17424 29765 18064
rect 29811 17424 29824 18064
rect 29752 17380 29824 17424
rect 28924 17308 29824 17380
rect 4672 15906 5572 15978
rect 4672 15862 4744 15906
rect 4672 15222 4685 15862
rect 4731 15222 4744 15862
rect 5500 15862 5572 15906
rect 4672 15178 4744 15222
rect 5500 15222 5513 15862
rect 5559 15222 5572 15862
rect 5500 15178 5572 15222
rect 4672 15106 5572 15178
rect 6158 15906 7058 15978
rect 6158 15862 6230 15906
rect 6158 15222 6171 15862
rect 6217 15222 6230 15862
rect 6986 15862 7058 15906
rect 6158 15178 6230 15222
rect 6986 15222 6999 15862
rect 7045 15222 7058 15862
rect 6986 15178 7058 15222
rect 6158 15106 7058 15178
rect 8714 15903 9614 15975
rect 8714 15859 8786 15903
rect 8714 15219 8727 15859
rect 8773 15219 8786 15859
rect 9542 15859 9614 15903
rect 8714 15175 8786 15219
rect 9542 15219 9555 15859
rect 9601 15219 9614 15859
rect 9542 15175 9614 15219
rect 8714 15103 9614 15175
rect 10200 15903 11100 15975
rect 10200 15859 10272 15903
rect 10200 15219 10213 15859
rect 10259 15219 10272 15859
rect 11028 15859 11100 15903
rect 10200 15175 10272 15219
rect 11028 15219 11041 15859
rect 11087 15219 11100 15859
rect 11028 15175 11100 15219
rect 10200 15103 11100 15175
rect 12756 15903 13656 15975
rect 12756 15859 12828 15903
rect 12756 15219 12769 15859
rect 12815 15219 12828 15859
rect 13584 15859 13656 15903
rect 12756 15175 12828 15219
rect 13584 15219 13597 15859
rect 13643 15219 13656 15859
rect 13584 15175 13656 15219
rect 12756 15103 13656 15175
rect 14242 15903 15142 15975
rect 14242 15859 14314 15903
rect 14242 15219 14255 15859
rect 14301 15219 14314 15859
rect 15070 15859 15142 15903
rect 14242 15175 14314 15219
rect 15070 15219 15083 15859
rect 15129 15219 15142 15859
rect 15070 15175 15142 15219
rect 14242 15103 15142 15175
rect 16798 15903 17698 15975
rect 16798 15859 16870 15903
rect 16798 15219 16811 15859
rect 16857 15219 16870 15859
rect 17626 15859 17698 15903
rect 16798 15175 16870 15219
rect 17626 15219 17639 15859
rect 17685 15219 17698 15859
rect 17626 15175 17698 15219
rect 16798 15103 17698 15175
rect 18284 15903 19184 15975
rect 18284 15859 18356 15903
rect 18284 15219 18297 15859
rect 18343 15219 18356 15859
rect 19112 15859 19184 15903
rect 18284 15175 18356 15219
rect 19112 15219 19125 15859
rect 19171 15219 19184 15859
rect 19112 15175 19184 15219
rect 18284 15103 19184 15175
rect 20840 15903 21740 15975
rect 20840 15859 20912 15903
rect 20840 15219 20853 15859
rect 20899 15219 20912 15859
rect 21668 15859 21740 15903
rect 20840 15175 20912 15219
rect 21668 15219 21681 15859
rect 21727 15219 21740 15859
rect 21668 15175 21740 15219
rect 20840 15103 21740 15175
rect 22326 15903 23226 15975
rect 22326 15859 22398 15903
rect 22326 15219 22339 15859
rect 22385 15219 22398 15859
rect 23154 15859 23226 15903
rect 22326 15175 22398 15219
rect 23154 15219 23167 15859
rect 23213 15219 23226 15859
rect 23154 15175 23226 15219
rect 22326 15103 23226 15175
rect 24882 15903 25782 15975
rect 24882 15859 24954 15903
rect 24882 15219 24895 15859
rect 24941 15219 24954 15859
rect 25710 15859 25782 15903
rect 24882 15175 24954 15219
rect 25710 15219 25723 15859
rect 25769 15219 25782 15859
rect 25710 15175 25782 15219
rect 24882 15103 25782 15175
rect 26368 15903 27268 15975
rect 26368 15859 26440 15903
rect 26368 15219 26381 15859
rect 26427 15219 26440 15859
rect 27196 15859 27268 15903
rect 26368 15175 26440 15219
rect 27196 15219 27209 15859
rect 27255 15219 27268 15859
rect 27196 15175 27268 15219
rect 26368 15103 27268 15175
rect 28924 15903 29824 15975
rect 28924 15859 28996 15903
rect 28924 15219 28937 15859
rect 28983 15219 28996 15859
rect 29752 15859 29824 15903
rect 28924 15175 28996 15219
rect 29752 15219 29765 15859
rect 29811 15219 29824 15859
rect 29752 15175 29824 15219
rect 28924 15103 29824 15175
rect 30410 15903 31310 15975
rect 30410 15859 30482 15903
rect 30410 15219 30423 15859
rect 30469 15219 30482 15859
rect 31238 15859 31310 15903
rect 30410 15175 30482 15219
rect 31238 15219 31251 15859
rect 31297 15219 31310 15859
rect 31238 15175 31310 15219
rect 30410 15103 31310 15175
rect 4672 13701 5572 13773
rect 4672 13657 4744 13701
rect 4672 13017 4685 13657
rect 4731 13017 4744 13657
rect 5500 13657 5572 13701
rect 4672 12973 4744 13017
rect 5500 13017 5513 13657
rect 5559 13017 5572 13657
rect 5500 12973 5572 13017
rect 4672 12901 5572 12973
rect 6158 13702 7058 13774
rect 6158 13658 6230 13702
rect 6158 13018 6171 13658
rect 6217 13018 6230 13658
rect 6986 13658 7058 13702
rect 6158 12974 6230 13018
rect 6986 13018 6999 13658
rect 7045 13018 7058 13658
rect 6986 12974 7058 13018
rect 6158 12902 7058 12974
rect 8714 13698 9614 13770
rect 8714 13654 8786 13698
rect 8714 13014 8727 13654
rect 8773 13014 8786 13654
rect 9542 13654 9614 13698
rect 8714 12970 8786 13014
rect 9542 13014 9555 13654
rect 9601 13014 9614 13654
rect 9542 12970 9614 13014
rect 8714 12898 9614 12970
rect 10200 13699 11100 13771
rect 10200 13655 10272 13699
rect 10200 13015 10213 13655
rect 10259 13015 10272 13655
rect 11028 13655 11100 13699
rect 10200 12971 10272 13015
rect 11028 13015 11041 13655
rect 11087 13015 11100 13655
rect 11028 12971 11100 13015
rect 10200 12899 11100 12971
rect 12756 13698 13656 13770
rect 12756 13654 12828 13698
rect 12756 13014 12769 13654
rect 12815 13014 12828 13654
rect 13584 13654 13656 13698
rect 12756 12970 12828 13014
rect 13584 13014 13597 13654
rect 13643 13014 13656 13654
rect 13584 12970 13656 13014
rect 12756 12898 13656 12970
rect 14242 13699 15142 13771
rect 14242 13655 14314 13699
rect 14242 13015 14255 13655
rect 14301 13015 14314 13655
rect 15070 13655 15142 13699
rect 14242 12971 14314 13015
rect 15070 13015 15083 13655
rect 15129 13015 15142 13655
rect 15070 12971 15142 13015
rect 14242 12899 15142 12971
rect 16798 13698 17698 13770
rect 16798 13654 16870 13698
rect 16798 13014 16811 13654
rect 16857 13014 16870 13654
rect 17626 13654 17698 13698
rect 16798 12970 16870 13014
rect 17626 13014 17639 13654
rect 17685 13014 17698 13654
rect 17626 12970 17698 13014
rect 16798 12898 17698 12970
rect 18284 13699 19184 13771
rect 18284 13655 18356 13699
rect 18284 13015 18297 13655
rect 18343 13015 18356 13655
rect 19112 13655 19184 13699
rect 18284 12971 18356 13015
rect 19112 13015 19125 13655
rect 19171 13015 19184 13655
rect 19112 12971 19184 13015
rect 18284 12899 19184 12971
rect 20840 13698 21740 13770
rect 20840 13654 20912 13698
rect 20840 13014 20853 13654
rect 20899 13014 20912 13654
rect 21668 13654 21740 13698
rect 20840 12970 20912 13014
rect 21668 13014 21681 13654
rect 21727 13014 21740 13654
rect 21668 12970 21740 13014
rect 20840 12898 21740 12970
rect 22326 13699 23226 13771
rect 22326 13655 22398 13699
rect 22326 13015 22339 13655
rect 22385 13015 22398 13655
rect 23154 13655 23226 13699
rect 22326 12971 22398 13015
rect 23154 13015 23167 13655
rect 23213 13015 23226 13655
rect 23154 12971 23226 13015
rect 22326 12899 23226 12971
rect 24882 13698 25782 13770
rect 24882 13654 24954 13698
rect 24882 13014 24895 13654
rect 24941 13014 24954 13654
rect 25710 13654 25782 13698
rect 24882 12970 24954 13014
rect 25710 13014 25723 13654
rect 25769 13014 25782 13654
rect 25710 12970 25782 13014
rect 24882 12898 25782 12970
rect 26368 13699 27268 13771
rect 26368 13655 26440 13699
rect 26368 13015 26381 13655
rect 26427 13015 26440 13655
rect 27196 13655 27268 13699
rect 26368 12971 26440 13015
rect 27196 13015 27209 13655
rect 27255 13015 27268 13655
rect 27196 12971 27268 13015
rect 26368 12899 27268 12971
rect 28924 13698 29824 13770
rect 28924 13654 28996 13698
rect 28924 13014 28937 13654
rect 28983 13014 28996 13654
rect 29752 13654 29824 13698
rect 28924 12970 28996 13014
rect 29752 13014 29765 13654
rect 29811 13014 29824 13654
rect 29752 12970 29824 13014
rect 28924 12898 29824 12970
rect 30410 13699 31310 13771
rect 30410 13655 30482 13699
rect 30410 13015 30423 13655
rect 30469 13015 30482 13655
rect 31238 13655 31310 13699
rect 30410 12971 30482 13015
rect 31238 13015 31251 13655
rect 31297 13015 31310 13655
rect 31238 12971 31310 13015
rect 30410 12899 31310 12971
rect 4672 11496 5572 11568
rect 4672 11452 4744 11496
rect 4672 10812 4685 11452
rect 4731 10812 4744 11452
rect 5500 11452 5572 11496
rect 4672 10768 4744 10812
rect 5500 10812 5513 11452
rect 5559 10812 5572 11452
rect 5500 10768 5572 10812
rect 4672 10696 5572 10768
rect 8714 11493 9614 11565
rect 8714 11449 8786 11493
rect 8714 10809 8727 11449
rect 8773 10809 8786 11449
rect 9542 11449 9614 11493
rect 8714 10765 8786 10809
rect 9542 10809 9555 11449
rect 9601 10809 9614 11449
rect 9542 10765 9614 10809
rect 8714 10693 9614 10765
rect 12756 11493 13656 11565
rect 12756 11449 12828 11493
rect 12756 10809 12769 11449
rect 12815 10809 12828 11449
rect 13584 11449 13656 11493
rect 12756 10765 12828 10809
rect 13584 10809 13597 11449
rect 13643 10809 13656 11449
rect 13584 10765 13656 10809
rect 12756 10693 13656 10765
rect 16798 11493 17698 11565
rect 16798 11449 16870 11493
rect 16798 10809 16811 11449
rect 16857 10809 16870 11449
rect 17626 11449 17698 11493
rect 16798 10765 16870 10809
rect 17626 10809 17639 11449
rect 17685 10809 17698 11449
rect 17626 10765 17698 10809
rect 16798 10693 17698 10765
rect 20840 11493 21740 11565
rect 20840 11449 20912 11493
rect 20840 10809 20853 11449
rect 20899 10809 20912 11449
rect 21668 11449 21740 11493
rect 20840 10765 20912 10809
rect 21668 10809 21681 11449
rect 21727 10809 21740 11449
rect 21668 10765 21740 10809
rect 20840 10693 21740 10765
rect 24882 11493 25782 11565
rect 24882 11449 24954 11493
rect 24882 10809 24895 11449
rect 24941 10809 24954 11449
rect 25710 11449 25782 11493
rect 24882 10765 24954 10809
rect 25710 10809 25723 11449
rect 25769 10809 25782 11449
rect 25710 10765 25782 10809
rect 24882 10693 25782 10765
rect 28924 11493 29824 11565
rect 28924 11449 28996 11493
rect 28924 10809 28937 11449
rect 28983 10809 28996 11449
rect 29752 11449 29824 11493
rect 28924 10765 28996 10809
rect 29752 10809 29765 11449
rect 29811 10809 29824 11449
rect 29752 10765 29824 10809
rect 28924 10693 29824 10765
rect 660 8532 1560 8604
rect 660 8488 732 8532
rect 660 7848 673 8488
rect 719 7848 732 8488
rect 1488 8488 1560 8532
rect 660 7804 732 7848
rect 1488 7848 1501 8488
rect 1547 7848 1560 8488
rect 1488 7804 1560 7848
rect 660 7732 1560 7804
rect 4672 8532 5572 8604
rect 4672 8488 4744 8532
rect 4672 7848 4685 8488
rect 4731 7848 4744 8488
rect 5500 8488 5572 8532
rect 4672 7804 4744 7848
rect 5500 7848 5513 8488
rect 5559 7848 5572 8488
rect 5500 7804 5572 7848
rect 4672 7732 5572 7804
rect 8714 8532 9614 8604
rect 8714 8488 8786 8532
rect 8714 7848 8727 8488
rect 8773 7848 8786 8488
rect 9542 8488 9614 8532
rect 8714 7804 8786 7848
rect 9542 7848 9555 8488
rect 9601 7848 9614 8488
rect 9542 7804 9614 7848
rect 8714 7732 9614 7804
rect 12756 8532 13656 8604
rect 12756 8488 12828 8532
rect 12756 7848 12769 8488
rect 12815 7848 12828 8488
rect 13584 8488 13656 8532
rect 12756 7804 12828 7848
rect 13584 7848 13597 8488
rect 13643 7848 13656 8488
rect 13584 7804 13656 7848
rect 12756 7732 13656 7804
rect 16798 8532 17698 8604
rect 16798 8488 16870 8532
rect 16798 7848 16811 8488
rect 16857 7848 16870 8488
rect 17626 8488 17698 8532
rect 16798 7804 16870 7848
rect 17626 7848 17639 8488
rect 17685 7848 17698 8488
rect 17626 7804 17698 7848
rect 16798 7732 17698 7804
rect 20840 8532 21740 8604
rect 20840 8488 20912 8532
rect 20840 7848 20853 8488
rect 20899 7848 20912 8488
rect 21668 8488 21740 8532
rect 20840 7804 20912 7848
rect 21668 7848 21681 8488
rect 21727 7848 21740 8488
rect 21668 7804 21740 7848
rect 20840 7732 21740 7804
rect 24882 8532 25782 8604
rect 24882 8488 24954 8532
rect 24882 7848 24895 8488
rect 24941 7848 24954 8488
rect 25710 8488 25782 8532
rect 24882 7804 24954 7848
rect 25710 7848 25723 8488
rect 25769 7848 25782 8488
rect 25710 7804 25782 7848
rect 24882 7732 25782 7804
rect 660 6327 1560 6399
rect 660 6283 732 6327
rect 660 5643 673 6283
rect 719 5643 732 6283
rect 1488 6283 1560 6327
rect 660 5599 732 5643
rect 1488 5643 1501 6283
rect 1547 5643 1560 6283
rect 1488 5599 1560 5643
rect 660 5527 1560 5599
rect 2146 6327 3046 6399
rect 2146 6283 2218 6327
rect 2146 5643 2159 6283
rect 2205 5643 2218 6283
rect 2974 6283 3046 6327
rect 2146 5599 2218 5643
rect 2974 5643 2987 6283
rect 3033 5643 3046 6283
rect 2974 5599 3046 5643
rect 2146 5527 3046 5599
rect 4672 6327 5572 6399
rect 4672 6283 4744 6327
rect 4672 5643 4685 6283
rect 4731 5643 4744 6283
rect 5500 6283 5572 6327
rect 4672 5599 4744 5643
rect 5500 5643 5513 6283
rect 5559 5643 5572 6283
rect 5500 5599 5572 5643
rect 4672 5527 5572 5599
rect 6158 6327 7058 6399
rect 6158 6283 6230 6327
rect 6158 5643 6171 6283
rect 6217 5643 6230 6283
rect 6986 6283 7058 6327
rect 6158 5599 6230 5643
rect 6986 5643 6999 6283
rect 7045 5643 7058 6283
rect 6986 5599 7058 5643
rect 6158 5527 7058 5599
rect 8714 6327 9614 6399
rect 8714 6283 8786 6327
rect 8714 5643 8727 6283
rect 8773 5643 8786 6283
rect 9542 6283 9614 6327
rect 8714 5599 8786 5643
rect 9542 5643 9555 6283
rect 9601 5643 9614 6283
rect 9542 5599 9614 5643
rect 8714 5527 9614 5599
rect 10200 6327 11100 6399
rect 10200 6283 10272 6327
rect 10200 5643 10213 6283
rect 10259 5643 10272 6283
rect 11028 6283 11100 6327
rect 10200 5599 10272 5643
rect 11028 5643 11041 6283
rect 11087 5643 11100 6283
rect 11028 5599 11100 5643
rect 10200 5527 11100 5599
rect 12756 6327 13656 6399
rect 12756 6283 12828 6327
rect 12756 5643 12769 6283
rect 12815 5643 12828 6283
rect 13584 6283 13656 6327
rect 12756 5599 12828 5643
rect 13584 5643 13597 6283
rect 13643 5643 13656 6283
rect 13584 5599 13656 5643
rect 12756 5527 13656 5599
rect 14242 6327 15142 6399
rect 14242 6283 14314 6327
rect 14242 5643 14255 6283
rect 14301 5643 14314 6283
rect 15070 6283 15142 6327
rect 14242 5599 14314 5643
rect 15070 5643 15083 6283
rect 15129 5643 15142 6283
rect 15070 5599 15142 5643
rect 14242 5527 15142 5599
rect 16798 6327 17698 6399
rect 16798 6283 16870 6327
rect 16798 5643 16811 6283
rect 16857 5643 16870 6283
rect 17626 6283 17698 6327
rect 16798 5599 16870 5643
rect 17626 5643 17639 6283
rect 17685 5643 17698 6283
rect 17626 5599 17698 5643
rect 16798 5527 17698 5599
rect 18284 6327 19184 6399
rect 18284 6283 18356 6327
rect 18284 5643 18297 6283
rect 18343 5643 18356 6283
rect 19112 6283 19184 6327
rect 18284 5599 18356 5643
rect 19112 5643 19125 6283
rect 19171 5643 19184 6283
rect 19112 5599 19184 5643
rect 18284 5527 19184 5599
rect 20840 6327 21740 6399
rect 20840 6283 20912 6327
rect 20840 5643 20853 6283
rect 20899 5643 20912 6283
rect 21668 6283 21740 6327
rect 20840 5599 20912 5643
rect 21668 5643 21681 6283
rect 21727 5643 21740 6283
rect 21668 5599 21740 5643
rect 20840 5527 21740 5599
rect 22326 6327 23226 6399
rect 22326 6283 22398 6327
rect 22326 5643 22339 6283
rect 22385 5643 22398 6283
rect 23154 6283 23226 6327
rect 22326 5599 22398 5643
rect 23154 5643 23167 6283
rect 23213 5643 23226 6283
rect 23154 5599 23226 5643
rect 22326 5527 23226 5599
rect 24882 6327 25782 6399
rect 24882 6283 24954 6327
rect 24882 5643 24895 6283
rect 24941 5643 24954 6283
rect 25710 6283 25782 6327
rect 24882 5599 24954 5643
rect 25710 5643 25723 6283
rect 25769 5643 25782 6283
rect 25710 5599 25782 5643
rect 24882 5527 25782 5599
rect 26368 6327 27268 6399
rect 26368 6283 26440 6327
rect 26368 5643 26381 6283
rect 26427 5643 26440 6283
rect 27196 6283 27268 6327
rect 26368 5599 26440 5643
rect 27196 5643 27209 6283
rect 27255 5643 27268 6283
rect 27196 5599 27268 5643
rect 26368 5527 27268 5599
rect 660 4122 1560 4194
rect 660 4078 732 4122
rect 660 3438 673 4078
rect 719 3438 732 4078
rect 1488 4078 1560 4122
rect 660 3394 732 3438
rect 1488 3438 1501 4078
rect 1547 3438 1560 4078
rect 1488 3394 1560 3438
rect 660 3322 1560 3394
rect 2146 4123 3046 4195
rect 2146 4079 2218 4123
rect 2146 3439 2159 4079
rect 2205 3439 2218 4079
rect 2974 4079 3046 4123
rect 2146 3395 2218 3439
rect 2974 3439 2987 4079
rect 3033 3439 3046 4079
rect 2974 3395 3046 3439
rect 2146 3323 3046 3395
rect 4672 4122 5572 4194
rect 4672 4078 4744 4122
rect 4672 3438 4685 4078
rect 4731 3438 4744 4078
rect 5500 4078 5572 4122
rect 4672 3394 4744 3438
rect 5500 3438 5513 4078
rect 5559 3438 5572 4078
rect 5500 3394 5572 3438
rect 4672 3322 5572 3394
rect 6158 4123 7058 4195
rect 6158 4079 6230 4123
rect 6158 3439 6171 4079
rect 6217 3439 6230 4079
rect 6986 4079 7058 4123
rect 6158 3395 6230 3439
rect 6986 3439 6999 4079
rect 7045 3439 7058 4079
rect 6986 3395 7058 3439
rect 6158 3323 7058 3395
rect 8714 4122 9614 4194
rect 8714 4078 8786 4122
rect 8714 3438 8727 4078
rect 8773 3438 8786 4078
rect 9542 4078 9614 4122
rect 8714 3394 8786 3438
rect 9542 3438 9555 4078
rect 9601 3438 9614 4078
rect 9542 3394 9614 3438
rect 8714 3322 9614 3394
rect 10200 4123 11100 4195
rect 10200 4079 10272 4123
rect 10200 3439 10213 4079
rect 10259 3439 10272 4079
rect 11028 4079 11100 4123
rect 10200 3395 10272 3439
rect 11028 3439 11041 4079
rect 11087 3439 11100 4079
rect 11028 3395 11100 3439
rect 10200 3323 11100 3395
rect 12756 4122 13656 4194
rect 12756 4078 12828 4122
rect 12756 3438 12769 4078
rect 12815 3438 12828 4078
rect 13584 4078 13656 4122
rect 12756 3394 12828 3438
rect 13584 3438 13597 4078
rect 13643 3438 13656 4078
rect 13584 3394 13656 3438
rect 12756 3322 13656 3394
rect 14242 4123 15142 4195
rect 14242 4079 14314 4123
rect 14242 3439 14255 4079
rect 14301 3439 14314 4079
rect 15070 4079 15142 4123
rect 14242 3395 14314 3439
rect 15070 3439 15083 4079
rect 15129 3439 15142 4079
rect 15070 3395 15142 3439
rect 14242 3323 15142 3395
rect 16798 4122 17698 4194
rect 16798 4078 16870 4122
rect 16798 3438 16811 4078
rect 16857 3438 16870 4078
rect 17626 4078 17698 4122
rect 16798 3394 16870 3438
rect 17626 3438 17639 4078
rect 17685 3438 17698 4078
rect 17626 3394 17698 3438
rect 16798 3322 17698 3394
rect 18284 4123 19184 4195
rect 18284 4079 18356 4123
rect 18284 3439 18297 4079
rect 18343 3439 18356 4079
rect 19112 4079 19184 4123
rect 18284 3395 18356 3439
rect 19112 3439 19125 4079
rect 19171 3439 19184 4079
rect 19112 3395 19184 3439
rect 18284 3323 19184 3395
rect 20840 4122 21740 4194
rect 20840 4078 20912 4122
rect 20840 3438 20853 4078
rect 20899 3438 20912 4078
rect 21668 4078 21740 4122
rect 20840 3394 20912 3438
rect 21668 3438 21681 4078
rect 21727 3438 21740 4078
rect 21668 3394 21740 3438
rect 20840 3322 21740 3394
rect 22326 4123 23226 4195
rect 22326 4079 22398 4123
rect 22326 3439 22339 4079
rect 22385 3439 22398 4079
rect 23154 4079 23226 4123
rect 22326 3395 22398 3439
rect 23154 3439 23167 4079
rect 23213 3439 23226 4079
rect 23154 3395 23226 3439
rect 22326 3323 23226 3395
rect 24882 4122 25782 4194
rect 24882 4078 24954 4122
rect 24882 3438 24895 4078
rect 24941 3438 24954 4078
rect 25710 4078 25782 4122
rect 24882 3394 24954 3438
rect 25710 3438 25723 4078
rect 25769 3438 25782 4078
rect 25710 3394 25782 3438
rect 24882 3322 25782 3394
rect 26368 4123 27268 4195
rect 26368 4079 26440 4123
rect 26368 3439 26381 4079
rect 26427 3439 26440 4079
rect 27196 4079 27268 4123
rect 26368 3395 26440 3439
rect 27196 3439 27209 4079
rect 27255 3439 27268 4079
rect 27196 3395 27268 3439
rect 26368 3323 27268 3395
rect 660 1917 1560 1989
rect 660 1873 732 1917
rect 660 1233 673 1873
rect 719 1233 732 1873
rect 1488 1873 1560 1917
rect 660 1189 732 1233
rect 1488 1233 1501 1873
rect 1547 1233 1560 1873
rect 1488 1189 1560 1233
rect 660 1117 1560 1189
rect 4672 1917 5572 1989
rect 4672 1873 4744 1917
rect 4672 1233 4685 1873
rect 4731 1233 4744 1873
rect 5500 1873 5572 1917
rect 4672 1189 4744 1233
rect 5500 1233 5513 1873
rect 5559 1233 5572 1873
rect 5500 1189 5572 1233
rect 4672 1117 5572 1189
rect 8714 1917 9614 1989
rect 8714 1873 8786 1917
rect 8714 1233 8727 1873
rect 8773 1233 8786 1873
rect 9542 1873 9614 1917
rect 8714 1189 8786 1233
rect 9542 1233 9555 1873
rect 9601 1233 9614 1873
rect 9542 1189 9614 1233
rect 8714 1117 9614 1189
rect 12756 1917 13656 1989
rect 12756 1873 12828 1917
rect 12756 1233 12769 1873
rect 12815 1233 12828 1873
rect 13584 1873 13656 1917
rect 12756 1189 12828 1233
rect 13584 1233 13597 1873
rect 13643 1233 13656 1873
rect 13584 1189 13656 1233
rect 12756 1117 13656 1189
rect 16798 1917 17698 1989
rect 16798 1873 16870 1917
rect 16798 1233 16811 1873
rect 16857 1233 16870 1873
rect 17626 1873 17698 1917
rect 16798 1189 16870 1233
rect 17626 1233 17639 1873
rect 17685 1233 17698 1873
rect 17626 1189 17698 1233
rect 16798 1117 17698 1189
rect 20840 1917 21740 1989
rect 20840 1873 20912 1917
rect 20840 1233 20853 1873
rect 20899 1233 20912 1873
rect 21668 1873 21740 1917
rect 20840 1189 20912 1233
rect 21668 1233 21681 1873
rect 21727 1233 21740 1873
rect 21668 1189 21740 1233
rect 20840 1117 21740 1189
rect 24882 1917 25782 1989
rect 24882 1873 24954 1917
rect 24882 1233 24895 1873
rect 24941 1233 24954 1873
rect 25710 1873 25782 1917
rect 24882 1189 24954 1233
rect 25710 1233 25723 1873
rect 25769 1233 25782 1873
rect 25710 1189 25782 1233
rect 24882 1117 25782 1189
<< psubdiffcont >>
rect 4685 16567 4731 16907
rect 5513 16567 5559 16907
rect 8727 16564 8773 16904
rect 9555 16564 9601 16904
rect 12769 16564 12815 16904
rect 13597 16564 13643 16904
rect 16811 16564 16857 16904
rect 17639 16564 17685 16904
rect 20853 16564 20899 16904
rect 21681 16564 21727 16904
rect 24895 16564 24941 16904
rect 25723 16564 25769 16904
rect 28937 16564 28983 16904
rect 29765 16564 29811 16904
rect 4685 14362 4731 14702
rect 5513 14362 5559 14702
rect 6171 14362 6217 14702
rect 6999 14362 7045 14702
rect 8727 14359 8773 14699
rect 9555 14359 9601 14699
rect 10213 14359 10259 14699
rect 11041 14359 11087 14699
rect 12769 14359 12815 14699
rect 13597 14359 13643 14699
rect 14255 14359 14301 14699
rect 15083 14359 15129 14699
rect 16811 14359 16857 14699
rect 17639 14359 17685 14699
rect 18297 14359 18343 14699
rect 19125 14359 19171 14699
rect 20853 14359 20899 14699
rect 21681 14359 21727 14699
rect 22339 14359 22385 14699
rect 23167 14359 23213 14699
rect 24895 14359 24941 14699
rect 25723 14359 25769 14699
rect 26381 14359 26427 14699
rect 27209 14359 27255 14699
rect 28937 14359 28983 14699
rect 29765 14359 29811 14699
rect 30423 14359 30469 14699
rect 31251 14359 31297 14699
rect 4685 12157 4731 12497
rect 5513 12157 5559 12497
rect 6171 12158 6217 12498
rect 6999 12158 7045 12498
rect 8727 12154 8773 12494
rect 9555 12154 9601 12494
rect 10213 12155 10259 12495
rect 11041 12155 11087 12495
rect 12769 12154 12815 12494
rect 13597 12154 13643 12494
rect 14255 12155 14301 12495
rect 15083 12155 15129 12495
rect 16811 12154 16857 12494
rect 17639 12154 17685 12494
rect 18297 12155 18343 12495
rect 19125 12155 19171 12495
rect 20853 12154 20899 12494
rect 21681 12154 21727 12494
rect 22339 12155 22385 12495
rect 23167 12155 23213 12495
rect 24895 12154 24941 12494
rect 25723 12154 25769 12494
rect 26381 12155 26427 12495
rect 27209 12155 27255 12495
rect 28937 12154 28983 12494
rect 29765 12154 29811 12494
rect 30423 12155 30469 12495
rect 31251 12155 31297 12495
rect 4685 9952 4731 10292
rect 5513 9952 5559 10292
rect 8727 9949 8773 10289
rect 9555 9949 9601 10289
rect 12769 9949 12815 10289
rect 13597 9949 13643 10289
rect 16811 9949 16857 10289
rect 17639 9949 17685 10289
rect 20853 9949 20899 10289
rect 21681 9949 21727 10289
rect 24895 9949 24941 10289
rect 25723 9949 25769 10289
rect 28937 9949 28983 10289
rect 29765 9949 29811 10289
rect 673 6988 719 7328
rect 1501 6988 1547 7328
rect 4685 6988 4731 7328
rect 5513 6988 5559 7328
rect 8727 6988 8773 7328
rect 9555 6988 9601 7328
rect 12769 6988 12815 7328
rect 13597 6988 13643 7328
rect 16811 6988 16857 7328
rect 17639 6988 17685 7328
rect 20853 6988 20899 7328
rect 21681 6988 21727 7328
rect 24895 6988 24941 7328
rect 25723 6988 25769 7328
rect 673 4783 719 5123
rect 1501 4783 1547 5123
rect 2159 4783 2205 5123
rect 2987 4783 3033 5123
rect 4685 4783 4731 5123
rect 5513 4783 5559 5123
rect 6171 4783 6217 5123
rect 6999 4783 7045 5123
rect 8727 4783 8773 5123
rect 9555 4783 9601 5123
rect 10213 4783 10259 5123
rect 11041 4783 11087 5123
rect 12769 4783 12815 5123
rect 13597 4783 13643 5123
rect 14255 4783 14301 5123
rect 15083 4783 15129 5123
rect 16811 4783 16857 5123
rect 17639 4783 17685 5123
rect 18297 4783 18343 5123
rect 19125 4783 19171 5123
rect 20853 4783 20899 5123
rect 21681 4783 21727 5123
rect 22339 4783 22385 5123
rect 23167 4783 23213 5123
rect 24895 4783 24941 5123
rect 25723 4783 25769 5123
rect 26381 4783 26427 5123
rect 27209 4783 27255 5123
rect 673 2578 719 2918
rect 1501 2578 1547 2918
rect 2159 2579 2205 2919
rect 2987 2579 3033 2919
rect 4685 2578 4731 2918
rect 5513 2578 5559 2918
rect 6171 2579 6217 2919
rect 6999 2579 7045 2919
rect 8727 2578 8773 2918
rect 9555 2578 9601 2918
rect 10213 2579 10259 2919
rect 11041 2579 11087 2919
rect 12769 2578 12815 2918
rect 13597 2578 13643 2918
rect 14255 2579 14301 2919
rect 15083 2579 15129 2919
rect 16811 2578 16857 2918
rect 17639 2578 17685 2918
rect 18297 2579 18343 2919
rect 19125 2579 19171 2919
rect 20853 2578 20899 2918
rect 21681 2578 21727 2918
rect 22339 2579 22385 2919
rect 23167 2579 23213 2919
rect 24895 2578 24941 2918
rect 25723 2578 25769 2918
rect 26381 2579 26427 2919
rect 27209 2579 27255 2919
rect 673 373 719 713
rect 1501 373 1547 713
rect 4685 373 4731 713
rect 5513 373 5559 713
rect 8727 373 8773 713
rect 9555 373 9601 713
rect 12769 373 12815 713
rect 13597 373 13643 713
rect 16811 373 16857 713
rect 17639 373 17685 713
rect 20853 373 20899 713
rect 21681 373 21727 713
rect 24895 373 24941 713
rect 25723 373 25769 713
<< nsubdiffcont >>
rect 4685 17427 4731 18067
rect 5513 17427 5559 18067
rect 8727 17424 8773 18064
rect 9555 17424 9601 18064
rect 12769 17424 12815 18064
rect 13597 17424 13643 18064
rect 16811 17424 16857 18064
rect 17639 17424 17685 18064
rect 20853 17424 20899 18064
rect 21681 17424 21727 18064
rect 24895 17424 24941 18064
rect 25723 17424 25769 18064
rect 28937 17424 28983 18064
rect 29765 17424 29811 18064
rect 4685 15222 4731 15862
rect 5513 15222 5559 15862
rect 6171 15222 6217 15862
rect 6999 15222 7045 15862
rect 8727 15219 8773 15859
rect 9555 15219 9601 15859
rect 10213 15219 10259 15859
rect 11041 15219 11087 15859
rect 12769 15219 12815 15859
rect 13597 15219 13643 15859
rect 14255 15219 14301 15859
rect 15083 15219 15129 15859
rect 16811 15219 16857 15859
rect 17639 15219 17685 15859
rect 18297 15219 18343 15859
rect 19125 15219 19171 15859
rect 20853 15219 20899 15859
rect 21681 15219 21727 15859
rect 22339 15219 22385 15859
rect 23167 15219 23213 15859
rect 24895 15219 24941 15859
rect 25723 15219 25769 15859
rect 26381 15219 26427 15859
rect 27209 15219 27255 15859
rect 28937 15219 28983 15859
rect 29765 15219 29811 15859
rect 30423 15219 30469 15859
rect 31251 15219 31297 15859
rect 4685 13017 4731 13657
rect 5513 13017 5559 13657
rect 6171 13018 6217 13658
rect 6999 13018 7045 13658
rect 8727 13014 8773 13654
rect 9555 13014 9601 13654
rect 10213 13015 10259 13655
rect 11041 13015 11087 13655
rect 12769 13014 12815 13654
rect 13597 13014 13643 13654
rect 14255 13015 14301 13655
rect 15083 13015 15129 13655
rect 16811 13014 16857 13654
rect 17639 13014 17685 13654
rect 18297 13015 18343 13655
rect 19125 13015 19171 13655
rect 20853 13014 20899 13654
rect 21681 13014 21727 13654
rect 22339 13015 22385 13655
rect 23167 13015 23213 13655
rect 24895 13014 24941 13654
rect 25723 13014 25769 13654
rect 26381 13015 26427 13655
rect 27209 13015 27255 13655
rect 28937 13014 28983 13654
rect 29765 13014 29811 13654
rect 30423 13015 30469 13655
rect 31251 13015 31297 13655
rect 4685 10812 4731 11452
rect 5513 10812 5559 11452
rect 8727 10809 8773 11449
rect 9555 10809 9601 11449
rect 12769 10809 12815 11449
rect 13597 10809 13643 11449
rect 16811 10809 16857 11449
rect 17639 10809 17685 11449
rect 20853 10809 20899 11449
rect 21681 10809 21727 11449
rect 24895 10809 24941 11449
rect 25723 10809 25769 11449
rect 28937 10809 28983 11449
rect 29765 10809 29811 11449
rect 673 7848 719 8488
rect 1501 7848 1547 8488
rect 4685 7848 4731 8488
rect 5513 7848 5559 8488
rect 8727 7848 8773 8488
rect 9555 7848 9601 8488
rect 12769 7848 12815 8488
rect 13597 7848 13643 8488
rect 16811 7848 16857 8488
rect 17639 7848 17685 8488
rect 20853 7848 20899 8488
rect 21681 7848 21727 8488
rect 24895 7848 24941 8488
rect 25723 7848 25769 8488
rect 673 5643 719 6283
rect 1501 5643 1547 6283
rect 2159 5643 2205 6283
rect 2987 5643 3033 6283
rect 4685 5643 4731 6283
rect 5513 5643 5559 6283
rect 6171 5643 6217 6283
rect 6999 5643 7045 6283
rect 8727 5643 8773 6283
rect 9555 5643 9601 6283
rect 10213 5643 10259 6283
rect 11041 5643 11087 6283
rect 12769 5643 12815 6283
rect 13597 5643 13643 6283
rect 14255 5643 14301 6283
rect 15083 5643 15129 6283
rect 16811 5643 16857 6283
rect 17639 5643 17685 6283
rect 18297 5643 18343 6283
rect 19125 5643 19171 6283
rect 20853 5643 20899 6283
rect 21681 5643 21727 6283
rect 22339 5643 22385 6283
rect 23167 5643 23213 6283
rect 24895 5643 24941 6283
rect 25723 5643 25769 6283
rect 26381 5643 26427 6283
rect 27209 5643 27255 6283
rect 673 3438 719 4078
rect 1501 3438 1547 4078
rect 2159 3439 2205 4079
rect 2987 3439 3033 4079
rect 4685 3438 4731 4078
rect 5513 3438 5559 4078
rect 6171 3439 6217 4079
rect 6999 3439 7045 4079
rect 8727 3438 8773 4078
rect 9555 3438 9601 4078
rect 10213 3439 10259 4079
rect 11041 3439 11087 4079
rect 12769 3438 12815 4078
rect 13597 3438 13643 4078
rect 14255 3439 14301 4079
rect 15083 3439 15129 4079
rect 16811 3438 16857 4078
rect 17639 3438 17685 4078
rect 18297 3439 18343 4079
rect 19125 3439 19171 4079
rect 20853 3438 20899 4078
rect 21681 3438 21727 4078
rect 22339 3439 22385 4079
rect 23167 3439 23213 4079
rect 24895 3438 24941 4078
rect 25723 3438 25769 4078
rect 26381 3439 26427 4079
rect 27209 3439 27255 4079
rect 673 1233 719 1873
rect 1501 1233 1547 1873
rect 4685 1233 4731 1873
rect 5513 1233 5559 1873
rect 8727 1233 8773 1873
rect 9555 1233 9601 1873
rect 12769 1233 12815 1873
rect 13597 1233 13643 1873
rect 16811 1233 16857 1873
rect 17639 1233 17685 1873
rect 20853 1233 20899 1873
rect 21681 1233 21727 1873
rect 24895 1233 24941 1873
rect 25723 1233 25769 1873
<< polysilicon >>
rect 4898 18076 4978 18089
rect 4898 18030 4911 18076
rect 4965 18030 4978 18076
rect 4898 17997 4978 18030
rect 5082 18076 5162 18089
rect 5082 18030 5095 18076
rect 5149 18030 5162 18076
rect 5082 17997 5162 18030
rect 5266 18076 5346 18089
rect 5266 18030 5279 18076
rect 5333 18030 5346 18076
rect 5266 17997 5346 18030
rect 4898 17464 4978 17497
rect 4898 17418 4911 17464
rect 4965 17418 4978 17464
rect 4898 17405 4978 17418
rect 5082 17464 5162 17497
rect 5082 17418 5095 17464
rect 5149 17418 5162 17464
rect 5082 17405 5162 17418
rect 5266 17464 5346 17497
rect 5266 17418 5279 17464
rect 5333 17418 5346 17464
rect 5266 17405 5346 17418
rect 8940 18073 9020 18086
rect 8940 18027 8953 18073
rect 9007 18027 9020 18073
rect 8940 17994 9020 18027
rect 9124 18073 9204 18086
rect 9124 18027 9137 18073
rect 9191 18027 9204 18073
rect 9124 17994 9204 18027
rect 9308 18073 9388 18086
rect 9308 18027 9321 18073
rect 9375 18027 9388 18073
rect 9308 17994 9388 18027
rect 8940 17461 9020 17494
rect 8940 17415 8953 17461
rect 9007 17415 9020 17461
rect 8940 17402 9020 17415
rect 9124 17461 9204 17494
rect 9124 17415 9137 17461
rect 9191 17415 9204 17461
rect 9124 17402 9204 17415
rect 9308 17461 9388 17494
rect 9308 17415 9321 17461
rect 9375 17415 9388 17461
rect 9308 17402 9388 17415
rect 12982 18073 13062 18086
rect 12982 18027 12995 18073
rect 13049 18027 13062 18073
rect 12982 17994 13062 18027
rect 13166 18073 13246 18086
rect 13166 18027 13179 18073
rect 13233 18027 13246 18073
rect 13166 17994 13246 18027
rect 13350 18073 13430 18086
rect 13350 18027 13363 18073
rect 13417 18027 13430 18073
rect 13350 17994 13430 18027
rect 12982 17461 13062 17494
rect 12982 17415 12995 17461
rect 13049 17415 13062 17461
rect 12982 17402 13062 17415
rect 13166 17461 13246 17494
rect 13166 17415 13179 17461
rect 13233 17415 13246 17461
rect 13166 17402 13246 17415
rect 13350 17461 13430 17494
rect 13350 17415 13363 17461
rect 13417 17415 13430 17461
rect 13350 17402 13430 17415
rect 17024 18073 17104 18086
rect 17024 18027 17037 18073
rect 17091 18027 17104 18073
rect 17024 17994 17104 18027
rect 17208 18073 17288 18086
rect 17208 18027 17221 18073
rect 17275 18027 17288 18073
rect 17208 17994 17288 18027
rect 17392 18073 17472 18086
rect 17392 18027 17405 18073
rect 17459 18027 17472 18073
rect 17392 17994 17472 18027
rect 17024 17461 17104 17494
rect 17024 17415 17037 17461
rect 17091 17415 17104 17461
rect 17024 17402 17104 17415
rect 17208 17461 17288 17494
rect 17208 17415 17221 17461
rect 17275 17415 17288 17461
rect 17208 17402 17288 17415
rect 17392 17461 17472 17494
rect 17392 17415 17405 17461
rect 17459 17415 17472 17461
rect 17392 17402 17472 17415
rect 21066 18073 21146 18086
rect 21066 18027 21079 18073
rect 21133 18027 21146 18073
rect 21066 17994 21146 18027
rect 21250 18073 21330 18086
rect 21250 18027 21263 18073
rect 21317 18027 21330 18073
rect 21250 17994 21330 18027
rect 21434 18073 21514 18086
rect 21434 18027 21447 18073
rect 21501 18027 21514 18073
rect 21434 17994 21514 18027
rect 21066 17461 21146 17494
rect 21066 17415 21079 17461
rect 21133 17415 21146 17461
rect 21066 17402 21146 17415
rect 21250 17461 21330 17494
rect 21250 17415 21263 17461
rect 21317 17415 21330 17461
rect 21250 17402 21330 17415
rect 21434 17461 21514 17494
rect 21434 17415 21447 17461
rect 21501 17415 21514 17461
rect 21434 17402 21514 17415
rect 25108 18073 25188 18086
rect 25108 18027 25121 18073
rect 25175 18027 25188 18073
rect 25108 17994 25188 18027
rect 25292 18073 25372 18086
rect 25292 18027 25305 18073
rect 25359 18027 25372 18073
rect 25292 17994 25372 18027
rect 25476 18073 25556 18086
rect 25476 18027 25489 18073
rect 25543 18027 25556 18073
rect 25476 17994 25556 18027
rect 25108 17461 25188 17494
rect 25108 17415 25121 17461
rect 25175 17415 25188 17461
rect 25108 17402 25188 17415
rect 25292 17461 25372 17494
rect 25292 17415 25305 17461
rect 25359 17415 25372 17461
rect 25292 17402 25372 17415
rect 25476 17461 25556 17494
rect 25476 17415 25489 17461
rect 25543 17415 25556 17461
rect 25476 17402 25556 17415
rect 29150 18073 29230 18086
rect 29150 18027 29163 18073
rect 29217 18027 29230 18073
rect 29150 17994 29230 18027
rect 29334 18073 29414 18086
rect 29334 18027 29347 18073
rect 29401 18027 29414 18073
rect 29334 17994 29414 18027
rect 29518 18073 29598 18086
rect 29518 18027 29531 18073
rect 29585 18027 29598 18073
rect 29518 17994 29598 18027
rect 29150 17461 29230 17494
rect 29150 17415 29163 17461
rect 29217 17415 29230 17461
rect 29150 17402 29230 17415
rect 29334 17461 29414 17494
rect 29334 17415 29347 17461
rect 29401 17415 29414 17461
rect 29334 17402 29414 17415
rect 29518 17461 29598 17494
rect 29518 17415 29531 17461
rect 29585 17415 29598 17461
rect 29518 17402 29598 17415
rect 4898 16916 4978 16929
rect 4898 16870 4911 16916
rect 4965 16870 4978 16916
rect 4898 16837 4978 16870
rect 5082 16916 5162 16929
rect 5082 16870 5095 16916
rect 5149 16870 5162 16916
rect 5082 16837 5162 16870
rect 5266 16916 5346 16929
rect 5266 16870 5279 16916
rect 5333 16870 5346 16916
rect 5266 16837 5346 16870
rect 4898 16604 4978 16637
rect 4898 16558 4911 16604
rect 4965 16558 4978 16604
rect 4898 16545 4978 16558
rect 5082 16604 5162 16637
rect 5082 16558 5095 16604
rect 5149 16558 5162 16604
rect 5082 16545 5162 16558
rect 5266 16604 5346 16637
rect 5266 16558 5279 16604
rect 5333 16558 5346 16604
rect 5266 16545 5346 16558
rect 8940 16913 9020 16926
rect 8940 16867 8953 16913
rect 9007 16867 9020 16913
rect 8940 16834 9020 16867
rect 9124 16913 9204 16926
rect 9124 16867 9137 16913
rect 9191 16867 9204 16913
rect 9124 16834 9204 16867
rect 9308 16913 9388 16926
rect 9308 16867 9321 16913
rect 9375 16867 9388 16913
rect 9308 16834 9388 16867
rect 8940 16601 9020 16634
rect 8940 16555 8953 16601
rect 9007 16555 9020 16601
rect 8940 16542 9020 16555
rect 9124 16601 9204 16634
rect 9124 16555 9137 16601
rect 9191 16555 9204 16601
rect 9124 16542 9204 16555
rect 9308 16601 9388 16634
rect 9308 16555 9321 16601
rect 9375 16555 9388 16601
rect 9308 16542 9388 16555
rect 12982 16913 13062 16926
rect 12982 16867 12995 16913
rect 13049 16867 13062 16913
rect 12982 16834 13062 16867
rect 13166 16913 13246 16926
rect 13166 16867 13179 16913
rect 13233 16867 13246 16913
rect 13166 16834 13246 16867
rect 13350 16913 13430 16926
rect 13350 16867 13363 16913
rect 13417 16867 13430 16913
rect 13350 16834 13430 16867
rect 12982 16601 13062 16634
rect 12982 16555 12995 16601
rect 13049 16555 13062 16601
rect 12982 16542 13062 16555
rect 13166 16601 13246 16634
rect 13166 16555 13179 16601
rect 13233 16555 13246 16601
rect 13166 16542 13246 16555
rect 13350 16601 13430 16634
rect 13350 16555 13363 16601
rect 13417 16555 13430 16601
rect 13350 16542 13430 16555
rect 17024 16913 17104 16926
rect 17024 16867 17037 16913
rect 17091 16867 17104 16913
rect 17024 16834 17104 16867
rect 17208 16913 17288 16926
rect 17208 16867 17221 16913
rect 17275 16867 17288 16913
rect 17208 16834 17288 16867
rect 17392 16913 17472 16926
rect 17392 16867 17405 16913
rect 17459 16867 17472 16913
rect 17392 16834 17472 16867
rect 17024 16601 17104 16634
rect 17024 16555 17037 16601
rect 17091 16555 17104 16601
rect 17024 16542 17104 16555
rect 17208 16601 17288 16634
rect 17208 16555 17221 16601
rect 17275 16555 17288 16601
rect 17208 16542 17288 16555
rect 17392 16601 17472 16634
rect 17392 16555 17405 16601
rect 17459 16555 17472 16601
rect 17392 16542 17472 16555
rect 21066 16913 21146 16926
rect 21066 16867 21079 16913
rect 21133 16867 21146 16913
rect 21066 16834 21146 16867
rect 21250 16913 21330 16926
rect 21250 16867 21263 16913
rect 21317 16867 21330 16913
rect 21250 16834 21330 16867
rect 21434 16913 21514 16926
rect 21434 16867 21447 16913
rect 21501 16867 21514 16913
rect 21434 16834 21514 16867
rect 21066 16601 21146 16634
rect 21066 16555 21079 16601
rect 21133 16555 21146 16601
rect 21066 16542 21146 16555
rect 21250 16601 21330 16634
rect 21250 16555 21263 16601
rect 21317 16555 21330 16601
rect 21250 16542 21330 16555
rect 21434 16601 21514 16634
rect 21434 16555 21447 16601
rect 21501 16555 21514 16601
rect 21434 16542 21514 16555
rect 25108 16913 25188 16926
rect 25108 16867 25121 16913
rect 25175 16867 25188 16913
rect 25108 16834 25188 16867
rect 25292 16913 25372 16926
rect 25292 16867 25305 16913
rect 25359 16867 25372 16913
rect 25292 16834 25372 16867
rect 25476 16913 25556 16926
rect 25476 16867 25489 16913
rect 25543 16867 25556 16913
rect 25476 16834 25556 16867
rect 25108 16601 25188 16634
rect 25108 16555 25121 16601
rect 25175 16555 25188 16601
rect 25108 16542 25188 16555
rect 25292 16601 25372 16634
rect 25292 16555 25305 16601
rect 25359 16555 25372 16601
rect 25292 16542 25372 16555
rect 25476 16601 25556 16634
rect 25476 16555 25489 16601
rect 25543 16555 25556 16601
rect 25476 16542 25556 16555
rect 29150 16913 29230 16926
rect 29150 16867 29163 16913
rect 29217 16867 29230 16913
rect 29150 16834 29230 16867
rect 29334 16913 29414 16926
rect 29334 16867 29347 16913
rect 29401 16867 29414 16913
rect 29334 16834 29414 16867
rect 29518 16913 29598 16926
rect 29518 16867 29531 16913
rect 29585 16867 29598 16913
rect 29518 16834 29598 16867
rect 29150 16601 29230 16634
rect 29150 16555 29163 16601
rect 29217 16555 29230 16601
rect 29150 16542 29230 16555
rect 29334 16601 29414 16634
rect 29334 16555 29347 16601
rect 29401 16555 29414 16601
rect 29334 16542 29414 16555
rect 29518 16601 29598 16634
rect 29518 16555 29531 16601
rect 29585 16555 29598 16601
rect 29518 16542 29598 16555
rect 4898 15871 4978 15884
rect 4898 15825 4911 15871
rect 4965 15825 4978 15871
rect 4898 15792 4978 15825
rect 5082 15871 5162 15884
rect 5082 15825 5095 15871
rect 5149 15825 5162 15871
rect 5082 15792 5162 15825
rect 5266 15871 5346 15884
rect 5266 15825 5279 15871
rect 5333 15825 5346 15871
rect 5266 15792 5346 15825
rect 4898 15259 4978 15292
rect 4898 15213 4911 15259
rect 4965 15213 4978 15259
rect 4898 15200 4978 15213
rect 5082 15259 5162 15292
rect 5082 15213 5095 15259
rect 5149 15213 5162 15259
rect 5082 15200 5162 15213
rect 5266 15259 5346 15292
rect 5266 15213 5279 15259
rect 5333 15213 5346 15259
rect 5266 15200 5346 15213
rect 6384 15871 6464 15884
rect 6384 15825 6397 15871
rect 6451 15825 6464 15871
rect 6384 15792 6464 15825
rect 6568 15871 6648 15884
rect 6568 15825 6581 15871
rect 6635 15825 6648 15871
rect 6568 15792 6648 15825
rect 6752 15871 6832 15884
rect 6752 15825 6765 15871
rect 6819 15825 6832 15871
rect 6752 15792 6832 15825
rect 6384 15259 6464 15292
rect 6384 15213 6397 15259
rect 6451 15213 6464 15259
rect 6384 15200 6464 15213
rect 6568 15259 6648 15292
rect 6568 15213 6581 15259
rect 6635 15213 6648 15259
rect 6568 15200 6648 15213
rect 6752 15259 6832 15292
rect 6752 15213 6765 15259
rect 6819 15213 6832 15259
rect 6752 15200 6832 15213
rect 8940 15868 9020 15881
rect 8940 15822 8953 15868
rect 9007 15822 9020 15868
rect 8940 15789 9020 15822
rect 9124 15868 9204 15881
rect 9124 15822 9137 15868
rect 9191 15822 9204 15868
rect 9124 15789 9204 15822
rect 9308 15868 9388 15881
rect 9308 15822 9321 15868
rect 9375 15822 9388 15868
rect 9308 15789 9388 15822
rect 8940 15256 9020 15289
rect 8940 15210 8953 15256
rect 9007 15210 9020 15256
rect 8940 15197 9020 15210
rect 9124 15256 9204 15289
rect 9124 15210 9137 15256
rect 9191 15210 9204 15256
rect 9124 15197 9204 15210
rect 9308 15256 9388 15289
rect 9308 15210 9321 15256
rect 9375 15210 9388 15256
rect 9308 15197 9388 15210
rect 10426 15868 10506 15881
rect 10426 15822 10439 15868
rect 10493 15822 10506 15868
rect 10426 15789 10506 15822
rect 10610 15868 10690 15881
rect 10610 15822 10623 15868
rect 10677 15822 10690 15868
rect 10610 15789 10690 15822
rect 10794 15868 10874 15881
rect 10794 15822 10807 15868
rect 10861 15822 10874 15868
rect 10794 15789 10874 15822
rect 10426 15256 10506 15289
rect 10426 15210 10439 15256
rect 10493 15210 10506 15256
rect 10426 15197 10506 15210
rect 10610 15256 10690 15289
rect 10610 15210 10623 15256
rect 10677 15210 10690 15256
rect 10610 15197 10690 15210
rect 10794 15256 10874 15289
rect 10794 15210 10807 15256
rect 10861 15210 10874 15256
rect 10794 15197 10874 15210
rect 12982 15868 13062 15881
rect 12982 15822 12995 15868
rect 13049 15822 13062 15868
rect 12982 15789 13062 15822
rect 13166 15868 13246 15881
rect 13166 15822 13179 15868
rect 13233 15822 13246 15868
rect 13166 15789 13246 15822
rect 13350 15868 13430 15881
rect 13350 15822 13363 15868
rect 13417 15822 13430 15868
rect 13350 15789 13430 15822
rect 12982 15256 13062 15289
rect 12982 15210 12995 15256
rect 13049 15210 13062 15256
rect 12982 15197 13062 15210
rect 13166 15256 13246 15289
rect 13166 15210 13179 15256
rect 13233 15210 13246 15256
rect 13166 15197 13246 15210
rect 13350 15256 13430 15289
rect 13350 15210 13363 15256
rect 13417 15210 13430 15256
rect 13350 15197 13430 15210
rect 14468 15868 14548 15881
rect 14468 15822 14481 15868
rect 14535 15822 14548 15868
rect 14468 15789 14548 15822
rect 14652 15868 14732 15881
rect 14652 15822 14665 15868
rect 14719 15822 14732 15868
rect 14652 15789 14732 15822
rect 14836 15868 14916 15881
rect 14836 15822 14849 15868
rect 14903 15822 14916 15868
rect 14836 15789 14916 15822
rect 14468 15256 14548 15289
rect 14468 15210 14481 15256
rect 14535 15210 14548 15256
rect 14468 15197 14548 15210
rect 14652 15256 14732 15289
rect 14652 15210 14665 15256
rect 14719 15210 14732 15256
rect 14652 15197 14732 15210
rect 14836 15256 14916 15289
rect 14836 15210 14849 15256
rect 14903 15210 14916 15256
rect 14836 15197 14916 15210
rect 17024 15868 17104 15881
rect 17024 15822 17037 15868
rect 17091 15822 17104 15868
rect 17024 15789 17104 15822
rect 17208 15868 17288 15881
rect 17208 15822 17221 15868
rect 17275 15822 17288 15868
rect 17208 15789 17288 15822
rect 17392 15868 17472 15881
rect 17392 15822 17405 15868
rect 17459 15822 17472 15868
rect 17392 15789 17472 15822
rect 17024 15256 17104 15289
rect 17024 15210 17037 15256
rect 17091 15210 17104 15256
rect 17024 15197 17104 15210
rect 17208 15256 17288 15289
rect 17208 15210 17221 15256
rect 17275 15210 17288 15256
rect 17208 15197 17288 15210
rect 17392 15256 17472 15289
rect 17392 15210 17405 15256
rect 17459 15210 17472 15256
rect 17392 15197 17472 15210
rect 18510 15868 18590 15881
rect 18510 15822 18523 15868
rect 18577 15822 18590 15868
rect 18510 15789 18590 15822
rect 18694 15868 18774 15881
rect 18694 15822 18707 15868
rect 18761 15822 18774 15868
rect 18694 15789 18774 15822
rect 18878 15868 18958 15881
rect 18878 15822 18891 15868
rect 18945 15822 18958 15868
rect 18878 15789 18958 15822
rect 18510 15256 18590 15289
rect 18510 15210 18523 15256
rect 18577 15210 18590 15256
rect 18510 15197 18590 15210
rect 18694 15256 18774 15289
rect 18694 15210 18707 15256
rect 18761 15210 18774 15256
rect 18694 15197 18774 15210
rect 18878 15256 18958 15289
rect 18878 15210 18891 15256
rect 18945 15210 18958 15256
rect 18878 15197 18958 15210
rect 21066 15868 21146 15881
rect 21066 15822 21079 15868
rect 21133 15822 21146 15868
rect 21066 15789 21146 15822
rect 21250 15868 21330 15881
rect 21250 15822 21263 15868
rect 21317 15822 21330 15868
rect 21250 15789 21330 15822
rect 21434 15868 21514 15881
rect 21434 15822 21447 15868
rect 21501 15822 21514 15868
rect 21434 15789 21514 15822
rect 21066 15256 21146 15289
rect 21066 15210 21079 15256
rect 21133 15210 21146 15256
rect 21066 15197 21146 15210
rect 21250 15256 21330 15289
rect 21250 15210 21263 15256
rect 21317 15210 21330 15256
rect 21250 15197 21330 15210
rect 21434 15256 21514 15289
rect 21434 15210 21447 15256
rect 21501 15210 21514 15256
rect 21434 15197 21514 15210
rect 22552 15868 22632 15881
rect 22552 15822 22565 15868
rect 22619 15822 22632 15868
rect 22552 15789 22632 15822
rect 22736 15868 22816 15881
rect 22736 15822 22749 15868
rect 22803 15822 22816 15868
rect 22736 15789 22816 15822
rect 22920 15868 23000 15881
rect 22920 15822 22933 15868
rect 22987 15822 23000 15868
rect 22920 15789 23000 15822
rect 22552 15256 22632 15289
rect 22552 15210 22565 15256
rect 22619 15210 22632 15256
rect 22552 15197 22632 15210
rect 22736 15256 22816 15289
rect 22736 15210 22749 15256
rect 22803 15210 22816 15256
rect 22736 15197 22816 15210
rect 22920 15256 23000 15289
rect 22920 15210 22933 15256
rect 22987 15210 23000 15256
rect 22920 15197 23000 15210
rect 25108 15868 25188 15881
rect 25108 15822 25121 15868
rect 25175 15822 25188 15868
rect 25108 15789 25188 15822
rect 25292 15868 25372 15881
rect 25292 15822 25305 15868
rect 25359 15822 25372 15868
rect 25292 15789 25372 15822
rect 25476 15868 25556 15881
rect 25476 15822 25489 15868
rect 25543 15822 25556 15868
rect 25476 15789 25556 15822
rect 25108 15256 25188 15289
rect 25108 15210 25121 15256
rect 25175 15210 25188 15256
rect 25108 15197 25188 15210
rect 25292 15256 25372 15289
rect 25292 15210 25305 15256
rect 25359 15210 25372 15256
rect 25292 15197 25372 15210
rect 25476 15256 25556 15289
rect 25476 15210 25489 15256
rect 25543 15210 25556 15256
rect 25476 15197 25556 15210
rect 26594 15868 26674 15881
rect 26594 15822 26607 15868
rect 26661 15822 26674 15868
rect 26594 15789 26674 15822
rect 26778 15868 26858 15881
rect 26778 15822 26791 15868
rect 26845 15822 26858 15868
rect 26778 15789 26858 15822
rect 26962 15868 27042 15881
rect 26962 15822 26975 15868
rect 27029 15822 27042 15868
rect 26962 15789 27042 15822
rect 26594 15256 26674 15289
rect 26594 15210 26607 15256
rect 26661 15210 26674 15256
rect 26594 15197 26674 15210
rect 26778 15256 26858 15289
rect 26778 15210 26791 15256
rect 26845 15210 26858 15256
rect 26778 15197 26858 15210
rect 26962 15256 27042 15289
rect 26962 15210 26975 15256
rect 27029 15210 27042 15256
rect 26962 15197 27042 15210
rect 29150 15868 29230 15881
rect 29150 15822 29163 15868
rect 29217 15822 29230 15868
rect 29150 15789 29230 15822
rect 29334 15868 29414 15881
rect 29334 15822 29347 15868
rect 29401 15822 29414 15868
rect 29334 15789 29414 15822
rect 29518 15868 29598 15881
rect 29518 15822 29531 15868
rect 29585 15822 29598 15868
rect 29518 15789 29598 15822
rect 29150 15256 29230 15289
rect 29150 15210 29163 15256
rect 29217 15210 29230 15256
rect 29150 15197 29230 15210
rect 29334 15256 29414 15289
rect 29334 15210 29347 15256
rect 29401 15210 29414 15256
rect 29334 15197 29414 15210
rect 29518 15256 29598 15289
rect 29518 15210 29531 15256
rect 29585 15210 29598 15256
rect 29518 15197 29598 15210
rect 30636 15868 30716 15881
rect 30636 15822 30649 15868
rect 30703 15822 30716 15868
rect 30636 15789 30716 15822
rect 30820 15868 30900 15881
rect 30820 15822 30833 15868
rect 30887 15822 30900 15868
rect 30820 15789 30900 15822
rect 31004 15868 31084 15881
rect 31004 15822 31017 15868
rect 31071 15822 31084 15868
rect 31004 15789 31084 15822
rect 30636 15256 30716 15289
rect 30636 15210 30649 15256
rect 30703 15210 30716 15256
rect 30636 15197 30716 15210
rect 30820 15256 30900 15289
rect 30820 15210 30833 15256
rect 30887 15210 30900 15256
rect 30820 15197 30900 15210
rect 31004 15256 31084 15289
rect 31004 15210 31017 15256
rect 31071 15210 31084 15256
rect 31004 15197 31084 15210
rect 4898 14711 4978 14724
rect 4898 14665 4911 14711
rect 4965 14665 4978 14711
rect 4898 14632 4978 14665
rect 5082 14711 5162 14724
rect 5082 14665 5095 14711
rect 5149 14665 5162 14711
rect 5082 14632 5162 14665
rect 5266 14711 5346 14724
rect 5266 14665 5279 14711
rect 5333 14665 5346 14711
rect 5266 14632 5346 14665
rect 4898 14399 4978 14432
rect 4898 14353 4911 14399
rect 4965 14353 4978 14399
rect 4898 14340 4978 14353
rect 5082 14399 5162 14432
rect 5082 14353 5095 14399
rect 5149 14353 5162 14399
rect 5082 14340 5162 14353
rect 5266 14399 5346 14432
rect 5266 14353 5279 14399
rect 5333 14353 5346 14399
rect 5266 14340 5346 14353
rect 6384 14711 6464 14724
rect 6384 14665 6397 14711
rect 6451 14665 6464 14711
rect 6384 14632 6464 14665
rect 6568 14711 6648 14724
rect 6568 14665 6581 14711
rect 6635 14665 6648 14711
rect 6568 14632 6648 14665
rect 6752 14711 6832 14724
rect 6752 14665 6765 14711
rect 6819 14665 6832 14711
rect 6752 14632 6832 14665
rect 6384 14399 6464 14432
rect 6384 14353 6397 14399
rect 6451 14353 6464 14399
rect 6384 14340 6464 14353
rect 6568 14399 6648 14432
rect 6568 14353 6581 14399
rect 6635 14353 6648 14399
rect 6568 14340 6648 14353
rect 6752 14399 6832 14432
rect 6752 14353 6765 14399
rect 6819 14353 6832 14399
rect 6752 14340 6832 14353
rect 8940 14708 9020 14721
rect 8940 14662 8953 14708
rect 9007 14662 9020 14708
rect 8940 14629 9020 14662
rect 9124 14708 9204 14721
rect 9124 14662 9137 14708
rect 9191 14662 9204 14708
rect 9124 14629 9204 14662
rect 9308 14708 9388 14721
rect 9308 14662 9321 14708
rect 9375 14662 9388 14708
rect 9308 14629 9388 14662
rect 8940 14396 9020 14429
rect 8940 14350 8953 14396
rect 9007 14350 9020 14396
rect 8940 14337 9020 14350
rect 9124 14396 9204 14429
rect 9124 14350 9137 14396
rect 9191 14350 9204 14396
rect 9124 14337 9204 14350
rect 9308 14396 9388 14429
rect 9308 14350 9321 14396
rect 9375 14350 9388 14396
rect 9308 14337 9388 14350
rect 10426 14708 10506 14721
rect 10426 14662 10439 14708
rect 10493 14662 10506 14708
rect 10426 14629 10506 14662
rect 10610 14708 10690 14721
rect 10610 14662 10623 14708
rect 10677 14662 10690 14708
rect 10610 14629 10690 14662
rect 10794 14708 10874 14721
rect 10794 14662 10807 14708
rect 10861 14662 10874 14708
rect 10794 14629 10874 14662
rect 10426 14396 10506 14429
rect 10426 14350 10439 14396
rect 10493 14350 10506 14396
rect 10426 14337 10506 14350
rect 10610 14396 10690 14429
rect 10610 14350 10623 14396
rect 10677 14350 10690 14396
rect 10610 14337 10690 14350
rect 10794 14396 10874 14429
rect 10794 14350 10807 14396
rect 10861 14350 10874 14396
rect 10794 14337 10874 14350
rect 12982 14708 13062 14721
rect 12982 14662 12995 14708
rect 13049 14662 13062 14708
rect 12982 14629 13062 14662
rect 13166 14708 13246 14721
rect 13166 14662 13179 14708
rect 13233 14662 13246 14708
rect 13166 14629 13246 14662
rect 13350 14708 13430 14721
rect 13350 14662 13363 14708
rect 13417 14662 13430 14708
rect 13350 14629 13430 14662
rect 12982 14396 13062 14429
rect 12982 14350 12995 14396
rect 13049 14350 13062 14396
rect 12982 14337 13062 14350
rect 13166 14396 13246 14429
rect 13166 14350 13179 14396
rect 13233 14350 13246 14396
rect 13166 14337 13246 14350
rect 13350 14396 13430 14429
rect 13350 14350 13363 14396
rect 13417 14350 13430 14396
rect 13350 14337 13430 14350
rect 14468 14708 14548 14721
rect 14468 14662 14481 14708
rect 14535 14662 14548 14708
rect 14468 14629 14548 14662
rect 14652 14708 14732 14721
rect 14652 14662 14665 14708
rect 14719 14662 14732 14708
rect 14652 14629 14732 14662
rect 14836 14708 14916 14721
rect 14836 14662 14849 14708
rect 14903 14662 14916 14708
rect 14836 14629 14916 14662
rect 14468 14396 14548 14429
rect 14468 14350 14481 14396
rect 14535 14350 14548 14396
rect 14468 14337 14548 14350
rect 14652 14396 14732 14429
rect 14652 14350 14665 14396
rect 14719 14350 14732 14396
rect 14652 14337 14732 14350
rect 14836 14396 14916 14429
rect 14836 14350 14849 14396
rect 14903 14350 14916 14396
rect 14836 14337 14916 14350
rect 17024 14708 17104 14721
rect 17024 14662 17037 14708
rect 17091 14662 17104 14708
rect 17024 14629 17104 14662
rect 17208 14708 17288 14721
rect 17208 14662 17221 14708
rect 17275 14662 17288 14708
rect 17208 14629 17288 14662
rect 17392 14708 17472 14721
rect 17392 14662 17405 14708
rect 17459 14662 17472 14708
rect 17392 14629 17472 14662
rect 17024 14396 17104 14429
rect 17024 14350 17037 14396
rect 17091 14350 17104 14396
rect 17024 14337 17104 14350
rect 17208 14396 17288 14429
rect 17208 14350 17221 14396
rect 17275 14350 17288 14396
rect 17208 14337 17288 14350
rect 17392 14396 17472 14429
rect 17392 14350 17405 14396
rect 17459 14350 17472 14396
rect 17392 14337 17472 14350
rect 18510 14708 18590 14721
rect 18510 14662 18523 14708
rect 18577 14662 18590 14708
rect 18510 14629 18590 14662
rect 18694 14708 18774 14721
rect 18694 14662 18707 14708
rect 18761 14662 18774 14708
rect 18694 14629 18774 14662
rect 18878 14708 18958 14721
rect 18878 14662 18891 14708
rect 18945 14662 18958 14708
rect 18878 14629 18958 14662
rect 18510 14396 18590 14429
rect 18510 14350 18523 14396
rect 18577 14350 18590 14396
rect 18510 14337 18590 14350
rect 18694 14396 18774 14429
rect 18694 14350 18707 14396
rect 18761 14350 18774 14396
rect 18694 14337 18774 14350
rect 18878 14396 18958 14429
rect 18878 14350 18891 14396
rect 18945 14350 18958 14396
rect 18878 14337 18958 14350
rect 21066 14708 21146 14721
rect 21066 14662 21079 14708
rect 21133 14662 21146 14708
rect 21066 14629 21146 14662
rect 21250 14708 21330 14721
rect 21250 14662 21263 14708
rect 21317 14662 21330 14708
rect 21250 14629 21330 14662
rect 21434 14708 21514 14721
rect 21434 14662 21447 14708
rect 21501 14662 21514 14708
rect 21434 14629 21514 14662
rect 21066 14396 21146 14429
rect 21066 14350 21079 14396
rect 21133 14350 21146 14396
rect 21066 14337 21146 14350
rect 21250 14396 21330 14429
rect 21250 14350 21263 14396
rect 21317 14350 21330 14396
rect 21250 14337 21330 14350
rect 21434 14396 21514 14429
rect 21434 14350 21447 14396
rect 21501 14350 21514 14396
rect 21434 14337 21514 14350
rect 22552 14708 22632 14721
rect 22552 14662 22565 14708
rect 22619 14662 22632 14708
rect 22552 14629 22632 14662
rect 22736 14708 22816 14721
rect 22736 14662 22749 14708
rect 22803 14662 22816 14708
rect 22736 14629 22816 14662
rect 22920 14708 23000 14721
rect 22920 14662 22933 14708
rect 22987 14662 23000 14708
rect 22920 14629 23000 14662
rect 22552 14396 22632 14429
rect 22552 14350 22565 14396
rect 22619 14350 22632 14396
rect 22552 14337 22632 14350
rect 22736 14396 22816 14429
rect 22736 14350 22749 14396
rect 22803 14350 22816 14396
rect 22736 14337 22816 14350
rect 22920 14396 23000 14429
rect 22920 14350 22933 14396
rect 22987 14350 23000 14396
rect 22920 14337 23000 14350
rect 25108 14708 25188 14721
rect 25108 14662 25121 14708
rect 25175 14662 25188 14708
rect 25108 14629 25188 14662
rect 25292 14708 25372 14721
rect 25292 14662 25305 14708
rect 25359 14662 25372 14708
rect 25292 14629 25372 14662
rect 25476 14708 25556 14721
rect 25476 14662 25489 14708
rect 25543 14662 25556 14708
rect 25476 14629 25556 14662
rect 25108 14396 25188 14429
rect 25108 14350 25121 14396
rect 25175 14350 25188 14396
rect 25108 14337 25188 14350
rect 25292 14396 25372 14429
rect 25292 14350 25305 14396
rect 25359 14350 25372 14396
rect 25292 14337 25372 14350
rect 25476 14396 25556 14429
rect 25476 14350 25489 14396
rect 25543 14350 25556 14396
rect 25476 14337 25556 14350
rect 26594 14708 26674 14721
rect 26594 14662 26607 14708
rect 26661 14662 26674 14708
rect 26594 14629 26674 14662
rect 26778 14708 26858 14721
rect 26778 14662 26791 14708
rect 26845 14662 26858 14708
rect 26778 14629 26858 14662
rect 26962 14708 27042 14721
rect 26962 14662 26975 14708
rect 27029 14662 27042 14708
rect 26962 14629 27042 14662
rect 26594 14396 26674 14429
rect 26594 14350 26607 14396
rect 26661 14350 26674 14396
rect 26594 14337 26674 14350
rect 26778 14396 26858 14429
rect 26778 14350 26791 14396
rect 26845 14350 26858 14396
rect 26778 14337 26858 14350
rect 26962 14396 27042 14429
rect 26962 14350 26975 14396
rect 27029 14350 27042 14396
rect 26962 14337 27042 14350
rect 29150 14708 29230 14721
rect 29150 14662 29163 14708
rect 29217 14662 29230 14708
rect 29150 14629 29230 14662
rect 29334 14708 29414 14721
rect 29334 14662 29347 14708
rect 29401 14662 29414 14708
rect 29334 14629 29414 14662
rect 29518 14708 29598 14721
rect 29518 14662 29531 14708
rect 29585 14662 29598 14708
rect 29518 14629 29598 14662
rect 29150 14396 29230 14429
rect 29150 14350 29163 14396
rect 29217 14350 29230 14396
rect 29150 14337 29230 14350
rect 29334 14396 29414 14429
rect 29334 14350 29347 14396
rect 29401 14350 29414 14396
rect 29334 14337 29414 14350
rect 29518 14396 29598 14429
rect 29518 14350 29531 14396
rect 29585 14350 29598 14396
rect 29518 14337 29598 14350
rect 30636 14708 30716 14721
rect 30636 14662 30649 14708
rect 30703 14662 30716 14708
rect 30636 14629 30716 14662
rect 30820 14708 30900 14721
rect 30820 14662 30833 14708
rect 30887 14662 30900 14708
rect 30820 14629 30900 14662
rect 31004 14708 31084 14721
rect 31004 14662 31017 14708
rect 31071 14662 31084 14708
rect 31004 14629 31084 14662
rect 30636 14396 30716 14429
rect 30636 14350 30649 14396
rect 30703 14350 30716 14396
rect 30636 14337 30716 14350
rect 30820 14396 30900 14429
rect 30820 14350 30833 14396
rect 30887 14350 30900 14396
rect 30820 14337 30900 14350
rect 31004 14396 31084 14429
rect 31004 14350 31017 14396
rect 31071 14350 31084 14396
rect 31004 14337 31084 14350
rect 4898 13666 4978 13679
rect 4898 13620 4911 13666
rect 4965 13620 4978 13666
rect 4898 13587 4978 13620
rect 5082 13666 5162 13679
rect 5082 13620 5095 13666
rect 5149 13620 5162 13666
rect 5082 13587 5162 13620
rect 5266 13666 5346 13679
rect 5266 13620 5279 13666
rect 5333 13620 5346 13666
rect 5266 13587 5346 13620
rect 4898 13054 4978 13087
rect 4898 13008 4911 13054
rect 4965 13008 4978 13054
rect 4898 12995 4978 13008
rect 5082 13054 5162 13087
rect 5082 13008 5095 13054
rect 5149 13008 5162 13054
rect 5082 12995 5162 13008
rect 5266 13054 5346 13087
rect 5266 13008 5279 13054
rect 5333 13008 5346 13054
rect 5266 12995 5346 13008
rect 6384 13667 6464 13680
rect 6384 13621 6397 13667
rect 6451 13621 6464 13667
rect 6384 13588 6464 13621
rect 6568 13667 6648 13680
rect 6568 13621 6581 13667
rect 6635 13621 6648 13667
rect 6568 13588 6648 13621
rect 6752 13667 6832 13680
rect 6752 13621 6765 13667
rect 6819 13621 6832 13667
rect 6752 13588 6832 13621
rect 6384 13055 6464 13088
rect 6384 13009 6397 13055
rect 6451 13009 6464 13055
rect 6384 12996 6464 13009
rect 6568 13055 6648 13088
rect 6568 13009 6581 13055
rect 6635 13009 6648 13055
rect 6568 12996 6648 13009
rect 6752 13055 6832 13088
rect 6752 13009 6765 13055
rect 6819 13009 6832 13055
rect 6752 12996 6832 13009
rect 8940 13663 9020 13676
rect 8940 13617 8953 13663
rect 9007 13617 9020 13663
rect 8940 13584 9020 13617
rect 9124 13663 9204 13676
rect 9124 13617 9137 13663
rect 9191 13617 9204 13663
rect 9124 13584 9204 13617
rect 9308 13663 9388 13676
rect 9308 13617 9321 13663
rect 9375 13617 9388 13663
rect 9308 13584 9388 13617
rect 8940 13051 9020 13084
rect 8940 13005 8953 13051
rect 9007 13005 9020 13051
rect 8940 12992 9020 13005
rect 9124 13051 9204 13084
rect 9124 13005 9137 13051
rect 9191 13005 9204 13051
rect 9124 12992 9204 13005
rect 9308 13051 9388 13084
rect 9308 13005 9321 13051
rect 9375 13005 9388 13051
rect 9308 12992 9388 13005
rect 10426 13664 10506 13677
rect 10426 13618 10439 13664
rect 10493 13618 10506 13664
rect 10426 13585 10506 13618
rect 10610 13664 10690 13677
rect 10610 13618 10623 13664
rect 10677 13618 10690 13664
rect 10610 13585 10690 13618
rect 10794 13664 10874 13677
rect 10794 13618 10807 13664
rect 10861 13618 10874 13664
rect 10794 13585 10874 13618
rect 10426 13052 10506 13085
rect 10426 13006 10439 13052
rect 10493 13006 10506 13052
rect 10426 12993 10506 13006
rect 10610 13052 10690 13085
rect 10610 13006 10623 13052
rect 10677 13006 10690 13052
rect 10610 12993 10690 13006
rect 10794 13052 10874 13085
rect 10794 13006 10807 13052
rect 10861 13006 10874 13052
rect 10794 12993 10874 13006
rect 12982 13663 13062 13676
rect 12982 13617 12995 13663
rect 13049 13617 13062 13663
rect 12982 13584 13062 13617
rect 13166 13663 13246 13676
rect 13166 13617 13179 13663
rect 13233 13617 13246 13663
rect 13166 13584 13246 13617
rect 13350 13663 13430 13676
rect 13350 13617 13363 13663
rect 13417 13617 13430 13663
rect 13350 13584 13430 13617
rect 12982 13051 13062 13084
rect 12982 13005 12995 13051
rect 13049 13005 13062 13051
rect 12982 12992 13062 13005
rect 13166 13051 13246 13084
rect 13166 13005 13179 13051
rect 13233 13005 13246 13051
rect 13166 12992 13246 13005
rect 13350 13051 13430 13084
rect 13350 13005 13363 13051
rect 13417 13005 13430 13051
rect 13350 12992 13430 13005
rect 14468 13664 14548 13677
rect 14468 13618 14481 13664
rect 14535 13618 14548 13664
rect 14468 13585 14548 13618
rect 14652 13664 14732 13677
rect 14652 13618 14665 13664
rect 14719 13618 14732 13664
rect 14652 13585 14732 13618
rect 14836 13664 14916 13677
rect 14836 13618 14849 13664
rect 14903 13618 14916 13664
rect 14836 13585 14916 13618
rect 14468 13052 14548 13085
rect 14468 13006 14481 13052
rect 14535 13006 14548 13052
rect 14468 12993 14548 13006
rect 14652 13052 14732 13085
rect 14652 13006 14665 13052
rect 14719 13006 14732 13052
rect 14652 12993 14732 13006
rect 14836 13052 14916 13085
rect 14836 13006 14849 13052
rect 14903 13006 14916 13052
rect 14836 12993 14916 13006
rect 17024 13663 17104 13676
rect 17024 13617 17037 13663
rect 17091 13617 17104 13663
rect 17024 13584 17104 13617
rect 17208 13663 17288 13676
rect 17208 13617 17221 13663
rect 17275 13617 17288 13663
rect 17208 13584 17288 13617
rect 17392 13663 17472 13676
rect 17392 13617 17405 13663
rect 17459 13617 17472 13663
rect 17392 13584 17472 13617
rect 17024 13051 17104 13084
rect 17024 13005 17037 13051
rect 17091 13005 17104 13051
rect 17024 12992 17104 13005
rect 17208 13051 17288 13084
rect 17208 13005 17221 13051
rect 17275 13005 17288 13051
rect 17208 12992 17288 13005
rect 17392 13051 17472 13084
rect 17392 13005 17405 13051
rect 17459 13005 17472 13051
rect 17392 12992 17472 13005
rect 18510 13664 18590 13677
rect 18510 13618 18523 13664
rect 18577 13618 18590 13664
rect 18510 13585 18590 13618
rect 18694 13664 18774 13677
rect 18694 13618 18707 13664
rect 18761 13618 18774 13664
rect 18694 13585 18774 13618
rect 18878 13664 18958 13677
rect 18878 13618 18891 13664
rect 18945 13618 18958 13664
rect 18878 13585 18958 13618
rect 18510 13052 18590 13085
rect 18510 13006 18523 13052
rect 18577 13006 18590 13052
rect 18510 12993 18590 13006
rect 18694 13052 18774 13085
rect 18694 13006 18707 13052
rect 18761 13006 18774 13052
rect 18694 12993 18774 13006
rect 18878 13052 18958 13085
rect 18878 13006 18891 13052
rect 18945 13006 18958 13052
rect 18878 12993 18958 13006
rect 21066 13663 21146 13676
rect 21066 13617 21079 13663
rect 21133 13617 21146 13663
rect 21066 13584 21146 13617
rect 21250 13663 21330 13676
rect 21250 13617 21263 13663
rect 21317 13617 21330 13663
rect 21250 13584 21330 13617
rect 21434 13663 21514 13676
rect 21434 13617 21447 13663
rect 21501 13617 21514 13663
rect 21434 13584 21514 13617
rect 21066 13051 21146 13084
rect 21066 13005 21079 13051
rect 21133 13005 21146 13051
rect 21066 12992 21146 13005
rect 21250 13051 21330 13084
rect 21250 13005 21263 13051
rect 21317 13005 21330 13051
rect 21250 12992 21330 13005
rect 21434 13051 21514 13084
rect 21434 13005 21447 13051
rect 21501 13005 21514 13051
rect 21434 12992 21514 13005
rect 22552 13664 22632 13677
rect 22552 13618 22565 13664
rect 22619 13618 22632 13664
rect 22552 13585 22632 13618
rect 22736 13664 22816 13677
rect 22736 13618 22749 13664
rect 22803 13618 22816 13664
rect 22736 13585 22816 13618
rect 22920 13664 23000 13677
rect 22920 13618 22933 13664
rect 22987 13618 23000 13664
rect 22920 13585 23000 13618
rect 22552 13052 22632 13085
rect 22552 13006 22565 13052
rect 22619 13006 22632 13052
rect 22552 12993 22632 13006
rect 22736 13052 22816 13085
rect 22736 13006 22749 13052
rect 22803 13006 22816 13052
rect 22736 12993 22816 13006
rect 22920 13052 23000 13085
rect 22920 13006 22933 13052
rect 22987 13006 23000 13052
rect 22920 12993 23000 13006
rect 25108 13663 25188 13676
rect 25108 13617 25121 13663
rect 25175 13617 25188 13663
rect 25108 13584 25188 13617
rect 25292 13663 25372 13676
rect 25292 13617 25305 13663
rect 25359 13617 25372 13663
rect 25292 13584 25372 13617
rect 25476 13663 25556 13676
rect 25476 13617 25489 13663
rect 25543 13617 25556 13663
rect 25476 13584 25556 13617
rect 25108 13051 25188 13084
rect 25108 13005 25121 13051
rect 25175 13005 25188 13051
rect 25108 12992 25188 13005
rect 25292 13051 25372 13084
rect 25292 13005 25305 13051
rect 25359 13005 25372 13051
rect 25292 12992 25372 13005
rect 25476 13051 25556 13084
rect 25476 13005 25489 13051
rect 25543 13005 25556 13051
rect 25476 12992 25556 13005
rect 26594 13664 26674 13677
rect 26594 13618 26607 13664
rect 26661 13618 26674 13664
rect 26594 13585 26674 13618
rect 26778 13664 26858 13677
rect 26778 13618 26791 13664
rect 26845 13618 26858 13664
rect 26778 13585 26858 13618
rect 26962 13664 27042 13677
rect 26962 13618 26975 13664
rect 27029 13618 27042 13664
rect 26962 13585 27042 13618
rect 26594 13052 26674 13085
rect 26594 13006 26607 13052
rect 26661 13006 26674 13052
rect 26594 12993 26674 13006
rect 26778 13052 26858 13085
rect 26778 13006 26791 13052
rect 26845 13006 26858 13052
rect 26778 12993 26858 13006
rect 26962 13052 27042 13085
rect 26962 13006 26975 13052
rect 27029 13006 27042 13052
rect 26962 12993 27042 13006
rect 29150 13663 29230 13676
rect 29150 13617 29163 13663
rect 29217 13617 29230 13663
rect 29150 13584 29230 13617
rect 29334 13663 29414 13676
rect 29334 13617 29347 13663
rect 29401 13617 29414 13663
rect 29334 13584 29414 13617
rect 29518 13663 29598 13676
rect 29518 13617 29531 13663
rect 29585 13617 29598 13663
rect 29518 13584 29598 13617
rect 29150 13051 29230 13084
rect 29150 13005 29163 13051
rect 29217 13005 29230 13051
rect 29150 12992 29230 13005
rect 29334 13051 29414 13084
rect 29334 13005 29347 13051
rect 29401 13005 29414 13051
rect 29334 12992 29414 13005
rect 29518 13051 29598 13084
rect 29518 13005 29531 13051
rect 29585 13005 29598 13051
rect 29518 12992 29598 13005
rect 30636 13664 30716 13677
rect 30636 13618 30649 13664
rect 30703 13618 30716 13664
rect 30636 13585 30716 13618
rect 30820 13664 30900 13677
rect 30820 13618 30833 13664
rect 30887 13618 30900 13664
rect 30820 13585 30900 13618
rect 31004 13664 31084 13677
rect 31004 13618 31017 13664
rect 31071 13618 31084 13664
rect 31004 13585 31084 13618
rect 30636 13052 30716 13085
rect 30636 13006 30649 13052
rect 30703 13006 30716 13052
rect 30636 12993 30716 13006
rect 30820 13052 30900 13085
rect 30820 13006 30833 13052
rect 30887 13006 30900 13052
rect 30820 12993 30900 13006
rect 31004 13052 31084 13085
rect 31004 13006 31017 13052
rect 31071 13006 31084 13052
rect 31004 12993 31084 13006
rect 4898 12506 4978 12519
rect 4898 12460 4911 12506
rect 4965 12460 4978 12506
rect 4898 12427 4978 12460
rect 5082 12506 5162 12519
rect 5082 12460 5095 12506
rect 5149 12460 5162 12506
rect 5082 12427 5162 12460
rect 5266 12506 5346 12519
rect 5266 12460 5279 12506
rect 5333 12460 5346 12506
rect 5266 12427 5346 12460
rect 4898 12194 4978 12227
rect 4898 12148 4911 12194
rect 4965 12148 4978 12194
rect 4898 12135 4978 12148
rect 5082 12194 5162 12227
rect 5082 12148 5095 12194
rect 5149 12148 5162 12194
rect 5082 12135 5162 12148
rect 5266 12194 5346 12227
rect 5266 12148 5279 12194
rect 5333 12148 5346 12194
rect 5266 12135 5346 12148
rect 6384 12507 6464 12520
rect 6384 12461 6397 12507
rect 6451 12461 6464 12507
rect 6384 12428 6464 12461
rect 6568 12507 6648 12520
rect 6568 12461 6581 12507
rect 6635 12461 6648 12507
rect 6568 12428 6648 12461
rect 6752 12507 6832 12520
rect 6752 12461 6765 12507
rect 6819 12461 6832 12507
rect 6752 12428 6832 12461
rect 6384 12195 6464 12228
rect 6384 12149 6397 12195
rect 6451 12149 6464 12195
rect 6384 12136 6464 12149
rect 6568 12195 6648 12228
rect 6568 12149 6581 12195
rect 6635 12149 6648 12195
rect 6568 12136 6648 12149
rect 6752 12195 6832 12228
rect 6752 12149 6765 12195
rect 6819 12149 6832 12195
rect 6752 12136 6832 12149
rect 8940 12503 9020 12516
rect 8940 12457 8953 12503
rect 9007 12457 9020 12503
rect 8940 12424 9020 12457
rect 9124 12503 9204 12516
rect 9124 12457 9137 12503
rect 9191 12457 9204 12503
rect 9124 12424 9204 12457
rect 9308 12503 9388 12516
rect 9308 12457 9321 12503
rect 9375 12457 9388 12503
rect 9308 12424 9388 12457
rect 8940 12191 9020 12224
rect 8940 12145 8953 12191
rect 9007 12145 9020 12191
rect 8940 12132 9020 12145
rect 9124 12191 9204 12224
rect 9124 12145 9137 12191
rect 9191 12145 9204 12191
rect 9124 12132 9204 12145
rect 9308 12191 9388 12224
rect 9308 12145 9321 12191
rect 9375 12145 9388 12191
rect 9308 12132 9388 12145
rect 10426 12504 10506 12517
rect 10426 12458 10439 12504
rect 10493 12458 10506 12504
rect 10426 12425 10506 12458
rect 10610 12504 10690 12517
rect 10610 12458 10623 12504
rect 10677 12458 10690 12504
rect 10610 12425 10690 12458
rect 10794 12504 10874 12517
rect 10794 12458 10807 12504
rect 10861 12458 10874 12504
rect 10794 12425 10874 12458
rect 10426 12192 10506 12225
rect 10426 12146 10439 12192
rect 10493 12146 10506 12192
rect 10426 12133 10506 12146
rect 10610 12192 10690 12225
rect 10610 12146 10623 12192
rect 10677 12146 10690 12192
rect 10610 12133 10690 12146
rect 10794 12192 10874 12225
rect 10794 12146 10807 12192
rect 10861 12146 10874 12192
rect 10794 12133 10874 12146
rect 12982 12503 13062 12516
rect 12982 12457 12995 12503
rect 13049 12457 13062 12503
rect 12982 12424 13062 12457
rect 13166 12503 13246 12516
rect 13166 12457 13179 12503
rect 13233 12457 13246 12503
rect 13166 12424 13246 12457
rect 13350 12503 13430 12516
rect 13350 12457 13363 12503
rect 13417 12457 13430 12503
rect 13350 12424 13430 12457
rect 12982 12191 13062 12224
rect 12982 12145 12995 12191
rect 13049 12145 13062 12191
rect 12982 12132 13062 12145
rect 13166 12191 13246 12224
rect 13166 12145 13179 12191
rect 13233 12145 13246 12191
rect 13166 12132 13246 12145
rect 13350 12191 13430 12224
rect 13350 12145 13363 12191
rect 13417 12145 13430 12191
rect 13350 12132 13430 12145
rect 14468 12504 14548 12517
rect 14468 12458 14481 12504
rect 14535 12458 14548 12504
rect 14468 12425 14548 12458
rect 14652 12504 14732 12517
rect 14652 12458 14665 12504
rect 14719 12458 14732 12504
rect 14652 12425 14732 12458
rect 14836 12504 14916 12517
rect 14836 12458 14849 12504
rect 14903 12458 14916 12504
rect 14836 12425 14916 12458
rect 14468 12192 14548 12225
rect 14468 12146 14481 12192
rect 14535 12146 14548 12192
rect 14468 12133 14548 12146
rect 14652 12192 14732 12225
rect 14652 12146 14665 12192
rect 14719 12146 14732 12192
rect 14652 12133 14732 12146
rect 14836 12192 14916 12225
rect 14836 12146 14849 12192
rect 14903 12146 14916 12192
rect 14836 12133 14916 12146
rect 17024 12503 17104 12516
rect 17024 12457 17037 12503
rect 17091 12457 17104 12503
rect 17024 12424 17104 12457
rect 17208 12503 17288 12516
rect 17208 12457 17221 12503
rect 17275 12457 17288 12503
rect 17208 12424 17288 12457
rect 17392 12503 17472 12516
rect 17392 12457 17405 12503
rect 17459 12457 17472 12503
rect 17392 12424 17472 12457
rect 17024 12191 17104 12224
rect 17024 12145 17037 12191
rect 17091 12145 17104 12191
rect 17024 12132 17104 12145
rect 17208 12191 17288 12224
rect 17208 12145 17221 12191
rect 17275 12145 17288 12191
rect 17208 12132 17288 12145
rect 17392 12191 17472 12224
rect 17392 12145 17405 12191
rect 17459 12145 17472 12191
rect 17392 12132 17472 12145
rect 18510 12504 18590 12517
rect 18510 12458 18523 12504
rect 18577 12458 18590 12504
rect 18510 12425 18590 12458
rect 18694 12504 18774 12517
rect 18694 12458 18707 12504
rect 18761 12458 18774 12504
rect 18694 12425 18774 12458
rect 18878 12504 18958 12517
rect 18878 12458 18891 12504
rect 18945 12458 18958 12504
rect 18878 12425 18958 12458
rect 18510 12192 18590 12225
rect 18510 12146 18523 12192
rect 18577 12146 18590 12192
rect 18510 12133 18590 12146
rect 18694 12192 18774 12225
rect 18694 12146 18707 12192
rect 18761 12146 18774 12192
rect 18694 12133 18774 12146
rect 18878 12192 18958 12225
rect 18878 12146 18891 12192
rect 18945 12146 18958 12192
rect 18878 12133 18958 12146
rect 21066 12503 21146 12516
rect 21066 12457 21079 12503
rect 21133 12457 21146 12503
rect 21066 12424 21146 12457
rect 21250 12503 21330 12516
rect 21250 12457 21263 12503
rect 21317 12457 21330 12503
rect 21250 12424 21330 12457
rect 21434 12503 21514 12516
rect 21434 12457 21447 12503
rect 21501 12457 21514 12503
rect 21434 12424 21514 12457
rect 21066 12191 21146 12224
rect 21066 12145 21079 12191
rect 21133 12145 21146 12191
rect 21066 12132 21146 12145
rect 21250 12191 21330 12224
rect 21250 12145 21263 12191
rect 21317 12145 21330 12191
rect 21250 12132 21330 12145
rect 21434 12191 21514 12224
rect 21434 12145 21447 12191
rect 21501 12145 21514 12191
rect 21434 12132 21514 12145
rect 22552 12504 22632 12517
rect 22552 12458 22565 12504
rect 22619 12458 22632 12504
rect 22552 12425 22632 12458
rect 22736 12504 22816 12517
rect 22736 12458 22749 12504
rect 22803 12458 22816 12504
rect 22736 12425 22816 12458
rect 22920 12504 23000 12517
rect 22920 12458 22933 12504
rect 22987 12458 23000 12504
rect 22920 12425 23000 12458
rect 22552 12192 22632 12225
rect 22552 12146 22565 12192
rect 22619 12146 22632 12192
rect 22552 12133 22632 12146
rect 22736 12192 22816 12225
rect 22736 12146 22749 12192
rect 22803 12146 22816 12192
rect 22736 12133 22816 12146
rect 22920 12192 23000 12225
rect 22920 12146 22933 12192
rect 22987 12146 23000 12192
rect 22920 12133 23000 12146
rect 25108 12503 25188 12516
rect 25108 12457 25121 12503
rect 25175 12457 25188 12503
rect 25108 12424 25188 12457
rect 25292 12503 25372 12516
rect 25292 12457 25305 12503
rect 25359 12457 25372 12503
rect 25292 12424 25372 12457
rect 25476 12503 25556 12516
rect 25476 12457 25489 12503
rect 25543 12457 25556 12503
rect 25476 12424 25556 12457
rect 25108 12191 25188 12224
rect 25108 12145 25121 12191
rect 25175 12145 25188 12191
rect 25108 12132 25188 12145
rect 25292 12191 25372 12224
rect 25292 12145 25305 12191
rect 25359 12145 25372 12191
rect 25292 12132 25372 12145
rect 25476 12191 25556 12224
rect 25476 12145 25489 12191
rect 25543 12145 25556 12191
rect 25476 12132 25556 12145
rect 26594 12504 26674 12517
rect 26594 12458 26607 12504
rect 26661 12458 26674 12504
rect 26594 12425 26674 12458
rect 26778 12504 26858 12517
rect 26778 12458 26791 12504
rect 26845 12458 26858 12504
rect 26778 12425 26858 12458
rect 26962 12504 27042 12517
rect 26962 12458 26975 12504
rect 27029 12458 27042 12504
rect 26962 12425 27042 12458
rect 26594 12192 26674 12225
rect 26594 12146 26607 12192
rect 26661 12146 26674 12192
rect 26594 12133 26674 12146
rect 26778 12192 26858 12225
rect 26778 12146 26791 12192
rect 26845 12146 26858 12192
rect 26778 12133 26858 12146
rect 26962 12192 27042 12225
rect 26962 12146 26975 12192
rect 27029 12146 27042 12192
rect 26962 12133 27042 12146
rect 29150 12503 29230 12516
rect 29150 12457 29163 12503
rect 29217 12457 29230 12503
rect 29150 12424 29230 12457
rect 29334 12503 29414 12516
rect 29334 12457 29347 12503
rect 29401 12457 29414 12503
rect 29334 12424 29414 12457
rect 29518 12503 29598 12516
rect 29518 12457 29531 12503
rect 29585 12457 29598 12503
rect 29518 12424 29598 12457
rect 29150 12191 29230 12224
rect 29150 12145 29163 12191
rect 29217 12145 29230 12191
rect 29150 12132 29230 12145
rect 29334 12191 29414 12224
rect 29334 12145 29347 12191
rect 29401 12145 29414 12191
rect 29334 12132 29414 12145
rect 29518 12191 29598 12224
rect 29518 12145 29531 12191
rect 29585 12145 29598 12191
rect 29518 12132 29598 12145
rect 30636 12504 30716 12517
rect 30636 12458 30649 12504
rect 30703 12458 30716 12504
rect 30636 12425 30716 12458
rect 30820 12504 30900 12517
rect 30820 12458 30833 12504
rect 30887 12458 30900 12504
rect 30820 12425 30900 12458
rect 31004 12504 31084 12517
rect 31004 12458 31017 12504
rect 31071 12458 31084 12504
rect 31004 12425 31084 12458
rect 30636 12192 30716 12225
rect 30636 12146 30649 12192
rect 30703 12146 30716 12192
rect 30636 12133 30716 12146
rect 30820 12192 30900 12225
rect 30820 12146 30833 12192
rect 30887 12146 30900 12192
rect 30820 12133 30900 12146
rect 31004 12192 31084 12225
rect 31004 12146 31017 12192
rect 31071 12146 31084 12192
rect 31004 12133 31084 12146
rect 4898 11461 4978 11474
rect 4898 11415 4911 11461
rect 4965 11415 4978 11461
rect 4898 11382 4978 11415
rect 5082 11461 5162 11474
rect 5082 11415 5095 11461
rect 5149 11415 5162 11461
rect 5082 11382 5162 11415
rect 5266 11461 5346 11474
rect 5266 11415 5279 11461
rect 5333 11415 5346 11461
rect 5266 11382 5346 11415
rect 4898 10849 4978 10882
rect 4898 10803 4911 10849
rect 4965 10803 4978 10849
rect 4898 10790 4978 10803
rect 5082 10849 5162 10882
rect 5082 10803 5095 10849
rect 5149 10803 5162 10849
rect 5082 10790 5162 10803
rect 5266 10849 5346 10882
rect 5266 10803 5279 10849
rect 5333 10803 5346 10849
rect 5266 10790 5346 10803
rect 8940 11458 9020 11471
rect 8940 11412 8953 11458
rect 9007 11412 9020 11458
rect 8940 11379 9020 11412
rect 9124 11458 9204 11471
rect 9124 11412 9137 11458
rect 9191 11412 9204 11458
rect 9124 11379 9204 11412
rect 9308 11458 9388 11471
rect 9308 11412 9321 11458
rect 9375 11412 9388 11458
rect 9308 11379 9388 11412
rect 8940 10846 9020 10879
rect 8940 10800 8953 10846
rect 9007 10800 9020 10846
rect 8940 10787 9020 10800
rect 9124 10846 9204 10879
rect 9124 10800 9137 10846
rect 9191 10800 9204 10846
rect 9124 10787 9204 10800
rect 9308 10846 9388 10879
rect 9308 10800 9321 10846
rect 9375 10800 9388 10846
rect 9308 10787 9388 10800
rect 12982 11458 13062 11471
rect 12982 11412 12995 11458
rect 13049 11412 13062 11458
rect 12982 11379 13062 11412
rect 13166 11458 13246 11471
rect 13166 11412 13179 11458
rect 13233 11412 13246 11458
rect 13166 11379 13246 11412
rect 13350 11458 13430 11471
rect 13350 11412 13363 11458
rect 13417 11412 13430 11458
rect 13350 11379 13430 11412
rect 12982 10846 13062 10879
rect 12982 10800 12995 10846
rect 13049 10800 13062 10846
rect 12982 10787 13062 10800
rect 13166 10846 13246 10879
rect 13166 10800 13179 10846
rect 13233 10800 13246 10846
rect 13166 10787 13246 10800
rect 13350 10846 13430 10879
rect 13350 10800 13363 10846
rect 13417 10800 13430 10846
rect 13350 10787 13430 10800
rect 17024 11458 17104 11471
rect 17024 11412 17037 11458
rect 17091 11412 17104 11458
rect 17024 11379 17104 11412
rect 17208 11458 17288 11471
rect 17208 11412 17221 11458
rect 17275 11412 17288 11458
rect 17208 11379 17288 11412
rect 17392 11458 17472 11471
rect 17392 11412 17405 11458
rect 17459 11412 17472 11458
rect 17392 11379 17472 11412
rect 17024 10846 17104 10879
rect 17024 10800 17037 10846
rect 17091 10800 17104 10846
rect 17024 10787 17104 10800
rect 17208 10846 17288 10879
rect 17208 10800 17221 10846
rect 17275 10800 17288 10846
rect 17208 10787 17288 10800
rect 17392 10846 17472 10879
rect 17392 10800 17405 10846
rect 17459 10800 17472 10846
rect 17392 10787 17472 10800
rect 21066 11458 21146 11471
rect 21066 11412 21079 11458
rect 21133 11412 21146 11458
rect 21066 11379 21146 11412
rect 21250 11458 21330 11471
rect 21250 11412 21263 11458
rect 21317 11412 21330 11458
rect 21250 11379 21330 11412
rect 21434 11458 21514 11471
rect 21434 11412 21447 11458
rect 21501 11412 21514 11458
rect 21434 11379 21514 11412
rect 21066 10846 21146 10879
rect 21066 10800 21079 10846
rect 21133 10800 21146 10846
rect 21066 10787 21146 10800
rect 21250 10846 21330 10879
rect 21250 10800 21263 10846
rect 21317 10800 21330 10846
rect 21250 10787 21330 10800
rect 21434 10846 21514 10879
rect 21434 10800 21447 10846
rect 21501 10800 21514 10846
rect 21434 10787 21514 10800
rect 25108 11458 25188 11471
rect 25108 11412 25121 11458
rect 25175 11412 25188 11458
rect 25108 11379 25188 11412
rect 25292 11458 25372 11471
rect 25292 11412 25305 11458
rect 25359 11412 25372 11458
rect 25292 11379 25372 11412
rect 25476 11458 25556 11471
rect 25476 11412 25489 11458
rect 25543 11412 25556 11458
rect 25476 11379 25556 11412
rect 25108 10846 25188 10879
rect 25108 10800 25121 10846
rect 25175 10800 25188 10846
rect 25108 10787 25188 10800
rect 25292 10846 25372 10879
rect 25292 10800 25305 10846
rect 25359 10800 25372 10846
rect 25292 10787 25372 10800
rect 25476 10846 25556 10879
rect 25476 10800 25489 10846
rect 25543 10800 25556 10846
rect 25476 10787 25556 10800
rect 29150 11458 29230 11471
rect 29150 11412 29163 11458
rect 29217 11412 29230 11458
rect 29150 11379 29230 11412
rect 29334 11458 29414 11471
rect 29334 11412 29347 11458
rect 29401 11412 29414 11458
rect 29334 11379 29414 11412
rect 29518 11458 29598 11471
rect 29518 11412 29531 11458
rect 29585 11412 29598 11458
rect 29518 11379 29598 11412
rect 29150 10846 29230 10879
rect 29150 10800 29163 10846
rect 29217 10800 29230 10846
rect 29150 10787 29230 10800
rect 29334 10846 29414 10879
rect 29334 10800 29347 10846
rect 29401 10800 29414 10846
rect 29334 10787 29414 10800
rect 29518 10846 29598 10879
rect 29518 10800 29531 10846
rect 29585 10800 29598 10846
rect 29518 10787 29598 10800
rect 4898 10301 4978 10314
rect 4898 10255 4911 10301
rect 4965 10255 4978 10301
rect 4898 10222 4978 10255
rect 5082 10301 5162 10314
rect 5082 10255 5095 10301
rect 5149 10255 5162 10301
rect 5082 10222 5162 10255
rect 5266 10301 5346 10314
rect 5266 10255 5279 10301
rect 5333 10255 5346 10301
rect 5266 10222 5346 10255
rect 4898 9989 4978 10022
rect 4898 9943 4911 9989
rect 4965 9943 4978 9989
rect 4898 9930 4978 9943
rect 5082 9989 5162 10022
rect 5082 9943 5095 9989
rect 5149 9943 5162 9989
rect 5082 9930 5162 9943
rect 5266 9989 5346 10022
rect 5266 9943 5279 9989
rect 5333 9943 5346 9989
rect 5266 9930 5346 9943
rect 8940 10298 9020 10311
rect 8940 10252 8953 10298
rect 9007 10252 9020 10298
rect 8940 10219 9020 10252
rect 9124 10298 9204 10311
rect 9124 10252 9137 10298
rect 9191 10252 9204 10298
rect 9124 10219 9204 10252
rect 9308 10298 9388 10311
rect 9308 10252 9321 10298
rect 9375 10252 9388 10298
rect 9308 10219 9388 10252
rect 8940 9986 9020 10019
rect 8940 9940 8953 9986
rect 9007 9940 9020 9986
rect 8940 9927 9020 9940
rect 9124 9986 9204 10019
rect 9124 9940 9137 9986
rect 9191 9940 9204 9986
rect 9124 9927 9204 9940
rect 9308 9986 9388 10019
rect 9308 9940 9321 9986
rect 9375 9940 9388 9986
rect 9308 9927 9388 9940
rect 12982 10298 13062 10311
rect 12982 10252 12995 10298
rect 13049 10252 13062 10298
rect 12982 10219 13062 10252
rect 13166 10298 13246 10311
rect 13166 10252 13179 10298
rect 13233 10252 13246 10298
rect 13166 10219 13246 10252
rect 13350 10298 13430 10311
rect 13350 10252 13363 10298
rect 13417 10252 13430 10298
rect 13350 10219 13430 10252
rect 12982 9986 13062 10019
rect 12982 9940 12995 9986
rect 13049 9940 13062 9986
rect 12982 9927 13062 9940
rect 13166 9986 13246 10019
rect 13166 9940 13179 9986
rect 13233 9940 13246 9986
rect 13166 9927 13246 9940
rect 13350 9986 13430 10019
rect 13350 9940 13363 9986
rect 13417 9940 13430 9986
rect 13350 9927 13430 9940
rect 17024 10298 17104 10311
rect 17024 10252 17037 10298
rect 17091 10252 17104 10298
rect 17024 10219 17104 10252
rect 17208 10298 17288 10311
rect 17208 10252 17221 10298
rect 17275 10252 17288 10298
rect 17208 10219 17288 10252
rect 17392 10298 17472 10311
rect 17392 10252 17405 10298
rect 17459 10252 17472 10298
rect 17392 10219 17472 10252
rect 17024 9986 17104 10019
rect 17024 9940 17037 9986
rect 17091 9940 17104 9986
rect 17024 9927 17104 9940
rect 17208 9986 17288 10019
rect 17208 9940 17221 9986
rect 17275 9940 17288 9986
rect 17208 9927 17288 9940
rect 17392 9986 17472 10019
rect 17392 9940 17405 9986
rect 17459 9940 17472 9986
rect 17392 9927 17472 9940
rect 21066 10298 21146 10311
rect 21066 10252 21079 10298
rect 21133 10252 21146 10298
rect 21066 10219 21146 10252
rect 21250 10298 21330 10311
rect 21250 10252 21263 10298
rect 21317 10252 21330 10298
rect 21250 10219 21330 10252
rect 21434 10298 21514 10311
rect 21434 10252 21447 10298
rect 21501 10252 21514 10298
rect 21434 10219 21514 10252
rect 21066 9986 21146 10019
rect 21066 9940 21079 9986
rect 21133 9940 21146 9986
rect 21066 9927 21146 9940
rect 21250 9986 21330 10019
rect 21250 9940 21263 9986
rect 21317 9940 21330 9986
rect 21250 9927 21330 9940
rect 21434 9986 21514 10019
rect 21434 9940 21447 9986
rect 21501 9940 21514 9986
rect 21434 9927 21514 9940
rect 25108 10298 25188 10311
rect 25108 10252 25121 10298
rect 25175 10252 25188 10298
rect 25108 10219 25188 10252
rect 25292 10298 25372 10311
rect 25292 10252 25305 10298
rect 25359 10252 25372 10298
rect 25292 10219 25372 10252
rect 25476 10298 25556 10311
rect 25476 10252 25489 10298
rect 25543 10252 25556 10298
rect 25476 10219 25556 10252
rect 25108 9986 25188 10019
rect 25108 9940 25121 9986
rect 25175 9940 25188 9986
rect 25108 9927 25188 9940
rect 25292 9986 25372 10019
rect 25292 9940 25305 9986
rect 25359 9940 25372 9986
rect 25292 9927 25372 9940
rect 25476 9986 25556 10019
rect 25476 9940 25489 9986
rect 25543 9940 25556 9986
rect 25476 9927 25556 9940
rect 29150 10298 29230 10311
rect 29150 10252 29163 10298
rect 29217 10252 29230 10298
rect 29150 10219 29230 10252
rect 29334 10298 29414 10311
rect 29334 10252 29347 10298
rect 29401 10252 29414 10298
rect 29334 10219 29414 10252
rect 29518 10298 29598 10311
rect 29518 10252 29531 10298
rect 29585 10252 29598 10298
rect 29518 10219 29598 10252
rect 29150 9986 29230 10019
rect 29150 9940 29163 9986
rect 29217 9940 29230 9986
rect 29150 9927 29230 9940
rect 29334 9986 29414 10019
rect 29334 9940 29347 9986
rect 29401 9940 29414 9986
rect 29334 9927 29414 9940
rect 29518 9986 29598 10019
rect 29518 9940 29531 9986
rect 29585 9940 29598 9986
rect 29518 9927 29598 9940
rect 886 8497 966 8510
rect 886 8451 899 8497
rect 953 8451 966 8497
rect 886 8418 966 8451
rect 1070 8497 1150 8510
rect 1070 8451 1083 8497
rect 1137 8451 1150 8497
rect 1070 8418 1150 8451
rect 1254 8497 1334 8510
rect 1254 8451 1267 8497
rect 1321 8451 1334 8497
rect 1254 8418 1334 8451
rect 886 7885 966 7918
rect 886 7839 899 7885
rect 953 7839 966 7885
rect 886 7826 966 7839
rect 1070 7885 1150 7918
rect 1070 7839 1083 7885
rect 1137 7839 1150 7885
rect 1070 7826 1150 7839
rect 1254 7885 1334 7918
rect 1254 7839 1267 7885
rect 1321 7839 1334 7885
rect 1254 7826 1334 7839
rect 4898 8497 4978 8510
rect 4898 8451 4911 8497
rect 4965 8451 4978 8497
rect 4898 8418 4978 8451
rect 5082 8497 5162 8510
rect 5082 8451 5095 8497
rect 5149 8451 5162 8497
rect 5082 8418 5162 8451
rect 5266 8497 5346 8510
rect 5266 8451 5279 8497
rect 5333 8451 5346 8497
rect 5266 8418 5346 8451
rect 4898 7885 4978 7918
rect 4898 7839 4911 7885
rect 4965 7839 4978 7885
rect 4898 7826 4978 7839
rect 5082 7885 5162 7918
rect 5082 7839 5095 7885
rect 5149 7839 5162 7885
rect 5082 7826 5162 7839
rect 5266 7885 5346 7918
rect 5266 7839 5279 7885
rect 5333 7839 5346 7885
rect 5266 7826 5346 7839
rect 8940 8497 9020 8510
rect 8940 8451 8953 8497
rect 9007 8451 9020 8497
rect 8940 8418 9020 8451
rect 9124 8497 9204 8510
rect 9124 8451 9137 8497
rect 9191 8451 9204 8497
rect 9124 8418 9204 8451
rect 9308 8497 9388 8510
rect 9308 8451 9321 8497
rect 9375 8451 9388 8497
rect 9308 8418 9388 8451
rect 8940 7885 9020 7918
rect 8940 7839 8953 7885
rect 9007 7839 9020 7885
rect 8940 7826 9020 7839
rect 9124 7885 9204 7918
rect 9124 7839 9137 7885
rect 9191 7839 9204 7885
rect 9124 7826 9204 7839
rect 9308 7885 9388 7918
rect 9308 7839 9321 7885
rect 9375 7839 9388 7885
rect 9308 7826 9388 7839
rect 12982 8497 13062 8510
rect 12982 8451 12995 8497
rect 13049 8451 13062 8497
rect 12982 8418 13062 8451
rect 13166 8497 13246 8510
rect 13166 8451 13179 8497
rect 13233 8451 13246 8497
rect 13166 8418 13246 8451
rect 13350 8497 13430 8510
rect 13350 8451 13363 8497
rect 13417 8451 13430 8497
rect 13350 8418 13430 8451
rect 12982 7885 13062 7918
rect 12982 7839 12995 7885
rect 13049 7839 13062 7885
rect 12982 7826 13062 7839
rect 13166 7885 13246 7918
rect 13166 7839 13179 7885
rect 13233 7839 13246 7885
rect 13166 7826 13246 7839
rect 13350 7885 13430 7918
rect 13350 7839 13363 7885
rect 13417 7839 13430 7885
rect 13350 7826 13430 7839
rect 17024 8497 17104 8510
rect 17024 8451 17037 8497
rect 17091 8451 17104 8497
rect 17024 8418 17104 8451
rect 17208 8497 17288 8510
rect 17208 8451 17221 8497
rect 17275 8451 17288 8497
rect 17208 8418 17288 8451
rect 17392 8497 17472 8510
rect 17392 8451 17405 8497
rect 17459 8451 17472 8497
rect 17392 8418 17472 8451
rect 17024 7885 17104 7918
rect 17024 7839 17037 7885
rect 17091 7839 17104 7885
rect 17024 7826 17104 7839
rect 17208 7885 17288 7918
rect 17208 7839 17221 7885
rect 17275 7839 17288 7885
rect 17208 7826 17288 7839
rect 17392 7885 17472 7918
rect 17392 7839 17405 7885
rect 17459 7839 17472 7885
rect 17392 7826 17472 7839
rect 21066 8497 21146 8510
rect 21066 8451 21079 8497
rect 21133 8451 21146 8497
rect 21066 8418 21146 8451
rect 21250 8497 21330 8510
rect 21250 8451 21263 8497
rect 21317 8451 21330 8497
rect 21250 8418 21330 8451
rect 21434 8497 21514 8510
rect 21434 8451 21447 8497
rect 21501 8451 21514 8497
rect 21434 8418 21514 8451
rect 21066 7885 21146 7918
rect 21066 7839 21079 7885
rect 21133 7839 21146 7885
rect 21066 7826 21146 7839
rect 21250 7885 21330 7918
rect 21250 7839 21263 7885
rect 21317 7839 21330 7885
rect 21250 7826 21330 7839
rect 21434 7885 21514 7918
rect 21434 7839 21447 7885
rect 21501 7839 21514 7885
rect 21434 7826 21514 7839
rect 25108 8497 25188 8510
rect 25108 8451 25121 8497
rect 25175 8451 25188 8497
rect 25108 8418 25188 8451
rect 25292 8497 25372 8510
rect 25292 8451 25305 8497
rect 25359 8451 25372 8497
rect 25292 8418 25372 8451
rect 25476 8497 25556 8510
rect 25476 8451 25489 8497
rect 25543 8451 25556 8497
rect 25476 8418 25556 8451
rect 25108 7885 25188 7918
rect 25108 7839 25121 7885
rect 25175 7839 25188 7885
rect 25108 7826 25188 7839
rect 25292 7885 25372 7918
rect 25292 7839 25305 7885
rect 25359 7839 25372 7885
rect 25292 7826 25372 7839
rect 25476 7885 25556 7918
rect 25476 7839 25489 7885
rect 25543 7839 25556 7885
rect 25476 7826 25556 7839
rect 886 7337 966 7350
rect 886 7291 899 7337
rect 953 7291 966 7337
rect 886 7258 966 7291
rect 1070 7337 1150 7350
rect 1070 7291 1083 7337
rect 1137 7291 1150 7337
rect 1070 7258 1150 7291
rect 1254 7337 1334 7350
rect 1254 7291 1267 7337
rect 1321 7291 1334 7337
rect 1254 7258 1334 7291
rect 886 7025 966 7058
rect 886 6979 899 7025
rect 953 6979 966 7025
rect 886 6966 966 6979
rect 1070 7025 1150 7058
rect 1070 6979 1083 7025
rect 1137 6979 1150 7025
rect 1070 6966 1150 6979
rect 1254 7025 1334 7058
rect 1254 6979 1267 7025
rect 1321 6979 1334 7025
rect 1254 6966 1334 6979
rect 4898 7337 4978 7350
rect 4898 7291 4911 7337
rect 4965 7291 4978 7337
rect 4898 7258 4978 7291
rect 5082 7337 5162 7350
rect 5082 7291 5095 7337
rect 5149 7291 5162 7337
rect 5082 7258 5162 7291
rect 5266 7337 5346 7350
rect 5266 7291 5279 7337
rect 5333 7291 5346 7337
rect 5266 7258 5346 7291
rect 4898 7025 4978 7058
rect 4898 6979 4911 7025
rect 4965 6979 4978 7025
rect 4898 6966 4978 6979
rect 5082 7025 5162 7058
rect 5082 6979 5095 7025
rect 5149 6979 5162 7025
rect 5082 6966 5162 6979
rect 5266 7025 5346 7058
rect 5266 6979 5279 7025
rect 5333 6979 5346 7025
rect 5266 6966 5346 6979
rect 8940 7337 9020 7350
rect 8940 7291 8953 7337
rect 9007 7291 9020 7337
rect 8940 7258 9020 7291
rect 9124 7337 9204 7350
rect 9124 7291 9137 7337
rect 9191 7291 9204 7337
rect 9124 7258 9204 7291
rect 9308 7337 9388 7350
rect 9308 7291 9321 7337
rect 9375 7291 9388 7337
rect 9308 7258 9388 7291
rect 8940 7025 9020 7058
rect 8940 6979 8953 7025
rect 9007 6979 9020 7025
rect 8940 6966 9020 6979
rect 9124 7025 9204 7058
rect 9124 6979 9137 7025
rect 9191 6979 9204 7025
rect 9124 6966 9204 6979
rect 9308 7025 9388 7058
rect 9308 6979 9321 7025
rect 9375 6979 9388 7025
rect 9308 6966 9388 6979
rect 12982 7337 13062 7350
rect 12982 7291 12995 7337
rect 13049 7291 13062 7337
rect 12982 7258 13062 7291
rect 13166 7337 13246 7350
rect 13166 7291 13179 7337
rect 13233 7291 13246 7337
rect 13166 7258 13246 7291
rect 13350 7337 13430 7350
rect 13350 7291 13363 7337
rect 13417 7291 13430 7337
rect 13350 7258 13430 7291
rect 12982 7025 13062 7058
rect 12982 6979 12995 7025
rect 13049 6979 13062 7025
rect 12982 6966 13062 6979
rect 13166 7025 13246 7058
rect 13166 6979 13179 7025
rect 13233 6979 13246 7025
rect 13166 6966 13246 6979
rect 13350 7025 13430 7058
rect 13350 6979 13363 7025
rect 13417 6979 13430 7025
rect 13350 6966 13430 6979
rect 17024 7337 17104 7350
rect 17024 7291 17037 7337
rect 17091 7291 17104 7337
rect 17024 7258 17104 7291
rect 17208 7337 17288 7350
rect 17208 7291 17221 7337
rect 17275 7291 17288 7337
rect 17208 7258 17288 7291
rect 17392 7337 17472 7350
rect 17392 7291 17405 7337
rect 17459 7291 17472 7337
rect 17392 7258 17472 7291
rect 17024 7025 17104 7058
rect 17024 6979 17037 7025
rect 17091 6979 17104 7025
rect 17024 6966 17104 6979
rect 17208 7025 17288 7058
rect 17208 6979 17221 7025
rect 17275 6979 17288 7025
rect 17208 6966 17288 6979
rect 17392 7025 17472 7058
rect 17392 6979 17405 7025
rect 17459 6979 17472 7025
rect 17392 6966 17472 6979
rect 21066 7337 21146 7350
rect 21066 7291 21079 7337
rect 21133 7291 21146 7337
rect 21066 7258 21146 7291
rect 21250 7337 21330 7350
rect 21250 7291 21263 7337
rect 21317 7291 21330 7337
rect 21250 7258 21330 7291
rect 21434 7337 21514 7350
rect 21434 7291 21447 7337
rect 21501 7291 21514 7337
rect 21434 7258 21514 7291
rect 21066 7025 21146 7058
rect 21066 6979 21079 7025
rect 21133 6979 21146 7025
rect 21066 6966 21146 6979
rect 21250 7025 21330 7058
rect 21250 6979 21263 7025
rect 21317 6979 21330 7025
rect 21250 6966 21330 6979
rect 21434 7025 21514 7058
rect 21434 6979 21447 7025
rect 21501 6979 21514 7025
rect 21434 6966 21514 6979
rect 25108 7337 25188 7350
rect 25108 7291 25121 7337
rect 25175 7291 25188 7337
rect 25108 7258 25188 7291
rect 25292 7337 25372 7350
rect 25292 7291 25305 7337
rect 25359 7291 25372 7337
rect 25292 7258 25372 7291
rect 25476 7337 25556 7350
rect 25476 7291 25489 7337
rect 25543 7291 25556 7337
rect 25476 7258 25556 7291
rect 25108 7025 25188 7058
rect 25108 6979 25121 7025
rect 25175 6979 25188 7025
rect 25108 6966 25188 6979
rect 25292 7025 25372 7058
rect 25292 6979 25305 7025
rect 25359 6979 25372 7025
rect 25292 6966 25372 6979
rect 25476 7025 25556 7058
rect 25476 6979 25489 7025
rect 25543 6979 25556 7025
rect 25476 6966 25556 6979
rect 886 6292 966 6305
rect 886 6246 899 6292
rect 953 6246 966 6292
rect 886 6213 966 6246
rect 1070 6292 1150 6305
rect 1070 6246 1083 6292
rect 1137 6246 1150 6292
rect 1070 6213 1150 6246
rect 1254 6292 1334 6305
rect 1254 6246 1267 6292
rect 1321 6246 1334 6292
rect 1254 6213 1334 6246
rect 886 5680 966 5713
rect 886 5634 899 5680
rect 953 5634 966 5680
rect 886 5621 966 5634
rect 1070 5680 1150 5713
rect 1070 5634 1083 5680
rect 1137 5634 1150 5680
rect 1070 5621 1150 5634
rect 1254 5680 1334 5713
rect 1254 5634 1267 5680
rect 1321 5634 1334 5680
rect 1254 5621 1334 5634
rect 2372 6292 2452 6305
rect 2372 6246 2385 6292
rect 2439 6246 2452 6292
rect 2372 6213 2452 6246
rect 2556 6292 2636 6305
rect 2556 6246 2569 6292
rect 2623 6246 2636 6292
rect 2556 6213 2636 6246
rect 2740 6292 2820 6305
rect 2740 6246 2753 6292
rect 2807 6246 2820 6292
rect 2740 6213 2820 6246
rect 2372 5680 2452 5713
rect 2372 5634 2385 5680
rect 2439 5634 2452 5680
rect 2372 5621 2452 5634
rect 2556 5680 2636 5713
rect 2556 5634 2569 5680
rect 2623 5634 2636 5680
rect 2556 5621 2636 5634
rect 2740 5680 2820 5713
rect 2740 5634 2753 5680
rect 2807 5634 2820 5680
rect 2740 5621 2820 5634
rect 4898 6292 4978 6305
rect 4898 6246 4911 6292
rect 4965 6246 4978 6292
rect 4898 6213 4978 6246
rect 5082 6292 5162 6305
rect 5082 6246 5095 6292
rect 5149 6246 5162 6292
rect 5082 6213 5162 6246
rect 5266 6292 5346 6305
rect 5266 6246 5279 6292
rect 5333 6246 5346 6292
rect 5266 6213 5346 6246
rect 4898 5680 4978 5713
rect 4898 5634 4911 5680
rect 4965 5634 4978 5680
rect 4898 5621 4978 5634
rect 5082 5680 5162 5713
rect 5082 5634 5095 5680
rect 5149 5634 5162 5680
rect 5082 5621 5162 5634
rect 5266 5680 5346 5713
rect 5266 5634 5279 5680
rect 5333 5634 5346 5680
rect 5266 5621 5346 5634
rect 6384 6292 6464 6305
rect 6384 6246 6397 6292
rect 6451 6246 6464 6292
rect 6384 6213 6464 6246
rect 6568 6292 6648 6305
rect 6568 6246 6581 6292
rect 6635 6246 6648 6292
rect 6568 6213 6648 6246
rect 6752 6292 6832 6305
rect 6752 6246 6765 6292
rect 6819 6246 6832 6292
rect 6752 6213 6832 6246
rect 6384 5680 6464 5713
rect 6384 5634 6397 5680
rect 6451 5634 6464 5680
rect 6384 5621 6464 5634
rect 6568 5680 6648 5713
rect 6568 5634 6581 5680
rect 6635 5634 6648 5680
rect 6568 5621 6648 5634
rect 6752 5680 6832 5713
rect 6752 5634 6765 5680
rect 6819 5634 6832 5680
rect 6752 5621 6832 5634
rect 8940 6292 9020 6305
rect 8940 6246 8953 6292
rect 9007 6246 9020 6292
rect 8940 6213 9020 6246
rect 9124 6292 9204 6305
rect 9124 6246 9137 6292
rect 9191 6246 9204 6292
rect 9124 6213 9204 6246
rect 9308 6292 9388 6305
rect 9308 6246 9321 6292
rect 9375 6246 9388 6292
rect 9308 6213 9388 6246
rect 8940 5680 9020 5713
rect 8940 5634 8953 5680
rect 9007 5634 9020 5680
rect 8940 5621 9020 5634
rect 9124 5680 9204 5713
rect 9124 5634 9137 5680
rect 9191 5634 9204 5680
rect 9124 5621 9204 5634
rect 9308 5680 9388 5713
rect 9308 5634 9321 5680
rect 9375 5634 9388 5680
rect 9308 5621 9388 5634
rect 10426 6292 10506 6305
rect 10426 6246 10439 6292
rect 10493 6246 10506 6292
rect 10426 6213 10506 6246
rect 10610 6292 10690 6305
rect 10610 6246 10623 6292
rect 10677 6246 10690 6292
rect 10610 6213 10690 6246
rect 10794 6292 10874 6305
rect 10794 6246 10807 6292
rect 10861 6246 10874 6292
rect 10794 6213 10874 6246
rect 10426 5680 10506 5713
rect 10426 5634 10439 5680
rect 10493 5634 10506 5680
rect 10426 5621 10506 5634
rect 10610 5680 10690 5713
rect 10610 5634 10623 5680
rect 10677 5634 10690 5680
rect 10610 5621 10690 5634
rect 10794 5680 10874 5713
rect 10794 5634 10807 5680
rect 10861 5634 10874 5680
rect 10794 5621 10874 5634
rect 12982 6292 13062 6305
rect 12982 6246 12995 6292
rect 13049 6246 13062 6292
rect 12982 6213 13062 6246
rect 13166 6292 13246 6305
rect 13166 6246 13179 6292
rect 13233 6246 13246 6292
rect 13166 6213 13246 6246
rect 13350 6292 13430 6305
rect 13350 6246 13363 6292
rect 13417 6246 13430 6292
rect 13350 6213 13430 6246
rect 12982 5680 13062 5713
rect 12982 5634 12995 5680
rect 13049 5634 13062 5680
rect 12982 5621 13062 5634
rect 13166 5680 13246 5713
rect 13166 5634 13179 5680
rect 13233 5634 13246 5680
rect 13166 5621 13246 5634
rect 13350 5680 13430 5713
rect 13350 5634 13363 5680
rect 13417 5634 13430 5680
rect 13350 5621 13430 5634
rect 14468 6292 14548 6305
rect 14468 6246 14481 6292
rect 14535 6246 14548 6292
rect 14468 6213 14548 6246
rect 14652 6292 14732 6305
rect 14652 6246 14665 6292
rect 14719 6246 14732 6292
rect 14652 6213 14732 6246
rect 14836 6292 14916 6305
rect 14836 6246 14849 6292
rect 14903 6246 14916 6292
rect 14836 6213 14916 6246
rect 14468 5680 14548 5713
rect 14468 5634 14481 5680
rect 14535 5634 14548 5680
rect 14468 5621 14548 5634
rect 14652 5680 14732 5713
rect 14652 5634 14665 5680
rect 14719 5634 14732 5680
rect 14652 5621 14732 5634
rect 14836 5680 14916 5713
rect 14836 5634 14849 5680
rect 14903 5634 14916 5680
rect 14836 5621 14916 5634
rect 17024 6292 17104 6305
rect 17024 6246 17037 6292
rect 17091 6246 17104 6292
rect 17024 6213 17104 6246
rect 17208 6292 17288 6305
rect 17208 6246 17221 6292
rect 17275 6246 17288 6292
rect 17208 6213 17288 6246
rect 17392 6292 17472 6305
rect 17392 6246 17405 6292
rect 17459 6246 17472 6292
rect 17392 6213 17472 6246
rect 17024 5680 17104 5713
rect 17024 5634 17037 5680
rect 17091 5634 17104 5680
rect 17024 5621 17104 5634
rect 17208 5680 17288 5713
rect 17208 5634 17221 5680
rect 17275 5634 17288 5680
rect 17208 5621 17288 5634
rect 17392 5680 17472 5713
rect 17392 5634 17405 5680
rect 17459 5634 17472 5680
rect 17392 5621 17472 5634
rect 18510 6292 18590 6305
rect 18510 6246 18523 6292
rect 18577 6246 18590 6292
rect 18510 6213 18590 6246
rect 18694 6292 18774 6305
rect 18694 6246 18707 6292
rect 18761 6246 18774 6292
rect 18694 6213 18774 6246
rect 18878 6292 18958 6305
rect 18878 6246 18891 6292
rect 18945 6246 18958 6292
rect 18878 6213 18958 6246
rect 18510 5680 18590 5713
rect 18510 5634 18523 5680
rect 18577 5634 18590 5680
rect 18510 5621 18590 5634
rect 18694 5680 18774 5713
rect 18694 5634 18707 5680
rect 18761 5634 18774 5680
rect 18694 5621 18774 5634
rect 18878 5680 18958 5713
rect 18878 5634 18891 5680
rect 18945 5634 18958 5680
rect 18878 5621 18958 5634
rect 21066 6292 21146 6305
rect 21066 6246 21079 6292
rect 21133 6246 21146 6292
rect 21066 6213 21146 6246
rect 21250 6292 21330 6305
rect 21250 6246 21263 6292
rect 21317 6246 21330 6292
rect 21250 6213 21330 6246
rect 21434 6292 21514 6305
rect 21434 6246 21447 6292
rect 21501 6246 21514 6292
rect 21434 6213 21514 6246
rect 21066 5680 21146 5713
rect 21066 5634 21079 5680
rect 21133 5634 21146 5680
rect 21066 5621 21146 5634
rect 21250 5680 21330 5713
rect 21250 5634 21263 5680
rect 21317 5634 21330 5680
rect 21250 5621 21330 5634
rect 21434 5680 21514 5713
rect 21434 5634 21447 5680
rect 21501 5634 21514 5680
rect 21434 5621 21514 5634
rect 22552 6292 22632 6305
rect 22552 6246 22565 6292
rect 22619 6246 22632 6292
rect 22552 6213 22632 6246
rect 22736 6292 22816 6305
rect 22736 6246 22749 6292
rect 22803 6246 22816 6292
rect 22736 6213 22816 6246
rect 22920 6292 23000 6305
rect 22920 6246 22933 6292
rect 22987 6246 23000 6292
rect 22920 6213 23000 6246
rect 22552 5680 22632 5713
rect 22552 5634 22565 5680
rect 22619 5634 22632 5680
rect 22552 5621 22632 5634
rect 22736 5680 22816 5713
rect 22736 5634 22749 5680
rect 22803 5634 22816 5680
rect 22736 5621 22816 5634
rect 22920 5680 23000 5713
rect 22920 5634 22933 5680
rect 22987 5634 23000 5680
rect 22920 5621 23000 5634
rect 25108 6292 25188 6305
rect 25108 6246 25121 6292
rect 25175 6246 25188 6292
rect 25108 6213 25188 6246
rect 25292 6292 25372 6305
rect 25292 6246 25305 6292
rect 25359 6246 25372 6292
rect 25292 6213 25372 6246
rect 25476 6292 25556 6305
rect 25476 6246 25489 6292
rect 25543 6246 25556 6292
rect 25476 6213 25556 6246
rect 25108 5680 25188 5713
rect 25108 5634 25121 5680
rect 25175 5634 25188 5680
rect 25108 5621 25188 5634
rect 25292 5680 25372 5713
rect 25292 5634 25305 5680
rect 25359 5634 25372 5680
rect 25292 5621 25372 5634
rect 25476 5680 25556 5713
rect 25476 5634 25489 5680
rect 25543 5634 25556 5680
rect 25476 5621 25556 5634
rect 26594 6292 26674 6305
rect 26594 6246 26607 6292
rect 26661 6246 26674 6292
rect 26594 6213 26674 6246
rect 26778 6292 26858 6305
rect 26778 6246 26791 6292
rect 26845 6246 26858 6292
rect 26778 6213 26858 6246
rect 26962 6292 27042 6305
rect 26962 6246 26975 6292
rect 27029 6246 27042 6292
rect 26962 6213 27042 6246
rect 26594 5680 26674 5713
rect 26594 5634 26607 5680
rect 26661 5634 26674 5680
rect 26594 5621 26674 5634
rect 26778 5680 26858 5713
rect 26778 5634 26791 5680
rect 26845 5634 26858 5680
rect 26778 5621 26858 5634
rect 26962 5680 27042 5713
rect 26962 5634 26975 5680
rect 27029 5634 27042 5680
rect 26962 5621 27042 5634
rect 886 5132 966 5145
rect 886 5086 899 5132
rect 953 5086 966 5132
rect 886 5053 966 5086
rect 1070 5132 1150 5145
rect 1070 5086 1083 5132
rect 1137 5086 1150 5132
rect 1070 5053 1150 5086
rect 1254 5132 1334 5145
rect 1254 5086 1267 5132
rect 1321 5086 1334 5132
rect 1254 5053 1334 5086
rect 886 4820 966 4853
rect 886 4774 899 4820
rect 953 4774 966 4820
rect 886 4761 966 4774
rect 1070 4820 1150 4853
rect 1070 4774 1083 4820
rect 1137 4774 1150 4820
rect 1070 4761 1150 4774
rect 1254 4820 1334 4853
rect 1254 4774 1267 4820
rect 1321 4774 1334 4820
rect 1254 4761 1334 4774
rect 2372 5132 2452 5145
rect 2372 5086 2385 5132
rect 2439 5086 2452 5132
rect 2372 5053 2452 5086
rect 2556 5132 2636 5145
rect 2556 5086 2569 5132
rect 2623 5086 2636 5132
rect 2556 5053 2636 5086
rect 2740 5132 2820 5145
rect 2740 5086 2753 5132
rect 2807 5086 2820 5132
rect 2740 5053 2820 5086
rect 2372 4820 2452 4853
rect 2372 4774 2385 4820
rect 2439 4774 2452 4820
rect 2372 4761 2452 4774
rect 2556 4820 2636 4853
rect 2556 4774 2569 4820
rect 2623 4774 2636 4820
rect 2556 4761 2636 4774
rect 2740 4820 2820 4853
rect 2740 4774 2753 4820
rect 2807 4774 2820 4820
rect 2740 4761 2820 4774
rect 4898 5132 4978 5145
rect 4898 5086 4911 5132
rect 4965 5086 4978 5132
rect 4898 5053 4978 5086
rect 5082 5132 5162 5145
rect 5082 5086 5095 5132
rect 5149 5086 5162 5132
rect 5082 5053 5162 5086
rect 5266 5132 5346 5145
rect 5266 5086 5279 5132
rect 5333 5086 5346 5132
rect 5266 5053 5346 5086
rect 4898 4820 4978 4853
rect 4898 4774 4911 4820
rect 4965 4774 4978 4820
rect 4898 4761 4978 4774
rect 5082 4820 5162 4853
rect 5082 4774 5095 4820
rect 5149 4774 5162 4820
rect 5082 4761 5162 4774
rect 5266 4820 5346 4853
rect 5266 4774 5279 4820
rect 5333 4774 5346 4820
rect 5266 4761 5346 4774
rect 6384 5132 6464 5145
rect 6384 5086 6397 5132
rect 6451 5086 6464 5132
rect 6384 5053 6464 5086
rect 6568 5132 6648 5145
rect 6568 5086 6581 5132
rect 6635 5086 6648 5132
rect 6568 5053 6648 5086
rect 6752 5132 6832 5145
rect 6752 5086 6765 5132
rect 6819 5086 6832 5132
rect 6752 5053 6832 5086
rect 6384 4820 6464 4853
rect 6384 4774 6397 4820
rect 6451 4774 6464 4820
rect 6384 4761 6464 4774
rect 6568 4820 6648 4853
rect 6568 4774 6581 4820
rect 6635 4774 6648 4820
rect 6568 4761 6648 4774
rect 6752 4820 6832 4853
rect 6752 4774 6765 4820
rect 6819 4774 6832 4820
rect 6752 4761 6832 4774
rect 8940 5132 9020 5145
rect 8940 5086 8953 5132
rect 9007 5086 9020 5132
rect 8940 5053 9020 5086
rect 9124 5132 9204 5145
rect 9124 5086 9137 5132
rect 9191 5086 9204 5132
rect 9124 5053 9204 5086
rect 9308 5132 9388 5145
rect 9308 5086 9321 5132
rect 9375 5086 9388 5132
rect 9308 5053 9388 5086
rect 8940 4820 9020 4853
rect 8940 4774 8953 4820
rect 9007 4774 9020 4820
rect 8940 4761 9020 4774
rect 9124 4820 9204 4853
rect 9124 4774 9137 4820
rect 9191 4774 9204 4820
rect 9124 4761 9204 4774
rect 9308 4820 9388 4853
rect 9308 4774 9321 4820
rect 9375 4774 9388 4820
rect 9308 4761 9388 4774
rect 10426 5132 10506 5145
rect 10426 5086 10439 5132
rect 10493 5086 10506 5132
rect 10426 5053 10506 5086
rect 10610 5132 10690 5145
rect 10610 5086 10623 5132
rect 10677 5086 10690 5132
rect 10610 5053 10690 5086
rect 10794 5132 10874 5145
rect 10794 5086 10807 5132
rect 10861 5086 10874 5132
rect 10794 5053 10874 5086
rect 10426 4820 10506 4853
rect 10426 4774 10439 4820
rect 10493 4774 10506 4820
rect 10426 4761 10506 4774
rect 10610 4820 10690 4853
rect 10610 4774 10623 4820
rect 10677 4774 10690 4820
rect 10610 4761 10690 4774
rect 10794 4820 10874 4853
rect 10794 4774 10807 4820
rect 10861 4774 10874 4820
rect 10794 4761 10874 4774
rect 12982 5132 13062 5145
rect 12982 5086 12995 5132
rect 13049 5086 13062 5132
rect 12982 5053 13062 5086
rect 13166 5132 13246 5145
rect 13166 5086 13179 5132
rect 13233 5086 13246 5132
rect 13166 5053 13246 5086
rect 13350 5132 13430 5145
rect 13350 5086 13363 5132
rect 13417 5086 13430 5132
rect 13350 5053 13430 5086
rect 12982 4820 13062 4853
rect 12982 4774 12995 4820
rect 13049 4774 13062 4820
rect 12982 4761 13062 4774
rect 13166 4820 13246 4853
rect 13166 4774 13179 4820
rect 13233 4774 13246 4820
rect 13166 4761 13246 4774
rect 13350 4820 13430 4853
rect 13350 4774 13363 4820
rect 13417 4774 13430 4820
rect 13350 4761 13430 4774
rect 14468 5132 14548 5145
rect 14468 5086 14481 5132
rect 14535 5086 14548 5132
rect 14468 5053 14548 5086
rect 14652 5132 14732 5145
rect 14652 5086 14665 5132
rect 14719 5086 14732 5132
rect 14652 5053 14732 5086
rect 14836 5132 14916 5145
rect 14836 5086 14849 5132
rect 14903 5086 14916 5132
rect 14836 5053 14916 5086
rect 14468 4820 14548 4853
rect 14468 4774 14481 4820
rect 14535 4774 14548 4820
rect 14468 4761 14548 4774
rect 14652 4820 14732 4853
rect 14652 4774 14665 4820
rect 14719 4774 14732 4820
rect 14652 4761 14732 4774
rect 14836 4820 14916 4853
rect 14836 4774 14849 4820
rect 14903 4774 14916 4820
rect 14836 4761 14916 4774
rect 17024 5132 17104 5145
rect 17024 5086 17037 5132
rect 17091 5086 17104 5132
rect 17024 5053 17104 5086
rect 17208 5132 17288 5145
rect 17208 5086 17221 5132
rect 17275 5086 17288 5132
rect 17208 5053 17288 5086
rect 17392 5132 17472 5145
rect 17392 5086 17405 5132
rect 17459 5086 17472 5132
rect 17392 5053 17472 5086
rect 17024 4820 17104 4853
rect 17024 4774 17037 4820
rect 17091 4774 17104 4820
rect 17024 4761 17104 4774
rect 17208 4820 17288 4853
rect 17208 4774 17221 4820
rect 17275 4774 17288 4820
rect 17208 4761 17288 4774
rect 17392 4820 17472 4853
rect 17392 4774 17405 4820
rect 17459 4774 17472 4820
rect 17392 4761 17472 4774
rect 18510 5132 18590 5145
rect 18510 5086 18523 5132
rect 18577 5086 18590 5132
rect 18510 5053 18590 5086
rect 18694 5132 18774 5145
rect 18694 5086 18707 5132
rect 18761 5086 18774 5132
rect 18694 5053 18774 5086
rect 18878 5132 18958 5145
rect 18878 5086 18891 5132
rect 18945 5086 18958 5132
rect 18878 5053 18958 5086
rect 18510 4820 18590 4853
rect 18510 4774 18523 4820
rect 18577 4774 18590 4820
rect 18510 4761 18590 4774
rect 18694 4820 18774 4853
rect 18694 4774 18707 4820
rect 18761 4774 18774 4820
rect 18694 4761 18774 4774
rect 18878 4820 18958 4853
rect 18878 4774 18891 4820
rect 18945 4774 18958 4820
rect 18878 4761 18958 4774
rect 21066 5132 21146 5145
rect 21066 5086 21079 5132
rect 21133 5086 21146 5132
rect 21066 5053 21146 5086
rect 21250 5132 21330 5145
rect 21250 5086 21263 5132
rect 21317 5086 21330 5132
rect 21250 5053 21330 5086
rect 21434 5132 21514 5145
rect 21434 5086 21447 5132
rect 21501 5086 21514 5132
rect 21434 5053 21514 5086
rect 21066 4820 21146 4853
rect 21066 4774 21079 4820
rect 21133 4774 21146 4820
rect 21066 4761 21146 4774
rect 21250 4820 21330 4853
rect 21250 4774 21263 4820
rect 21317 4774 21330 4820
rect 21250 4761 21330 4774
rect 21434 4820 21514 4853
rect 21434 4774 21447 4820
rect 21501 4774 21514 4820
rect 21434 4761 21514 4774
rect 22552 5132 22632 5145
rect 22552 5086 22565 5132
rect 22619 5086 22632 5132
rect 22552 5053 22632 5086
rect 22736 5132 22816 5145
rect 22736 5086 22749 5132
rect 22803 5086 22816 5132
rect 22736 5053 22816 5086
rect 22920 5132 23000 5145
rect 22920 5086 22933 5132
rect 22987 5086 23000 5132
rect 22920 5053 23000 5086
rect 22552 4820 22632 4853
rect 22552 4774 22565 4820
rect 22619 4774 22632 4820
rect 22552 4761 22632 4774
rect 22736 4820 22816 4853
rect 22736 4774 22749 4820
rect 22803 4774 22816 4820
rect 22736 4761 22816 4774
rect 22920 4820 23000 4853
rect 22920 4774 22933 4820
rect 22987 4774 23000 4820
rect 22920 4761 23000 4774
rect 25108 5132 25188 5145
rect 25108 5086 25121 5132
rect 25175 5086 25188 5132
rect 25108 5053 25188 5086
rect 25292 5132 25372 5145
rect 25292 5086 25305 5132
rect 25359 5086 25372 5132
rect 25292 5053 25372 5086
rect 25476 5132 25556 5145
rect 25476 5086 25489 5132
rect 25543 5086 25556 5132
rect 25476 5053 25556 5086
rect 25108 4820 25188 4853
rect 25108 4774 25121 4820
rect 25175 4774 25188 4820
rect 25108 4761 25188 4774
rect 25292 4820 25372 4853
rect 25292 4774 25305 4820
rect 25359 4774 25372 4820
rect 25292 4761 25372 4774
rect 25476 4820 25556 4853
rect 25476 4774 25489 4820
rect 25543 4774 25556 4820
rect 25476 4761 25556 4774
rect 26594 5132 26674 5145
rect 26594 5086 26607 5132
rect 26661 5086 26674 5132
rect 26594 5053 26674 5086
rect 26778 5132 26858 5145
rect 26778 5086 26791 5132
rect 26845 5086 26858 5132
rect 26778 5053 26858 5086
rect 26962 5132 27042 5145
rect 26962 5086 26975 5132
rect 27029 5086 27042 5132
rect 26962 5053 27042 5086
rect 26594 4820 26674 4853
rect 26594 4774 26607 4820
rect 26661 4774 26674 4820
rect 26594 4761 26674 4774
rect 26778 4820 26858 4853
rect 26778 4774 26791 4820
rect 26845 4774 26858 4820
rect 26778 4761 26858 4774
rect 26962 4820 27042 4853
rect 26962 4774 26975 4820
rect 27029 4774 27042 4820
rect 26962 4761 27042 4774
rect 886 4087 966 4100
rect 886 4041 899 4087
rect 953 4041 966 4087
rect 886 4008 966 4041
rect 1070 4087 1150 4100
rect 1070 4041 1083 4087
rect 1137 4041 1150 4087
rect 1070 4008 1150 4041
rect 1254 4087 1334 4100
rect 1254 4041 1267 4087
rect 1321 4041 1334 4087
rect 1254 4008 1334 4041
rect 886 3475 966 3508
rect 886 3429 899 3475
rect 953 3429 966 3475
rect 886 3416 966 3429
rect 1070 3475 1150 3508
rect 1070 3429 1083 3475
rect 1137 3429 1150 3475
rect 1070 3416 1150 3429
rect 1254 3475 1334 3508
rect 1254 3429 1267 3475
rect 1321 3429 1334 3475
rect 1254 3416 1334 3429
rect 2372 4088 2452 4101
rect 2372 4042 2385 4088
rect 2439 4042 2452 4088
rect 2372 4009 2452 4042
rect 2556 4088 2636 4101
rect 2556 4042 2569 4088
rect 2623 4042 2636 4088
rect 2556 4009 2636 4042
rect 2740 4088 2820 4101
rect 2740 4042 2753 4088
rect 2807 4042 2820 4088
rect 2740 4009 2820 4042
rect 2372 3476 2452 3509
rect 2372 3430 2385 3476
rect 2439 3430 2452 3476
rect 2372 3417 2452 3430
rect 2556 3476 2636 3509
rect 2556 3430 2569 3476
rect 2623 3430 2636 3476
rect 2556 3417 2636 3430
rect 2740 3476 2820 3509
rect 2740 3430 2753 3476
rect 2807 3430 2820 3476
rect 2740 3417 2820 3430
rect 4898 4087 4978 4100
rect 4898 4041 4911 4087
rect 4965 4041 4978 4087
rect 4898 4008 4978 4041
rect 5082 4087 5162 4100
rect 5082 4041 5095 4087
rect 5149 4041 5162 4087
rect 5082 4008 5162 4041
rect 5266 4087 5346 4100
rect 5266 4041 5279 4087
rect 5333 4041 5346 4087
rect 5266 4008 5346 4041
rect 4898 3475 4978 3508
rect 4898 3429 4911 3475
rect 4965 3429 4978 3475
rect 4898 3416 4978 3429
rect 5082 3475 5162 3508
rect 5082 3429 5095 3475
rect 5149 3429 5162 3475
rect 5082 3416 5162 3429
rect 5266 3475 5346 3508
rect 5266 3429 5279 3475
rect 5333 3429 5346 3475
rect 5266 3416 5346 3429
rect 6384 4088 6464 4101
rect 6384 4042 6397 4088
rect 6451 4042 6464 4088
rect 6384 4009 6464 4042
rect 6568 4088 6648 4101
rect 6568 4042 6581 4088
rect 6635 4042 6648 4088
rect 6568 4009 6648 4042
rect 6752 4088 6832 4101
rect 6752 4042 6765 4088
rect 6819 4042 6832 4088
rect 6752 4009 6832 4042
rect 6384 3476 6464 3509
rect 6384 3430 6397 3476
rect 6451 3430 6464 3476
rect 6384 3417 6464 3430
rect 6568 3476 6648 3509
rect 6568 3430 6581 3476
rect 6635 3430 6648 3476
rect 6568 3417 6648 3430
rect 6752 3476 6832 3509
rect 6752 3430 6765 3476
rect 6819 3430 6832 3476
rect 6752 3417 6832 3430
rect 8940 4087 9020 4100
rect 8940 4041 8953 4087
rect 9007 4041 9020 4087
rect 8940 4008 9020 4041
rect 9124 4087 9204 4100
rect 9124 4041 9137 4087
rect 9191 4041 9204 4087
rect 9124 4008 9204 4041
rect 9308 4087 9388 4100
rect 9308 4041 9321 4087
rect 9375 4041 9388 4087
rect 9308 4008 9388 4041
rect 8940 3475 9020 3508
rect 8940 3429 8953 3475
rect 9007 3429 9020 3475
rect 8940 3416 9020 3429
rect 9124 3475 9204 3508
rect 9124 3429 9137 3475
rect 9191 3429 9204 3475
rect 9124 3416 9204 3429
rect 9308 3475 9388 3508
rect 9308 3429 9321 3475
rect 9375 3429 9388 3475
rect 9308 3416 9388 3429
rect 10426 4088 10506 4101
rect 10426 4042 10439 4088
rect 10493 4042 10506 4088
rect 10426 4009 10506 4042
rect 10610 4088 10690 4101
rect 10610 4042 10623 4088
rect 10677 4042 10690 4088
rect 10610 4009 10690 4042
rect 10794 4088 10874 4101
rect 10794 4042 10807 4088
rect 10861 4042 10874 4088
rect 10794 4009 10874 4042
rect 10426 3476 10506 3509
rect 10426 3430 10439 3476
rect 10493 3430 10506 3476
rect 10426 3417 10506 3430
rect 10610 3476 10690 3509
rect 10610 3430 10623 3476
rect 10677 3430 10690 3476
rect 10610 3417 10690 3430
rect 10794 3476 10874 3509
rect 10794 3430 10807 3476
rect 10861 3430 10874 3476
rect 10794 3417 10874 3430
rect 12982 4087 13062 4100
rect 12982 4041 12995 4087
rect 13049 4041 13062 4087
rect 12982 4008 13062 4041
rect 13166 4087 13246 4100
rect 13166 4041 13179 4087
rect 13233 4041 13246 4087
rect 13166 4008 13246 4041
rect 13350 4087 13430 4100
rect 13350 4041 13363 4087
rect 13417 4041 13430 4087
rect 13350 4008 13430 4041
rect 12982 3475 13062 3508
rect 12982 3429 12995 3475
rect 13049 3429 13062 3475
rect 12982 3416 13062 3429
rect 13166 3475 13246 3508
rect 13166 3429 13179 3475
rect 13233 3429 13246 3475
rect 13166 3416 13246 3429
rect 13350 3475 13430 3508
rect 13350 3429 13363 3475
rect 13417 3429 13430 3475
rect 13350 3416 13430 3429
rect 14468 4088 14548 4101
rect 14468 4042 14481 4088
rect 14535 4042 14548 4088
rect 14468 4009 14548 4042
rect 14652 4088 14732 4101
rect 14652 4042 14665 4088
rect 14719 4042 14732 4088
rect 14652 4009 14732 4042
rect 14836 4088 14916 4101
rect 14836 4042 14849 4088
rect 14903 4042 14916 4088
rect 14836 4009 14916 4042
rect 14468 3476 14548 3509
rect 14468 3430 14481 3476
rect 14535 3430 14548 3476
rect 14468 3417 14548 3430
rect 14652 3476 14732 3509
rect 14652 3430 14665 3476
rect 14719 3430 14732 3476
rect 14652 3417 14732 3430
rect 14836 3476 14916 3509
rect 14836 3430 14849 3476
rect 14903 3430 14916 3476
rect 14836 3417 14916 3430
rect 17024 4087 17104 4100
rect 17024 4041 17037 4087
rect 17091 4041 17104 4087
rect 17024 4008 17104 4041
rect 17208 4087 17288 4100
rect 17208 4041 17221 4087
rect 17275 4041 17288 4087
rect 17208 4008 17288 4041
rect 17392 4087 17472 4100
rect 17392 4041 17405 4087
rect 17459 4041 17472 4087
rect 17392 4008 17472 4041
rect 17024 3475 17104 3508
rect 17024 3429 17037 3475
rect 17091 3429 17104 3475
rect 17024 3416 17104 3429
rect 17208 3475 17288 3508
rect 17208 3429 17221 3475
rect 17275 3429 17288 3475
rect 17208 3416 17288 3429
rect 17392 3475 17472 3508
rect 17392 3429 17405 3475
rect 17459 3429 17472 3475
rect 17392 3416 17472 3429
rect 18510 4088 18590 4101
rect 18510 4042 18523 4088
rect 18577 4042 18590 4088
rect 18510 4009 18590 4042
rect 18694 4088 18774 4101
rect 18694 4042 18707 4088
rect 18761 4042 18774 4088
rect 18694 4009 18774 4042
rect 18878 4088 18958 4101
rect 18878 4042 18891 4088
rect 18945 4042 18958 4088
rect 18878 4009 18958 4042
rect 18510 3476 18590 3509
rect 18510 3430 18523 3476
rect 18577 3430 18590 3476
rect 18510 3417 18590 3430
rect 18694 3476 18774 3509
rect 18694 3430 18707 3476
rect 18761 3430 18774 3476
rect 18694 3417 18774 3430
rect 18878 3476 18958 3509
rect 18878 3430 18891 3476
rect 18945 3430 18958 3476
rect 18878 3417 18958 3430
rect 21066 4087 21146 4100
rect 21066 4041 21079 4087
rect 21133 4041 21146 4087
rect 21066 4008 21146 4041
rect 21250 4087 21330 4100
rect 21250 4041 21263 4087
rect 21317 4041 21330 4087
rect 21250 4008 21330 4041
rect 21434 4087 21514 4100
rect 21434 4041 21447 4087
rect 21501 4041 21514 4087
rect 21434 4008 21514 4041
rect 21066 3475 21146 3508
rect 21066 3429 21079 3475
rect 21133 3429 21146 3475
rect 21066 3416 21146 3429
rect 21250 3475 21330 3508
rect 21250 3429 21263 3475
rect 21317 3429 21330 3475
rect 21250 3416 21330 3429
rect 21434 3475 21514 3508
rect 21434 3429 21447 3475
rect 21501 3429 21514 3475
rect 21434 3416 21514 3429
rect 22552 4088 22632 4101
rect 22552 4042 22565 4088
rect 22619 4042 22632 4088
rect 22552 4009 22632 4042
rect 22736 4088 22816 4101
rect 22736 4042 22749 4088
rect 22803 4042 22816 4088
rect 22736 4009 22816 4042
rect 22920 4088 23000 4101
rect 22920 4042 22933 4088
rect 22987 4042 23000 4088
rect 22920 4009 23000 4042
rect 22552 3476 22632 3509
rect 22552 3430 22565 3476
rect 22619 3430 22632 3476
rect 22552 3417 22632 3430
rect 22736 3476 22816 3509
rect 22736 3430 22749 3476
rect 22803 3430 22816 3476
rect 22736 3417 22816 3430
rect 22920 3476 23000 3509
rect 22920 3430 22933 3476
rect 22987 3430 23000 3476
rect 22920 3417 23000 3430
rect 25108 4087 25188 4100
rect 25108 4041 25121 4087
rect 25175 4041 25188 4087
rect 25108 4008 25188 4041
rect 25292 4087 25372 4100
rect 25292 4041 25305 4087
rect 25359 4041 25372 4087
rect 25292 4008 25372 4041
rect 25476 4087 25556 4100
rect 25476 4041 25489 4087
rect 25543 4041 25556 4087
rect 25476 4008 25556 4041
rect 25108 3475 25188 3508
rect 25108 3429 25121 3475
rect 25175 3429 25188 3475
rect 25108 3416 25188 3429
rect 25292 3475 25372 3508
rect 25292 3429 25305 3475
rect 25359 3429 25372 3475
rect 25292 3416 25372 3429
rect 25476 3475 25556 3508
rect 25476 3429 25489 3475
rect 25543 3429 25556 3475
rect 25476 3416 25556 3429
rect 26594 4088 26674 4101
rect 26594 4042 26607 4088
rect 26661 4042 26674 4088
rect 26594 4009 26674 4042
rect 26778 4088 26858 4101
rect 26778 4042 26791 4088
rect 26845 4042 26858 4088
rect 26778 4009 26858 4042
rect 26962 4088 27042 4101
rect 26962 4042 26975 4088
rect 27029 4042 27042 4088
rect 26962 4009 27042 4042
rect 26594 3476 26674 3509
rect 26594 3430 26607 3476
rect 26661 3430 26674 3476
rect 26594 3417 26674 3430
rect 26778 3476 26858 3509
rect 26778 3430 26791 3476
rect 26845 3430 26858 3476
rect 26778 3417 26858 3430
rect 26962 3476 27042 3509
rect 26962 3430 26975 3476
rect 27029 3430 27042 3476
rect 26962 3417 27042 3430
rect 886 2927 966 2940
rect 886 2881 899 2927
rect 953 2881 966 2927
rect 886 2848 966 2881
rect 1070 2927 1150 2940
rect 1070 2881 1083 2927
rect 1137 2881 1150 2927
rect 1070 2848 1150 2881
rect 1254 2927 1334 2940
rect 1254 2881 1267 2927
rect 1321 2881 1334 2927
rect 1254 2848 1334 2881
rect 886 2615 966 2648
rect 886 2569 899 2615
rect 953 2569 966 2615
rect 886 2556 966 2569
rect 1070 2615 1150 2648
rect 1070 2569 1083 2615
rect 1137 2569 1150 2615
rect 1070 2556 1150 2569
rect 1254 2615 1334 2648
rect 1254 2569 1267 2615
rect 1321 2569 1334 2615
rect 1254 2556 1334 2569
rect 2372 2928 2452 2941
rect 2372 2882 2385 2928
rect 2439 2882 2452 2928
rect 2372 2849 2452 2882
rect 2556 2928 2636 2941
rect 2556 2882 2569 2928
rect 2623 2882 2636 2928
rect 2556 2849 2636 2882
rect 2740 2928 2820 2941
rect 2740 2882 2753 2928
rect 2807 2882 2820 2928
rect 2740 2849 2820 2882
rect 2372 2616 2452 2649
rect 2372 2570 2385 2616
rect 2439 2570 2452 2616
rect 2372 2557 2452 2570
rect 2556 2616 2636 2649
rect 2556 2570 2569 2616
rect 2623 2570 2636 2616
rect 2556 2557 2636 2570
rect 2740 2616 2820 2649
rect 2740 2570 2753 2616
rect 2807 2570 2820 2616
rect 2740 2557 2820 2570
rect 4898 2927 4978 2940
rect 4898 2881 4911 2927
rect 4965 2881 4978 2927
rect 4898 2848 4978 2881
rect 5082 2927 5162 2940
rect 5082 2881 5095 2927
rect 5149 2881 5162 2927
rect 5082 2848 5162 2881
rect 5266 2927 5346 2940
rect 5266 2881 5279 2927
rect 5333 2881 5346 2927
rect 5266 2848 5346 2881
rect 4898 2615 4978 2648
rect 4898 2569 4911 2615
rect 4965 2569 4978 2615
rect 4898 2556 4978 2569
rect 5082 2615 5162 2648
rect 5082 2569 5095 2615
rect 5149 2569 5162 2615
rect 5082 2556 5162 2569
rect 5266 2615 5346 2648
rect 5266 2569 5279 2615
rect 5333 2569 5346 2615
rect 5266 2556 5346 2569
rect 6384 2928 6464 2941
rect 6384 2882 6397 2928
rect 6451 2882 6464 2928
rect 6384 2849 6464 2882
rect 6568 2928 6648 2941
rect 6568 2882 6581 2928
rect 6635 2882 6648 2928
rect 6568 2849 6648 2882
rect 6752 2928 6832 2941
rect 6752 2882 6765 2928
rect 6819 2882 6832 2928
rect 6752 2849 6832 2882
rect 6384 2616 6464 2649
rect 6384 2570 6397 2616
rect 6451 2570 6464 2616
rect 6384 2557 6464 2570
rect 6568 2616 6648 2649
rect 6568 2570 6581 2616
rect 6635 2570 6648 2616
rect 6568 2557 6648 2570
rect 6752 2616 6832 2649
rect 6752 2570 6765 2616
rect 6819 2570 6832 2616
rect 6752 2557 6832 2570
rect 8940 2927 9020 2940
rect 8940 2881 8953 2927
rect 9007 2881 9020 2927
rect 8940 2848 9020 2881
rect 9124 2927 9204 2940
rect 9124 2881 9137 2927
rect 9191 2881 9204 2927
rect 9124 2848 9204 2881
rect 9308 2927 9388 2940
rect 9308 2881 9321 2927
rect 9375 2881 9388 2927
rect 9308 2848 9388 2881
rect 8940 2615 9020 2648
rect 8940 2569 8953 2615
rect 9007 2569 9020 2615
rect 8940 2556 9020 2569
rect 9124 2615 9204 2648
rect 9124 2569 9137 2615
rect 9191 2569 9204 2615
rect 9124 2556 9204 2569
rect 9308 2615 9388 2648
rect 9308 2569 9321 2615
rect 9375 2569 9388 2615
rect 9308 2556 9388 2569
rect 10426 2928 10506 2941
rect 10426 2882 10439 2928
rect 10493 2882 10506 2928
rect 10426 2849 10506 2882
rect 10610 2928 10690 2941
rect 10610 2882 10623 2928
rect 10677 2882 10690 2928
rect 10610 2849 10690 2882
rect 10794 2928 10874 2941
rect 10794 2882 10807 2928
rect 10861 2882 10874 2928
rect 10794 2849 10874 2882
rect 10426 2616 10506 2649
rect 10426 2570 10439 2616
rect 10493 2570 10506 2616
rect 10426 2557 10506 2570
rect 10610 2616 10690 2649
rect 10610 2570 10623 2616
rect 10677 2570 10690 2616
rect 10610 2557 10690 2570
rect 10794 2616 10874 2649
rect 10794 2570 10807 2616
rect 10861 2570 10874 2616
rect 10794 2557 10874 2570
rect 12982 2927 13062 2940
rect 12982 2881 12995 2927
rect 13049 2881 13062 2927
rect 12982 2848 13062 2881
rect 13166 2927 13246 2940
rect 13166 2881 13179 2927
rect 13233 2881 13246 2927
rect 13166 2848 13246 2881
rect 13350 2927 13430 2940
rect 13350 2881 13363 2927
rect 13417 2881 13430 2927
rect 13350 2848 13430 2881
rect 12982 2615 13062 2648
rect 12982 2569 12995 2615
rect 13049 2569 13062 2615
rect 12982 2556 13062 2569
rect 13166 2615 13246 2648
rect 13166 2569 13179 2615
rect 13233 2569 13246 2615
rect 13166 2556 13246 2569
rect 13350 2615 13430 2648
rect 13350 2569 13363 2615
rect 13417 2569 13430 2615
rect 13350 2556 13430 2569
rect 14468 2928 14548 2941
rect 14468 2882 14481 2928
rect 14535 2882 14548 2928
rect 14468 2849 14548 2882
rect 14652 2928 14732 2941
rect 14652 2882 14665 2928
rect 14719 2882 14732 2928
rect 14652 2849 14732 2882
rect 14836 2928 14916 2941
rect 14836 2882 14849 2928
rect 14903 2882 14916 2928
rect 14836 2849 14916 2882
rect 14468 2616 14548 2649
rect 14468 2570 14481 2616
rect 14535 2570 14548 2616
rect 14468 2557 14548 2570
rect 14652 2616 14732 2649
rect 14652 2570 14665 2616
rect 14719 2570 14732 2616
rect 14652 2557 14732 2570
rect 14836 2616 14916 2649
rect 14836 2570 14849 2616
rect 14903 2570 14916 2616
rect 14836 2557 14916 2570
rect 17024 2927 17104 2940
rect 17024 2881 17037 2927
rect 17091 2881 17104 2927
rect 17024 2848 17104 2881
rect 17208 2927 17288 2940
rect 17208 2881 17221 2927
rect 17275 2881 17288 2927
rect 17208 2848 17288 2881
rect 17392 2927 17472 2940
rect 17392 2881 17405 2927
rect 17459 2881 17472 2927
rect 17392 2848 17472 2881
rect 17024 2615 17104 2648
rect 17024 2569 17037 2615
rect 17091 2569 17104 2615
rect 17024 2556 17104 2569
rect 17208 2615 17288 2648
rect 17208 2569 17221 2615
rect 17275 2569 17288 2615
rect 17208 2556 17288 2569
rect 17392 2615 17472 2648
rect 17392 2569 17405 2615
rect 17459 2569 17472 2615
rect 17392 2556 17472 2569
rect 18510 2928 18590 2941
rect 18510 2882 18523 2928
rect 18577 2882 18590 2928
rect 18510 2849 18590 2882
rect 18694 2928 18774 2941
rect 18694 2882 18707 2928
rect 18761 2882 18774 2928
rect 18694 2849 18774 2882
rect 18878 2928 18958 2941
rect 18878 2882 18891 2928
rect 18945 2882 18958 2928
rect 18878 2849 18958 2882
rect 18510 2616 18590 2649
rect 18510 2570 18523 2616
rect 18577 2570 18590 2616
rect 18510 2557 18590 2570
rect 18694 2616 18774 2649
rect 18694 2570 18707 2616
rect 18761 2570 18774 2616
rect 18694 2557 18774 2570
rect 18878 2616 18958 2649
rect 18878 2570 18891 2616
rect 18945 2570 18958 2616
rect 18878 2557 18958 2570
rect 21066 2927 21146 2940
rect 21066 2881 21079 2927
rect 21133 2881 21146 2927
rect 21066 2848 21146 2881
rect 21250 2927 21330 2940
rect 21250 2881 21263 2927
rect 21317 2881 21330 2927
rect 21250 2848 21330 2881
rect 21434 2927 21514 2940
rect 21434 2881 21447 2927
rect 21501 2881 21514 2927
rect 21434 2848 21514 2881
rect 21066 2615 21146 2648
rect 21066 2569 21079 2615
rect 21133 2569 21146 2615
rect 21066 2556 21146 2569
rect 21250 2615 21330 2648
rect 21250 2569 21263 2615
rect 21317 2569 21330 2615
rect 21250 2556 21330 2569
rect 21434 2615 21514 2648
rect 21434 2569 21447 2615
rect 21501 2569 21514 2615
rect 21434 2556 21514 2569
rect 22552 2928 22632 2941
rect 22552 2882 22565 2928
rect 22619 2882 22632 2928
rect 22552 2849 22632 2882
rect 22736 2928 22816 2941
rect 22736 2882 22749 2928
rect 22803 2882 22816 2928
rect 22736 2849 22816 2882
rect 22920 2928 23000 2941
rect 22920 2882 22933 2928
rect 22987 2882 23000 2928
rect 22920 2849 23000 2882
rect 22552 2616 22632 2649
rect 22552 2570 22565 2616
rect 22619 2570 22632 2616
rect 22552 2557 22632 2570
rect 22736 2616 22816 2649
rect 22736 2570 22749 2616
rect 22803 2570 22816 2616
rect 22736 2557 22816 2570
rect 22920 2616 23000 2649
rect 22920 2570 22933 2616
rect 22987 2570 23000 2616
rect 22920 2557 23000 2570
rect 25108 2927 25188 2940
rect 25108 2881 25121 2927
rect 25175 2881 25188 2927
rect 25108 2848 25188 2881
rect 25292 2927 25372 2940
rect 25292 2881 25305 2927
rect 25359 2881 25372 2927
rect 25292 2848 25372 2881
rect 25476 2927 25556 2940
rect 25476 2881 25489 2927
rect 25543 2881 25556 2927
rect 25476 2848 25556 2881
rect 25108 2615 25188 2648
rect 25108 2569 25121 2615
rect 25175 2569 25188 2615
rect 25108 2556 25188 2569
rect 25292 2615 25372 2648
rect 25292 2569 25305 2615
rect 25359 2569 25372 2615
rect 25292 2556 25372 2569
rect 25476 2615 25556 2648
rect 25476 2569 25489 2615
rect 25543 2569 25556 2615
rect 25476 2556 25556 2569
rect 26594 2928 26674 2941
rect 26594 2882 26607 2928
rect 26661 2882 26674 2928
rect 26594 2849 26674 2882
rect 26778 2928 26858 2941
rect 26778 2882 26791 2928
rect 26845 2882 26858 2928
rect 26778 2849 26858 2882
rect 26962 2928 27042 2941
rect 26962 2882 26975 2928
rect 27029 2882 27042 2928
rect 26962 2849 27042 2882
rect 26594 2616 26674 2649
rect 26594 2570 26607 2616
rect 26661 2570 26674 2616
rect 26594 2557 26674 2570
rect 26778 2616 26858 2649
rect 26778 2570 26791 2616
rect 26845 2570 26858 2616
rect 26778 2557 26858 2570
rect 26962 2616 27042 2649
rect 26962 2570 26975 2616
rect 27029 2570 27042 2616
rect 26962 2557 27042 2570
rect 886 1882 966 1895
rect 886 1836 899 1882
rect 953 1836 966 1882
rect 886 1803 966 1836
rect 1070 1882 1150 1895
rect 1070 1836 1083 1882
rect 1137 1836 1150 1882
rect 1070 1803 1150 1836
rect 1254 1882 1334 1895
rect 1254 1836 1267 1882
rect 1321 1836 1334 1882
rect 1254 1803 1334 1836
rect 886 1270 966 1303
rect 886 1224 899 1270
rect 953 1224 966 1270
rect 886 1211 966 1224
rect 1070 1270 1150 1303
rect 1070 1224 1083 1270
rect 1137 1224 1150 1270
rect 1070 1211 1150 1224
rect 1254 1270 1334 1303
rect 1254 1224 1267 1270
rect 1321 1224 1334 1270
rect 1254 1211 1334 1224
rect 4898 1882 4978 1895
rect 4898 1836 4911 1882
rect 4965 1836 4978 1882
rect 4898 1803 4978 1836
rect 5082 1882 5162 1895
rect 5082 1836 5095 1882
rect 5149 1836 5162 1882
rect 5082 1803 5162 1836
rect 5266 1882 5346 1895
rect 5266 1836 5279 1882
rect 5333 1836 5346 1882
rect 5266 1803 5346 1836
rect 4898 1270 4978 1303
rect 4898 1224 4911 1270
rect 4965 1224 4978 1270
rect 4898 1211 4978 1224
rect 5082 1270 5162 1303
rect 5082 1224 5095 1270
rect 5149 1224 5162 1270
rect 5082 1211 5162 1224
rect 5266 1270 5346 1303
rect 5266 1224 5279 1270
rect 5333 1224 5346 1270
rect 5266 1211 5346 1224
rect 8940 1882 9020 1895
rect 8940 1836 8953 1882
rect 9007 1836 9020 1882
rect 8940 1803 9020 1836
rect 9124 1882 9204 1895
rect 9124 1836 9137 1882
rect 9191 1836 9204 1882
rect 9124 1803 9204 1836
rect 9308 1882 9388 1895
rect 9308 1836 9321 1882
rect 9375 1836 9388 1882
rect 9308 1803 9388 1836
rect 8940 1270 9020 1303
rect 8940 1224 8953 1270
rect 9007 1224 9020 1270
rect 8940 1211 9020 1224
rect 9124 1270 9204 1303
rect 9124 1224 9137 1270
rect 9191 1224 9204 1270
rect 9124 1211 9204 1224
rect 9308 1270 9388 1303
rect 9308 1224 9321 1270
rect 9375 1224 9388 1270
rect 9308 1211 9388 1224
rect 12982 1882 13062 1895
rect 12982 1836 12995 1882
rect 13049 1836 13062 1882
rect 12982 1803 13062 1836
rect 13166 1882 13246 1895
rect 13166 1836 13179 1882
rect 13233 1836 13246 1882
rect 13166 1803 13246 1836
rect 13350 1882 13430 1895
rect 13350 1836 13363 1882
rect 13417 1836 13430 1882
rect 13350 1803 13430 1836
rect 12982 1270 13062 1303
rect 12982 1224 12995 1270
rect 13049 1224 13062 1270
rect 12982 1211 13062 1224
rect 13166 1270 13246 1303
rect 13166 1224 13179 1270
rect 13233 1224 13246 1270
rect 13166 1211 13246 1224
rect 13350 1270 13430 1303
rect 13350 1224 13363 1270
rect 13417 1224 13430 1270
rect 13350 1211 13430 1224
rect 17024 1882 17104 1895
rect 17024 1836 17037 1882
rect 17091 1836 17104 1882
rect 17024 1803 17104 1836
rect 17208 1882 17288 1895
rect 17208 1836 17221 1882
rect 17275 1836 17288 1882
rect 17208 1803 17288 1836
rect 17392 1882 17472 1895
rect 17392 1836 17405 1882
rect 17459 1836 17472 1882
rect 17392 1803 17472 1836
rect 17024 1270 17104 1303
rect 17024 1224 17037 1270
rect 17091 1224 17104 1270
rect 17024 1211 17104 1224
rect 17208 1270 17288 1303
rect 17208 1224 17221 1270
rect 17275 1224 17288 1270
rect 17208 1211 17288 1224
rect 17392 1270 17472 1303
rect 17392 1224 17405 1270
rect 17459 1224 17472 1270
rect 17392 1211 17472 1224
rect 21066 1882 21146 1895
rect 21066 1836 21079 1882
rect 21133 1836 21146 1882
rect 21066 1803 21146 1836
rect 21250 1882 21330 1895
rect 21250 1836 21263 1882
rect 21317 1836 21330 1882
rect 21250 1803 21330 1836
rect 21434 1882 21514 1895
rect 21434 1836 21447 1882
rect 21501 1836 21514 1882
rect 21434 1803 21514 1836
rect 21066 1270 21146 1303
rect 21066 1224 21079 1270
rect 21133 1224 21146 1270
rect 21066 1211 21146 1224
rect 21250 1270 21330 1303
rect 21250 1224 21263 1270
rect 21317 1224 21330 1270
rect 21250 1211 21330 1224
rect 21434 1270 21514 1303
rect 21434 1224 21447 1270
rect 21501 1224 21514 1270
rect 21434 1211 21514 1224
rect 25108 1882 25188 1895
rect 25108 1836 25121 1882
rect 25175 1836 25188 1882
rect 25108 1803 25188 1836
rect 25292 1882 25372 1895
rect 25292 1836 25305 1882
rect 25359 1836 25372 1882
rect 25292 1803 25372 1836
rect 25476 1882 25556 1895
rect 25476 1836 25489 1882
rect 25543 1836 25556 1882
rect 25476 1803 25556 1836
rect 25108 1270 25188 1303
rect 25108 1224 25121 1270
rect 25175 1224 25188 1270
rect 25108 1211 25188 1224
rect 25292 1270 25372 1303
rect 25292 1224 25305 1270
rect 25359 1224 25372 1270
rect 25292 1211 25372 1224
rect 25476 1270 25556 1303
rect 25476 1224 25489 1270
rect 25543 1224 25556 1270
rect 25476 1211 25556 1224
rect 886 722 966 735
rect 886 676 899 722
rect 953 676 966 722
rect 886 643 966 676
rect 1070 722 1150 735
rect 1070 676 1083 722
rect 1137 676 1150 722
rect 1070 643 1150 676
rect 1254 722 1334 735
rect 1254 676 1267 722
rect 1321 676 1334 722
rect 1254 643 1334 676
rect 886 410 966 443
rect 886 364 899 410
rect 953 364 966 410
rect 886 351 966 364
rect 1070 410 1150 443
rect 1070 364 1083 410
rect 1137 364 1150 410
rect 1070 351 1150 364
rect 1254 410 1334 443
rect 1254 364 1267 410
rect 1321 364 1334 410
rect 1254 351 1334 364
rect 4898 722 4978 735
rect 4898 676 4911 722
rect 4965 676 4978 722
rect 4898 643 4978 676
rect 5082 722 5162 735
rect 5082 676 5095 722
rect 5149 676 5162 722
rect 5082 643 5162 676
rect 5266 722 5346 735
rect 5266 676 5279 722
rect 5333 676 5346 722
rect 5266 643 5346 676
rect 4898 410 4978 443
rect 4898 364 4911 410
rect 4965 364 4978 410
rect 4898 351 4978 364
rect 5082 410 5162 443
rect 5082 364 5095 410
rect 5149 364 5162 410
rect 5082 351 5162 364
rect 5266 410 5346 443
rect 5266 364 5279 410
rect 5333 364 5346 410
rect 5266 351 5346 364
rect 8940 722 9020 735
rect 8940 676 8953 722
rect 9007 676 9020 722
rect 8940 643 9020 676
rect 9124 722 9204 735
rect 9124 676 9137 722
rect 9191 676 9204 722
rect 9124 643 9204 676
rect 9308 722 9388 735
rect 9308 676 9321 722
rect 9375 676 9388 722
rect 9308 643 9388 676
rect 8940 410 9020 443
rect 8940 364 8953 410
rect 9007 364 9020 410
rect 8940 351 9020 364
rect 9124 410 9204 443
rect 9124 364 9137 410
rect 9191 364 9204 410
rect 9124 351 9204 364
rect 9308 410 9388 443
rect 9308 364 9321 410
rect 9375 364 9388 410
rect 9308 351 9388 364
rect 12982 722 13062 735
rect 12982 676 12995 722
rect 13049 676 13062 722
rect 12982 643 13062 676
rect 13166 722 13246 735
rect 13166 676 13179 722
rect 13233 676 13246 722
rect 13166 643 13246 676
rect 13350 722 13430 735
rect 13350 676 13363 722
rect 13417 676 13430 722
rect 13350 643 13430 676
rect 12982 410 13062 443
rect 12982 364 12995 410
rect 13049 364 13062 410
rect 12982 351 13062 364
rect 13166 410 13246 443
rect 13166 364 13179 410
rect 13233 364 13246 410
rect 13166 351 13246 364
rect 13350 410 13430 443
rect 13350 364 13363 410
rect 13417 364 13430 410
rect 13350 351 13430 364
rect 17024 722 17104 735
rect 17024 676 17037 722
rect 17091 676 17104 722
rect 17024 643 17104 676
rect 17208 722 17288 735
rect 17208 676 17221 722
rect 17275 676 17288 722
rect 17208 643 17288 676
rect 17392 722 17472 735
rect 17392 676 17405 722
rect 17459 676 17472 722
rect 17392 643 17472 676
rect 17024 410 17104 443
rect 17024 364 17037 410
rect 17091 364 17104 410
rect 17024 351 17104 364
rect 17208 410 17288 443
rect 17208 364 17221 410
rect 17275 364 17288 410
rect 17208 351 17288 364
rect 17392 410 17472 443
rect 17392 364 17405 410
rect 17459 364 17472 410
rect 17392 351 17472 364
rect 21066 722 21146 735
rect 21066 676 21079 722
rect 21133 676 21146 722
rect 21066 643 21146 676
rect 21250 722 21330 735
rect 21250 676 21263 722
rect 21317 676 21330 722
rect 21250 643 21330 676
rect 21434 722 21514 735
rect 21434 676 21447 722
rect 21501 676 21514 722
rect 21434 643 21514 676
rect 21066 410 21146 443
rect 21066 364 21079 410
rect 21133 364 21146 410
rect 21066 351 21146 364
rect 21250 410 21330 443
rect 21250 364 21263 410
rect 21317 364 21330 410
rect 21250 351 21330 364
rect 21434 410 21514 443
rect 21434 364 21447 410
rect 21501 364 21514 410
rect 21434 351 21514 364
rect 25108 722 25188 735
rect 25108 676 25121 722
rect 25175 676 25188 722
rect 25108 643 25188 676
rect 25292 722 25372 735
rect 25292 676 25305 722
rect 25359 676 25372 722
rect 25292 643 25372 676
rect 25476 722 25556 735
rect 25476 676 25489 722
rect 25543 676 25556 722
rect 25476 643 25556 676
rect 25108 410 25188 443
rect 25108 364 25121 410
rect 25175 364 25188 410
rect 25108 351 25188 364
rect 25292 410 25372 443
rect 25292 364 25305 410
rect 25359 364 25372 410
rect 25292 351 25372 364
rect 25476 410 25556 443
rect 25476 364 25489 410
rect 25543 364 25556 410
rect 25476 351 25556 364
<< polycontact >>
rect 4911 18030 4965 18076
rect 5095 18030 5149 18076
rect 5279 18030 5333 18076
rect 4911 17418 4965 17464
rect 5095 17418 5149 17464
rect 5279 17418 5333 17464
rect 8953 18027 9007 18073
rect 9137 18027 9191 18073
rect 9321 18027 9375 18073
rect 8953 17415 9007 17461
rect 9137 17415 9191 17461
rect 9321 17415 9375 17461
rect 12995 18027 13049 18073
rect 13179 18027 13233 18073
rect 13363 18027 13417 18073
rect 12995 17415 13049 17461
rect 13179 17415 13233 17461
rect 13363 17415 13417 17461
rect 17037 18027 17091 18073
rect 17221 18027 17275 18073
rect 17405 18027 17459 18073
rect 17037 17415 17091 17461
rect 17221 17415 17275 17461
rect 17405 17415 17459 17461
rect 21079 18027 21133 18073
rect 21263 18027 21317 18073
rect 21447 18027 21501 18073
rect 21079 17415 21133 17461
rect 21263 17415 21317 17461
rect 21447 17415 21501 17461
rect 25121 18027 25175 18073
rect 25305 18027 25359 18073
rect 25489 18027 25543 18073
rect 25121 17415 25175 17461
rect 25305 17415 25359 17461
rect 25489 17415 25543 17461
rect 29163 18027 29217 18073
rect 29347 18027 29401 18073
rect 29531 18027 29585 18073
rect 29163 17415 29217 17461
rect 29347 17415 29401 17461
rect 29531 17415 29585 17461
rect 4911 16870 4965 16916
rect 5095 16870 5149 16916
rect 5279 16870 5333 16916
rect 4911 16558 4965 16604
rect 5095 16558 5149 16604
rect 5279 16558 5333 16604
rect 8953 16867 9007 16913
rect 9137 16867 9191 16913
rect 9321 16867 9375 16913
rect 8953 16555 9007 16601
rect 9137 16555 9191 16601
rect 9321 16555 9375 16601
rect 12995 16867 13049 16913
rect 13179 16867 13233 16913
rect 13363 16867 13417 16913
rect 12995 16555 13049 16601
rect 13179 16555 13233 16601
rect 13363 16555 13417 16601
rect 17037 16867 17091 16913
rect 17221 16867 17275 16913
rect 17405 16867 17459 16913
rect 17037 16555 17091 16601
rect 17221 16555 17275 16601
rect 17405 16555 17459 16601
rect 21079 16867 21133 16913
rect 21263 16867 21317 16913
rect 21447 16867 21501 16913
rect 21079 16555 21133 16601
rect 21263 16555 21317 16601
rect 21447 16555 21501 16601
rect 25121 16867 25175 16913
rect 25305 16867 25359 16913
rect 25489 16867 25543 16913
rect 25121 16555 25175 16601
rect 25305 16555 25359 16601
rect 25489 16555 25543 16601
rect 29163 16867 29217 16913
rect 29347 16867 29401 16913
rect 29531 16867 29585 16913
rect 29163 16555 29217 16601
rect 29347 16555 29401 16601
rect 29531 16555 29585 16601
rect 4911 15825 4965 15871
rect 5095 15825 5149 15871
rect 5279 15825 5333 15871
rect 4911 15213 4965 15259
rect 5095 15213 5149 15259
rect 5279 15213 5333 15259
rect 6397 15825 6451 15871
rect 6581 15825 6635 15871
rect 6765 15825 6819 15871
rect 6397 15213 6451 15259
rect 6581 15213 6635 15259
rect 6765 15213 6819 15259
rect 8953 15822 9007 15868
rect 9137 15822 9191 15868
rect 9321 15822 9375 15868
rect 8953 15210 9007 15256
rect 9137 15210 9191 15256
rect 9321 15210 9375 15256
rect 10439 15822 10493 15868
rect 10623 15822 10677 15868
rect 10807 15822 10861 15868
rect 10439 15210 10493 15256
rect 10623 15210 10677 15256
rect 10807 15210 10861 15256
rect 12995 15822 13049 15868
rect 13179 15822 13233 15868
rect 13363 15822 13417 15868
rect 12995 15210 13049 15256
rect 13179 15210 13233 15256
rect 13363 15210 13417 15256
rect 14481 15822 14535 15868
rect 14665 15822 14719 15868
rect 14849 15822 14903 15868
rect 14481 15210 14535 15256
rect 14665 15210 14719 15256
rect 14849 15210 14903 15256
rect 17037 15822 17091 15868
rect 17221 15822 17275 15868
rect 17405 15822 17459 15868
rect 17037 15210 17091 15256
rect 17221 15210 17275 15256
rect 17405 15210 17459 15256
rect 18523 15822 18577 15868
rect 18707 15822 18761 15868
rect 18891 15822 18945 15868
rect 18523 15210 18577 15256
rect 18707 15210 18761 15256
rect 18891 15210 18945 15256
rect 21079 15822 21133 15868
rect 21263 15822 21317 15868
rect 21447 15822 21501 15868
rect 21079 15210 21133 15256
rect 21263 15210 21317 15256
rect 21447 15210 21501 15256
rect 22565 15822 22619 15868
rect 22749 15822 22803 15868
rect 22933 15822 22987 15868
rect 22565 15210 22619 15256
rect 22749 15210 22803 15256
rect 22933 15210 22987 15256
rect 25121 15822 25175 15868
rect 25305 15822 25359 15868
rect 25489 15822 25543 15868
rect 25121 15210 25175 15256
rect 25305 15210 25359 15256
rect 25489 15210 25543 15256
rect 26607 15822 26661 15868
rect 26791 15822 26845 15868
rect 26975 15822 27029 15868
rect 26607 15210 26661 15256
rect 26791 15210 26845 15256
rect 26975 15210 27029 15256
rect 29163 15822 29217 15868
rect 29347 15822 29401 15868
rect 29531 15822 29585 15868
rect 29163 15210 29217 15256
rect 29347 15210 29401 15256
rect 29531 15210 29585 15256
rect 30649 15822 30703 15868
rect 30833 15822 30887 15868
rect 31017 15822 31071 15868
rect 30649 15210 30703 15256
rect 30833 15210 30887 15256
rect 31017 15210 31071 15256
rect 4911 14665 4965 14711
rect 5095 14665 5149 14711
rect 5279 14665 5333 14711
rect 4911 14353 4965 14399
rect 5095 14353 5149 14399
rect 5279 14353 5333 14399
rect 6397 14665 6451 14711
rect 6581 14665 6635 14711
rect 6765 14665 6819 14711
rect 6397 14353 6451 14399
rect 6581 14353 6635 14399
rect 6765 14353 6819 14399
rect 8953 14662 9007 14708
rect 9137 14662 9191 14708
rect 9321 14662 9375 14708
rect 8953 14350 9007 14396
rect 9137 14350 9191 14396
rect 9321 14350 9375 14396
rect 10439 14662 10493 14708
rect 10623 14662 10677 14708
rect 10807 14662 10861 14708
rect 10439 14350 10493 14396
rect 10623 14350 10677 14396
rect 10807 14350 10861 14396
rect 12995 14662 13049 14708
rect 13179 14662 13233 14708
rect 13363 14662 13417 14708
rect 12995 14350 13049 14396
rect 13179 14350 13233 14396
rect 13363 14350 13417 14396
rect 14481 14662 14535 14708
rect 14665 14662 14719 14708
rect 14849 14662 14903 14708
rect 14481 14350 14535 14396
rect 14665 14350 14719 14396
rect 14849 14350 14903 14396
rect 17037 14662 17091 14708
rect 17221 14662 17275 14708
rect 17405 14662 17459 14708
rect 17037 14350 17091 14396
rect 17221 14350 17275 14396
rect 17405 14350 17459 14396
rect 18523 14662 18577 14708
rect 18707 14662 18761 14708
rect 18891 14662 18945 14708
rect 18523 14350 18577 14396
rect 18707 14350 18761 14396
rect 18891 14350 18945 14396
rect 21079 14662 21133 14708
rect 21263 14662 21317 14708
rect 21447 14662 21501 14708
rect 21079 14350 21133 14396
rect 21263 14350 21317 14396
rect 21447 14350 21501 14396
rect 22565 14662 22619 14708
rect 22749 14662 22803 14708
rect 22933 14662 22987 14708
rect 22565 14350 22619 14396
rect 22749 14350 22803 14396
rect 22933 14350 22987 14396
rect 25121 14662 25175 14708
rect 25305 14662 25359 14708
rect 25489 14662 25543 14708
rect 25121 14350 25175 14396
rect 25305 14350 25359 14396
rect 25489 14350 25543 14396
rect 26607 14662 26661 14708
rect 26791 14662 26845 14708
rect 26975 14662 27029 14708
rect 26607 14350 26661 14396
rect 26791 14350 26845 14396
rect 26975 14350 27029 14396
rect 29163 14662 29217 14708
rect 29347 14662 29401 14708
rect 29531 14662 29585 14708
rect 29163 14350 29217 14396
rect 29347 14350 29401 14396
rect 29531 14350 29585 14396
rect 30649 14662 30703 14708
rect 30833 14662 30887 14708
rect 31017 14662 31071 14708
rect 30649 14350 30703 14396
rect 30833 14350 30887 14396
rect 31017 14350 31071 14396
rect 4911 13620 4965 13666
rect 5095 13620 5149 13666
rect 5279 13620 5333 13666
rect 4911 13008 4965 13054
rect 5095 13008 5149 13054
rect 5279 13008 5333 13054
rect 6397 13621 6451 13667
rect 6581 13621 6635 13667
rect 6765 13621 6819 13667
rect 6397 13009 6451 13055
rect 6581 13009 6635 13055
rect 6765 13009 6819 13055
rect 8953 13617 9007 13663
rect 9137 13617 9191 13663
rect 9321 13617 9375 13663
rect 8953 13005 9007 13051
rect 9137 13005 9191 13051
rect 9321 13005 9375 13051
rect 10439 13618 10493 13664
rect 10623 13618 10677 13664
rect 10807 13618 10861 13664
rect 10439 13006 10493 13052
rect 10623 13006 10677 13052
rect 10807 13006 10861 13052
rect 12995 13617 13049 13663
rect 13179 13617 13233 13663
rect 13363 13617 13417 13663
rect 12995 13005 13049 13051
rect 13179 13005 13233 13051
rect 13363 13005 13417 13051
rect 14481 13618 14535 13664
rect 14665 13618 14719 13664
rect 14849 13618 14903 13664
rect 14481 13006 14535 13052
rect 14665 13006 14719 13052
rect 14849 13006 14903 13052
rect 17037 13617 17091 13663
rect 17221 13617 17275 13663
rect 17405 13617 17459 13663
rect 17037 13005 17091 13051
rect 17221 13005 17275 13051
rect 17405 13005 17459 13051
rect 18523 13618 18577 13664
rect 18707 13618 18761 13664
rect 18891 13618 18945 13664
rect 18523 13006 18577 13052
rect 18707 13006 18761 13052
rect 18891 13006 18945 13052
rect 21079 13617 21133 13663
rect 21263 13617 21317 13663
rect 21447 13617 21501 13663
rect 21079 13005 21133 13051
rect 21263 13005 21317 13051
rect 21447 13005 21501 13051
rect 22565 13618 22619 13664
rect 22749 13618 22803 13664
rect 22933 13618 22987 13664
rect 22565 13006 22619 13052
rect 22749 13006 22803 13052
rect 22933 13006 22987 13052
rect 25121 13617 25175 13663
rect 25305 13617 25359 13663
rect 25489 13617 25543 13663
rect 25121 13005 25175 13051
rect 25305 13005 25359 13051
rect 25489 13005 25543 13051
rect 26607 13618 26661 13664
rect 26791 13618 26845 13664
rect 26975 13618 27029 13664
rect 26607 13006 26661 13052
rect 26791 13006 26845 13052
rect 26975 13006 27029 13052
rect 29163 13617 29217 13663
rect 29347 13617 29401 13663
rect 29531 13617 29585 13663
rect 29163 13005 29217 13051
rect 29347 13005 29401 13051
rect 29531 13005 29585 13051
rect 30649 13618 30703 13664
rect 30833 13618 30887 13664
rect 31017 13618 31071 13664
rect 30649 13006 30703 13052
rect 30833 13006 30887 13052
rect 31017 13006 31071 13052
rect 4911 12460 4965 12506
rect 5095 12460 5149 12506
rect 5279 12460 5333 12506
rect 4911 12148 4965 12194
rect 5095 12148 5149 12194
rect 5279 12148 5333 12194
rect 6397 12461 6451 12507
rect 6581 12461 6635 12507
rect 6765 12461 6819 12507
rect 6397 12149 6451 12195
rect 6581 12149 6635 12195
rect 6765 12149 6819 12195
rect 8953 12457 9007 12503
rect 9137 12457 9191 12503
rect 9321 12457 9375 12503
rect 8953 12145 9007 12191
rect 9137 12145 9191 12191
rect 9321 12145 9375 12191
rect 10439 12458 10493 12504
rect 10623 12458 10677 12504
rect 10807 12458 10861 12504
rect 10439 12146 10493 12192
rect 10623 12146 10677 12192
rect 10807 12146 10861 12192
rect 12995 12457 13049 12503
rect 13179 12457 13233 12503
rect 13363 12457 13417 12503
rect 12995 12145 13049 12191
rect 13179 12145 13233 12191
rect 13363 12145 13417 12191
rect 14481 12458 14535 12504
rect 14665 12458 14719 12504
rect 14849 12458 14903 12504
rect 14481 12146 14535 12192
rect 14665 12146 14719 12192
rect 14849 12146 14903 12192
rect 17037 12457 17091 12503
rect 17221 12457 17275 12503
rect 17405 12457 17459 12503
rect 17037 12145 17091 12191
rect 17221 12145 17275 12191
rect 17405 12145 17459 12191
rect 18523 12458 18577 12504
rect 18707 12458 18761 12504
rect 18891 12458 18945 12504
rect 18523 12146 18577 12192
rect 18707 12146 18761 12192
rect 18891 12146 18945 12192
rect 21079 12457 21133 12503
rect 21263 12457 21317 12503
rect 21447 12457 21501 12503
rect 21079 12145 21133 12191
rect 21263 12145 21317 12191
rect 21447 12145 21501 12191
rect 22565 12458 22619 12504
rect 22749 12458 22803 12504
rect 22933 12458 22987 12504
rect 22565 12146 22619 12192
rect 22749 12146 22803 12192
rect 22933 12146 22987 12192
rect 25121 12457 25175 12503
rect 25305 12457 25359 12503
rect 25489 12457 25543 12503
rect 25121 12145 25175 12191
rect 25305 12145 25359 12191
rect 25489 12145 25543 12191
rect 26607 12458 26661 12504
rect 26791 12458 26845 12504
rect 26975 12458 27029 12504
rect 26607 12146 26661 12192
rect 26791 12146 26845 12192
rect 26975 12146 27029 12192
rect 29163 12457 29217 12503
rect 29347 12457 29401 12503
rect 29531 12457 29585 12503
rect 29163 12145 29217 12191
rect 29347 12145 29401 12191
rect 29531 12145 29585 12191
rect 30649 12458 30703 12504
rect 30833 12458 30887 12504
rect 31017 12458 31071 12504
rect 30649 12146 30703 12192
rect 30833 12146 30887 12192
rect 31017 12146 31071 12192
rect 4911 11415 4965 11461
rect 5095 11415 5149 11461
rect 5279 11415 5333 11461
rect 4911 10803 4965 10849
rect 5095 10803 5149 10849
rect 5279 10803 5333 10849
rect 8953 11412 9007 11458
rect 9137 11412 9191 11458
rect 9321 11412 9375 11458
rect 8953 10800 9007 10846
rect 9137 10800 9191 10846
rect 9321 10800 9375 10846
rect 12995 11412 13049 11458
rect 13179 11412 13233 11458
rect 13363 11412 13417 11458
rect 12995 10800 13049 10846
rect 13179 10800 13233 10846
rect 13363 10800 13417 10846
rect 17037 11412 17091 11458
rect 17221 11412 17275 11458
rect 17405 11412 17459 11458
rect 17037 10800 17091 10846
rect 17221 10800 17275 10846
rect 17405 10800 17459 10846
rect 21079 11412 21133 11458
rect 21263 11412 21317 11458
rect 21447 11412 21501 11458
rect 21079 10800 21133 10846
rect 21263 10800 21317 10846
rect 21447 10800 21501 10846
rect 25121 11412 25175 11458
rect 25305 11412 25359 11458
rect 25489 11412 25543 11458
rect 25121 10800 25175 10846
rect 25305 10800 25359 10846
rect 25489 10800 25543 10846
rect 29163 11412 29217 11458
rect 29347 11412 29401 11458
rect 29531 11412 29585 11458
rect 29163 10800 29217 10846
rect 29347 10800 29401 10846
rect 29531 10800 29585 10846
rect 4911 10255 4965 10301
rect 5095 10255 5149 10301
rect 5279 10255 5333 10301
rect 4911 9943 4965 9989
rect 5095 9943 5149 9989
rect 5279 9943 5333 9989
rect 8953 10252 9007 10298
rect 9137 10252 9191 10298
rect 9321 10252 9375 10298
rect 8953 9940 9007 9986
rect 9137 9940 9191 9986
rect 9321 9940 9375 9986
rect 12995 10252 13049 10298
rect 13179 10252 13233 10298
rect 13363 10252 13417 10298
rect 12995 9940 13049 9986
rect 13179 9940 13233 9986
rect 13363 9940 13417 9986
rect 17037 10252 17091 10298
rect 17221 10252 17275 10298
rect 17405 10252 17459 10298
rect 17037 9940 17091 9986
rect 17221 9940 17275 9986
rect 17405 9940 17459 9986
rect 21079 10252 21133 10298
rect 21263 10252 21317 10298
rect 21447 10252 21501 10298
rect 21079 9940 21133 9986
rect 21263 9940 21317 9986
rect 21447 9940 21501 9986
rect 25121 10252 25175 10298
rect 25305 10252 25359 10298
rect 25489 10252 25543 10298
rect 25121 9940 25175 9986
rect 25305 9940 25359 9986
rect 25489 9940 25543 9986
rect 29163 10252 29217 10298
rect 29347 10252 29401 10298
rect 29531 10252 29585 10298
rect 29163 9940 29217 9986
rect 29347 9940 29401 9986
rect 29531 9940 29585 9986
rect 899 8451 953 8497
rect 1083 8451 1137 8497
rect 1267 8451 1321 8497
rect 899 7839 953 7885
rect 1083 7839 1137 7885
rect 1267 7839 1321 7885
rect 4911 8451 4965 8497
rect 5095 8451 5149 8497
rect 5279 8451 5333 8497
rect 4911 7839 4965 7885
rect 5095 7839 5149 7885
rect 5279 7839 5333 7885
rect 8953 8451 9007 8497
rect 9137 8451 9191 8497
rect 9321 8451 9375 8497
rect 8953 7839 9007 7885
rect 9137 7839 9191 7885
rect 9321 7839 9375 7885
rect 12995 8451 13049 8497
rect 13179 8451 13233 8497
rect 13363 8451 13417 8497
rect 12995 7839 13049 7885
rect 13179 7839 13233 7885
rect 13363 7839 13417 7885
rect 17037 8451 17091 8497
rect 17221 8451 17275 8497
rect 17405 8451 17459 8497
rect 17037 7839 17091 7885
rect 17221 7839 17275 7885
rect 17405 7839 17459 7885
rect 21079 8451 21133 8497
rect 21263 8451 21317 8497
rect 21447 8451 21501 8497
rect 21079 7839 21133 7885
rect 21263 7839 21317 7885
rect 21447 7839 21501 7885
rect 25121 8451 25175 8497
rect 25305 8451 25359 8497
rect 25489 8451 25543 8497
rect 25121 7839 25175 7885
rect 25305 7839 25359 7885
rect 25489 7839 25543 7885
rect 899 7291 953 7337
rect 1083 7291 1137 7337
rect 1267 7291 1321 7337
rect 899 6979 953 7025
rect 1083 6979 1137 7025
rect 1267 6979 1321 7025
rect 4911 7291 4965 7337
rect 5095 7291 5149 7337
rect 5279 7291 5333 7337
rect 4911 6979 4965 7025
rect 5095 6979 5149 7025
rect 5279 6979 5333 7025
rect 8953 7291 9007 7337
rect 9137 7291 9191 7337
rect 9321 7291 9375 7337
rect 8953 6979 9007 7025
rect 9137 6979 9191 7025
rect 9321 6979 9375 7025
rect 12995 7291 13049 7337
rect 13179 7291 13233 7337
rect 13363 7291 13417 7337
rect 12995 6979 13049 7025
rect 13179 6979 13233 7025
rect 13363 6979 13417 7025
rect 17037 7291 17091 7337
rect 17221 7291 17275 7337
rect 17405 7291 17459 7337
rect 17037 6979 17091 7025
rect 17221 6979 17275 7025
rect 17405 6979 17459 7025
rect 21079 7291 21133 7337
rect 21263 7291 21317 7337
rect 21447 7291 21501 7337
rect 21079 6979 21133 7025
rect 21263 6979 21317 7025
rect 21447 6979 21501 7025
rect 25121 7291 25175 7337
rect 25305 7291 25359 7337
rect 25489 7291 25543 7337
rect 25121 6979 25175 7025
rect 25305 6979 25359 7025
rect 25489 6979 25543 7025
rect 899 6246 953 6292
rect 1083 6246 1137 6292
rect 1267 6246 1321 6292
rect 899 5634 953 5680
rect 1083 5634 1137 5680
rect 1267 5634 1321 5680
rect 2385 6246 2439 6292
rect 2569 6246 2623 6292
rect 2753 6246 2807 6292
rect 2385 5634 2439 5680
rect 2569 5634 2623 5680
rect 2753 5634 2807 5680
rect 4911 6246 4965 6292
rect 5095 6246 5149 6292
rect 5279 6246 5333 6292
rect 4911 5634 4965 5680
rect 5095 5634 5149 5680
rect 5279 5634 5333 5680
rect 6397 6246 6451 6292
rect 6581 6246 6635 6292
rect 6765 6246 6819 6292
rect 6397 5634 6451 5680
rect 6581 5634 6635 5680
rect 6765 5634 6819 5680
rect 8953 6246 9007 6292
rect 9137 6246 9191 6292
rect 9321 6246 9375 6292
rect 8953 5634 9007 5680
rect 9137 5634 9191 5680
rect 9321 5634 9375 5680
rect 10439 6246 10493 6292
rect 10623 6246 10677 6292
rect 10807 6246 10861 6292
rect 10439 5634 10493 5680
rect 10623 5634 10677 5680
rect 10807 5634 10861 5680
rect 12995 6246 13049 6292
rect 13179 6246 13233 6292
rect 13363 6246 13417 6292
rect 12995 5634 13049 5680
rect 13179 5634 13233 5680
rect 13363 5634 13417 5680
rect 14481 6246 14535 6292
rect 14665 6246 14719 6292
rect 14849 6246 14903 6292
rect 14481 5634 14535 5680
rect 14665 5634 14719 5680
rect 14849 5634 14903 5680
rect 17037 6246 17091 6292
rect 17221 6246 17275 6292
rect 17405 6246 17459 6292
rect 17037 5634 17091 5680
rect 17221 5634 17275 5680
rect 17405 5634 17459 5680
rect 18523 6246 18577 6292
rect 18707 6246 18761 6292
rect 18891 6246 18945 6292
rect 18523 5634 18577 5680
rect 18707 5634 18761 5680
rect 18891 5634 18945 5680
rect 21079 6246 21133 6292
rect 21263 6246 21317 6292
rect 21447 6246 21501 6292
rect 21079 5634 21133 5680
rect 21263 5634 21317 5680
rect 21447 5634 21501 5680
rect 22565 6246 22619 6292
rect 22749 6246 22803 6292
rect 22933 6246 22987 6292
rect 22565 5634 22619 5680
rect 22749 5634 22803 5680
rect 22933 5634 22987 5680
rect 25121 6246 25175 6292
rect 25305 6246 25359 6292
rect 25489 6246 25543 6292
rect 25121 5634 25175 5680
rect 25305 5634 25359 5680
rect 25489 5634 25543 5680
rect 26607 6246 26661 6292
rect 26791 6246 26845 6292
rect 26975 6246 27029 6292
rect 26607 5634 26661 5680
rect 26791 5634 26845 5680
rect 26975 5634 27029 5680
rect 899 5086 953 5132
rect 1083 5086 1137 5132
rect 1267 5086 1321 5132
rect 899 4774 953 4820
rect 1083 4774 1137 4820
rect 1267 4774 1321 4820
rect 2385 5086 2439 5132
rect 2569 5086 2623 5132
rect 2753 5086 2807 5132
rect 2385 4774 2439 4820
rect 2569 4774 2623 4820
rect 2753 4774 2807 4820
rect 4911 5086 4965 5132
rect 5095 5086 5149 5132
rect 5279 5086 5333 5132
rect 4911 4774 4965 4820
rect 5095 4774 5149 4820
rect 5279 4774 5333 4820
rect 6397 5086 6451 5132
rect 6581 5086 6635 5132
rect 6765 5086 6819 5132
rect 6397 4774 6451 4820
rect 6581 4774 6635 4820
rect 6765 4774 6819 4820
rect 8953 5086 9007 5132
rect 9137 5086 9191 5132
rect 9321 5086 9375 5132
rect 8953 4774 9007 4820
rect 9137 4774 9191 4820
rect 9321 4774 9375 4820
rect 10439 5086 10493 5132
rect 10623 5086 10677 5132
rect 10807 5086 10861 5132
rect 10439 4774 10493 4820
rect 10623 4774 10677 4820
rect 10807 4774 10861 4820
rect 12995 5086 13049 5132
rect 13179 5086 13233 5132
rect 13363 5086 13417 5132
rect 12995 4774 13049 4820
rect 13179 4774 13233 4820
rect 13363 4774 13417 4820
rect 14481 5086 14535 5132
rect 14665 5086 14719 5132
rect 14849 5086 14903 5132
rect 14481 4774 14535 4820
rect 14665 4774 14719 4820
rect 14849 4774 14903 4820
rect 17037 5086 17091 5132
rect 17221 5086 17275 5132
rect 17405 5086 17459 5132
rect 17037 4774 17091 4820
rect 17221 4774 17275 4820
rect 17405 4774 17459 4820
rect 18523 5086 18577 5132
rect 18707 5086 18761 5132
rect 18891 5086 18945 5132
rect 18523 4774 18577 4820
rect 18707 4774 18761 4820
rect 18891 4774 18945 4820
rect 21079 5086 21133 5132
rect 21263 5086 21317 5132
rect 21447 5086 21501 5132
rect 21079 4774 21133 4820
rect 21263 4774 21317 4820
rect 21447 4774 21501 4820
rect 22565 5086 22619 5132
rect 22749 5086 22803 5132
rect 22933 5086 22987 5132
rect 22565 4774 22619 4820
rect 22749 4774 22803 4820
rect 22933 4774 22987 4820
rect 25121 5086 25175 5132
rect 25305 5086 25359 5132
rect 25489 5086 25543 5132
rect 25121 4774 25175 4820
rect 25305 4774 25359 4820
rect 25489 4774 25543 4820
rect 26607 5086 26661 5132
rect 26791 5086 26845 5132
rect 26975 5086 27029 5132
rect 26607 4774 26661 4820
rect 26791 4774 26845 4820
rect 26975 4774 27029 4820
rect 899 4041 953 4087
rect 1083 4041 1137 4087
rect 1267 4041 1321 4087
rect 899 3429 953 3475
rect 1083 3429 1137 3475
rect 1267 3429 1321 3475
rect 2385 4042 2439 4088
rect 2569 4042 2623 4088
rect 2753 4042 2807 4088
rect 2385 3430 2439 3476
rect 2569 3430 2623 3476
rect 2753 3430 2807 3476
rect 4911 4041 4965 4087
rect 5095 4041 5149 4087
rect 5279 4041 5333 4087
rect 4911 3429 4965 3475
rect 5095 3429 5149 3475
rect 5279 3429 5333 3475
rect 6397 4042 6451 4088
rect 6581 4042 6635 4088
rect 6765 4042 6819 4088
rect 6397 3430 6451 3476
rect 6581 3430 6635 3476
rect 6765 3430 6819 3476
rect 8953 4041 9007 4087
rect 9137 4041 9191 4087
rect 9321 4041 9375 4087
rect 8953 3429 9007 3475
rect 9137 3429 9191 3475
rect 9321 3429 9375 3475
rect 10439 4042 10493 4088
rect 10623 4042 10677 4088
rect 10807 4042 10861 4088
rect 10439 3430 10493 3476
rect 10623 3430 10677 3476
rect 10807 3430 10861 3476
rect 12995 4041 13049 4087
rect 13179 4041 13233 4087
rect 13363 4041 13417 4087
rect 12995 3429 13049 3475
rect 13179 3429 13233 3475
rect 13363 3429 13417 3475
rect 14481 4042 14535 4088
rect 14665 4042 14719 4088
rect 14849 4042 14903 4088
rect 14481 3430 14535 3476
rect 14665 3430 14719 3476
rect 14849 3430 14903 3476
rect 17037 4041 17091 4087
rect 17221 4041 17275 4087
rect 17405 4041 17459 4087
rect 17037 3429 17091 3475
rect 17221 3429 17275 3475
rect 17405 3429 17459 3475
rect 18523 4042 18577 4088
rect 18707 4042 18761 4088
rect 18891 4042 18945 4088
rect 18523 3430 18577 3476
rect 18707 3430 18761 3476
rect 18891 3430 18945 3476
rect 21079 4041 21133 4087
rect 21263 4041 21317 4087
rect 21447 4041 21501 4087
rect 21079 3429 21133 3475
rect 21263 3429 21317 3475
rect 21447 3429 21501 3475
rect 22565 4042 22619 4088
rect 22749 4042 22803 4088
rect 22933 4042 22987 4088
rect 22565 3430 22619 3476
rect 22749 3430 22803 3476
rect 22933 3430 22987 3476
rect 25121 4041 25175 4087
rect 25305 4041 25359 4087
rect 25489 4041 25543 4087
rect 25121 3429 25175 3475
rect 25305 3429 25359 3475
rect 25489 3429 25543 3475
rect 26607 4042 26661 4088
rect 26791 4042 26845 4088
rect 26975 4042 27029 4088
rect 26607 3430 26661 3476
rect 26791 3430 26845 3476
rect 26975 3430 27029 3476
rect 899 2881 953 2927
rect 1083 2881 1137 2927
rect 1267 2881 1321 2927
rect 899 2569 953 2615
rect 1083 2569 1137 2615
rect 1267 2569 1321 2615
rect 2385 2882 2439 2928
rect 2569 2882 2623 2928
rect 2753 2882 2807 2928
rect 2385 2570 2439 2616
rect 2569 2570 2623 2616
rect 2753 2570 2807 2616
rect 4911 2881 4965 2927
rect 5095 2881 5149 2927
rect 5279 2881 5333 2927
rect 4911 2569 4965 2615
rect 5095 2569 5149 2615
rect 5279 2569 5333 2615
rect 6397 2882 6451 2928
rect 6581 2882 6635 2928
rect 6765 2882 6819 2928
rect 6397 2570 6451 2616
rect 6581 2570 6635 2616
rect 6765 2570 6819 2616
rect 8953 2881 9007 2927
rect 9137 2881 9191 2927
rect 9321 2881 9375 2927
rect 8953 2569 9007 2615
rect 9137 2569 9191 2615
rect 9321 2569 9375 2615
rect 10439 2882 10493 2928
rect 10623 2882 10677 2928
rect 10807 2882 10861 2928
rect 10439 2570 10493 2616
rect 10623 2570 10677 2616
rect 10807 2570 10861 2616
rect 12995 2881 13049 2927
rect 13179 2881 13233 2927
rect 13363 2881 13417 2927
rect 12995 2569 13049 2615
rect 13179 2569 13233 2615
rect 13363 2569 13417 2615
rect 14481 2882 14535 2928
rect 14665 2882 14719 2928
rect 14849 2882 14903 2928
rect 14481 2570 14535 2616
rect 14665 2570 14719 2616
rect 14849 2570 14903 2616
rect 17037 2881 17091 2927
rect 17221 2881 17275 2927
rect 17405 2881 17459 2927
rect 17037 2569 17091 2615
rect 17221 2569 17275 2615
rect 17405 2569 17459 2615
rect 18523 2882 18577 2928
rect 18707 2882 18761 2928
rect 18891 2882 18945 2928
rect 18523 2570 18577 2616
rect 18707 2570 18761 2616
rect 18891 2570 18945 2616
rect 21079 2881 21133 2927
rect 21263 2881 21317 2927
rect 21447 2881 21501 2927
rect 21079 2569 21133 2615
rect 21263 2569 21317 2615
rect 21447 2569 21501 2615
rect 22565 2882 22619 2928
rect 22749 2882 22803 2928
rect 22933 2882 22987 2928
rect 22565 2570 22619 2616
rect 22749 2570 22803 2616
rect 22933 2570 22987 2616
rect 25121 2881 25175 2927
rect 25305 2881 25359 2927
rect 25489 2881 25543 2927
rect 25121 2569 25175 2615
rect 25305 2569 25359 2615
rect 25489 2569 25543 2615
rect 26607 2882 26661 2928
rect 26791 2882 26845 2928
rect 26975 2882 27029 2928
rect 26607 2570 26661 2616
rect 26791 2570 26845 2616
rect 26975 2570 27029 2616
rect 899 1836 953 1882
rect 1083 1836 1137 1882
rect 1267 1836 1321 1882
rect 899 1224 953 1270
rect 1083 1224 1137 1270
rect 1267 1224 1321 1270
rect 4911 1836 4965 1882
rect 5095 1836 5149 1882
rect 5279 1836 5333 1882
rect 4911 1224 4965 1270
rect 5095 1224 5149 1270
rect 5279 1224 5333 1270
rect 8953 1836 9007 1882
rect 9137 1836 9191 1882
rect 9321 1836 9375 1882
rect 8953 1224 9007 1270
rect 9137 1224 9191 1270
rect 9321 1224 9375 1270
rect 12995 1836 13049 1882
rect 13179 1836 13233 1882
rect 13363 1836 13417 1882
rect 12995 1224 13049 1270
rect 13179 1224 13233 1270
rect 13363 1224 13417 1270
rect 17037 1836 17091 1882
rect 17221 1836 17275 1882
rect 17405 1836 17459 1882
rect 17037 1224 17091 1270
rect 17221 1224 17275 1270
rect 17405 1224 17459 1270
rect 21079 1836 21133 1882
rect 21263 1836 21317 1882
rect 21447 1836 21501 1882
rect 21079 1224 21133 1270
rect 21263 1224 21317 1270
rect 21447 1224 21501 1270
rect 25121 1836 25175 1882
rect 25305 1836 25359 1882
rect 25489 1836 25543 1882
rect 25121 1224 25175 1270
rect 25305 1224 25359 1270
rect 25489 1224 25543 1270
rect 899 676 953 722
rect 1083 676 1137 722
rect 1267 676 1321 722
rect 899 364 953 410
rect 1083 364 1137 410
rect 1267 364 1321 410
rect 4911 676 4965 722
rect 5095 676 5149 722
rect 5279 676 5333 722
rect 4911 364 4965 410
rect 5095 364 5149 410
rect 5279 364 5333 410
rect 8953 676 9007 722
rect 9137 676 9191 722
rect 9321 676 9375 722
rect 8953 364 9007 410
rect 9137 364 9191 410
rect 9321 364 9375 410
rect 12995 676 13049 722
rect 13179 676 13233 722
rect 13363 676 13417 722
rect 12995 364 13049 410
rect 13179 364 13233 410
rect 13363 364 13417 410
rect 17037 676 17091 722
rect 17221 676 17275 722
rect 17405 676 17459 722
rect 17037 364 17091 410
rect 17221 364 17275 410
rect 17405 364 17459 410
rect 21079 676 21133 722
rect 21263 676 21317 722
rect 21447 676 21501 722
rect 21079 364 21133 410
rect 21263 364 21317 410
rect 21447 364 21501 410
rect 25121 676 25175 722
rect 25305 676 25359 722
rect 25489 676 25543 722
rect 25121 364 25175 410
rect 25305 364 25359 410
rect 25489 364 25543 410
<< metal1 >>
rect 12038 19089 12108 19101
rect 19896 19089 19966 19091
rect 12038 19033 12050 19089
rect 12106 19033 19898 19089
rect 19954 19033 19966 19089
rect 12038 19031 12108 19033
rect 19896 19031 19966 19033
rect 16080 18913 16150 18925
rect 23938 18913 24008 18915
rect 16080 18857 16092 18913
rect 16148 18857 23940 18913
rect 23996 18857 24008 18913
rect 16080 18855 16150 18857
rect 23938 18855 24008 18857
rect 3900 18737 3970 18749
rect 11758 18737 11828 18739
rect 3900 18681 3912 18737
rect 3968 18681 11760 18737
rect 11816 18681 11828 18737
rect 3900 18679 3970 18681
rect 11758 18679 11828 18681
rect 20122 18737 20192 18749
rect 27980 18737 28050 18739
rect 20122 18681 20134 18737
rect 20190 18681 27982 18737
rect 28038 18681 28050 18737
rect 20122 18679 20192 18681
rect 27980 18679 28050 18681
rect 7996 18561 8066 18573
rect 15854 18561 15924 18563
rect 7996 18505 8008 18561
rect 8064 18505 15856 18561
rect 15912 18505 15924 18561
rect 7996 18503 8066 18505
rect 15854 18503 15924 18505
rect 24164 18561 24234 18573
rect 32022 18561 32092 18573
rect 24164 18505 24176 18561
rect 24232 18505 32024 18561
rect 32080 18505 32092 18561
rect 24164 18503 24234 18505
rect 32022 18503 32092 18505
rect 4505 18332 6052 18388
rect 3546 17311 3616 17323
rect 4505 17311 4561 18332
rect 5174 18280 5260 18284
rect 5174 18224 5186 18280
rect 5242 18224 5260 18280
rect 5174 18212 5260 18224
rect 4685 18067 4731 18078
rect 4900 18076 4976 18109
rect 4900 18030 4911 18076
rect 4965 18030 4976 18076
rect 5084 18076 5160 18109
rect 5084 18030 5095 18076
rect 5149 18030 5160 18076
rect 5268 18076 5344 18109
rect 5268 18030 5279 18076
rect 5333 18030 5344 18076
rect 5513 18067 5559 18078
rect 4823 17984 4869 17995
rect 4806 17957 4823 17959
rect 5007 17984 5053 17995
rect 4869 17957 4886 17959
rect 4731 17837 4818 17957
rect 4874 17837 4886 17957
rect 4806 17835 4823 17837
rect 4731 17537 4823 17657
rect 4869 17835 4886 17837
rect 4990 17657 5007 17659
rect 5191 17984 5237 17995
rect 5174 17957 5191 17959
rect 5375 17984 5421 17995
rect 5237 17957 5254 17959
rect 5174 17837 5186 17957
rect 5242 17837 5254 17957
rect 5174 17835 5191 17837
rect 5053 17657 5070 17659
rect 4990 17537 5002 17657
rect 5058 17537 5070 17657
rect 4990 17535 5007 17537
rect 4823 17499 4869 17510
rect 5053 17535 5070 17537
rect 5007 17499 5053 17510
rect 5237 17835 5254 17837
rect 5358 17657 5375 17659
rect 5496 17957 5513 17959
rect 5559 17957 5576 17959
rect 5496 17836 5508 17957
rect 5564 17836 5576 17957
rect 5496 17834 5513 17836
rect 5421 17657 5438 17659
rect 5358 17537 5370 17657
rect 5426 17537 5438 17657
rect 5358 17535 5375 17537
rect 5191 17499 5237 17510
rect 5421 17535 5438 17537
rect 5375 17499 5421 17510
rect 4900 17461 4911 17464
rect 4965 17461 4976 17464
rect 5084 17461 5095 17464
rect 5149 17461 5160 17464
rect 5268 17461 5279 17464
rect 5333 17461 5344 17464
rect 4685 17416 4731 17427
rect 4898 17405 4910 17461
rect 4966 17405 4978 17461
rect 4898 17391 4978 17405
rect 5082 17405 5094 17461
rect 5150 17405 5162 17461
rect 5082 17391 5162 17405
rect 5266 17405 5278 17461
rect 5334 17405 5346 17461
rect 5559 17834 5576 17836
rect 5513 17416 5559 17427
rect 5266 17391 5346 17405
rect 4898 17311 4978 17313
rect 3546 17255 3558 17311
rect 3614 17255 4910 17311
rect 4966 17255 4978 17311
rect 3546 17253 3616 17255
rect 4898 17253 4978 17255
rect 4226 17195 4296 17207
rect 5082 17195 5162 17197
rect 4226 17139 4238 17195
rect 4294 17139 5094 17195
rect 5150 17139 5162 17195
rect 4226 17127 4296 17139
rect 5082 17137 5162 17139
rect 5411 17195 5491 17197
rect 5678 17195 5748 17207
rect 5411 17139 5423 17195
rect 5479 17139 5680 17195
rect 5736 17139 5748 17195
rect 5411 17137 5491 17139
rect 5678 17129 5748 17139
rect 5266 17079 5346 17081
rect 4510 17023 5278 17079
rect 5334 17023 5346 17079
rect 4510 16292 4566 17023
rect 5266 17021 5346 17023
rect 4898 16929 4978 16943
rect 4685 16907 4731 16918
rect 4898 16873 4910 16929
rect 4966 16873 4978 16929
rect 5082 16929 5162 16943
rect 5082 16873 5094 16929
rect 5150 16873 5162 16929
rect 5266 16929 5346 16943
rect 5266 16873 5278 16929
rect 5334 16873 5346 16929
rect 5513 16907 5559 16918
rect 4900 16870 4911 16873
rect 4965 16870 4976 16873
rect 5084 16870 5095 16873
rect 5149 16870 5160 16873
rect 5268 16870 5279 16873
rect 5333 16870 5344 16873
rect 4823 16824 4869 16835
rect 4731 16650 4823 16824
rect 4823 16639 4869 16650
rect 5007 16824 5053 16835
rect 5007 16639 5053 16650
rect 5191 16824 5237 16835
rect 5375 16824 5421 16835
rect 5358 16797 5375 16799
rect 5421 16797 5438 16799
rect 5358 16677 5370 16797
rect 5426 16677 5438 16797
rect 5358 16675 5375 16677
rect 5191 16639 5237 16650
rect 5421 16675 5438 16677
rect 5375 16639 5421 16650
rect 4685 16422 4731 16567
rect 4900 16558 4911 16604
rect 4965 16558 4976 16604
rect 4900 16525 4976 16558
rect 5084 16558 5095 16604
rect 5149 16558 5160 16604
rect 5084 16525 5160 16558
rect 5268 16558 5279 16604
rect 5333 16558 5344 16604
rect 5268 16525 5344 16558
rect 5513 16422 5559 16567
rect 4673 16410 4753 16422
rect 4673 16354 4685 16410
rect 4741 16354 4753 16410
rect 4673 16342 4753 16354
rect 5491 16410 5571 16422
rect 5491 16354 5503 16410
rect 5559 16354 5571 16410
rect 5491 16342 5571 16354
rect 5844 16292 5924 16302
rect 4510 16236 5856 16292
rect 5912 16236 5924 16292
rect 5844 16234 5924 16236
rect 5678 16183 5748 16185
rect 4510 16182 5748 16183
rect 4510 16128 5680 16182
rect 5736 16128 5748 16182
rect 4510 16127 5748 16128
rect 4510 15106 4566 16127
rect 5678 16119 5748 16127
rect 5174 16075 5260 16079
rect 5174 16019 5186 16075
rect 5242 16019 5260 16075
rect 5174 16007 5260 16019
rect 4685 15862 4731 15873
rect 4900 15871 4976 15904
rect 4900 15825 4911 15871
rect 4965 15825 4976 15871
rect 5084 15871 5160 15904
rect 5084 15825 5095 15871
rect 5149 15825 5160 15871
rect 5268 15871 5344 15904
rect 5268 15825 5279 15871
rect 5333 15825 5344 15871
rect 5513 15862 5559 15873
rect 4823 15779 4869 15790
rect 4806 15752 4823 15754
rect 5007 15779 5053 15790
rect 4869 15752 4886 15754
rect 4731 15632 4818 15752
rect 4874 15632 4886 15752
rect 4806 15630 4823 15632
rect 4731 15332 4823 15452
rect 4869 15630 4886 15632
rect 4990 15452 5007 15454
rect 5191 15779 5237 15790
rect 5174 15752 5191 15754
rect 5375 15779 5421 15790
rect 5237 15752 5254 15754
rect 5174 15632 5186 15752
rect 5242 15632 5254 15752
rect 5174 15630 5191 15632
rect 5053 15452 5070 15454
rect 4990 15332 5002 15452
rect 5058 15332 5070 15452
rect 4990 15330 5007 15332
rect 4823 15294 4869 15305
rect 5053 15330 5070 15332
rect 5007 15294 5053 15305
rect 5237 15630 5254 15632
rect 5358 15452 5375 15454
rect 5496 15752 5513 15754
rect 5559 15752 5576 15754
rect 5496 15631 5508 15752
rect 5564 15631 5576 15752
rect 5496 15629 5513 15631
rect 5421 15452 5438 15454
rect 5358 15332 5370 15452
rect 5426 15332 5438 15452
rect 5358 15330 5375 15332
rect 5191 15294 5237 15305
rect 5421 15330 5438 15332
rect 5375 15294 5421 15305
rect 4900 15256 4911 15259
rect 4965 15256 4976 15259
rect 5084 15256 5095 15259
rect 5149 15256 5160 15259
rect 5268 15256 5279 15259
rect 5333 15256 5344 15259
rect 4685 15211 4731 15222
rect 4898 15200 4910 15256
rect 4966 15200 4978 15256
rect 4898 15186 4978 15200
rect 5082 15200 5094 15256
rect 5150 15200 5162 15256
rect 5082 15186 5162 15200
rect 5266 15200 5278 15256
rect 5334 15200 5346 15256
rect 5559 15629 5576 15631
rect 5513 15211 5559 15222
rect 5266 15186 5346 15200
rect 4898 15106 4978 15108
rect 4510 15050 4910 15106
rect 4966 15050 4978 15106
rect 5996 15106 6052 18332
rect 8547 18329 10094 18385
rect 7558 17308 7628 17320
rect 8547 17308 8603 18329
rect 9216 18277 9302 18281
rect 9216 18221 9228 18277
rect 9284 18221 9302 18277
rect 9216 18209 9302 18221
rect 8727 18064 8773 18075
rect 8942 18073 9018 18106
rect 8942 18027 8953 18073
rect 9007 18027 9018 18073
rect 9126 18073 9202 18106
rect 9126 18027 9137 18073
rect 9191 18027 9202 18073
rect 9310 18073 9386 18106
rect 9310 18027 9321 18073
rect 9375 18027 9386 18073
rect 9555 18064 9601 18075
rect 8865 17981 8911 17992
rect 8848 17954 8865 17956
rect 9049 17981 9095 17992
rect 8911 17954 8928 17956
rect 8773 17834 8860 17954
rect 8916 17834 8928 17954
rect 8848 17832 8865 17834
rect 8773 17534 8865 17654
rect 8911 17832 8928 17834
rect 9032 17654 9049 17656
rect 9233 17981 9279 17992
rect 9216 17954 9233 17956
rect 9417 17981 9463 17992
rect 9279 17954 9296 17956
rect 9216 17834 9228 17954
rect 9284 17834 9296 17954
rect 9216 17832 9233 17834
rect 9095 17654 9112 17656
rect 9032 17534 9044 17654
rect 9100 17534 9112 17654
rect 9032 17532 9049 17534
rect 8865 17496 8911 17507
rect 9095 17532 9112 17534
rect 9049 17496 9095 17507
rect 9279 17832 9296 17834
rect 9400 17654 9417 17656
rect 9538 17954 9555 17956
rect 9601 17954 9618 17956
rect 9538 17833 9550 17954
rect 9606 17833 9618 17954
rect 9538 17831 9555 17833
rect 9463 17654 9480 17656
rect 9400 17534 9412 17654
rect 9468 17534 9480 17654
rect 9400 17532 9417 17534
rect 9233 17496 9279 17507
rect 9463 17532 9480 17534
rect 9417 17496 9463 17507
rect 8942 17458 8953 17461
rect 9007 17458 9018 17461
rect 9126 17458 9137 17461
rect 9191 17458 9202 17461
rect 9310 17458 9321 17461
rect 9375 17458 9386 17461
rect 8727 17413 8773 17424
rect 8940 17402 8952 17458
rect 9008 17402 9020 17458
rect 8940 17388 9020 17402
rect 9124 17402 9136 17458
rect 9192 17402 9204 17458
rect 9124 17388 9204 17402
rect 9308 17402 9320 17458
rect 9376 17402 9388 17458
rect 9601 17831 9618 17833
rect 9555 17413 9601 17424
rect 9308 17388 9388 17402
rect 8940 17308 9020 17310
rect 7558 17252 7570 17308
rect 7626 17252 8952 17308
rect 9008 17252 9020 17308
rect 7558 17250 7628 17252
rect 8940 17250 9020 17252
rect 8268 17192 8338 17204
rect 9124 17192 9204 17194
rect 8268 17136 8280 17192
rect 8336 17136 9136 17192
rect 9192 17136 9204 17192
rect 8268 17124 8338 17136
rect 9124 17134 9204 17136
rect 9453 17192 9533 17194
rect 9720 17192 9790 17204
rect 9453 17136 9465 17192
rect 9521 17136 9722 17192
rect 9778 17136 9790 17192
rect 9453 17134 9533 17136
rect 9720 17126 9790 17136
rect 9308 17076 9388 17078
rect 8552 17020 9320 17076
rect 9376 17020 9388 17076
rect 8552 16289 8608 17020
rect 9308 17018 9388 17020
rect 8940 16926 9020 16940
rect 8727 16904 8773 16915
rect 8940 16870 8952 16926
rect 9008 16870 9020 16926
rect 9124 16926 9204 16940
rect 9124 16870 9136 16926
rect 9192 16870 9204 16926
rect 9308 16926 9388 16940
rect 9308 16870 9320 16926
rect 9376 16870 9388 16926
rect 9555 16904 9601 16915
rect 8942 16867 8953 16870
rect 9007 16867 9018 16870
rect 9126 16867 9137 16870
rect 9191 16867 9202 16870
rect 9310 16867 9321 16870
rect 9375 16867 9386 16870
rect 8865 16821 8911 16832
rect 8773 16647 8865 16821
rect 8865 16636 8911 16647
rect 9049 16821 9095 16832
rect 9049 16636 9095 16647
rect 9233 16821 9279 16832
rect 9417 16821 9463 16832
rect 9400 16794 9417 16796
rect 9463 16794 9480 16796
rect 9400 16674 9412 16794
rect 9468 16674 9480 16794
rect 9400 16672 9417 16674
rect 9233 16636 9279 16647
rect 9463 16672 9480 16674
rect 9417 16636 9463 16647
rect 8727 16419 8773 16564
rect 8942 16555 8953 16601
rect 9007 16555 9018 16601
rect 8942 16522 9018 16555
rect 9126 16555 9137 16601
rect 9191 16555 9202 16601
rect 9126 16522 9202 16555
rect 9310 16555 9321 16601
rect 9375 16555 9386 16601
rect 9310 16522 9386 16555
rect 9555 16419 9601 16564
rect 8715 16407 8795 16419
rect 8715 16351 8727 16407
rect 8783 16351 8795 16407
rect 8715 16339 8795 16351
rect 9533 16407 9613 16419
rect 9533 16351 9545 16407
rect 9601 16351 9613 16407
rect 9533 16339 9613 16351
rect 9886 16289 9966 16299
rect 8552 16233 9898 16289
rect 9954 16233 9966 16289
rect 9886 16231 9966 16233
rect 9720 16180 9790 16182
rect 8552 16179 9790 16180
rect 8552 16125 9722 16179
rect 9778 16125 9790 16179
rect 8552 16124 9790 16125
rect 6660 16075 6746 16079
rect 6660 16019 6672 16075
rect 6728 16019 6746 16075
rect 6660 16007 6746 16019
rect 6171 15862 6217 15873
rect 6386 15871 6462 15904
rect 6386 15825 6397 15871
rect 6451 15825 6462 15871
rect 6570 15871 6646 15904
rect 6570 15825 6581 15871
rect 6635 15825 6646 15871
rect 6754 15871 6830 15904
rect 6754 15825 6765 15871
rect 6819 15825 6830 15871
rect 6999 15862 7045 15873
rect 6309 15779 6355 15790
rect 6292 15752 6309 15754
rect 6493 15779 6539 15790
rect 6355 15752 6372 15754
rect 6217 15632 6304 15752
rect 6360 15632 6372 15752
rect 6292 15630 6309 15632
rect 6217 15332 6309 15452
rect 6355 15630 6372 15632
rect 6476 15452 6493 15454
rect 6677 15779 6723 15790
rect 6660 15752 6677 15754
rect 6861 15779 6907 15790
rect 6723 15752 6740 15754
rect 6660 15632 6672 15752
rect 6728 15632 6740 15752
rect 6660 15630 6677 15632
rect 6539 15452 6556 15454
rect 6476 15332 6488 15452
rect 6544 15332 6556 15452
rect 6476 15330 6493 15332
rect 6309 15294 6355 15305
rect 6539 15330 6556 15332
rect 6493 15294 6539 15305
rect 6723 15630 6740 15632
rect 6844 15452 6861 15454
rect 6982 15752 6999 15754
rect 7045 15752 7062 15754
rect 6982 15631 6994 15752
rect 7050 15631 7062 15752
rect 6982 15629 6999 15631
rect 6907 15452 6924 15454
rect 6844 15332 6856 15452
rect 6912 15332 6924 15452
rect 6844 15330 6861 15332
rect 6677 15294 6723 15305
rect 6907 15330 6924 15332
rect 6861 15294 6907 15305
rect 6386 15256 6397 15259
rect 6451 15256 6462 15259
rect 6570 15256 6581 15259
rect 6635 15256 6646 15259
rect 6754 15256 6765 15259
rect 6819 15256 6830 15259
rect 6171 15211 6217 15222
rect 6384 15200 6396 15256
rect 6452 15200 6464 15256
rect 6384 15186 6464 15200
rect 6568 15200 6580 15256
rect 6636 15200 6648 15256
rect 6568 15186 6648 15200
rect 6752 15200 6764 15256
rect 6820 15200 6832 15256
rect 7045 15629 7062 15631
rect 6999 15211 7045 15222
rect 6752 15186 6832 15200
rect 6384 15106 6464 15108
rect 5996 15050 6396 15106
rect 6452 15050 6464 15106
rect 4898 15048 4978 15050
rect 6384 15048 6464 15050
rect 8552 15103 8608 16124
rect 9720 16116 9790 16124
rect 9216 16072 9302 16076
rect 9216 16016 9228 16072
rect 9284 16016 9302 16072
rect 9216 16004 9302 16016
rect 8727 15859 8773 15870
rect 8942 15868 9018 15901
rect 8942 15822 8953 15868
rect 9007 15822 9018 15868
rect 9126 15868 9202 15901
rect 9126 15822 9137 15868
rect 9191 15822 9202 15868
rect 9310 15868 9386 15901
rect 9310 15822 9321 15868
rect 9375 15822 9386 15868
rect 9555 15859 9601 15870
rect 8865 15776 8911 15787
rect 8848 15749 8865 15751
rect 9049 15776 9095 15787
rect 8911 15749 8928 15751
rect 8773 15629 8860 15749
rect 8916 15629 8928 15749
rect 8848 15627 8865 15629
rect 8773 15329 8865 15449
rect 8911 15627 8928 15629
rect 9032 15449 9049 15451
rect 9233 15776 9279 15787
rect 9216 15749 9233 15751
rect 9417 15776 9463 15787
rect 9279 15749 9296 15751
rect 9216 15629 9228 15749
rect 9284 15629 9296 15749
rect 9216 15627 9233 15629
rect 9095 15449 9112 15451
rect 9032 15329 9044 15449
rect 9100 15329 9112 15449
rect 9032 15327 9049 15329
rect 8865 15291 8911 15302
rect 9095 15327 9112 15329
rect 9049 15291 9095 15302
rect 9279 15627 9296 15629
rect 9400 15449 9417 15451
rect 9538 15749 9555 15751
rect 9601 15749 9618 15751
rect 9538 15628 9550 15749
rect 9606 15628 9618 15749
rect 9538 15626 9555 15628
rect 9463 15449 9480 15451
rect 9400 15329 9412 15449
rect 9468 15329 9480 15449
rect 9400 15327 9417 15329
rect 9233 15291 9279 15302
rect 9463 15327 9480 15329
rect 9417 15291 9463 15302
rect 8942 15253 8953 15256
rect 9007 15253 9018 15256
rect 9126 15253 9137 15256
rect 9191 15253 9202 15256
rect 9310 15253 9321 15256
rect 9375 15253 9386 15256
rect 8727 15208 8773 15219
rect 8940 15197 8952 15253
rect 9008 15197 9020 15253
rect 8940 15183 9020 15197
rect 9124 15197 9136 15253
rect 9192 15197 9204 15253
rect 9124 15183 9204 15197
rect 9308 15197 9320 15253
rect 9376 15197 9388 15253
rect 9601 15626 9618 15628
rect 9555 15208 9601 15219
rect 9308 15183 9388 15197
rect 8940 15103 9020 15105
rect 8552 15047 8952 15103
rect 9008 15047 9020 15103
rect 10038 15103 10094 18329
rect 12589 18329 14136 18385
rect 11600 17308 11670 17320
rect 12589 17308 12645 18329
rect 13258 18277 13344 18281
rect 13258 18221 13270 18277
rect 13326 18221 13344 18277
rect 13258 18209 13344 18221
rect 12769 18064 12815 18075
rect 12984 18073 13060 18106
rect 12984 18027 12995 18073
rect 13049 18027 13060 18073
rect 13168 18073 13244 18106
rect 13168 18027 13179 18073
rect 13233 18027 13244 18073
rect 13352 18073 13428 18106
rect 13352 18027 13363 18073
rect 13417 18027 13428 18073
rect 13597 18064 13643 18075
rect 12907 17981 12953 17992
rect 12890 17954 12907 17956
rect 13091 17981 13137 17992
rect 12953 17954 12970 17956
rect 12815 17834 12902 17954
rect 12958 17834 12970 17954
rect 12890 17832 12907 17834
rect 12815 17534 12907 17654
rect 12953 17832 12970 17834
rect 13074 17654 13091 17656
rect 13275 17981 13321 17992
rect 13258 17954 13275 17956
rect 13459 17981 13505 17992
rect 13321 17954 13338 17956
rect 13258 17834 13270 17954
rect 13326 17834 13338 17954
rect 13258 17832 13275 17834
rect 13137 17654 13154 17656
rect 13074 17534 13086 17654
rect 13142 17534 13154 17654
rect 13074 17532 13091 17534
rect 12907 17496 12953 17507
rect 13137 17532 13154 17534
rect 13091 17496 13137 17507
rect 13321 17832 13338 17834
rect 13442 17654 13459 17656
rect 13580 17954 13597 17956
rect 13643 17954 13660 17956
rect 13580 17833 13592 17954
rect 13648 17833 13660 17954
rect 13580 17831 13597 17833
rect 13505 17654 13522 17656
rect 13442 17534 13454 17654
rect 13510 17534 13522 17654
rect 13442 17532 13459 17534
rect 13275 17496 13321 17507
rect 13505 17532 13522 17534
rect 13459 17496 13505 17507
rect 12984 17458 12995 17461
rect 13049 17458 13060 17461
rect 13168 17458 13179 17461
rect 13233 17458 13244 17461
rect 13352 17458 13363 17461
rect 13417 17458 13428 17461
rect 12769 17413 12815 17424
rect 12982 17402 12994 17458
rect 13050 17402 13062 17458
rect 12982 17388 13062 17402
rect 13166 17402 13178 17458
rect 13234 17402 13246 17458
rect 13166 17388 13246 17402
rect 13350 17402 13362 17458
rect 13418 17402 13430 17458
rect 13643 17831 13660 17833
rect 13597 17413 13643 17424
rect 13350 17388 13430 17402
rect 12982 17308 13062 17310
rect 11600 17252 11612 17308
rect 11668 17252 12994 17308
rect 13050 17252 13062 17308
rect 11600 17250 11670 17252
rect 12982 17250 13062 17252
rect 12310 17192 12380 17204
rect 13166 17192 13246 17194
rect 12310 17136 12322 17192
rect 12378 17136 13178 17192
rect 13234 17136 13246 17192
rect 12310 17124 12380 17136
rect 13166 17134 13246 17136
rect 13495 17192 13575 17194
rect 13762 17192 13832 17204
rect 13495 17136 13507 17192
rect 13563 17136 13764 17192
rect 13820 17136 13832 17192
rect 13495 17134 13575 17136
rect 13762 17126 13832 17136
rect 13350 17076 13430 17078
rect 12594 17020 13362 17076
rect 13418 17020 13430 17076
rect 12594 16289 12650 17020
rect 13350 17018 13430 17020
rect 12982 16926 13062 16940
rect 12769 16904 12815 16915
rect 12982 16870 12994 16926
rect 13050 16870 13062 16926
rect 13166 16926 13246 16940
rect 13166 16870 13178 16926
rect 13234 16870 13246 16926
rect 13350 16926 13430 16940
rect 13350 16870 13362 16926
rect 13418 16870 13430 16926
rect 13597 16904 13643 16915
rect 12984 16867 12995 16870
rect 13049 16867 13060 16870
rect 13168 16867 13179 16870
rect 13233 16867 13244 16870
rect 13352 16867 13363 16870
rect 13417 16867 13428 16870
rect 12907 16821 12953 16832
rect 12815 16647 12907 16821
rect 12907 16636 12953 16647
rect 13091 16821 13137 16832
rect 13091 16636 13137 16647
rect 13275 16821 13321 16832
rect 13459 16821 13505 16832
rect 13442 16794 13459 16796
rect 13505 16794 13522 16796
rect 13442 16674 13454 16794
rect 13510 16674 13522 16794
rect 13442 16672 13459 16674
rect 13275 16636 13321 16647
rect 13505 16672 13522 16674
rect 13459 16636 13505 16647
rect 12769 16419 12815 16564
rect 12984 16555 12995 16601
rect 13049 16555 13060 16601
rect 12984 16522 13060 16555
rect 13168 16555 13179 16601
rect 13233 16555 13244 16601
rect 13168 16522 13244 16555
rect 13352 16555 13363 16601
rect 13417 16555 13428 16601
rect 13352 16522 13428 16555
rect 13597 16419 13643 16564
rect 12757 16407 12837 16419
rect 12757 16351 12769 16407
rect 12825 16351 12837 16407
rect 12757 16339 12837 16351
rect 13575 16407 13655 16419
rect 13575 16351 13587 16407
rect 13643 16351 13655 16407
rect 13575 16339 13655 16351
rect 13928 16289 14008 16299
rect 12594 16233 13940 16289
rect 13996 16233 14008 16289
rect 13928 16231 14008 16233
rect 13762 16180 13832 16182
rect 12594 16179 13832 16180
rect 12594 16125 13764 16179
rect 13820 16125 13832 16179
rect 12594 16124 13832 16125
rect 10702 16072 10788 16076
rect 10702 16016 10714 16072
rect 10770 16016 10788 16072
rect 10702 16004 10788 16016
rect 10213 15859 10259 15870
rect 10428 15868 10504 15901
rect 10428 15822 10439 15868
rect 10493 15822 10504 15868
rect 10612 15868 10688 15901
rect 10612 15822 10623 15868
rect 10677 15822 10688 15868
rect 10796 15868 10872 15901
rect 10796 15822 10807 15868
rect 10861 15822 10872 15868
rect 11041 15859 11087 15870
rect 10351 15776 10397 15787
rect 10334 15749 10351 15751
rect 10535 15776 10581 15787
rect 10397 15749 10414 15751
rect 10259 15629 10346 15749
rect 10402 15629 10414 15749
rect 10334 15627 10351 15629
rect 10259 15329 10351 15449
rect 10397 15627 10414 15629
rect 10518 15449 10535 15451
rect 10719 15776 10765 15787
rect 10702 15749 10719 15751
rect 10903 15776 10949 15787
rect 10765 15749 10782 15751
rect 10702 15629 10714 15749
rect 10770 15629 10782 15749
rect 10702 15627 10719 15629
rect 10581 15449 10598 15451
rect 10518 15329 10530 15449
rect 10586 15329 10598 15449
rect 10518 15327 10535 15329
rect 10351 15291 10397 15302
rect 10581 15327 10598 15329
rect 10535 15291 10581 15302
rect 10765 15627 10782 15629
rect 10886 15449 10903 15451
rect 11024 15749 11041 15751
rect 11087 15749 11104 15751
rect 11024 15628 11036 15749
rect 11092 15628 11104 15749
rect 11024 15626 11041 15628
rect 10949 15449 10966 15451
rect 10886 15329 10898 15449
rect 10954 15329 10966 15449
rect 10886 15327 10903 15329
rect 10719 15291 10765 15302
rect 10949 15327 10966 15329
rect 10903 15291 10949 15302
rect 10428 15253 10439 15256
rect 10493 15253 10504 15256
rect 10612 15253 10623 15256
rect 10677 15253 10688 15256
rect 10796 15253 10807 15256
rect 10861 15253 10872 15256
rect 10213 15208 10259 15219
rect 10426 15197 10438 15253
rect 10494 15197 10506 15253
rect 10426 15183 10506 15197
rect 10610 15197 10622 15253
rect 10678 15197 10690 15253
rect 10610 15183 10690 15197
rect 10794 15197 10806 15253
rect 10862 15197 10874 15253
rect 11087 15626 11104 15628
rect 11041 15208 11087 15219
rect 10794 15183 10874 15197
rect 10426 15103 10506 15105
rect 10038 15047 10438 15103
rect 10494 15047 10506 15103
rect 12594 15103 12650 16124
rect 13762 16116 13832 16124
rect 13258 16072 13344 16076
rect 13258 16016 13270 16072
rect 13326 16016 13344 16072
rect 13258 16004 13344 16016
rect 12769 15859 12815 15870
rect 12984 15868 13060 15901
rect 12984 15822 12995 15868
rect 13049 15822 13060 15868
rect 13168 15868 13244 15901
rect 13168 15822 13179 15868
rect 13233 15822 13244 15868
rect 13352 15868 13428 15901
rect 13352 15822 13363 15868
rect 13417 15822 13428 15868
rect 13597 15859 13643 15870
rect 12907 15776 12953 15787
rect 12890 15749 12907 15751
rect 13091 15776 13137 15787
rect 12953 15749 12970 15751
rect 12815 15629 12902 15749
rect 12958 15629 12970 15749
rect 12890 15627 12907 15629
rect 12815 15329 12907 15449
rect 12953 15627 12970 15629
rect 13074 15449 13091 15451
rect 13275 15776 13321 15787
rect 13258 15749 13275 15751
rect 13459 15776 13505 15787
rect 13321 15749 13338 15751
rect 13258 15629 13270 15749
rect 13326 15629 13338 15749
rect 13258 15627 13275 15629
rect 13137 15449 13154 15451
rect 13074 15329 13086 15449
rect 13142 15329 13154 15449
rect 13074 15327 13091 15329
rect 12907 15291 12953 15302
rect 13137 15327 13154 15329
rect 13091 15291 13137 15302
rect 13321 15627 13338 15629
rect 13442 15449 13459 15451
rect 13580 15749 13597 15751
rect 13643 15749 13660 15751
rect 13580 15628 13592 15749
rect 13648 15628 13660 15749
rect 13580 15626 13597 15628
rect 13505 15449 13522 15451
rect 13442 15329 13454 15449
rect 13510 15329 13522 15449
rect 13442 15327 13459 15329
rect 13275 15291 13321 15302
rect 13505 15327 13522 15329
rect 13459 15291 13505 15302
rect 12984 15253 12995 15256
rect 13049 15253 13060 15256
rect 13168 15253 13179 15256
rect 13233 15253 13244 15256
rect 13352 15253 13363 15256
rect 13417 15253 13428 15256
rect 12769 15208 12815 15219
rect 12982 15197 12994 15253
rect 13050 15197 13062 15253
rect 12982 15183 13062 15197
rect 13166 15197 13178 15253
rect 13234 15197 13246 15253
rect 13166 15183 13246 15197
rect 13350 15197 13362 15253
rect 13418 15197 13430 15253
rect 13643 15626 13660 15628
rect 13597 15208 13643 15219
rect 13350 15183 13430 15197
rect 12982 15103 13062 15105
rect 12594 15047 12994 15103
rect 13050 15047 13062 15103
rect 14080 15103 14136 18329
rect 16631 18329 18178 18385
rect 15642 17308 15712 17320
rect 16631 17308 16687 18329
rect 17300 18277 17386 18281
rect 17300 18221 17312 18277
rect 17368 18221 17386 18277
rect 17300 18209 17386 18221
rect 16811 18064 16857 18075
rect 17026 18073 17102 18106
rect 17026 18027 17037 18073
rect 17091 18027 17102 18073
rect 17210 18073 17286 18106
rect 17210 18027 17221 18073
rect 17275 18027 17286 18073
rect 17394 18073 17470 18106
rect 17394 18027 17405 18073
rect 17459 18027 17470 18073
rect 17639 18064 17685 18075
rect 16949 17981 16995 17992
rect 16932 17954 16949 17956
rect 17133 17981 17179 17992
rect 16995 17954 17012 17956
rect 16857 17834 16944 17954
rect 17000 17834 17012 17954
rect 16932 17832 16949 17834
rect 16857 17534 16949 17654
rect 16995 17832 17012 17834
rect 17116 17654 17133 17656
rect 17317 17981 17363 17992
rect 17300 17954 17317 17956
rect 17501 17981 17547 17992
rect 17363 17954 17380 17956
rect 17300 17834 17312 17954
rect 17368 17834 17380 17954
rect 17300 17832 17317 17834
rect 17179 17654 17196 17656
rect 17116 17534 17128 17654
rect 17184 17534 17196 17654
rect 17116 17532 17133 17534
rect 16949 17496 16995 17507
rect 17179 17532 17196 17534
rect 17133 17496 17179 17507
rect 17363 17832 17380 17834
rect 17484 17654 17501 17656
rect 17622 17954 17639 17956
rect 17685 17954 17702 17956
rect 17622 17833 17634 17954
rect 17690 17833 17702 17954
rect 17622 17831 17639 17833
rect 17547 17654 17564 17656
rect 17484 17534 17496 17654
rect 17552 17534 17564 17654
rect 17484 17532 17501 17534
rect 17317 17496 17363 17507
rect 17547 17532 17564 17534
rect 17501 17496 17547 17507
rect 17026 17458 17037 17461
rect 17091 17458 17102 17461
rect 17210 17458 17221 17461
rect 17275 17458 17286 17461
rect 17394 17458 17405 17461
rect 17459 17458 17470 17461
rect 16811 17413 16857 17424
rect 17024 17402 17036 17458
rect 17092 17402 17104 17458
rect 17024 17388 17104 17402
rect 17208 17402 17220 17458
rect 17276 17402 17288 17458
rect 17208 17388 17288 17402
rect 17392 17402 17404 17458
rect 17460 17402 17472 17458
rect 17685 17831 17702 17833
rect 17639 17413 17685 17424
rect 17392 17388 17472 17402
rect 17024 17308 17104 17310
rect 15642 17252 15654 17308
rect 15710 17252 17036 17308
rect 17092 17252 17104 17308
rect 15642 17250 15712 17252
rect 17024 17250 17104 17252
rect 16352 17192 16422 17204
rect 17208 17192 17288 17194
rect 16352 17136 16364 17192
rect 16420 17136 17220 17192
rect 17276 17136 17288 17192
rect 16352 17124 16422 17136
rect 17208 17134 17288 17136
rect 17537 17192 17617 17194
rect 17804 17192 17874 17204
rect 17537 17136 17549 17192
rect 17605 17136 17806 17192
rect 17862 17136 17874 17192
rect 17537 17134 17617 17136
rect 17804 17126 17874 17136
rect 17392 17076 17472 17078
rect 16636 17020 17404 17076
rect 17460 17020 17472 17076
rect 16636 16289 16692 17020
rect 17392 17018 17472 17020
rect 17024 16926 17104 16940
rect 16811 16904 16857 16915
rect 17024 16870 17036 16926
rect 17092 16870 17104 16926
rect 17208 16926 17288 16940
rect 17208 16870 17220 16926
rect 17276 16870 17288 16926
rect 17392 16926 17472 16940
rect 17392 16870 17404 16926
rect 17460 16870 17472 16926
rect 17639 16904 17685 16915
rect 17026 16867 17037 16870
rect 17091 16867 17102 16870
rect 17210 16867 17221 16870
rect 17275 16867 17286 16870
rect 17394 16867 17405 16870
rect 17459 16867 17470 16870
rect 16949 16821 16995 16832
rect 16857 16647 16949 16821
rect 16949 16636 16995 16647
rect 17133 16821 17179 16832
rect 17133 16636 17179 16647
rect 17317 16821 17363 16832
rect 17501 16821 17547 16832
rect 17484 16794 17501 16796
rect 17547 16794 17564 16796
rect 17484 16674 17496 16794
rect 17552 16674 17564 16794
rect 17484 16672 17501 16674
rect 17317 16636 17363 16647
rect 17547 16672 17564 16674
rect 17501 16636 17547 16647
rect 16811 16419 16857 16564
rect 17026 16555 17037 16601
rect 17091 16555 17102 16601
rect 17026 16522 17102 16555
rect 17210 16555 17221 16601
rect 17275 16555 17286 16601
rect 17210 16522 17286 16555
rect 17394 16555 17405 16601
rect 17459 16555 17470 16601
rect 17394 16522 17470 16555
rect 17639 16419 17685 16564
rect 16799 16407 16879 16419
rect 16799 16351 16811 16407
rect 16867 16351 16879 16407
rect 16799 16339 16879 16351
rect 17617 16407 17697 16419
rect 17617 16351 17629 16407
rect 17685 16351 17697 16407
rect 17617 16339 17697 16351
rect 17970 16289 18050 16299
rect 16636 16233 17982 16289
rect 18038 16233 18050 16289
rect 17970 16231 18050 16233
rect 17804 16180 17874 16182
rect 16636 16179 17874 16180
rect 16636 16125 17806 16179
rect 17862 16125 17874 16179
rect 16636 16124 17874 16125
rect 14744 16072 14830 16076
rect 14744 16016 14756 16072
rect 14812 16016 14830 16072
rect 14744 16004 14830 16016
rect 14255 15859 14301 15870
rect 14470 15868 14546 15901
rect 14470 15822 14481 15868
rect 14535 15822 14546 15868
rect 14654 15868 14730 15901
rect 14654 15822 14665 15868
rect 14719 15822 14730 15868
rect 14838 15868 14914 15901
rect 14838 15822 14849 15868
rect 14903 15822 14914 15868
rect 15083 15859 15129 15870
rect 14393 15776 14439 15787
rect 14376 15749 14393 15751
rect 14577 15776 14623 15787
rect 14439 15749 14456 15751
rect 14301 15629 14388 15749
rect 14444 15629 14456 15749
rect 14376 15627 14393 15629
rect 14301 15329 14393 15449
rect 14439 15627 14456 15629
rect 14560 15449 14577 15451
rect 14761 15776 14807 15787
rect 14744 15749 14761 15751
rect 14945 15776 14991 15787
rect 14807 15749 14824 15751
rect 14744 15629 14756 15749
rect 14812 15629 14824 15749
rect 14744 15627 14761 15629
rect 14623 15449 14640 15451
rect 14560 15329 14572 15449
rect 14628 15329 14640 15449
rect 14560 15327 14577 15329
rect 14393 15291 14439 15302
rect 14623 15327 14640 15329
rect 14577 15291 14623 15302
rect 14807 15627 14824 15629
rect 14928 15449 14945 15451
rect 15066 15749 15083 15751
rect 15129 15749 15146 15751
rect 15066 15628 15078 15749
rect 15134 15628 15146 15749
rect 15066 15626 15083 15628
rect 14991 15449 15008 15451
rect 14928 15329 14940 15449
rect 14996 15329 15008 15449
rect 14928 15327 14945 15329
rect 14761 15291 14807 15302
rect 14991 15327 15008 15329
rect 14945 15291 14991 15302
rect 14470 15253 14481 15256
rect 14535 15253 14546 15256
rect 14654 15253 14665 15256
rect 14719 15253 14730 15256
rect 14838 15253 14849 15256
rect 14903 15253 14914 15256
rect 14255 15208 14301 15219
rect 14468 15197 14480 15253
rect 14536 15197 14548 15253
rect 14468 15183 14548 15197
rect 14652 15197 14664 15253
rect 14720 15197 14732 15253
rect 14652 15183 14732 15197
rect 14836 15197 14848 15253
rect 14904 15197 14916 15253
rect 15129 15626 15146 15628
rect 15083 15208 15129 15219
rect 14836 15183 14916 15197
rect 14468 15103 14548 15105
rect 14080 15047 14480 15103
rect 14536 15047 14548 15103
rect 16636 15103 16692 16124
rect 17804 16116 17874 16124
rect 17300 16072 17386 16076
rect 17300 16016 17312 16072
rect 17368 16016 17386 16072
rect 17300 16004 17386 16016
rect 16811 15859 16857 15870
rect 17026 15868 17102 15901
rect 17026 15822 17037 15868
rect 17091 15822 17102 15868
rect 17210 15868 17286 15901
rect 17210 15822 17221 15868
rect 17275 15822 17286 15868
rect 17394 15868 17470 15901
rect 17394 15822 17405 15868
rect 17459 15822 17470 15868
rect 17639 15859 17685 15870
rect 16949 15776 16995 15787
rect 16932 15749 16949 15751
rect 17133 15776 17179 15787
rect 16995 15749 17012 15751
rect 16857 15629 16944 15749
rect 17000 15629 17012 15749
rect 16932 15627 16949 15629
rect 16857 15329 16949 15449
rect 16995 15627 17012 15629
rect 17116 15449 17133 15451
rect 17317 15776 17363 15787
rect 17300 15749 17317 15751
rect 17501 15776 17547 15787
rect 17363 15749 17380 15751
rect 17300 15629 17312 15749
rect 17368 15629 17380 15749
rect 17300 15627 17317 15629
rect 17179 15449 17196 15451
rect 17116 15329 17128 15449
rect 17184 15329 17196 15449
rect 17116 15327 17133 15329
rect 16949 15291 16995 15302
rect 17179 15327 17196 15329
rect 17133 15291 17179 15302
rect 17363 15627 17380 15629
rect 17484 15449 17501 15451
rect 17622 15749 17639 15751
rect 17685 15749 17702 15751
rect 17622 15628 17634 15749
rect 17690 15628 17702 15749
rect 17622 15626 17639 15628
rect 17547 15449 17564 15451
rect 17484 15329 17496 15449
rect 17552 15329 17564 15449
rect 17484 15327 17501 15329
rect 17317 15291 17363 15302
rect 17547 15327 17564 15329
rect 17501 15291 17547 15302
rect 17026 15253 17037 15256
rect 17091 15253 17102 15256
rect 17210 15253 17221 15256
rect 17275 15253 17286 15256
rect 17394 15253 17405 15256
rect 17459 15253 17470 15256
rect 16811 15208 16857 15219
rect 17024 15197 17036 15253
rect 17092 15197 17104 15253
rect 17024 15183 17104 15197
rect 17208 15197 17220 15253
rect 17276 15197 17288 15253
rect 17208 15183 17288 15197
rect 17392 15197 17404 15253
rect 17460 15197 17472 15253
rect 17685 15626 17702 15628
rect 17639 15208 17685 15219
rect 17392 15183 17472 15197
rect 17024 15103 17104 15105
rect 16636 15047 17036 15103
rect 17092 15047 17104 15103
rect 18122 15103 18178 18329
rect 20673 18329 22220 18385
rect 19684 17308 19754 17320
rect 20673 17308 20729 18329
rect 21342 18277 21428 18281
rect 21342 18221 21354 18277
rect 21410 18221 21428 18277
rect 21342 18209 21428 18221
rect 20853 18064 20899 18075
rect 21068 18073 21144 18106
rect 21068 18027 21079 18073
rect 21133 18027 21144 18073
rect 21252 18073 21328 18106
rect 21252 18027 21263 18073
rect 21317 18027 21328 18073
rect 21436 18073 21512 18106
rect 21436 18027 21447 18073
rect 21501 18027 21512 18073
rect 21681 18064 21727 18075
rect 20991 17981 21037 17992
rect 20974 17954 20991 17956
rect 21175 17981 21221 17992
rect 21037 17954 21054 17956
rect 20899 17834 20986 17954
rect 21042 17834 21054 17954
rect 20974 17832 20991 17834
rect 20899 17534 20991 17654
rect 21037 17832 21054 17834
rect 21158 17654 21175 17656
rect 21359 17981 21405 17992
rect 21342 17954 21359 17956
rect 21543 17981 21589 17992
rect 21405 17954 21422 17956
rect 21342 17834 21354 17954
rect 21410 17834 21422 17954
rect 21342 17832 21359 17834
rect 21221 17654 21238 17656
rect 21158 17534 21170 17654
rect 21226 17534 21238 17654
rect 21158 17532 21175 17534
rect 20991 17496 21037 17507
rect 21221 17532 21238 17534
rect 21175 17496 21221 17507
rect 21405 17832 21422 17834
rect 21526 17654 21543 17656
rect 21664 17954 21681 17956
rect 21727 17954 21744 17956
rect 21664 17833 21676 17954
rect 21732 17833 21744 17954
rect 21664 17831 21681 17833
rect 21589 17654 21606 17656
rect 21526 17534 21538 17654
rect 21594 17534 21606 17654
rect 21526 17532 21543 17534
rect 21359 17496 21405 17507
rect 21589 17532 21606 17534
rect 21543 17496 21589 17507
rect 21068 17458 21079 17461
rect 21133 17458 21144 17461
rect 21252 17458 21263 17461
rect 21317 17458 21328 17461
rect 21436 17458 21447 17461
rect 21501 17458 21512 17461
rect 20853 17413 20899 17424
rect 21066 17402 21078 17458
rect 21134 17402 21146 17458
rect 21066 17388 21146 17402
rect 21250 17402 21262 17458
rect 21318 17402 21330 17458
rect 21250 17388 21330 17402
rect 21434 17402 21446 17458
rect 21502 17402 21514 17458
rect 21727 17831 21744 17833
rect 21681 17413 21727 17424
rect 21434 17388 21514 17402
rect 21066 17308 21146 17310
rect 19684 17252 19696 17308
rect 19752 17252 21078 17308
rect 21134 17252 21146 17308
rect 19684 17250 19754 17252
rect 21066 17250 21146 17252
rect 20394 17192 20464 17204
rect 21250 17192 21330 17194
rect 20394 17136 20406 17192
rect 20462 17136 21262 17192
rect 21318 17136 21330 17192
rect 20394 17124 20464 17136
rect 21250 17134 21330 17136
rect 21579 17192 21659 17194
rect 21846 17192 21916 17204
rect 21579 17136 21591 17192
rect 21647 17136 21848 17192
rect 21904 17136 21916 17192
rect 21579 17134 21659 17136
rect 21846 17126 21916 17136
rect 21434 17076 21514 17078
rect 20678 17020 21446 17076
rect 21502 17020 21514 17076
rect 20678 16289 20734 17020
rect 21434 17018 21514 17020
rect 21066 16926 21146 16940
rect 20853 16904 20899 16915
rect 21066 16870 21078 16926
rect 21134 16870 21146 16926
rect 21250 16926 21330 16940
rect 21250 16870 21262 16926
rect 21318 16870 21330 16926
rect 21434 16926 21514 16940
rect 21434 16870 21446 16926
rect 21502 16870 21514 16926
rect 21681 16904 21727 16915
rect 21068 16867 21079 16870
rect 21133 16867 21144 16870
rect 21252 16867 21263 16870
rect 21317 16867 21328 16870
rect 21436 16867 21447 16870
rect 21501 16867 21512 16870
rect 20991 16821 21037 16832
rect 20899 16647 20991 16821
rect 20991 16636 21037 16647
rect 21175 16821 21221 16832
rect 21175 16636 21221 16647
rect 21359 16821 21405 16832
rect 21543 16821 21589 16832
rect 21526 16794 21543 16796
rect 21589 16794 21606 16796
rect 21526 16674 21538 16794
rect 21594 16674 21606 16794
rect 21526 16672 21543 16674
rect 21359 16636 21405 16647
rect 21589 16672 21606 16674
rect 21543 16636 21589 16647
rect 20853 16419 20899 16564
rect 21068 16555 21079 16601
rect 21133 16555 21144 16601
rect 21068 16522 21144 16555
rect 21252 16555 21263 16601
rect 21317 16555 21328 16601
rect 21252 16522 21328 16555
rect 21436 16555 21447 16601
rect 21501 16555 21512 16601
rect 21436 16522 21512 16555
rect 21681 16419 21727 16564
rect 20841 16407 20921 16419
rect 20841 16351 20853 16407
rect 20909 16351 20921 16407
rect 20841 16339 20921 16351
rect 21659 16407 21739 16419
rect 21659 16351 21671 16407
rect 21727 16351 21739 16407
rect 21659 16339 21739 16351
rect 22012 16289 22092 16299
rect 20678 16233 22024 16289
rect 22080 16233 22092 16289
rect 22012 16231 22092 16233
rect 21846 16180 21916 16182
rect 20678 16179 21916 16180
rect 20678 16125 21848 16179
rect 21904 16125 21916 16179
rect 20678 16124 21916 16125
rect 18786 16072 18872 16076
rect 18786 16016 18798 16072
rect 18854 16016 18872 16072
rect 18786 16004 18872 16016
rect 18297 15859 18343 15870
rect 18512 15868 18588 15901
rect 18512 15822 18523 15868
rect 18577 15822 18588 15868
rect 18696 15868 18772 15901
rect 18696 15822 18707 15868
rect 18761 15822 18772 15868
rect 18880 15868 18956 15901
rect 18880 15822 18891 15868
rect 18945 15822 18956 15868
rect 19125 15859 19171 15870
rect 18435 15776 18481 15787
rect 18418 15749 18435 15751
rect 18619 15776 18665 15787
rect 18481 15749 18498 15751
rect 18343 15629 18430 15749
rect 18486 15629 18498 15749
rect 18418 15627 18435 15629
rect 18343 15329 18435 15449
rect 18481 15627 18498 15629
rect 18602 15449 18619 15451
rect 18803 15776 18849 15787
rect 18786 15749 18803 15751
rect 18987 15776 19033 15787
rect 18849 15749 18866 15751
rect 18786 15629 18798 15749
rect 18854 15629 18866 15749
rect 18786 15627 18803 15629
rect 18665 15449 18682 15451
rect 18602 15329 18614 15449
rect 18670 15329 18682 15449
rect 18602 15327 18619 15329
rect 18435 15291 18481 15302
rect 18665 15327 18682 15329
rect 18619 15291 18665 15302
rect 18849 15627 18866 15629
rect 18970 15449 18987 15451
rect 19108 15749 19125 15751
rect 19171 15749 19188 15751
rect 19108 15628 19120 15749
rect 19176 15628 19188 15749
rect 19108 15626 19125 15628
rect 19033 15449 19050 15451
rect 18970 15329 18982 15449
rect 19038 15329 19050 15449
rect 18970 15327 18987 15329
rect 18803 15291 18849 15302
rect 19033 15327 19050 15329
rect 18987 15291 19033 15302
rect 18512 15253 18523 15256
rect 18577 15253 18588 15256
rect 18696 15253 18707 15256
rect 18761 15253 18772 15256
rect 18880 15253 18891 15256
rect 18945 15253 18956 15256
rect 18297 15208 18343 15219
rect 18510 15197 18522 15253
rect 18578 15197 18590 15253
rect 18510 15183 18590 15197
rect 18694 15197 18706 15253
rect 18762 15197 18774 15253
rect 18694 15183 18774 15197
rect 18878 15197 18890 15253
rect 18946 15197 18958 15253
rect 19171 15626 19188 15628
rect 19125 15208 19171 15219
rect 18878 15183 18958 15197
rect 18510 15103 18590 15105
rect 18122 15047 18522 15103
rect 18578 15047 18590 15103
rect 20678 15103 20734 16124
rect 21846 16116 21916 16124
rect 21342 16072 21428 16076
rect 21342 16016 21354 16072
rect 21410 16016 21428 16072
rect 21342 16004 21428 16016
rect 20853 15859 20899 15870
rect 21068 15868 21144 15901
rect 21068 15822 21079 15868
rect 21133 15822 21144 15868
rect 21252 15868 21328 15901
rect 21252 15822 21263 15868
rect 21317 15822 21328 15868
rect 21436 15868 21512 15901
rect 21436 15822 21447 15868
rect 21501 15822 21512 15868
rect 21681 15859 21727 15870
rect 20991 15776 21037 15787
rect 20974 15749 20991 15751
rect 21175 15776 21221 15787
rect 21037 15749 21054 15751
rect 20899 15629 20986 15749
rect 21042 15629 21054 15749
rect 20974 15627 20991 15629
rect 20899 15329 20991 15449
rect 21037 15627 21054 15629
rect 21158 15449 21175 15451
rect 21359 15776 21405 15787
rect 21342 15749 21359 15751
rect 21543 15776 21589 15787
rect 21405 15749 21422 15751
rect 21342 15629 21354 15749
rect 21410 15629 21422 15749
rect 21342 15627 21359 15629
rect 21221 15449 21238 15451
rect 21158 15329 21170 15449
rect 21226 15329 21238 15449
rect 21158 15327 21175 15329
rect 20991 15291 21037 15302
rect 21221 15327 21238 15329
rect 21175 15291 21221 15302
rect 21405 15627 21422 15629
rect 21526 15449 21543 15451
rect 21664 15749 21681 15751
rect 21727 15749 21744 15751
rect 21664 15628 21676 15749
rect 21732 15628 21744 15749
rect 21664 15626 21681 15628
rect 21589 15449 21606 15451
rect 21526 15329 21538 15449
rect 21594 15329 21606 15449
rect 21526 15327 21543 15329
rect 21359 15291 21405 15302
rect 21589 15327 21606 15329
rect 21543 15291 21589 15302
rect 21068 15253 21079 15256
rect 21133 15253 21144 15256
rect 21252 15253 21263 15256
rect 21317 15253 21328 15256
rect 21436 15253 21447 15256
rect 21501 15253 21512 15256
rect 20853 15208 20899 15219
rect 21066 15197 21078 15253
rect 21134 15197 21146 15253
rect 21066 15183 21146 15197
rect 21250 15197 21262 15253
rect 21318 15197 21330 15253
rect 21250 15183 21330 15197
rect 21434 15197 21446 15253
rect 21502 15197 21514 15253
rect 21727 15626 21744 15628
rect 21681 15208 21727 15219
rect 21434 15183 21514 15197
rect 21066 15103 21146 15105
rect 20678 15047 21078 15103
rect 21134 15047 21146 15103
rect 22164 15103 22220 18329
rect 24715 18329 26262 18385
rect 23726 17308 23796 17320
rect 24715 17308 24771 18329
rect 25384 18277 25470 18281
rect 25384 18221 25396 18277
rect 25452 18221 25470 18277
rect 25384 18209 25470 18221
rect 24895 18064 24941 18075
rect 25110 18073 25186 18106
rect 25110 18027 25121 18073
rect 25175 18027 25186 18073
rect 25294 18073 25370 18106
rect 25294 18027 25305 18073
rect 25359 18027 25370 18073
rect 25478 18073 25554 18106
rect 25478 18027 25489 18073
rect 25543 18027 25554 18073
rect 25723 18064 25769 18075
rect 25033 17981 25079 17992
rect 25016 17954 25033 17956
rect 25217 17981 25263 17992
rect 25079 17954 25096 17956
rect 24941 17834 25028 17954
rect 25084 17834 25096 17954
rect 25016 17832 25033 17834
rect 24941 17534 25033 17654
rect 25079 17832 25096 17834
rect 25200 17654 25217 17656
rect 25401 17981 25447 17992
rect 25384 17954 25401 17956
rect 25585 17981 25631 17992
rect 25447 17954 25464 17956
rect 25384 17834 25396 17954
rect 25452 17834 25464 17954
rect 25384 17832 25401 17834
rect 25263 17654 25280 17656
rect 25200 17534 25212 17654
rect 25268 17534 25280 17654
rect 25200 17532 25217 17534
rect 25033 17496 25079 17507
rect 25263 17532 25280 17534
rect 25217 17496 25263 17507
rect 25447 17832 25464 17834
rect 25568 17654 25585 17656
rect 25706 17954 25723 17956
rect 25769 17954 25786 17956
rect 25706 17833 25718 17954
rect 25774 17833 25786 17954
rect 25706 17831 25723 17833
rect 25631 17654 25648 17656
rect 25568 17534 25580 17654
rect 25636 17534 25648 17654
rect 25568 17532 25585 17534
rect 25401 17496 25447 17507
rect 25631 17532 25648 17534
rect 25585 17496 25631 17507
rect 25110 17458 25121 17461
rect 25175 17458 25186 17461
rect 25294 17458 25305 17461
rect 25359 17458 25370 17461
rect 25478 17458 25489 17461
rect 25543 17458 25554 17461
rect 24895 17413 24941 17424
rect 25108 17402 25120 17458
rect 25176 17402 25188 17458
rect 25108 17388 25188 17402
rect 25292 17402 25304 17458
rect 25360 17402 25372 17458
rect 25292 17388 25372 17402
rect 25476 17402 25488 17458
rect 25544 17402 25556 17458
rect 25769 17831 25786 17833
rect 25723 17413 25769 17424
rect 25476 17388 25556 17402
rect 25108 17308 25188 17310
rect 23726 17252 23738 17308
rect 23794 17252 25120 17308
rect 25176 17252 25188 17308
rect 23726 17250 23796 17252
rect 25108 17250 25188 17252
rect 24436 17192 24506 17204
rect 25292 17192 25372 17194
rect 24436 17136 24448 17192
rect 24504 17136 25304 17192
rect 25360 17136 25372 17192
rect 24436 17124 24506 17136
rect 25292 17134 25372 17136
rect 25621 17192 25701 17194
rect 25888 17192 25958 17204
rect 25621 17136 25633 17192
rect 25689 17136 25890 17192
rect 25946 17136 25958 17192
rect 25621 17134 25701 17136
rect 25888 17126 25958 17136
rect 25476 17076 25556 17078
rect 24720 17020 25488 17076
rect 25544 17020 25556 17076
rect 24720 16289 24776 17020
rect 25476 17018 25556 17020
rect 25108 16926 25188 16940
rect 24895 16904 24941 16915
rect 25108 16870 25120 16926
rect 25176 16870 25188 16926
rect 25292 16926 25372 16940
rect 25292 16870 25304 16926
rect 25360 16870 25372 16926
rect 25476 16926 25556 16940
rect 25476 16870 25488 16926
rect 25544 16870 25556 16926
rect 25723 16904 25769 16915
rect 25110 16867 25121 16870
rect 25175 16867 25186 16870
rect 25294 16867 25305 16870
rect 25359 16867 25370 16870
rect 25478 16867 25489 16870
rect 25543 16867 25554 16870
rect 25033 16821 25079 16832
rect 24941 16647 25033 16821
rect 25033 16636 25079 16647
rect 25217 16821 25263 16832
rect 25217 16636 25263 16647
rect 25401 16821 25447 16832
rect 25585 16821 25631 16832
rect 25568 16794 25585 16796
rect 25631 16794 25648 16796
rect 25568 16674 25580 16794
rect 25636 16674 25648 16794
rect 25568 16672 25585 16674
rect 25401 16636 25447 16647
rect 25631 16672 25648 16674
rect 25585 16636 25631 16647
rect 24895 16419 24941 16564
rect 25110 16555 25121 16601
rect 25175 16555 25186 16601
rect 25110 16522 25186 16555
rect 25294 16555 25305 16601
rect 25359 16555 25370 16601
rect 25294 16522 25370 16555
rect 25478 16555 25489 16601
rect 25543 16555 25554 16601
rect 25478 16522 25554 16555
rect 25723 16419 25769 16564
rect 24883 16407 24963 16419
rect 24883 16351 24895 16407
rect 24951 16351 24963 16407
rect 24883 16339 24963 16351
rect 25701 16407 25781 16419
rect 25701 16351 25713 16407
rect 25769 16351 25781 16407
rect 25701 16339 25781 16351
rect 26054 16289 26134 16299
rect 24720 16233 26066 16289
rect 26122 16233 26134 16289
rect 26054 16231 26134 16233
rect 25888 16180 25958 16182
rect 24720 16179 25958 16180
rect 24720 16125 25890 16179
rect 25946 16125 25958 16179
rect 24720 16124 25958 16125
rect 22828 16072 22914 16076
rect 22828 16016 22840 16072
rect 22896 16016 22914 16072
rect 22828 16004 22914 16016
rect 22339 15859 22385 15870
rect 22554 15868 22630 15901
rect 22554 15822 22565 15868
rect 22619 15822 22630 15868
rect 22738 15868 22814 15901
rect 22738 15822 22749 15868
rect 22803 15822 22814 15868
rect 22922 15868 22998 15901
rect 22922 15822 22933 15868
rect 22987 15822 22998 15868
rect 23167 15859 23213 15870
rect 22477 15776 22523 15787
rect 22460 15749 22477 15751
rect 22661 15776 22707 15787
rect 22523 15749 22540 15751
rect 22385 15629 22472 15749
rect 22528 15629 22540 15749
rect 22460 15627 22477 15629
rect 22385 15329 22477 15449
rect 22523 15627 22540 15629
rect 22644 15449 22661 15451
rect 22845 15776 22891 15787
rect 22828 15749 22845 15751
rect 23029 15776 23075 15787
rect 22891 15749 22908 15751
rect 22828 15629 22840 15749
rect 22896 15629 22908 15749
rect 22828 15627 22845 15629
rect 22707 15449 22724 15451
rect 22644 15329 22656 15449
rect 22712 15329 22724 15449
rect 22644 15327 22661 15329
rect 22477 15291 22523 15302
rect 22707 15327 22724 15329
rect 22661 15291 22707 15302
rect 22891 15627 22908 15629
rect 23012 15449 23029 15451
rect 23150 15749 23167 15751
rect 23213 15749 23230 15751
rect 23150 15628 23162 15749
rect 23218 15628 23230 15749
rect 23150 15626 23167 15628
rect 23075 15449 23092 15451
rect 23012 15329 23024 15449
rect 23080 15329 23092 15449
rect 23012 15327 23029 15329
rect 22845 15291 22891 15302
rect 23075 15327 23092 15329
rect 23029 15291 23075 15302
rect 22554 15253 22565 15256
rect 22619 15253 22630 15256
rect 22738 15253 22749 15256
rect 22803 15253 22814 15256
rect 22922 15253 22933 15256
rect 22987 15253 22998 15256
rect 22339 15208 22385 15219
rect 22552 15197 22564 15253
rect 22620 15197 22632 15253
rect 22552 15183 22632 15197
rect 22736 15197 22748 15253
rect 22804 15197 22816 15253
rect 22736 15183 22816 15197
rect 22920 15197 22932 15253
rect 22988 15197 23000 15253
rect 23213 15626 23230 15628
rect 23167 15208 23213 15219
rect 22920 15183 23000 15197
rect 22552 15103 22632 15105
rect 22164 15047 22564 15103
rect 22620 15047 22632 15103
rect 24720 15103 24776 16124
rect 25888 16116 25958 16124
rect 25384 16072 25470 16076
rect 25384 16016 25396 16072
rect 25452 16016 25470 16072
rect 25384 16004 25470 16016
rect 24895 15859 24941 15870
rect 25110 15868 25186 15901
rect 25110 15822 25121 15868
rect 25175 15822 25186 15868
rect 25294 15868 25370 15901
rect 25294 15822 25305 15868
rect 25359 15822 25370 15868
rect 25478 15868 25554 15901
rect 25478 15822 25489 15868
rect 25543 15822 25554 15868
rect 25723 15859 25769 15870
rect 25033 15776 25079 15787
rect 25016 15749 25033 15751
rect 25217 15776 25263 15787
rect 25079 15749 25096 15751
rect 24941 15629 25028 15749
rect 25084 15629 25096 15749
rect 25016 15627 25033 15629
rect 24941 15329 25033 15449
rect 25079 15627 25096 15629
rect 25200 15449 25217 15451
rect 25401 15776 25447 15787
rect 25384 15749 25401 15751
rect 25585 15776 25631 15787
rect 25447 15749 25464 15751
rect 25384 15629 25396 15749
rect 25452 15629 25464 15749
rect 25384 15627 25401 15629
rect 25263 15449 25280 15451
rect 25200 15329 25212 15449
rect 25268 15329 25280 15449
rect 25200 15327 25217 15329
rect 25033 15291 25079 15302
rect 25263 15327 25280 15329
rect 25217 15291 25263 15302
rect 25447 15627 25464 15629
rect 25568 15449 25585 15451
rect 25706 15749 25723 15751
rect 25769 15749 25786 15751
rect 25706 15628 25718 15749
rect 25774 15628 25786 15749
rect 25706 15626 25723 15628
rect 25631 15449 25648 15451
rect 25568 15329 25580 15449
rect 25636 15329 25648 15449
rect 25568 15327 25585 15329
rect 25401 15291 25447 15302
rect 25631 15327 25648 15329
rect 25585 15291 25631 15302
rect 25110 15253 25121 15256
rect 25175 15253 25186 15256
rect 25294 15253 25305 15256
rect 25359 15253 25370 15256
rect 25478 15253 25489 15256
rect 25543 15253 25554 15256
rect 24895 15208 24941 15219
rect 25108 15197 25120 15253
rect 25176 15197 25188 15253
rect 25108 15183 25188 15197
rect 25292 15197 25304 15253
rect 25360 15197 25372 15253
rect 25292 15183 25372 15197
rect 25476 15197 25488 15253
rect 25544 15197 25556 15253
rect 25769 15626 25786 15628
rect 25723 15208 25769 15219
rect 25476 15183 25556 15197
rect 25108 15103 25188 15105
rect 24720 15047 25120 15103
rect 25176 15047 25188 15103
rect 26206 15103 26262 18329
rect 28757 18329 30304 18385
rect 27768 17308 27848 17320
rect 28757 17308 28813 18329
rect 29426 18277 29512 18281
rect 29426 18221 29438 18277
rect 29494 18221 29512 18277
rect 29426 18209 29512 18221
rect 28937 18064 28983 18075
rect 29152 18073 29228 18106
rect 29152 18027 29163 18073
rect 29217 18027 29228 18073
rect 29336 18073 29412 18106
rect 29336 18027 29347 18073
rect 29401 18027 29412 18073
rect 29520 18073 29596 18106
rect 29520 18027 29531 18073
rect 29585 18027 29596 18073
rect 29765 18064 29811 18075
rect 29075 17981 29121 17992
rect 29058 17954 29075 17956
rect 29259 17981 29305 17992
rect 29121 17954 29138 17956
rect 28983 17834 29070 17954
rect 29126 17834 29138 17954
rect 29058 17832 29075 17834
rect 28983 17534 29075 17654
rect 29121 17832 29138 17834
rect 29242 17654 29259 17656
rect 29443 17981 29489 17992
rect 29426 17954 29443 17956
rect 29627 17981 29673 17992
rect 29489 17954 29506 17956
rect 29426 17834 29438 17954
rect 29494 17834 29506 17954
rect 29426 17832 29443 17834
rect 29305 17654 29322 17656
rect 29242 17534 29254 17654
rect 29310 17534 29322 17654
rect 29242 17532 29259 17534
rect 29075 17496 29121 17507
rect 29305 17532 29322 17534
rect 29259 17496 29305 17507
rect 29489 17832 29506 17834
rect 29610 17654 29627 17656
rect 29748 17954 29765 17956
rect 29811 17954 29828 17956
rect 29748 17833 29760 17954
rect 29816 17833 29828 17954
rect 29748 17831 29765 17833
rect 29673 17654 29690 17656
rect 29610 17534 29622 17654
rect 29678 17534 29690 17654
rect 29610 17532 29627 17534
rect 29443 17496 29489 17507
rect 29673 17532 29690 17534
rect 29627 17496 29673 17507
rect 29152 17458 29163 17461
rect 29217 17458 29228 17461
rect 29336 17458 29347 17461
rect 29401 17458 29412 17461
rect 29520 17458 29531 17461
rect 29585 17458 29596 17461
rect 28937 17413 28983 17424
rect 29150 17402 29162 17458
rect 29218 17402 29230 17458
rect 29150 17388 29230 17402
rect 29334 17402 29346 17458
rect 29402 17402 29414 17458
rect 29334 17388 29414 17402
rect 29518 17402 29530 17458
rect 29586 17402 29598 17458
rect 29811 17831 29828 17833
rect 29765 17413 29811 17424
rect 29518 17388 29598 17402
rect 29150 17308 29230 17310
rect 27768 17252 27780 17308
rect 27836 17252 29162 17308
rect 29218 17252 29230 17308
rect 27768 17250 27848 17252
rect 29150 17250 29230 17252
rect 28478 17192 28548 17204
rect 29334 17192 29414 17194
rect 28478 17136 28490 17192
rect 28546 17136 29346 17192
rect 29402 17136 29414 17192
rect 28478 17124 28548 17136
rect 29334 17134 29414 17136
rect 29663 17192 29743 17194
rect 29930 17192 30000 17204
rect 29663 17136 29675 17192
rect 29731 17136 29932 17192
rect 29988 17136 30000 17192
rect 29663 17134 29743 17136
rect 29930 17126 30000 17136
rect 29518 17076 29598 17078
rect 28762 17020 29530 17076
rect 29586 17020 29598 17076
rect 28762 16289 28818 17020
rect 29518 17018 29598 17020
rect 29150 16926 29230 16940
rect 28937 16904 28983 16915
rect 29150 16870 29162 16926
rect 29218 16870 29230 16926
rect 29334 16926 29414 16940
rect 29334 16870 29346 16926
rect 29402 16870 29414 16926
rect 29518 16926 29598 16940
rect 29518 16870 29530 16926
rect 29586 16870 29598 16926
rect 29765 16904 29811 16915
rect 29152 16867 29163 16870
rect 29217 16867 29228 16870
rect 29336 16867 29347 16870
rect 29401 16867 29412 16870
rect 29520 16867 29531 16870
rect 29585 16867 29596 16870
rect 29075 16821 29121 16832
rect 28983 16647 29075 16821
rect 29075 16636 29121 16647
rect 29259 16821 29305 16832
rect 29259 16636 29305 16647
rect 29443 16821 29489 16832
rect 29627 16821 29673 16832
rect 29610 16794 29627 16796
rect 29673 16794 29690 16796
rect 29610 16674 29622 16794
rect 29678 16674 29690 16794
rect 29610 16672 29627 16674
rect 29443 16636 29489 16647
rect 29673 16672 29690 16674
rect 29627 16636 29673 16647
rect 28937 16419 28983 16564
rect 29152 16555 29163 16601
rect 29217 16555 29228 16601
rect 29152 16522 29228 16555
rect 29336 16555 29347 16601
rect 29401 16555 29412 16601
rect 29336 16522 29412 16555
rect 29520 16555 29531 16601
rect 29585 16555 29596 16601
rect 29520 16522 29596 16555
rect 29765 16419 29811 16564
rect 28925 16407 29005 16419
rect 28925 16351 28937 16407
rect 28993 16351 29005 16407
rect 28925 16339 29005 16351
rect 29743 16407 29823 16419
rect 29743 16351 29755 16407
rect 29811 16351 29823 16407
rect 29743 16339 29823 16351
rect 30096 16289 30176 16299
rect 28762 16233 30108 16289
rect 30164 16233 30176 16289
rect 30096 16231 30176 16233
rect 29930 16180 30000 16182
rect 28762 16179 30000 16180
rect 28762 16125 29932 16179
rect 29988 16125 30000 16179
rect 28762 16124 30000 16125
rect 26870 16072 26956 16076
rect 26870 16016 26882 16072
rect 26938 16016 26956 16072
rect 26870 16004 26956 16016
rect 26381 15859 26427 15870
rect 26596 15868 26672 15901
rect 26596 15822 26607 15868
rect 26661 15822 26672 15868
rect 26780 15868 26856 15901
rect 26780 15822 26791 15868
rect 26845 15822 26856 15868
rect 26964 15868 27040 15901
rect 26964 15822 26975 15868
rect 27029 15822 27040 15868
rect 27209 15859 27255 15870
rect 26519 15776 26565 15787
rect 26502 15749 26519 15751
rect 26703 15776 26749 15787
rect 26565 15749 26582 15751
rect 26427 15629 26514 15749
rect 26570 15629 26582 15749
rect 26502 15627 26519 15629
rect 26427 15329 26519 15449
rect 26565 15627 26582 15629
rect 26686 15449 26703 15451
rect 26887 15776 26933 15787
rect 26870 15749 26887 15751
rect 27071 15776 27117 15787
rect 26933 15749 26950 15751
rect 26870 15629 26882 15749
rect 26938 15629 26950 15749
rect 26870 15627 26887 15629
rect 26749 15449 26766 15451
rect 26686 15329 26698 15449
rect 26754 15329 26766 15449
rect 26686 15327 26703 15329
rect 26519 15291 26565 15302
rect 26749 15327 26766 15329
rect 26703 15291 26749 15302
rect 26933 15627 26950 15629
rect 27054 15449 27071 15451
rect 27192 15749 27209 15751
rect 27255 15749 27272 15751
rect 27192 15628 27204 15749
rect 27260 15628 27272 15749
rect 27192 15626 27209 15628
rect 27117 15449 27134 15451
rect 27054 15329 27066 15449
rect 27122 15329 27134 15449
rect 27054 15327 27071 15329
rect 26887 15291 26933 15302
rect 27117 15327 27134 15329
rect 27071 15291 27117 15302
rect 26596 15253 26607 15256
rect 26661 15253 26672 15256
rect 26780 15253 26791 15256
rect 26845 15253 26856 15256
rect 26964 15253 26975 15256
rect 27029 15253 27040 15256
rect 26381 15208 26427 15219
rect 26594 15197 26606 15253
rect 26662 15197 26674 15253
rect 26594 15183 26674 15197
rect 26778 15197 26790 15253
rect 26846 15197 26858 15253
rect 26778 15183 26858 15197
rect 26962 15197 26974 15253
rect 27030 15197 27042 15253
rect 27255 15626 27272 15628
rect 27209 15208 27255 15219
rect 26962 15183 27042 15197
rect 26594 15103 26674 15105
rect 26206 15047 26606 15103
rect 26662 15047 26674 15103
rect 28762 15103 28818 16124
rect 29930 16116 30000 16124
rect 29426 16072 29512 16076
rect 29426 16016 29438 16072
rect 29494 16016 29512 16072
rect 29426 16004 29512 16016
rect 28937 15859 28983 15870
rect 29152 15868 29228 15901
rect 29152 15822 29163 15868
rect 29217 15822 29228 15868
rect 29336 15868 29412 15901
rect 29336 15822 29347 15868
rect 29401 15822 29412 15868
rect 29520 15868 29596 15901
rect 29520 15822 29531 15868
rect 29585 15822 29596 15868
rect 29765 15859 29811 15870
rect 29075 15776 29121 15787
rect 29058 15749 29075 15751
rect 29259 15776 29305 15787
rect 29121 15749 29138 15751
rect 28983 15629 29070 15749
rect 29126 15629 29138 15749
rect 29058 15627 29075 15629
rect 28983 15329 29075 15449
rect 29121 15627 29138 15629
rect 29242 15449 29259 15451
rect 29443 15776 29489 15787
rect 29426 15749 29443 15751
rect 29627 15776 29673 15787
rect 29489 15749 29506 15751
rect 29426 15629 29438 15749
rect 29494 15629 29506 15749
rect 29426 15627 29443 15629
rect 29305 15449 29322 15451
rect 29242 15329 29254 15449
rect 29310 15329 29322 15449
rect 29242 15327 29259 15329
rect 29075 15291 29121 15302
rect 29305 15327 29322 15329
rect 29259 15291 29305 15302
rect 29489 15627 29506 15629
rect 29610 15449 29627 15451
rect 29748 15749 29765 15751
rect 29811 15749 29828 15751
rect 29748 15628 29760 15749
rect 29816 15628 29828 15749
rect 29748 15626 29765 15628
rect 29673 15449 29690 15451
rect 29610 15329 29622 15449
rect 29678 15329 29690 15449
rect 29610 15327 29627 15329
rect 29443 15291 29489 15302
rect 29673 15327 29690 15329
rect 29627 15291 29673 15302
rect 29152 15253 29163 15256
rect 29217 15253 29228 15256
rect 29336 15253 29347 15256
rect 29401 15253 29412 15256
rect 29520 15253 29531 15256
rect 29585 15253 29596 15256
rect 28937 15208 28983 15219
rect 29150 15197 29162 15253
rect 29218 15197 29230 15253
rect 29150 15183 29230 15197
rect 29334 15197 29346 15253
rect 29402 15197 29414 15253
rect 29334 15183 29414 15197
rect 29518 15197 29530 15253
rect 29586 15197 29598 15253
rect 29811 15626 29828 15628
rect 29765 15208 29811 15219
rect 29518 15183 29598 15197
rect 29150 15103 29230 15105
rect 28762 15047 29162 15103
rect 29218 15047 29230 15103
rect 30248 15103 30304 18329
rect 30912 16072 30998 16076
rect 30912 16016 30924 16072
rect 30980 16016 30998 16072
rect 30912 16004 30998 16016
rect 30423 15859 30469 15870
rect 30638 15868 30714 15901
rect 30638 15822 30649 15868
rect 30703 15822 30714 15868
rect 30822 15868 30898 15901
rect 30822 15822 30833 15868
rect 30887 15822 30898 15868
rect 31006 15868 31082 15901
rect 31006 15822 31017 15868
rect 31071 15822 31082 15868
rect 31251 15859 31297 15870
rect 30561 15776 30607 15787
rect 30544 15749 30561 15751
rect 30745 15776 30791 15787
rect 30607 15749 30624 15751
rect 30469 15629 30556 15749
rect 30612 15629 30624 15749
rect 30544 15627 30561 15629
rect 30469 15329 30561 15449
rect 30607 15627 30624 15629
rect 30728 15449 30745 15451
rect 30929 15776 30975 15787
rect 30912 15749 30929 15751
rect 31113 15776 31159 15787
rect 30975 15749 30992 15751
rect 30912 15629 30924 15749
rect 30980 15629 30992 15749
rect 30912 15627 30929 15629
rect 30791 15449 30808 15451
rect 30728 15329 30740 15449
rect 30796 15329 30808 15449
rect 30728 15327 30745 15329
rect 30561 15291 30607 15302
rect 30791 15327 30808 15329
rect 30745 15291 30791 15302
rect 30975 15627 30992 15629
rect 31096 15449 31113 15451
rect 31234 15749 31251 15751
rect 31297 15749 31314 15751
rect 31234 15628 31246 15749
rect 31302 15628 31314 15749
rect 31234 15626 31251 15628
rect 31159 15449 31176 15451
rect 31096 15329 31108 15449
rect 31164 15329 31176 15449
rect 31096 15327 31113 15329
rect 30929 15291 30975 15302
rect 31159 15327 31176 15329
rect 31113 15291 31159 15302
rect 30638 15253 30649 15256
rect 30703 15253 30714 15256
rect 30822 15253 30833 15256
rect 30887 15253 30898 15256
rect 31006 15253 31017 15256
rect 31071 15253 31082 15256
rect 30423 15208 30469 15219
rect 30636 15197 30648 15253
rect 30704 15197 30716 15253
rect 30636 15183 30716 15197
rect 30820 15197 30832 15253
rect 30888 15197 30900 15253
rect 30820 15183 30900 15197
rect 31004 15197 31016 15253
rect 31072 15197 31084 15253
rect 31297 15626 31314 15628
rect 31251 15208 31297 15219
rect 31004 15183 31084 15197
rect 30636 15103 30716 15105
rect 30248 15047 30648 15103
rect 30704 15047 30716 15103
rect 8940 15045 9020 15047
rect 10426 15045 10506 15047
rect 12982 15045 13062 15047
rect 14468 15045 14548 15047
rect 17024 15045 17104 15047
rect 18510 15045 18590 15047
rect 21066 15045 21146 15047
rect 22552 15045 22632 15047
rect 25108 15045 25188 15047
rect 26594 15045 26674 15047
rect 29150 15045 29230 15047
rect 30636 15045 30716 15047
rect 4090 14990 4160 15004
rect 5082 14990 5162 14992
rect 4090 14934 4102 14990
rect 4158 14934 5094 14990
rect 5150 14934 5162 14990
rect 4090 14922 4160 14934
rect 5082 14932 5162 14934
rect 5411 14990 5491 14992
rect 5854 14990 5914 15000
rect 6568 14990 6648 14992
rect 5411 14934 5423 14990
rect 5479 14934 5856 14990
rect 5912 14934 6580 14990
rect 6636 14934 6648 14990
rect 5411 14932 5491 14934
rect 5854 14922 5914 14934
rect 6568 14932 6648 14934
rect 6897 14990 6977 14992
rect 7164 14990 7234 15002
rect 7704 14990 7774 14992
rect 6897 14934 6909 14990
rect 6965 14934 7166 14990
rect 7222 14934 7706 14990
rect 7762 14934 7774 14990
rect 6897 14932 6977 14934
rect 7164 14924 7234 14934
rect 7704 14922 7774 14934
rect 8132 14987 8202 15001
rect 9124 14987 9204 14989
rect 8132 14931 8144 14987
rect 8200 14931 9136 14987
rect 9192 14931 9204 14987
rect 8132 14919 8202 14931
rect 9124 14929 9204 14931
rect 9453 14987 9533 14989
rect 9896 14987 9956 14997
rect 10610 14987 10690 14989
rect 9453 14931 9465 14987
rect 9521 14931 9898 14987
rect 9954 14931 10622 14987
rect 10678 14931 10690 14987
rect 9453 14929 9533 14931
rect 9896 14919 9956 14931
rect 10610 14929 10690 14931
rect 10939 14987 11019 14989
rect 11206 14987 11276 14999
rect 11758 14987 11828 14999
rect 10939 14931 10951 14987
rect 11007 14931 11208 14987
rect 11264 14931 11760 14987
rect 11816 14931 11828 14987
rect 10939 14929 11019 14931
rect 11206 14921 11276 14931
rect 11758 14919 11828 14931
rect 12174 14987 12244 15001
rect 13166 14987 13246 14989
rect 12174 14931 12186 14987
rect 12242 14931 13178 14987
rect 13234 14931 13246 14987
rect 12174 14919 12244 14931
rect 13166 14929 13246 14931
rect 13495 14987 13575 14989
rect 13938 14987 13998 14997
rect 14652 14987 14732 14989
rect 13495 14931 13507 14987
rect 13563 14931 13940 14987
rect 13996 14931 14664 14987
rect 14720 14931 14732 14987
rect 13495 14929 13575 14931
rect 13938 14919 13998 14931
rect 14652 14929 14732 14931
rect 14981 14987 15061 14989
rect 15248 14987 15318 14999
rect 15854 14987 15924 14999
rect 14981 14931 14993 14987
rect 15049 14931 15250 14987
rect 15306 14931 15856 14987
rect 15912 14931 15924 14987
rect 14981 14929 15061 14931
rect 15248 14921 15318 14931
rect 15854 14919 15924 14931
rect 16216 14987 16286 15001
rect 17208 14987 17288 14989
rect 16216 14931 16228 14987
rect 16284 14931 17220 14987
rect 17276 14931 17288 14987
rect 16216 14919 16286 14931
rect 17208 14929 17288 14931
rect 17537 14987 17617 14989
rect 17980 14987 18040 14997
rect 18694 14987 18774 14989
rect 17537 14931 17549 14987
rect 17605 14931 17982 14987
rect 18038 14931 18706 14987
rect 18762 14931 18774 14987
rect 17537 14929 17617 14931
rect 17980 14919 18040 14931
rect 18694 14929 18774 14931
rect 19023 14987 19103 14989
rect 19290 14987 19360 14999
rect 19896 14987 19966 14999
rect 19023 14931 19035 14987
rect 19091 14931 19292 14987
rect 19348 14931 19898 14987
rect 19954 14931 19966 14987
rect 19023 14929 19103 14931
rect 19290 14921 19360 14931
rect 19896 14919 19966 14931
rect 20258 14987 20328 15001
rect 21250 14987 21330 14989
rect 20258 14931 20270 14987
rect 20326 14931 21262 14987
rect 21318 14931 21330 14987
rect 20258 14919 20328 14931
rect 21250 14929 21330 14931
rect 21579 14987 21659 14989
rect 22022 14987 22082 14997
rect 22736 14987 22816 14989
rect 21579 14931 21591 14987
rect 21647 14931 22024 14987
rect 22080 14931 22748 14987
rect 22804 14931 22816 14987
rect 21579 14929 21659 14931
rect 22022 14919 22082 14931
rect 22736 14929 22816 14931
rect 23065 14987 23145 14989
rect 23332 14987 23402 14999
rect 23938 14987 24008 14999
rect 23065 14931 23077 14987
rect 23133 14931 23334 14987
rect 23390 14931 23940 14987
rect 23996 14931 24008 14987
rect 23065 14929 23145 14931
rect 23332 14921 23402 14931
rect 23938 14919 24008 14931
rect 24300 14987 24370 15001
rect 25292 14987 25372 14989
rect 24300 14931 24312 14987
rect 24368 14931 25304 14987
rect 25360 14931 25372 14987
rect 24300 14919 24370 14931
rect 25292 14929 25372 14931
rect 25621 14987 25701 14989
rect 26064 14987 26124 14997
rect 26778 14987 26858 14989
rect 25621 14931 25633 14987
rect 25689 14931 26066 14987
rect 26122 14931 26790 14987
rect 26846 14931 26858 14987
rect 25621 14929 25701 14931
rect 26064 14919 26124 14931
rect 26778 14929 26858 14931
rect 27107 14987 27187 14989
rect 27374 14987 27444 14999
rect 27980 14987 28050 14999
rect 27107 14931 27119 14987
rect 27175 14931 27376 14987
rect 27432 14931 27982 14987
rect 28038 14931 28050 14987
rect 27107 14929 27187 14931
rect 27374 14921 27444 14931
rect 27980 14919 28050 14931
rect 28342 14987 28412 15001
rect 29334 14987 29414 14989
rect 28342 14931 28354 14987
rect 28410 14931 29346 14987
rect 29402 14931 29414 14987
rect 28342 14919 28412 14931
rect 29334 14929 29414 14931
rect 29663 14987 29743 14989
rect 30106 14987 30166 14997
rect 30820 14987 30900 14989
rect 29663 14931 29675 14987
rect 29731 14931 30108 14987
rect 30164 14931 30832 14987
rect 30888 14931 30900 14987
rect 29663 14929 29743 14931
rect 30106 14919 30166 14931
rect 30820 14929 30900 14931
rect 31149 14987 31229 14989
rect 31416 14987 31486 14999
rect 32022 14987 32092 14999
rect 31149 14931 31161 14987
rect 31217 14931 31418 14987
rect 31474 14931 32024 14987
rect 32080 14931 32092 14987
rect 31149 14929 31229 14931
rect 31416 14921 31486 14931
rect 32022 14919 32092 14931
rect 5266 14874 5346 14876
rect 6752 14874 6832 14876
rect 4374 14818 5278 14874
rect 5334 14818 5346 14874
rect 3900 14088 3970 14090
rect 4374 14088 4430 14818
rect 5266 14816 5346 14818
rect 5996 14818 6764 14874
rect 6820 14818 6832 14874
rect 9308 14871 9388 14873
rect 10794 14871 10874 14873
rect 13350 14871 13430 14873
rect 14836 14871 14916 14873
rect 17392 14871 17472 14873
rect 18878 14871 18958 14873
rect 21434 14871 21514 14873
rect 22920 14871 23000 14873
rect 25476 14871 25556 14873
rect 26962 14871 27042 14873
rect 29518 14871 29598 14873
rect 31004 14871 31084 14873
rect 4898 14724 4978 14738
rect 4685 14702 4731 14713
rect 4898 14668 4910 14724
rect 4966 14668 4978 14724
rect 5082 14724 5162 14738
rect 5082 14668 5094 14724
rect 5150 14668 5162 14724
rect 5266 14724 5346 14738
rect 5266 14668 5278 14724
rect 5334 14668 5346 14724
rect 5513 14702 5559 14713
rect 4900 14665 4911 14668
rect 4965 14665 4976 14668
rect 5084 14665 5095 14668
rect 5149 14665 5160 14668
rect 5268 14665 5279 14668
rect 5333 14665 5344 14668
rect 4823 14619 4869 14630
rect 4731 14445 4823 14619
rect 4823 14434 4869 14445
rect 5007 14619 5053 14630
rect 5007 14434 5053 14445
rect 5191 14619 5237 14630
rect 5375 14619 5421 14630
rect 5358 14592 5375 14594
rect 5421 14592 5438 14594
rect 5358 14472 5370 14592
rect 5426 14472 5438 14592
rect 5358 14470 5375 14472
rect 5191 14434 5237 14445
rect 5421 14470 5438 14472
rect 5375 14434 5421 14445
rect 4685 14217 4731 14362
rect 4900 14353 4911 14399
rect 4965 14353 4976 14399
rect 4900 14320 4976 14353
rect 5084 14353 5095 14399
rect 5149 14353 5160 14399
rect 5084 14320 5160 14353
rect 5268 14353 5279 14399
rect 5333 14353 5344 14399
rect 5268 14320 5344 14353
rect 5513 14217 5559 14362
rect 4673 14205 4753 14217
rect 4673 14149 4685 14205
rect 4741 14149 4753 14205
rect 4673 14137 4753 14149
rect 5491 14205 5569 14217
rect 5491 14149 5503 14205
rect 5559 14149 5569 14205
rect 5491 14137 5569 14149
rect 3900 14032 3912 14088
rect 3968 14032 4430 14088
rect 5996 14088 6052 14818
rect 6752 14816 6832 14818
rect 8416 14815 9320 14871
rect 9376 14815 9388 14871
rect 6384 14724 6464 14738
rect 6171 14702 6217 14713
rect 6384 14668 6396 14724
rect 6452 14668 6464 14724
rect 6568 14724 6648 14738
rect 6568 14668 6580 14724
rect 6636 14668 6648 14724
rect 6752 14724 6832 14738
rect 6752 14668 6764 14724
rect 6820 14668 6832 14724
rect 6999 14702 7045 14713
rect 6386 14665 6397 14668
rect 6451 14665 6462 14668
rect 6570 14665 6581 14668
rect 6635 14665 6646 14668
rect 6754 14665 6765 14668
rect 6819 14665 6830 14668
rect 6309 14619 6355 14630
rect 6217 14445 6309 14619
rect 6309 14434 6355 14445
rect 6493 14619 6539 14630
rect 6493 14434 6539 14445
rect 6677 14619 6723 14630
rect 6861 14619 6907 14630
rect 6844 14592 6861 14594
rect 6907 14592 6924 14594
rect 6844 14472 6856 14592
rect 6912 14472 6924 14592
rect 6844 14470 6861 14472
rect 6677 14434 6723 14445
rect 6907 14470 6924 14472
rect 6861 14434 6907 14445
rect 6171 14217 6217 14362
rect 6386 14353 6397 14399
rect 6451 14353 6462 14399
rect 6386 14320 6462 14353
rect 6570 14353 6581 14399
rect 6635 14353 6646 14399
rect 6570 14320 6646 14353
rect 6754 14353 6765 14399
rect 6819 14353 6830 14399
rect 6754 14320 6830 14353
rect 6999 14217 7045 14362
rect 6159 14205 6239 14217
rect 6159 14149 6171 14205
rect 6227 14149 6239 14205
rect 6159 14137 6239 14149
rect 6977 14205 7055 14217
rect 6977 14149 6989 14205
rect 7045 14149 7055 14205
rect 6977 14137 7055 14149
rect 7330 14088 7410 14098
rect 5996 14032 7342 14088
rect 7398 14032 7410 14088
rect 3900 14020 3970 14032
rect 4374 12785 4430 14032
rect 7330 14030 7410 14032
rect 7996 14085 8066 14087
rect 8416 14085 8472 14815
rect 9308 14813 9388 14815
rect 10038 14815 10806 14871
rect 10862 14815 10874 14871
rect 8940 14721 9020 14735
rect 8727 14699 8773 14710
rect 8940 14665 8952 14721
rect 9008 14665 9020 14721
rect 9124 14721 9204 14735
rect 9124 14665 9136 14721
rect 9192 14665 9204 14721
rect 9308 14721 9388 14735
rect 9308 14665 9320 14721
rect 9376 14665 9388 14721
rect 9555 14699 9601 14710
rect 8942 14662 8953 14665
rect 9007 14662 9018 14665
rect 9126 14662 9137 14665
rect 9191 14662 9202 14665
rect 9310 14662 9321 14665
rect 9375 14662 9386 14665
rect 8865 14616 8911 14627
rect 8773 14442 8865 14616
rect 8865 14431 8911 14442
rect 9049 14616 9095 14627
rect 9049 14431 9095 14442
rect 9233 14616 9279 14627
rect 9417 14616 9463 14627
rect 9400 14589 9417 14591
rect 9463 14589 9480 14591
rect 9400 14469 9412 14589
rect 9468 14469 9480 14589
rect 9400 14467 9417 14469
rect 9233 14431 9279 14442
rect 9463 14467 9480 14469
rect 9417 14431 9463 14442
rect 8727 14214 8773 14359
rect 8942 14350 8953 14396
rect 9007 14350 9018 14396
rect 8942 14317 9018 14350
rect 9126 14350 9137 14396
rect 9191 14350 9202 14396
rect 9126 14317 9202 14350
rect 9310 14350 9321 14396
rect 9375 14350 9386 14396
rect 9310 14317 9386 14350
rect 9555 14214 9601 14359
rect 8715 14202 8795 14214
rect 8715 14146 8727 14202
rect 8783 14146 8795 14202
rect 8715 14134 8795 14146
rect 9533 14202 9611 14214
rect 9533 14146 9545 14202
rect 9601 14146 9611 14202
rect 9533 14134 9611 14146
rect 7996 14029 8008 14085
rect 8064 14029 8472 14085
rect 10038 14085 10094 14815
rect 10794 14813 10874 14815
rect 12458 14815 13362 14871
rect 13418 14815 13430 14871
rect 10426 14721 10506 14735
rect 10213 14699 10259 14710
rect 10426 14665 10438 14721
rect 10494 14665 10506 14721
rect 10610 14721 10690 14735
rect 10610 14665 10622 14721
rect 10678 14665 10690 14721
rect 10794 14721 10874 14735
rect 10794 14665 10806 14721
rect 10862 14665 10874 14721
rect 11041 14699 11087 14710
rect 10428 14662 10439 14665
rect 10493 14662 10504 14665
rect 10612 14662 10623 14665
rect 10677 14662 10688 14665
rect 10796 14662 10807 14665
rect 10861 14662 10872 14665
rect 10351 14616 10397 14627
rect 10259 14442 10351 14616
rect 10351 14431 10397 14442
rect 10535 14616 10581 14627
rect 10535 14431 10581 14442
rect 10719 14616 10765 14627
rect 10903 14616 10949 14627
rect 10886 14589 10903 14591
rect 10949 14589 10966 14591
rect 10886 14469 10898 14589
rect 10954 14469 10966 14589
rect 10886 14467 10903 14469
rect 10719 14431 10765 14442
rect 10949 14467 10966 14469
rect 10903 14431 10949 14442
rect 10213 14214 10259 14359
rect 10428 14350 10439 14396
rect 10493 14350 10504 14396
rect 10428 14317 10504 14350
rect 10612 14350 10623 14396
rect 10677 14350 10688 14396
rect 10612 14317 10688 14350
rect 10796 14350 10807 14396
rect 10861 14350 10872 14396
rect 10796 14317 10872 14350
rect 11041 14214 11087 14359
rect 10201 14202 10281 14214
rect 10201 14146 10213 14202
rect 10269 14146 10281 14202
rect 10201 14134 10281 14146
rect 11019 14202 11097 14214
rect 11019 14146 11031 14202
rect 11087 14146 11097 14202
rect 11019 14134 11097 14146
rect 11372 14085 11452 14095
rect 10038 14029 11384 14085
rect 11440 14029 11452 14085
rect 7996 14017 8066 14029
rect 5854 13977 5924 13979
rect 7154 13978 7234 13980
rect 4510 13921 5856 13977
rect 5912 13921 5924 13977
rect 4510 12901 4566 13921
rect 5854 13909 5924 13921
rect 5996 13922 7166 13978
rect 7222 13922 7234 13978
rect 5174 13870 5260 13874
rect 5174 13814 5186 13870
rect 5242 13814 5260 13870
rect 5174 13802 5260 13814
rect 4685 13657 4731 13668
rect 4900 13666 4976 13699
rect 4900 13620 4911 13666
rect 4965 13620 4976 13666
rect 5084 13666 5160 13699
rect 5084 13620 5095 13666
rect 5149 13620 5160 13666
rect 5268 13666 5344 13699
rect 5268 13620 5279 13666
rect 5333 13620 5344 13666
rect 5513 13657 5559 13668
rect 4823 13574 4869 13585
rect 4806 13547 4823 13549
rect 5007 13574 5053 13585
rect 4869 13547 4886 13549
rect 4731 13427 4818 13547
rect 4874 13427 4886 13547
rect 4806 13425 4823 13427
rect 4731 13127 4823 13247
rect 4869 13425 4886 13427
rect 4990 13247 5007 13249
rect 5191 13574 5237 13585
rect 5174 13547 5191 13549
rect 5375 13574 5421 13585
rect 5237 13547 5254 13549
rect 5174 13427 5186 13547
rect 5242 13427 5254 13547
rect 5174 13425 5191 13427
rect 5053 13247 5070 13249
rect 4990 13127 5002 13247
rect 5058 13127 5070 13247
rect 4990 13125 5007 13127
rect 4823 13089 4869 13100
rect 5053 13125 5070 13127
rect 5007 13089 5053 13100
rect 5237 13425 5254 13427
rect 5358 13247 5375 13249
rect 5496 13547 5513 13549
rect 5559 13547 5576 13549
rect 5496 13426 5508 13547
rect 5564 13426 5576 13547
rect 5496 13424 5513 13426
rect 5421 13247 5438 13249
rect 5358 13127 5370 13247
rect 5426 13127 5438 13247
rect 5358 13125 5375 13127
rect 5191 13089 5237 13100
rect 5421 13125 5438 13127
rect 5375 13089 5421 13100
rect 4900 13051 4911 13054
rect 4965 13051 4976 13054
rect 5084 13051 5095 13054
rect 5149 13051 5160 13054
rect 5268 13051 5279 13054
rect 5333 13051 5344 13054
rect 4685 13006 4731 13017
rect 4898 12995 4910 13051
rect 4966 12995 4978 13051
rect 4898 12981 4978 12995
rect 5082 12995 5094 13051
rect 5150 12995 5162 13051
rect 5082 12981 5162 12995
rect 5266 12995 5278 13051
rect 5334 12995 5346 13051
rect 5559 13424 5576 13426
rect 5513 13006 5559 13017
rect 5266 12981 5346 12995
rect 4898 12901 4978 12903
rect 4510 12845 4910 12901
rect 4966 12845 4978 12901
rect 5996 12902 6052 13922
rect 7154 13910 7234 13922
rect 6660 13871 6746 13875
rect 6660 13815 6672 13871
rect 6728 13815 6746 13871
rect 6660 13803 6746 13815
rect 6171 13658 6217 13669
rect 6386 13667 6462 13700
rect 6386 13621 6397 13667
rect 6451 13621 6462 13667
rect 6570 13667 6646 13700
rect 6570 13621 6581 13667
rect 6635 13621 6646 13667
rect 6754 13667 6830 13700
rect 6754 13621 6765 13667
rect 6819 13621 6830 13667
rect 6999 13658 7045 13669
rect 6309 13575 6355 13586
rect 6292 13548 6309 13550
rect 6493 13575 6539 13586
rect 6355 13548 6372 13550
rect 6217 13428 6304 13548
rect 6360 13428 6372 13548
rect 6292 13426 6309 13428
rect 6217 13128 6309 13248
rect 6355 13426 6372 13428
rect 6476 13248 6493 13250
rect 6677 13575 6723 13586
rect 6660 13548 6677 13550
rect 6861 13575 6907 13586
rect 6723 13548 6740 13550
rect 6660 13428 6672 13548
rect 6728 13428 6740 13548
rect 6660 13426 6677 13428
rect 6539 13248 6556 13250
rect 6476 13128 6488 13248
rect 6544 13128 6556 13248
rect 6476 13126 6493 13128
rect 6309 13090 6355 13101
rect 6539 13126 6556 13128
rect 6493 13090 6539 13101
rect 6723 13426 6740 13428
rect 6844 13248 6861 13250
rect 6982 13548 6999 13550
rect 7045 13548 7062 13550
rect 6982 13427 6994 13548
rect 7050 13427 7062 13548
rect 6982 13425 6999 13427
rect 6907 13248 6924 13250
rect 6844 13128 6856 13248
rect 6912 13128 6924 13248
rect 6844 13126 6861 13128
rect 6677 13090 6723 13101
rect 6907 13126 6924 13128
rect 6861 13090 6907 13101
rect 6386 13052 6397 13055
rect 6451 13052 6462 13055
rect 6570 13052 6581 13055
rect 6635 13052 6646 13055
rect 6754 13052 6765 13055
rect 6819 13052 6830 13055
rect 6171 13007 6217 13018
rect 6384 12996 6396 13052
rect 6452 12996 6464 13052
rect 6384 12982 6464 12996
rect 6568 12996 6580 13052
rect 6636 12996 6648 13052
rect 6568 12982 6648 12996
rect 6752 12996 6764 13052
rect 6820 12996 6832 13052
rect 7045 13425 7062 13427
rect 6999 13007 7045 13018
rect 6752 12982 6832 12996
rect 6384 12902 6464 12904
rect 5996 12846 6396 12902
rect 6452 12846 6464 12902
rect 4898 12843 4978 12845
rect 6384 12844 6464 12846
rect 5082 12785 5162 12787
rect 4374 12729 5094 12785
rect 5150 12729 5162 12785
rect 5082 12727 5162 12729
rect 5411 12785 5491 12787
rect 5678 12786 5748 12797
rect 6568 12786 6648 12788
rect 5678 12785 6580 12786
rect 5411 12729 5423 12785
rect 5479 12729 5680 12785
rect 5736 12730 6580 12785
rect 6636 12730 6648 12786
rect 5736 12729 5996 12730
rect 5411 12727 5491 12729
rect 5678 12719 5748 12729
rect 6568 12728 6648 12730
rect 6897 12786 6977 12788
rect 7340 12786 7410 12796
rect 6897 12730 6909 12786
rect 6965 12730 7342 12786
rect 7398 12730 7410 12786
rect 6897 12728 6977 12730
rect 7340 12718 7410 12730
rect 8416 12782 8472 14029
rect 11372 14027 11452 14029
rect 12038 14085 12108 14087
rect 12458 14085 12514 14815
rect 13350 14813 13430 14815
rect 14080 14815 14848 14871
rect 14904 14815 14916 14871
rect 12982 14721 13062 14735
rect 12769 14699 12815 14710
rect 12982 14665 12994 14721
rect 13050 14665 13062 14721
rect 13166 14721 13246 14735
rect 13166 14665 13178 14721
rect 13234 14665 13246 14721
rect 13350 14721 13430 14735
rect 13350 14665 13362 14721
rect 13418 14665 13430 14721
rect 13597 14699 13643 14710
rect 12984 14662 12995 14665
rect 13049 14662 13060 14665
rect 13168 14662 13179 14665
rect 13233 14662 13244 14665
rect 13352 14662 13363 14665
rect 13417 14662 13428 14665
rect 12907 14616 12953 14627
rect 12815 14442 12907 14616
rect 12907 14431 12953 14442
rect 13091 14616 13137 14627
rect 13091 14431 13137 14442
rect 13275 14616 13321 14627
rect 13459 14616 13505 14627
rect 13442 14589 13459 14591
rect 13505 14589 13522 14591
rect 13442 14469 13454 14589
rect 13510 14469 13522 14589
rect 13442 14467 13459 14469
rect 13275 14431 13321 14442
rect 13505 14467 13522 14469
rect 13459 14431 13505 14442
rect 12769 14214 12815 14359
rect 12984 14350 12995 14396
rect 13049 14350 13060 14396
rect 12984 14317 13060 14350
rect 13168 14350 13179 14396
rect 13233 14350 13244 14396
rect 13168 14317 13244 14350
rect 13352 14350 13363 14396
rect 13417 14350 13428 14396
rect 13352 14317 13428 14350
rect 13597 14214 13643 14359
rect 12757 14202 12837 14214
rect 12757 14146 12769 14202
rect 12825 14146 12837 14202
rect 12757 14134 12837 14146
rect 13575 14202 13653 14214
rect 13575 14146 13587 14202
rect 13643 14146 13653 14202
rect 13575 14134 13653 14146
rect 12038 14029 12050 14085
rect 12106 14029 12514 14085
rect 14080 14085 14136 14815
rect 14836 14813 14916 14815
rect 16500 14815 17404 14871
rect 17460 14815 17472 14871
rect 14468 14721 14548 14735
rect 14255 14699 14301 14710
rect 14468 14665 14480 14721
rect 14536 14665 14548 14721
rect 14652 14721 14732 14735
rect 14652 14665 14664 14721
rect 14720 14665 14732 14721
rect 14836 14721 14916 14735
rect 14836 14665 14848 14721
rect 14904 14665 14916 14721
rect 15083 14699 15129 14710
rect 14470 14662 14481 14665
rect 14535 14662 14546 14665
rect 14654 14662 14665 14665
rect 14719 14662 14730 14665
rect 14838 14662 14849 14665
rect 14903 14662 14914 14665
rect 14393 14616 14439 14627
rect 14301 14442 14393 14616
rect 14393 14431 14439 14442
rect 14577 14616 14623 14627
rect 14577 14431 14623 14442
rect 14761 14616 14807 14627
rect 14945 14616 14991 14627
rect 14928 14589 14945 14591
rect 14991 14589 15008 14591
rect 14928 14469 14940 14589
rect 14996 14469 15008 14589
rect 14928 14467 14945 14469
rect 14761 14431 14807 14442
rect 14991 14467 15008 14469
rect 14945 14431 14991 14442
rect 14255 14214 14301 14359
rect 14470 14350 14481 14396
rect 14535 14350 14546 14396
rect 14470 14317 14546 14350
rect 14654 14350 14665 14396
rect 14719 14350 14730 14396
rect 14654 14317 14730 14350
rect 14838 14350 14849 14396
rect 14903 14350 14914 14396
rect 14838 14317 14914 14350
rect 15083 14214 15129 14359
rect 14243 14202 14323 14214
rect 14243 14146 14255 14202
rect 14311 14146 14323 14202
rect 14243 14134 14323 14146
rect 15061 14202 15139 14214
rect 15061 14146 15073 14202
rect 15129 14146 15139 14202
rect 15061 14134 15139 14146
rect 15414 14085 15494 14095
rect 14080 14029 15426 14085
rect 15482 14029 15494 14085
rect 12038 14017 12108 14029
rect 9896 13974 9966 13976
rect 11196 13975 11276 13977
rect 8552 13918 9898 13974
rect 9954 13918 9966 13974
rect 8552 12898 8608 13918
rect 9896 13906 9966 13918
rect 10038 13919 11208 13975
rect 11264 13919 11276 13975
rect 9216 13867 9302 13871
rect 9216 13811 9228 13867
rect 9284 13811 9302 13867
rect 9216 13799 9302 13811
rect 8727 13654 8773 13665
rect 8942 13663 9018 13696
rect 8942 13617 8953 13663
rect 9007 13617 9018 13663
rect 9126 13663 9202 13696
rect 9126 13617 9137 13663
rect 9191 13617 9202 13663
rect 9310 13663 9386 13696
rect 9310 13617 9321 13663
rect 9375 13617 9386 13663
rect 9555 13654 9601 13665
rect 8865 13571 8911 13582
rect 8848 13544 8865 13546
rect 9049 13571 9095 13582
rect 8911 13544 8928 13546
rect 8773 13424 8860 13544
rect 8916 13424 8928 13544
rect 8848 13422 8865 13424
rect 8773 13124 8865 13244
rect 8911 13422 8928 13424
rect 9032 13244 9049 13246
rect 9233 13571 9279 13582
rect 9216 13544 9233 13546
rect 9417 13571 9463 13582
rect 9279 13544 9296 13546
rect 9216 13424 9228 13544
rect 9284 13424 9296 13544
rect 9216 13422 9233 13424
rect 9095 13244 9112 13246
rect 9032 13124 9044 13244
rect 9100 13124 9112 13244
rect 9032 13122 9049 13124
rect 8865 13086 8911 13097
rect 9095 13122 9112 13124
rect 9049 13086 9095 13097
rect 9279 13422 9296 13424
rect 9400 13244 9417 13246
rect 9538 13544 9555 13546
rect 9601 13544 9618 13546
rect 9538 13423 9550 13544
rect 9606 13423 9618 13544
rect 9538 13421 9555 13423
rect 9463 13244 9480 13246
rect 9400 13124 9412 13244
rect 9468 13124 9480 13244
rect 9400 13122 9417 13124
rect 9233 13086 9279 13097
rect 9463 13122 9480 13124
rect 9417 13086 9463 13097
rect 8942 13048 8953 13051
rect 9007 13048 9018 13051
rect 9126 13048 9137 13051
rect 9191 13048 9202 13051
rect 9310 13048 9321 13051
rect 9375 13048 9386 13051
rect 8727 13003 8773 13014
rect 8940 12992 8952 13048
rect 9008 12992 9020 13048
rect 8940 12978 9020 12992
rect 9124 12992 9136 13048
rect 9192 12992 9204 13048
rect 9124 12978 9204 12992
rect 9308 12992 9320 13048
rect 9376 12992 9388 13048
rect 9601 13421 9618 13423
rect 9555 13003 9601 13014
rect 9308 12978 9388 12992
rect 8940 12898 9020 12900
rect 8552 12842 8952 12898
rect 9008 12842 9020 12898
rect 10038 12899 10094 13919
rect 11196 13907 11276 13919
rect 10702 13868 10788 13872
rect 10702 13812 10714 13868
rect 10770 13812 10788 13868
rect 10702 13800 10788 13812
rect 10213 13655 10259 13666
rect 10428 13664 10504 13697
rect 10428 13618 10439 13664
rect 10493 13618 10504 13664
rect 10612 13664 10688 13697
rect 10612 13618 10623 13664
rect 10677 13618 10688 13664
rect 10796 13664 10872 13697
rect 10796 13618 10807 13664
rect 10861 13618 10872 13664
rect 11041 13655 11087 13666
rect 10351 13572 10397 13583
rect 10334 13545 10351 13547
rect 10535 13572 10581 13583
rect 10397 13545 10414 13547
rect 10259 13425 10346 13545
rect 10402 13425 10414 13545
rect 10334 13423 10351 13425
rect 10259 13125 10351 13245
rect 10397 13423 10414 13425
rect 10518 13245 10535 13247
rect 10719 13572 10765 13583
rect 10702 13545 10719 13547
rect 10903 13572 10949 13583
rect 10765 13545 10782 13547
rect 10702 13425 10714 13545
rect 10770 13425 10782 13545
rect 10702 13423 10719 13425
rect 10581 13245 10598 13247
rect 10518 13125 10530 13245
rect 10586 13125 10598 13245
rect 10518 13123 10535 13125
rect 10351 13087 10397 13098
rect 10581 13123 10598 13125
rect 10535 13087 10581 13098
rect 10765 13423 10782 13425
rect 10886 13245 10903 13247
rect 11024 13545 11041 13547
rect 11087 13545 11104 13547
rect 11024 13424 11036 13545
rect 11092 13424 11104 13545
rect 11024 13422 11041 13424
rect 10949 13245 10966 13247
rect 10886 13125 10898 13245
rect 10954 13125 10966 13245
rect 10886 13123 10903 13125
rect 10719 13087 10765 13098
rect 10949 13123 10966 13125
rect 10903 13087 10949 13098
rect 10428 13049 10439 13052
rect 10493 13049 10504 13052
rect 10612 13049 10623 13052
rect 10677 13049 10688 13052
rect 10796 13049 10807 13052
rect 10861 13049 10872 13052
rect 10213 13004 10259 13015
rect 10426 12993 10438 13049
rect 10494 12993 10506 13049
rect 10426 12979 10506 12993
rect 10610 12993 10622 13049
rect 10678 12993 10690 13049
rect 10610 12979 10690 12993
rect 10794 12993 10806 13049
rect 10862 12993 10874 13049
rect 11087 13422 11104 13424
rect 11041 13004 11087 13015
rect 10794 12979 10874 12993
rect 10426 12899 10506 12901
rect 10038 12843 10438 12899
rect 10494 12843 10506 12899
rect 8940 12840 9020 12842
rect 10426 12841 10506 12843
rect 9124 12782 9204 12784
rect 8416 12726 9136 12782
rect 9192 12726 9204 12782
rect 9124 12724 9204 12726
rect 9453 12782 9533 12784
rect 9720 12783 9790 12794
rect 10610 12783 10690 12785
rect 9720 12782 10622 12783
rect 9453 12726 9465 12782
rect 9521 12726 9722 12782
rect 9778 12727 10622 12782
rect 10678 12727 10690 12783
rect 9778 12726 10038 12727
rect 9453 12724 9533 12726
rect 9720 12716 9790 12726
rect 10610 12725 10690 12727
rect 10939 12783 11019 12785
rect 11382 12783 11452 12793
rect 10939 12727 10951 12783
rect 11007 12727 11384 12783
rect 11440 12727 11452 12783
rect 10939 12725 11019 12727
rect 11382 12715 11452 12727
rect 12458 12782 12514 14029
rect 15414 14027 15494 14029
rect 16080 14085 16150 14087
rect 16500 14085 16556 14815
rect 17392 14813 17472 14815
rect 18122 14815 18890 14871
rect 18946 14815 18958 14871
rect 17024 14721 17104 14735
rect 16811 14699 16857 14710
rect 17024 14665 17036 14721
rect 17092 14665 17104 14721
rect 17208 14721 17288 14735
rect 17208 14665 17220 14721
rect 17276 14665 17288 14721
rect 17392 14721 17472 14735
rect 17392 14665 17404 14721
rect 17460 14665 17472 14721
rect 17639 14699 17685 14710
rect 17026 14662 17037 14665
rect 17091 14662 17102 14665
rect 17210 14662 17221 14665
rect 17275 14662 17286 14665
rect 17394 14662 17405 14665
rect 17459 14662 17470 14665
rect 16949 14616 16995 14627
rect 16857 14442 16949 14616
rect 16949 14431 16995 14442
rect 17133 14616 17179 14627
rect 17133 14431 17179 14442
rect 17317 14616 17363 14627
rect 17501 14616 17547 14627
rect 17484 14589 17501 14591
rect 17547 14589 17564 14591
rect 17484 14469 17496 14589
rect 17552 14469 17564 14589
rect 17484 14467 17501 14469
rect 17317 14431 17363 14442
rect 17547 14467 17564 14469
rect 17501 14431 17547 14442
rect 16811 14214 16857 14359
rect 17026 14350 17037 14396
rect 17091 14350 17102 14396
rect 17026 14317 17102 14350
rect 17210 14350 17221 14396
rect 17275 14350 17286 14396
rect 17210 14317 17286 14350
rect 17394 14350 17405 14396
rect 17459 14350 17470 14396
rect 17394 14317 17470 14350
rect 17639 14214 17685 14359
rect 16799 14202 16879 14214
rect 16799 14146 16811 14202
rect 16867 14146 16879 14202
rect 16799 14134 16879 14146
rect 17617 14202 17695 14214
rect 17617 14146 17629 14202
rect 17685 14146 17695 14202
rect 17617 14134 17695 14146
rect 16080 14029 16092 14085
rect 16148 14029 16556 14085
rect 18122 14085 18178 14815
rect 18878 14813 18958 14815
rect 20542 14815 21446 14871
rect 21502 14815 21514 14871
rect 18510 14721 18590 14735
rect 18297 14699 18343 14710
rect 18510 14665 18522 14721
rect 18578 14665 18590 14721
rect 18694 14721 18774 14735
rect 18694 14665 18706 14721
rect 18762 14665 18774 14721
rect 18878 14721 18958 14735
rect 18878 14665 18890 14721
rect 18946 14665 18958 14721
rect 19125 14699 19171 14710
rect 18512 14662 18523 14665
rect 18577 14662 18588 14665
rect 18696 14662 18707 14665
rect 18761 14662 18772 14665
rect 18880 14662 18891 14665
rect 18945 14662 18956 14665
rect 18435 14616 18481 14627
rect 18343 14442 18435 14616
rect 18435 14431 18481 14442
rect 18619 14616 18665 14627
rect 18619 14431 18665 14442
rect 18803 14616 18849 14627
rect 18987 14616 19033 14627
rect 18970 14589 18987 14591
rect 19033 14589 19050 14591
rect 18970 14469 18982 14589
rect 19038 14469 19050 14589
rect 18970 14467 18987 14469
rect 18803 14431 18849 14442
rect 19033 14467 19050 14469
rect 18987 14431 19033 14442
rect 18297 14214 18343 14359
rect 18512 14350 18523 14396
rect 18577 14350 18588 14396
rect 18512 14317 18588 14350
rect 18696 14350 18707 14396
rect 18761 14350 18772 14396
rect 18696 14317 18772 14350
rect 18880 14350 18891 14396
rect 18945 14350 18956 14396
rect 18880 14317 18956 14350
rect 19125 14214 19171 14359
rect 18285 14202 18365 14214
rect 18285 14146 18297 14202
rect 18353 14146 18365 14202
rect 18285 14134 18365 14146
rect 19103 14202 19181 14214
rect 19103 14146 19115 14202
rect 19171 14146 19181 14202
rect 19103 14134 19181 14146
rect 19456 14085 19536 14095
rect 18122 14029 19468 14085
rect 19524 14029 19536 14085
rect 16080 14017 16150 14029
rect 13938 13974 14008 13976
rect 15238 13975 15318 13977
rect 12594 13918 13940 13974
rect 13996 13918 14008 13974
rect 12594 12898 12650 13918
rect 13938 13906 14008 13918
rect 14080 13919 15250 13975
rect 15306 13919 15318 13975
rect 13258 13867 13344 13871
rect 13258 13811 13270 13867
rect 13326 13811 13344 13867
rect 13258 13799 13344 13811
rect 12769 13654 12815 13665
rect 12984 13663 13060 13696
rect 12984 13617 12995 13663
rect 13049 13617 13060 13663
rect 13168 13663 13244 13696
rect 13168 13617 13179 13663
rect 13233 13617 13244 13663
rect 13352 13663 13428 13696
rect 13352 13617 13363 13663
rect 13417 13617 13428 13663
rect 13597 13654 13643 13665
rect 12907 13571 12953 13582
rect 12890 13544 12907 13546
rect 13091 13571 13137 13582
rect 12953 13544 12970 13546
rect 12815 13424 12902 13544
rect 12958 13424 12970 13544
rect 12890 13422 12907 13424
rect 12815 13124 12907 13244
rect 12953 13422 12970 13424
rect 13074 13244 13091 13246
rect 13275 13571 13321 13582
rect 13258 13544 13275 13546
rect 13459 13571 13505 13582
rect 13321 13544 13338 13546
rect 13258 13424 13270 13544
rect 13326 13424 13338 13544
rect 13258 13422 13275 13424
rect 13137 13244 13154 13246
rect 13074 13124 13086 13244
rect 13142 13124 13154 13244
rect 13074 13122 13091 13124
rect 12907 13086 12953 13097
rect 13137 13122 13154 13124
rect 13091 13086 13137 13097
rect 13321 13422 13338 13424
rect 13442 13244 13459 13246
rect 13580 13544 13597 13546
rect 13643 13544 13660 13546
rect 13580 13423 13592 13544
rect 13648 13423 13660 13544
rect 13580 13421 13597 13423
rect 13505 13244 13522 13246
rect 13442 13124 13454 13244
rect 13510 13124 13522 13244
rect 13442 13122 13459 13124
rect 13275 13086 13321 13097
rect 13505 13122 13522 13124
rect 13459 13086 13505 13097
rect 12984 13048 12995 13051
rect 13049 13048 13060 13051
rect 13168 13048 13179 13051
rect 13233 13048 13244 13051
rect 13352 13048 13363 13051
rect 13417 13048 13428 13051
rect 12769 13003 12815 13014
rect 12982 12992 12994 13048
rect 13050 12992 13062 13048
rect 12982 12978 13062 12992
rect 13166 12992 13178 13048
rect 13234 12992 13246 13048
rect 13166 12978 13246 12992
rect 13350 12992 13362 13048
rect 13418 12992 13430 13048
rect 13643 13421 13660 13423
rect 13597 13003 13643 13014
rect 13350 12978 13430 12992
rect 12982 12898 13062 12900
rect 12594 12842 12994 12898
rect 13050 12842 13062 12898
rect 14080 12899 14136 13919
rect 15238 13907 15318 13919
rect 14744 13868 14830 13872
rect 14744 13812 14756 13868
rect 14812 13812 14830 13868
rect 14744 13800 14830 13812
rect 14255 13655 14301 13666
rect 14470 13664 14546 13697
rect 14470 13618 14481 13664
rect 14535 13618 14546 13664
rect 14654 13664 14730 13697
rect 14654 13618 14665 13664
rect 14719 13618 14730 13664
rect 14838 13664 14914 13697
rect 14838 13618 14849 13664
rect 14903 13618 14914 13664
rect 15083 13655 15129 13666
rect 14393 13572 14439 13583
rect 14376 13545 14393 13547
rect 14577 13572 14623 13583
rect 14439 13545 14456 13547
rect 14301 13425 14388 13545
rect 14444 13425 14456 13545
rect 14376 13423 14393 13425
rect 14301 13125 14393 13245
rect 14439 13423 14456 13425
rect 14560 13245 14577 13247
rect 14761 13572 14807 13583
rect 14744 13545 14761 13547
rect 14945 13572 14991 13583
rect 14807 13545 14824 13547
rect 14744 13425 14756 13545
rect 14812 13425 14824 13545
rect 14744 13423 14761 13425
rect 14623 13245 14640 13247
rect 14560 13125 14572 13245
rect 14628 13125 14640 13245
rect 14560 13123 14577 13125
rect 14393 13087 14439 13098
rect 14623 13123 14640 13125
rect 14577 13087 14623 13098
rect 14807 13423 14824 13425
rect 14928 13245 14945 13247
rect 15066 13545 15083 13547
rect 15129 13545 15146 13547
rect 15066 13424 15078 13545
rect 15134 13424 15146 13545
rect 15066 13422 15083 13424
rect 14991 13245 15008 13247
rect 14928 13125 14940 13245
rect 14996 13125 15008 13245
rect 14928 13123 14945 13125
rect 14761 13087 14807 13098
rect 14991 13123 15008 13125
rect 14945 13087 14991 13098
rect 14470 13049 14481 13052
rect 14535 13049 14546 13052
rect 14654 13049 14665 13052
rect 14719 13049 14730 13052
rect 14838 13049 14849 13052
rect 14903 13049 14914 13052
rect 14255 13004 14301 13015
rect 14468 12993 14480 13049
rect 14536 12993 14548 13049
rect 14468 12979 14548 12993
rect 14652 12993 14664 13049
rect 14720 12993 14732 13049
rect 14652 12979 14732 12993
rect 14836 12993 14848 13049
rect 14904 12993 14916 13049
rect 15129 13422 15146 13424
rect 15083 13004 15129 13015
rect 14836 12979 14916 12993
rect 14468 12899 14548 12901
rect 14080 12843 14480 12899
rect 14536 12843 14548 12899
rect 12982 12840 13062 12842
rect 14468 12841 14548 12843
rect 13166 12782 13246 12784
rect 12458 12726 13178 12782
rect 13234 12726 13246 12782
rect 13166 12724 13246 12726
rect 13495 12782 13575 12784
rect 13762 12783 13832 12794
rect 14652 12783 14732 12785
rect 13762 12782 14664 12783
rect 13495 12726 13507 12782
rect 13563 12726 13764 12782
rect 13820 12727 14664 12782
rect 14720 12727 14732 12783
rect 13820 12726 14080 12727
rect 13495 12724 13575 12726
rect 13762 12716 13832 12726
rect 14652 12725 14732 12727
rect 14981 12783 15061 12785
rect 15424 12783 15494 12793
rect 14981 12727 14993 12783
rect 15049 12727 15426 12783
rect 15482 12727 15494 12783
rect 14981 12725 15061 12727
rect 15424 12715 15494 12727
rect 16500 12782 16556 14029
rect 19456 14027 19536 14029
rect 20122 14085 20192 14087
rect 20542 14085 20598 14815
rect 21434 14813 21514 14815
rect 22164 14815 22932 14871
rect 22988 14815 23000 14871
rect 21066 14721 21146 14735
rect 20853 14699 20899 14710
rect 21066 14665 21078 14721
rect 21134 14665 21146 14721
rect 21250 14721 21330 14735
rect 21250 14665 21262 14721
rect 21318 14665 21330 14721
rect 21434 14721 21514 14735
rect 21434 14665 21446 14721
rect 21502 14665 21514 14721
rect 21681 14699 21727 14710
rect 21068 14662 21079 14665
rect 21133 14662 21144 14665
rect 21252 14662 21263 14665
rect 21317 14662 21328 14665
rect 21436 14662 21447 14665
rect 21501 14662 21512 14665
rect 20991 14616 21037 14627
rect 20899 14442 20991 14616
rect 20991 14431 21037 14442
rect 21175 14616 21221 14627
rect 21175 14431 21221 14442
rect 21359 14616 21405 14627
rect 21543 14616 21589 14627
rect 21526 14589 21543 14591
rect 21589 14589 21606 14591
rect 21526 14469 21538 14589
rect 21594 14469 21606 14589
rect 21526 14467 21543 14469
rect 21359 14431 21405 14442
rect 21589 14467 21606 14469
rect 21543 14431 21589 14442
rect 20853 14214 20899 14359
rect 21068 14350 21079 14396
rect 21133 14350 21144 14396
rect 21068 14317 21144 14350
rect 21252 14350 21263 14396
rect 21317 14350 21328 14396
rect 21252 14317 21328 14350
rect 21436 14350 21447 14396
rect 21501 14350 21512 14396
rect 21436 14317 21512 14350
rect 21681 14214 21727 14359
rect 20841 14202 20921 14214
rect 20841 14146 20853 14202
rect 20909 14146 20921 14202
rect 20841 14134 20921 14146
rect 21659 14202 21737 14214
rect 21659 14146 21671 14202
rect 21727 14146 21737 14202
rect 21659 14134 21737 14146
rect 20122 14029 20134 14085
rect 20190 14029 20598 14085
rect 22164 14085 22220 14815
rect 22920 14813 23000 14815
rect 24584 14815 25488 14871
rect 25544 14815 25556 14871
rect 22552 14721 22632 14735
rect 22339 14699 22385 14710
rect 22552 14665 22564 14721
rect 22620 14665 22632 14721
rect 22736 14721 22816 14735
rect 22736 14665 22748 14721
rect 22804 14665 22816 14721
rect 22920 14721 23000 14735
rect 22920 14665 22932 14721
rect 22988 14665 23000 14721
rect 23167 14699 23213 14710
rect 22554 14662 22565 14665
rect 22619 14662 22630 14665
rect 22738 14662 22749 14665
rect 22803 14662 22814 14665
rect 22922 14662 22933 14665
rect 22987 14662 22998 14665
rect 22477 14616 22523 14627
rect 22385 14442 22477 14616
rect 22477 14431 22523 14442
rect 22661 14616 22707 14627
rect 22661 14431 22707 14442
rect 22845 14616 22891 14627
rect 23029 14616 23075 14627
rect 23012 14589 23029 14591
rect 23075 14589 23092 14591
rect 23012 14469 23024 14589
rect 23080 14469 23092 14589
rect 23012 14467 23029 14469
rect 22845 14431 22891 14442
rect 23075 14467 23092 14469
rect 23029 14431 23075 14442
rect 22339 14214 22385 14359
rect 22554 14350 22565 14396
rect 22619 14350 22630 14396
rect 22554 14317 22630 14350
rect 22738 14350 22749 14396
rect 22803 14350 22814 14396
rect 22738 14317 22814 14350
rect 22922 14350 22933 14396
rect 22987 14350 22998 14396
rect 22922 14317 22998 14350
rect 23167 14214 23213 14359
rect 22327 14202 22407 14214
rect 22327 14146 22339 14202
rect 22395 14146 22407 14202
rect 22327 14134 22407 14146
rect 23145 14202 23223 14214
rect 23145 14146 23157 14202
rect 23213 14146 23223 14202
rect 23145 14134 23223 14146
rect 23498 14085 23578 14095
rect 22164 14029 23510 14085
rect 23566 14029 23578 14085
rect 20122 14017 20192 14029
rect 17980 13974 18050 13976
rect 19280 13975 19360 13977
rect 16636 13918 17982 13974
rect 18038 13918 18050 13974
rect 16636 12898 16692 13918
rect 17980 13906 18050 13918
rect 18122 13919 19292 13975
rect 19348 13919 19360 13975
rect 17300 13867 17386 13871
rect 17300 13811 17312 13867
rect 17368 13811 17386 13867
rect 17300 13799 17386 13811
rect 16811 13654 16857 13665
rect 17026 13663 17102 13696
rect 17026 13617 17037 13663
rect 17091 13617 17102 13663
rect 17210 13663 17286 13696
rect 17210 13617 17221 13663
rect 17275 13617 17286 13663
rect 17394 13663 17470 13696
rect 17394 13617 17405 13663
rect 17459 13617 17470 13663
rect 17639 13654 17685 13665
rect 16949 13571 16995 13582
rect 16932 13544 16949 13546
rect 17133 13571 17179 13582
rect 16995 13544 17012 13546
rect 16857 13424 16944 13544
rect 17000 13424 17012 13544
rect 16932 13422 16949 13424
rect 16857 13124 16949 13244
rect 16995 13422 17012 13424
rect 17116 13244 17133 13246
rect 17317 13571 17363 13582
rect 17300 13544 17317 13546
rect 17501 13571 17547 13582
rect 17363 13544 17380 13546
rect 17300 13424 17312 13544
rect 17368 13424 17380 13544
rect 17300 13422 17317 13424
rect 17179 13244 17196 13246
rect 17116 13124 17128 13244
rect 17184 13124 17196 13244
rect 17116 13122 17133 13124
rect 16949 13086 16995 13097
rect 17179 13122 17196 13124
rect 17133 13086 17179 13097
rect 17363 13422 17380 13424
rect 17484 13244 17501 13246
rect 17622 13544 17639 13546
rect 17685 13544 17702 13546
rect 17622 13423 17634 13544
rect 17690 13423 17702 13544
rect 17622 13421 17639 13423
rect 17547 13244 17564 13246
rect 17484 13124 17496 13244
rect 17552 13124 17564 13244
rect 17484 13122 17501 13124
rect 17317 13086 17363 13097
rect 17547 13122 17564 13124
rect 17501 13086 17547 13097
rect 17026 13048 17037 13051
rect 17091 13048 17102 13051
rect 17210 13048 17221 13051
rect 17275 13048 17286 13051
rect 17394 13048 17405 13051
rect 17459 13048 17470 13051
rect 16811 13003 16857 13014
rect 17024 12992 17036 13048
rect 17092 12992 17104 13048
rect 17024 12978 17104 12992
rect 17208 12992 17220 13048
rect 17276 12992 17288 13048
rect 17208 12978 17288 12992
rect 17392 12992 17404 13048
rect 17460 12992 17472 13048
rect 17685 13421 17702 13423
rect 17639 13003 17685 13014
rect 17392 12978 17472 12992
rect 17024 12898 17104 12900
rect 16636 12842 17036 12898
rect 17092 12842 17104 12898
rect 18122 12899 18178 13919
rect 19280 13907 19360 13919
rect 18786 13868 18872 13872
rect 18786 13812 18798 13868
rect 18854 13812 18872 13868
rect 18786 13800 18872 13812
rect 18297 13655 18343 13666
rect 18512 13664 18588 13697
rect 18512 13618 18523 13664
rect 18577 13618 18588 13664
rect 18696 13664 18772 13697
rect 18696 13618 18707 13664
rect 18761 13618 18772 13664
rect 18880 13664 18956 13697
rect 18880 13618 18891 13664
rect 18945 13618 18956 13664
rect 19125 13655 19171 13666
rect 18435 13572 18481 13583
rect 18418 13545 18435 13547
rect 18619 13572 18665 13583
rect 18481 13545 18498 13547
rect 18343 13425 18430 13545
rect 18486 13425 18498 13545
rect 18418 13423 18435 13425
rect 18343 13125 18435 13245
rect 18481 13423 18498 13425
rect 18602 13245 18619 13247
rect 18803 13572 18849 13583
rect 18786 13545 18803 13547
rect 18987 13572 19033 13583
rect 18849 13545 18866 13547
rect 18786 13425 18798 13545
rect 18854 13425 18866 13545
rect 18786 13423 18803 13425
rect 18665 13245 18682 13247
rect 18602 13125 18614 13245
rect 18670 13125 18682 13245
rect 18602 13123 18619 13125
rect 18435 13087 18481 13098
rect 18665 13123 18682 13125
rect 18619 13087 18665 13098
rect 18849 13423 18866 13425
rect 18970 13245 18987 13247
rect 19108 13545 19125 13547
rect 19171 13545 19188 13547
rect 19108 13424 19120 13545
rect 19176 13424 19188 13545
rect 19108 13422 19125 13424
rect 19033 13245 19050 13247
rect 18970 13125 18982 13245
rect 19038 13125 19050 13245
rect 18970 13123 18987 13125
rect 18803 13087 18849 13098
rect 19033 13123 19050 13125
rect 18987 13087 19033 13098
rect 18512 13049 18523 13052
rect 18577 13049 18588 13052
rect 18696 13049 18707 13052
rect 18761 13049 18772 13052
rect 18880 13049 18891 13052
rect 18945 13049 18956 13052
rect 18297 13004 18343 13015
rect 18510 12993 18522 13049
rect 18578 12993 18590 13049
rect 18510 12979 18590 12993
rect 18694 12993 18706 13049
rect 18762 12993 18774 13049
rect 18694 12979 18774 12993
rect 18878 12993 18890 13049
rect 18946 12993 18958 13049
rect 19171 13422 19188 13424
rect 19125 13004 19171 13015
rect 18878 12979 18958 12993
rect 18510 12899 18590 12901
rect 18122 12843 18522 12899
rect 18578 12843 18590 12899
rect 17024 12840 17104 12842
rect 18510 12841 18590 12843
rect 17208 12782 17288 12784
rect 16500 12726 17220 12782
rect 17276 12726 17288 12782
rect 17208 12724 17288 12726
rect 17537 12782 17617 12784
rect 17804 12783 17874 12794
rect 18694 12783 18774 12785
rect 17804 12782 18706 12783
rect 17537 12726 17549 12782
rect 17605 12726 17806 12782
rect 17862 12727 18706 12782
rect 18762 12727 18774 12783
rect 17862 12726 18122 12727
rect 17537 12724 17617 12726
rect 17804 12716 17874 12726
rect 18694 12725 18774 12727
rect 19023 12783 19103 12785
rect 19466 12783 19536 12793
rect 19023 12727 19035 12783
rect 19091 12727 19468 12783
rect 19524 12727 19536 12783
rect 19023 12725 19103 12727
rect 19466 12715 19536 12727
rect 20542 12782 20598 14029
rect 23498 14027 23578 14029
rect 24164 14085 24234 14087
rect 24584 14085 24640 14815
rect 25476 14813 25556 14815
rect 26206 14815 26974 14871
rect 27030 14815 27042 14871
rect 25108 14721 25188 14735
rect 24895 14699 24941 14710
rect 25108 14665 25120 14721
rect 25176 14665 25188 14721
rect 25292 14721 25372 14735
rect 25292 14665 25304 14721
rect 25360 14665 25372 14721
rect 25476 14721 25556 14735
rect 25476 14665 25488 14721
rect 25544 14665 25556 14721
rect 25723 14699 25769 14710
rect 25110 14662 25121 14665
rect 25175 14662 25186 14665
rect 25294 14662 25305 14665
rect 25359 14662 25370 14665
rect 25478 14662 25489 14665
rect 25543 14662 25554 14665
rect 25033 14616 25079 14627
rect 24941 14442 25033 14616
rect 25033 14431 25079 14442
rect 25217 14616 25263 14627
rect 25217 14431 25263 14442
rect 25401 14616 25447 14627
rect 25585 14616 25631 14627
rect 25568 14589 25585 14591
rect 25631 14589 25648 14591
rect 25568 14469 25580 14589
rect 25636 14469 25648 14589
rect 25568 14467 25585 14469
rect 25401 14431 25447 14442
rect 25631 14467 25648 14469
rect 25585 14431 25631 14442
rect 24895 14214 24941 14359
rect 25110 14350 25121 14396
rect 25175 14350 25186 14396
rect 25110 14317 25186 14350
rect 25294 14350 25305 14396
rect 25359 14350 25370 14396
rect 25294 14317 25370 14350
rect 25478 14350 25489 14396
rect 25543 14350 25554 14396
rect 25478 14317 25554 14350
rect 25723 14214 25769 14359
rect 24883 14202 24963 14214
rect 24883 14146 24895 14202
rect 24951 14146 24963 14202
rect 24883 14134 24963 14146
rect 25701 14202 25779 14214
rect 25701 14146 25713 14202
rect 25769 14146 25779 14202
rect 25701 14134 25779 14146
rect 24164 14029 24176 14085
rect 24232 14029 24640 14085
rect 26206 14085 26262 14815
rect 26962 14813 27042 14815
rect 28626 14815 29530 14871
rect 29586 14815 29598 14871
rect 26594 14721 26674 14735
rect 26381 14699 26427 14710
rect 26594 14665 26606 14721
rect 26662 14665 26674 14721
rect 26778 14721 26858 14735
rect 26778 14665 26790 14721
rect 26846 14665 26858 14721
rect 26962 14721 27042 14735
rect 26962 14665 26974 14721
rect 27030 14665 27042 14721
rect 27209 14699 27255 14710
rect 26596 14662 26607 14665
rect 26661 14662 26672 14665
rect 26780 14662 26791 14665
rect 26845 14662 26856 14665
rect 26964 14662 26975 14665
rect 27029 14662 27040 14665
rect 26519 14616 26565 14627
rect 26427 14442 26519 14616
rect 26519 14431 26565 14442
rect 26703 14616 26749 14627
rect 26703 14431 26749 14442
rect 26887 14616 26933 14627
rect 27071 14616 27117 14627
rect 27054 14589 27071 14591
rect 27117 14589 27134 14591
rect 27054 14469 27066 14589
rect 27122 14469 27134 14589
rect 27054 14467 27071 14469
rect 26887 14431 26933 14442
rect 27117 14467 27134 14469
rect 27071 14431 27117 14442
rect 26381 14214 26427 14359
rect 26596 14350 26607 14396
rect 26661 14350 26672 14396
rect 26596 14317 26672 14350
rect 26780 14350 26791 14396
rect 26845 14350 26856 14396
rect 26780 14317 26856 14350
rect 26964 14350 26975 14396
rect 27029 14350 27040 14396
rect 26964 14317 27040 14350
rect 27209 14214 27255 14359
rect 26369 14202 26449 14214
rect 26369 14146 26381 14202
rect 26437 14146 26449 14202
rect 26369 14134 26449 14146
rect 27187 14202 27265 14214
rect 27187 14146 27199 14202
rect 27255 14146 27265 14202
rect 27187 14134 27265 14146
rect 27540 14085 27620 14095
rect 26206 14029 27552 14085
rect 27608 14029 27620 14085
rect 24164 14017 24234 14029
rect 22022 13974 22092 13976
rect 23322 13975 23402 13977
rect 20678 13918 22024 13974
rect 22080 13918 22092 13974
rect 20678 12898 20734 13918
rect 22022 13906 22092 13918
rect 22164 13919 23334 13975
rect 23390 13919 23402 13975
rect 21342 13867 21428 13871
rect 21342 13811 21354 13867
rect 21410 13811 21428 13867
rect 21342 13799 21428 13811
rect 20853 13654 20899 13665
rect 21068 13663 21144 13696
rect 21068 13617 21079 13663
rect 21133 13617 21144 13663
rect 21252 13663 21328 13696
rect 21252 13617 21263 13663
rect 21317 13617 21328 13663
rect 21436 13663 21512 13696
rect 21436 13617 21447 13663
rect 21501 13617 21512 13663
rect 21681 13654 21727 13665
rect 20991 13571 21037 13582
rect 20974 13544 20991 13546
rect 21175 13571 21221 13582
rect 21037 13544 21054 13546
rect 20899 13424 20986 13544
rect 21042 13424 21054 13544
rect 20974 13422 20991 13424
rect 20899 13124 20991 13244
rect 21037 13422 21054 13424
rect 21158 13244 21175 13246
rect 21359 13571 21405 13582
rect 21342 13544 21359 13546
rect 21543 13571 21589 13582
rect 21405 13544 21422 13546
rect 21342 13424 21354 13544
rect 21410 13424 21422 13544
rect 21342 13422 21359 13424
rect 21221 13244 21238 13246
rect 21158 13124 21170 13244
rect 21226 13124 21238 13244
rect 21158 13122 21175 13124
rect 20991 13086 21037 13097
rect 21221 13122 21238 13124
rect 21175 13086 21221 13097
rect 21405 13422 21422 13424
rect 21526 13244 21543 13246
rect 21664 13544 21681 13546
rect 21727 13544 21744 13546
rect 21664 13423 21676 13544
rect 21732 13423 21744 13544
rect 21664 13421 21681 13423
rect 21589 13244 21606 13246
rect 21526 13124 21538 13244
rect 21594 13124 21606 13244
rect 21526 13122 21543 13124
rect 21359 13086 21405 13097
rect 21589 13122 21606 13124
rect 21543 13086 21589 13097
rect 21068 13048 21079 13051
rect 21133 13048 21144 13051
rect 21252 13048 21263 13051
rect 21317 13048 21328 13051
rect 21436 13048 21447 13051
rect 21501 13048 21512 13051
rect 20853 13003 20899 13014
rect 21066 12992 21078 13048
rect 21134 12992 21146 13048
rect 21066 12978 21146 12992
rect 21250 12992 21262 13048
rect 21318 12992 21330 13048
rect 21250 12978 21330 12992
rect 21434 12992 21446 13048
rect 21502 12992 21514 13048
rect 21727 13421 21744 13423
rect 21681 13003 21727 13014
rect 21434 12978 21514 12992
rect 21066 12898 21146 12900
rect 20678 12842 21078 12898
rect 21134 12842 21146 12898
rect 22164 12899 22220 13919
rect 23322 13907 23402 13919
rect 22828 13868 22914 13872
rect 22828 13812 22840 13868
rect 22896 13812 22914 13868
rect 22828 13800 22914 13812
rect 22339 13655 22385 13666
rect 22554 13664 22630 13697
rect 22554 13618 22565 13664
rect 22619 13618 22630 13664
rect 22738 13664 22814 13697
rect 22738 13618 22749 13664
rect 22803 13618 22814 13664
rect 22922 13664 22998 13697
rect 22922 13618 22933 13664
rect 22987 13618 22998 13664
rect 23167 13655 23213 13666
rect 22477 13572 22523 13583
rect 22460 13545 22477 13547
rect 22661 13572 22707 13583
rect 22523 13545 22540 13547
rect 22385 13425 22472 13545
rect 22528 13425 22540 13545
rect 22460 13423 22477 13425
rect 22385 13125 22477 13245
rect 22523 13423 22540 13425
rect 22644 13245 22661 13247
rect 22845 13572 22891 13583
rect 22828 13545 22845 13547
rect 23029 13572 23075 13583
rect 22891 13545 22908 13547
rect 22828 13425 22840 13545
rect 22896 13425 22908 13545
rect 22828 13423 22845 13425
rect 22707 13245 22724 13247
rect 22644 13125 22656 13245
rect 22712 13125 22724 13245
rect 22644 13123 22661 13125
rect 22477 13087 22523 13098
rect 22707 13123 22724 13125
rect 22661 13087 22707 13098
rect 22891 13423 22908 13425
rect 23012 13245 23029 13247
rect 23150 13545 23167 13547
rect 23213 13545 23230 13547
rect 23150 13424 23162 13545
rect 23218 13424 23230 13545
rect 23150 13422 23167 13424
rect 23075 13245 23092 13247
rect 23012 13125 23024 13245
rect 23080 13125 23092 13245
rect 23012 13123 23029 13125
rect 22845 13087 22891 13098
rect 23075 13123 23092 13125
rect 23029 13087 23075 13098
rect 22554 13049 22565 13052
rect 22619 13049 22630 13052
rect 22738 13049 22749 13052
rect 22803 13049 22814 13052
rect 22922 13049 22933 13052
rect 22987 13049 22998 13052
rect 22339 13004 22385 13015
rect 22552 12993 22564 13049
rect 22620 12993 22632 13049
rect 22552 12979 22632 12993
rect 22736 12993 22748 13049
rect 22804 12993 22816 13049
rect 22736 12979 22816 12993
rect 22920 12993 22932 13049
rect 22988 12993 23000 13049
rect 23213 13422 23230 13424
rect 23167 13004 23213 13015
rect 22920 12979 23000 12993
rect 22552 12899 22632 12901
rect 22164 12843 22564 12899
rect 22620 12843 22632 12899
rect 21066 12840 21146 12842
rect 22552 12841 22632 12843
rect 21250 12782 21330 12784
rect 20542 12726 21262 12782
rect 21318 12726 21330 12782
rect 21250 12724 21330 12726
rect 21579 12782 21659 12784
rect 21846 12783 21916 12794
rect 22736 12783 22816 12785
rect 21846 12782 22748 12783
rect 21579 12726 21591 12782
rect 21647 12726 21848 12782
rect 21904 12727 22748 12782
rect 22804 12727 22816 12783
rect 21904 12726 22164 12727
rect 21579 12724 21659 12726
rect 21846 12716 21916 12726
rect 22736 12725 22816 12727
rect 23065 12783 23145 12785
rect 23508 12783 23578 12793
rect 23065 12727 23077 12783
rect 23133 12727 23510 12783
rect 23566 12727 23578 12783
rect 23065 12725 23145 12727
rect 23508 12715 23578 12727
rect 24584 12782 24640 14029
rect 27540 14027 27620 14029
rect 28162 14085 28240 14097
rect 28626 14085 28682 14815
rect 29518 14813 29598 14815
rect 30248 14815 31016 14871
rect 31072 14815 31084 14871
rect 29150 14721 29230 14735
rect 28937 14699 28983 14710
rect 29150 14665 29162 14721
rect 29218 14665 29230 14721
rect 29334 14721 29414 14735
rect 29334 14665 29346 14721
rect 29402 14665 29414 14721
rect 29518 14721 29598 14735
rect 29518 14665 29530 14721
rect 29586 14665 29598 14721
rect 29765 14699 29811 14710
rect 29152 14662 29163 14665
rect 29217 14662 29228 14665
rect 29336 14662 29347 14665
rect 29401 14662 29412 14665
rect 29520 14662 29531 14665
rect 29585 14662 29596 14665
rect 29075 14616 29121 14627
rect 28983 14442 29075 14616
rect 29075 14431 29121 14442
rect 29259 14616 29305 14627
rect 29259 14431 29305 14442
rect 29443 14616 29489 14627
rect 29627 14616 29673 14627
rect 29610 14589 29627 14591
rect 29673 14589 29690 14591
rect 29610 14469 29622 14589
rect 29678 14469 29690 14589
rect 29610 14467 29627 14469
rect 29443 14431 29489 14442
rect 29673 14467 29690 14469
rect 29627 14431 29673 14442
rect 28937 14214 28983 14359
rect 29152 14350 29163 14396
rect 29217 14350 29228 14396
rect 29152 14317 29228 14350
rect 29336 14350 29347 14396
rect 29401 14350 29412 14396
rect 29336 14317 29412 14350
rect 29520 14350 29531 14396
rect 29585 14350 29596 14396
rect 29520 14317 29596 14350
rect 29765 14214 29811 14359
rect 28925 14202 29005 14214
rect 28925 14146 28937 14202
rect 28993 14146 29005 14202
rect 28925 14134 29005 14146
rect 29743 14202 29821 14214
rect 29743 14146 29755 14202
rect 29811 14146 29821 14202
rect 29743 14134 29821 14146
rect 28162 14029 28173 14085
rect 28229 14029 28682 14085
rect 30248 14085 30304 14815
rect 31004 14813 31084 14815
rect 30636 14721 30716 14735
rect 30423 14699 30469 14710
rect 30636 14665 30648 14721
rect 30704 14665 30716 14721
rect 30820 14721 30900 14735
rect 30820 14665 30832 14721
rect 30888 14665 30900 14721
rect 31004 14721 31084 14735
rect 31004 14665 31016 14721
rect 31072 14665 31084 14721
rect 31251 14699 31297 14710
rect 30638 14662 30649 14665
rect 30703 14662 30714 14665
rect 30822 14662 30833 14665
rect 30887 14662 30898 14665
rect 31006 14662 31017 14665
rect 31071 14662 31082 14665
rect 30561 14616 30607 14627
rect 30469 14442 30561 14616
rect 30561 14431 30607 14442
rect 30745 14616 30791 14627
rect 30745 14431 30791 14442
rect 30929 14616 30975 14627
rect 31113 14616 31159 14627
rect 31096 14589 31113 14591
rect 31159 14589 31176 14591
rect 31096 14469 31108 14589
rect 31164 14469 31176 14589
rect 31096 14467 31113 14469
rect 30929 14431 30975 14442
rect 31159 14467 31176 14469
rect 31113 14431 31159 14442
rect 30423 14214 30469 14359
rect 30638 14350 30649 14396
rect 30703 14350 30714 14396
rect 30638 14317 30714 14350
rect 30822 14350 30833 14396
rect 30887 14350 30898 14396
rect 30822 14317 30898 14350
rect 31006 14350 31017 14396
rect 31071 14350 31082 14396
rect 31006 14317 31082 14350
rect 31251 14214 31297 14359
rect 30411 14202 30491 14214
rect 30411 14146 30423 14202
rect 30479 14146 30491 14202
rect 30411 14134 30491 14146
rect 31229 14202 31307 14214
rect 31229 14146 31241 14202
rect 31297 14146 31307 14202
rect 31229 14134 31307 14146
rect 31582 14085 31662 14095
rect 30248 14029 31594 14085
rect 31650 14029 31662 14085
rect 28162 14017 28240 14029
rect 26064 13974 26134 13976
rect 27364 13975 27444 13977
rect 24720 13918 26066 13974
rect 26122 13918 26134 13974
rect 24720 12898 24776 13918
rect 26064 13906 26134 13918
rect 26206 13919 27376 13975
rect 27432 13919 27444 13975
rect 25384 13867 25470 13871
rect 25384 13811 25396 13867
rect 25452 13811 25470 13867
rect 25384 13799 25470 13811
rect 24895 13654 24941 13665
rect 25110 13663 25186 13696
rect 25110 13617 25121 13663
rect 25175 13617 25186 13663
rect 25294 13663 25370 13696
rect 25294 13617 25305 13663
rect 25359 13617 25370 13663
rect 25478 13663 25554 13696
rect 25478 13617 25489 13663
rect 25543 13617 25554 13663
rect 25723 13654 25769 13665
rect 25033 13571 25079 13582
rect 25016 13544 25033 13546
rect 25217 13571 25263 13582
rect 25079 13544 25096 13546
rect 24941 13424 25028 13544
rect 25084 13424 25096 13544
rect 25016 13422 25033 13424
rect 24941 13124 25033 13244
rect 25079 13422 25096 13424
rect 25200 13244 25217 13246
rect 25401 13571 25447 13582
rect 25384 13544 25401 13546
rect 25585 13571 25631 13582
rect 25447 13544 25464 13546
rect 25384 13424 25396 13544
rect 25452 13424 25464 13544
rect 25384 13422 25401 13424
rect 25263 13244 25280 13246
rect 25200 13124 25212 13244
rect 25268 13124 25280 13244
rect 25200 13122 25217 13124
rect 25033 13086 25079 13097
rect 25263 13122 25280 13124
rect 25217 13086 25263 13097
rect 25447 13422 25464 13424
rect 25568 13244 25585 13246
rect 25706 13544 25723 13546
rect 25769 13544 25786 13546
rect 25706 13423 25718 13544
rect 25774 13423 25786 13544
rect 25706 13421 25723 13423
rect 25631 13244 25648 13246
rect 25568 13124 25580 13244
rect 25636 13124 25648 13244
rect 25568 13122 25585 13124
rect 25401 13086 25447 13097
rect 25631 13122 25648 13124
rect 25585 13086 25631 13097
rect 25110 13048 25121 13051
rect 25175 13048 25186 13051
rect 25294 13048 25305 13051
rect 25359 13048 25370 13051
rect 25478 13048 25489 13051
rect 25543 13048 25554 13051
rect 24895 13003 24941 13014
rect 25108 12992 25120 13048
rect 25176 12992 25188 13048
rect 25108 12978 25188 12992
rect 25292 12992 25304 13048
rect 25360 12992 25372 13048
rect 25292 12978 25372 12992
rect 25476 12992 25488 13048
rect 25544 12992 25556 13048
rect 25769 13421 25786 13423
rect 25723 13003 25769 13014
rect 25476 12978 25556 12992
rect 25108 12898 25188 12900
rect 24720 12842 25120 12898
rect 25176 12842 25188 12898
rect 26206 12899 26262 13919
rect 27364 13907 27444 13919
rect 26870 13868 26956 13872
rect 26870 13812 26882 13868
rect 26938 13812 26956 13868
rect 26870 13800 26956 13812
rect 26381 13655 26427 13666
rect 26596 13664 26672 13697
rect 26596 13618 26607 13664
rect 26661 13618 26672 13664
rect 26780 13664 26856 13697
rect 26780 13618 26791 13664
rect 26845 13618 26856 13664
rect 26964 13664 27040 13697
rect 26964 13618 26975 13664
rect 27029 13618 27040 13664
rect 27209 13655 27255 13666
rect 26519 13572 26565 13583
rect 26502 13545 26519 13547
rect 26703 13572 26749 13583
rect 26565 13545 26582 13547
rect 26427 13425 26514 13545
rect 26570 13425 26582 13545
rect 26502 13423 26519 13425
rect 26427 13125 26519 13245
rect 26565 13423 26582 13425
rect 26686 13245 26703 13247
rect 26887 13572 26933 13583
rect 26870 13545 26887 13547
rect 27071 13572 27117 13583
rect 26933 13545 26950 13547
rect 26870 13425 26882 13545
rect 26938 13425 26950 13545
rect 26870 13423 26887 13425
rect 26749 13245 26766 13247
rect 26686 13125 26698 13245
rect 26754 13125 26766 13245
rect 26686 13123 26703 13125
rect 26519 13087 26565 13098
rect 26749 13123 26766 13125
rect 26703 13087 26749 13098
rect 26933 13423 26950 13425
rect 27054 13245 27071 13247
rect 27192 13545 27209 13547
rect 27255 13545 27272 13547
rect 27192 13424 27204 13545
rect 27260 13424 27272 13545
rect 27192 13422 27209 13424
rect 27117 13245 27134 13247
rect 27054 13125 27066 13245
rect 27122 13125 27134 13245
rect 27054 13123 27071 13125
rect 26887 13087 26933 13098
rect 27117 13123 27134 13125
rect 27071 13087 27117 13098
rect 26596 13049 26607 13052
rect 26661 13049 26672 13052
rect 26780 13049 26791 13052
rect 26845 13049 26856 13052
rect 26964 13049 26975 13052
rect 27029 13049 27040 13052
rect 26381 13004 26427 13015
rect 26594 12993 26606 13049
rect 26662 12993 26674 13049
rect 26594 12979 26674 12993
rect 26778 12993 26790 13049
rect 26846 12993 26858 13049
rect 26778 12979 26858 12993
rect 26962 12993 26974 13049
rect 27030 12993 27042 13049
rect 27255 13422 27272 13424
rect 27209 13004 27255 13015
rect 26962 12979 27042 12993
rect 26594 12899 26674 12901
rect 26206 12843 26606 12899
rect 26662 12843 26674 12899
rect 25108 12840 25188 12842
rect 26594 12841 26674 12843
rect 25292 12782 25372 12784
rect 24584 12726 25304 12782
rect 25360 12726 25372 12782
rect 25292 12724 25372 12726
rect 25621 12782 25701 12784
rect 25888 12783 25958 12794
rect 26778 12783 26858 12785
rect 25888 12782 26790 12783
rect 25621 12726 25633 12782
rect 25689 12726 25890 12782
rect 25946 12727 26790 12782
rect 26846 12727 26858 12783
rect 25946 12726 26206 12727
rect 25621 12724 25701 12726
rect 25888 12716 25958 12726
rect 26778 12725 26858 12727
rect 27107 12783 27187 12785
rect 27550 12783 27620 12793
rect 27107 12727 27119 12783
rect 27175 12727 27552 12783
rect 27608 12727 27620 12783
rect 27107 12725 27187 12727
rect 27550 12715 27620 12727
rect 28626 12782 28682 14029
rect 31582 14027 31662 14029
rect 30106 13974 30176 13976
rect 31406 13975 31486 13977
rect 28762 13918 30108 13974
rect 30164 13918 30176 13974
rect 28762 12898 28818 13918
rect 30106 13906 30176 13918
rect 30248 13919 31418 13975
rect 31474 13919 31486 13975
rect 29426 13867 29512 13871
rect 29426 13811 29438 13867
rect 29494 13811 29512 13867
rect 29426 13799 29512 13811
rect 28937 13654 28983 13665
rect 29152 13663 29228 13696
rect 29152 13617 29163 13663
rect 29217 13617 29228 13663
rect 29336 13663 29412 13696
rect 29336 13617 29347 13663
rect 29401 13617 29412 13663
rect 29520 13663 29596 13696
rect 29520 13617 29531 13663
rect 29585 13617 29596 13663
rect 29765 13654 29811 13665
rect 29075 13571 29121 13582
rect 29058 13544 29075 13546
rect 29259 13571 29305 13582
rect 29121 13544 29138 13546
rect 28983 13424 29070 13544
rect 29126 13424 29138 13544
rect 29058 13422 29075 13424
rect 28983 13124 29075 13244
rect 29121 13422 29138 13424
rect 29242 13244 29259 13246
rect 29443 13571 29489 13582
rect 29426 13544 29443 13546
rect 29627 13571 29673 13582
rect 29489 13544 29506 13546
rect 29426 13424 29438 13544
rect 29494 13424 29506 13544
rect 29426 13422 29443 13424
rect 29305 13244 29322 13246
rect 29242 13124 29254 13244
rect 29310 13124 29322 13244
rect 29242 13122 29259 13124
rect 29075 13086 29121 13097
rect 29305 13122 29322 13124
rect 29259 13086 29305 13097
rect 29489 13422 29506 13424
rect 29610 13244 29627 13246
rect 29748 13544 29765 13546
rect 29811 13544 29828 13546
rect 29748 13423 29760 13544
rect 29816 13423 29828 13544
rect 29748 13421 29765 13423
rect 29673 13244 29690 13246
rect 29610 13124 29622 13244
rect 29678 13124 29690 13244
rect 29610 13122 29627 13124
rect 29443 13086 29489 13097
rect 29673 13122 29690 13124
rect 29627 13086 29673 13097
rect 29152 13048 29163 13051
rect 29217 13048 29228 13051
rect 29336 13048 29347 13051
rect 29401 13048 29412 13051
rect 29520 13048 29531 13051
rect 29585 13048 29596 13051
rect 28937 13003 28983 13014
rect 29150 12992 29162 13048
rect 29218 12992 29230 13048
rect 29150 12978 29230 12992
rect 29334 12992 29346 13048
rect 29402 12992 29414 13048
rect 29334 12978 29414 12992
rect 29518 12992 29530 13048
rect 29586 12992 29598 13048
rect 29811 13421 29828 13423
rect 29765 13003 29811 13014
rect 29518 12978 29598 12992
rect 29150 12898 29230 12900
rect 28762 12842 29162 12898
rect 29218 12842 29230 12898
rect 30248 12899 30304 13919
rect 31406 13907 31486 13919
rect 30912 13868 30998 13872
rect 30912 13812 30924 13868
rect 30980 13812 30998 13868
rect 30912 13800 30998 13812
rect 30423 13655 30469 13666
rect 30638 13664 30714 13697
rect 30638 13618 30649 13664
rect 30703 13618 30714 13664
rect 30822 13664 30898 13697
rect 30822 13618 30833 13664
rect 30887 13618 30898 13664
rect 31006 13664 31082 13697
rect 31006 13618 31017 13664
rect 31071 13618 31082 13664
rect 31251 13655 31297 13666
rect 30561 13572 30607 13583
rect 30544 13545 30561 13547
rect 30745 13572 30791 13583
rect 30607 13545 30624 13547
rect 30469 13425 30556 13545
rect 30612 13425 30624 13545
rect 30544 13423 30561 13425
rect 30469 13125 30561 13245
rect 30607 13423 30624 13425
rect 30728 13245 30745 13247
rect 30929 13572 30975 13583
rect 30912 13545 30929 13547
rect 31113 13572 31159 13583
rect 30975 13545 30992 13547
rect 30912 13425 30924 13545
rect 30980 13425 30992 13545
rect 30912 13423 30929 13425
rect 30791 13245 30808 13247
rect 30728 13125 30740 13245
rect 30796 13125 30808 13245
rect 30728 13123 30745 13125
rect 30561 13087 30607 13098
rect 30791 13123 30808 13125
rect 30745 13087 30791 13098
rect 30975 13423 30992 13425
rect 31096 13245 31113 13247
rect 31234 13545 31251 13547
rect 31297 13545 31314 13547
rect 31234 13424 31246 13545
rect 31302 13424 31314 13545
rect 31234 13422 31251 13424
rect 31159 13245 31176 13247
rect 31096 13125 31108 13245
rect 31164 13125 31176 13245
rect 31096 13123 31113 13125
rect 30929 13087 30975 13098
rect 31159 13123 31176 13125
rect 31113 13087 31159 13098
rect 30638 13049 30649 13052
rect 30703 13049 30714 13052
rect 30822 13049 30833 13052
rect 30887 13049 30898 13052
rect 31006 13049 31017 13052
rect 31071 13049 31082 13052
rect 30423 13004 30469 13015
rect 30636 12993 30648 13049
rect 30704 12993 30716 13049
rect 30636 12979 30716 12993
rect 30820 12993 30832 13049
rect 30888 12993 30900 13049
rect 30820 12979 30900 12993
rect 31004 12993 31016 13049
rect 31072 12993 31084 13049
rect 31297 13422 31314 13424
rect 31251 13004 31297 13015
rect 31004 12979 31084 12993
rect 30636 12899 30716 12901
rect 30248 12843 30648 12899
rect 30704 12843 30716 12899
rect 29150 12840 29230 12842
rect 30636 12841 30716 12843
rect 29334 12782 29414 12784
rect 28626 12726 29346 12782
rect 29402 12726 29414 12782
rect 29334 12724 29414 12726
rect 29663 12782 29743 12784
rect 29930 12783 30000 12794
rect 30820 12783 30900 12785
rect 29930 12782 30832 12783
rect 29663 12726 29675 12782
rect 29731 12726 29932 12782
rect 29988 12727 30832 12782
rect 30888 12727 30900 12783
rect 29988 12726 30248 12727
rect 29663 12724 29743 12726
rect 29930 12716 30000 12726
rect 30820 12725 30900 12727
rect 31149 12783 31229 12785
rect 31592 12783 31662 12793
rect 31149 12727 31161 12783
rect 31217 12727 31594 12783
rect 31650 12727 31662 12783
rect 31149 12725 31229 12727
rect 31592 12715 31662 12727
rect 4226 12669 4296 12681
rect 5266 12669 5346 12671
rect 6752 12670 6832 12672
rect 4226 12613 4238 12669
rect 4294 12613 5278 12669
rect 5334 12613 5346 12669
rect 4226 12601 4296 12613
rect 4510 11882 4566 12613
rect 5266 12611 5346 12613
rect 5996 12614 6764 12670
rect 6820 12614 6832 12670
rect 4898 12519 4978 12533
rect 4685 12497 4731 12508
rect 4898 12463 4910 12519
rect 4966 12463 4978 12519
rect 5082 12519 5162 12533
rect 5082 12463 5094 12519
rect 5150 12463 5162 12519
rect 5266 12519 5346 12533
rect 5266 12463 5278 12519
rect 5334 12463 5346 12519
rect 5513 12497 5559 12508
rect 4900 12460 4911 12463
rect 4965 12460 4976 12463
rect 5084 12460 5095 12463
rect 5149 12460 5160 12463
rect 5268 12460 5279 12463
rect 5333 12460 5344 12463
rect 4823 12414 4869 12425
rect 4731 12240 4823 12414
rect 4823 12229 4869 12240
rect 5007 12414 5053 12425
rect 5007 12229 5053 12240
rect 5191 12414 5237 12425
rect 5375 12414 5421 12425
rect 5358 12387 5375 12389
rect 5421 12387 5438 12389
rect 5358 12267 5370 12387
rect 5426 12267 5438 12387
rect 5358 12265 5375 12267
rect 5191 12229 5237 12240
rect 5421 12265 5438 12267
rect 5375 12229 5421 12240
rect 4685 12012 4731 12157
rect 4900 12148 4911 12194
rect 4965 12148 4976 12194
rect 4900 12115 4976 12148
rect 5084 12148 5095 12194
rect 5149 12148 5160 12194
rect 5084 12115 5160 12148
rect 5268 12148 5279 12194
rect 5333 12148 5344 12194
rect 5268 12115 5344 12148
rect 5513 12012 5559 12157
rect 4673 12000 4753 12012
rect 4673 11944 4685 12000
rect 4741 11944 4753 12000
rect 4673 11932 4753 11944
rect 5491 12000 5569 12012
rect 5491 11944 5503 12000
rect 5559 11944 5569 12000
rect 5491 11932 5569 11944
rect 5844 11882 5924 11892
rect 4510 11826 5856 11882
rect 5912 11826 5924 11882
rect 5844 11824 5924 11826
rect 5678 11773 5748 11775
rect 4510 11772 5748 11773
rect 4510 11718 5680 11772
rect 5736 11718 5748 11772
rect 4510 11717 5748 11718
rect 4510 10696 4566 11717
rect 5678 11709 5748 11717
rect 5174 11665 5260 11669
rect 5174 11609 5186 11665
rect 5242 11609 5260 11665
rect 5174 11597 5260 11609
rect 4685 11452 4731 11463
rect 4900 11461 4976 11494
rect 4900 11415 4911 11461
rect 4965 11415 4976 11461
rect 5084 11461 5160 11494
rect 5084 11415 5095 11461
rect 5149 11415 5160 11461
rect 5268 11461 5344 11494
rect 5268 11415 5279 11461
rect 5333 11415 5344 11461
rect 5513 11452 5559 11463
rect 4823 11369 4869 11380
rect 4806 11342 4823 11344
rect 5007 11369 5053 11380
rect 4869 11342 4886 11344
rect 4731 11222 4818 11342
rect 4874 11222 4886 11342
rect 4806 11220 4823 11222
rect 4731 10922 4823 11042
rect 4869 11220 4886 11222
rect 4990 11042 5007 11044
rect 5191 11369 5237 11380
rect 5174 11342 5191 11344
rect 5375 11369 5421 11380
rect 5237 11342 5254 11344
rect 5174 11222 5186 11342
rect 5242 11222 5254 11342
rect 5174 11220 5191 11222
rect 5053 11042 5070 11044
rect 4990 10922 5002 11042
rect 5058 10922 5070 11042
rect 4990 10920 5007 10922
rect 4823 10884 4869 10895
rect 5053 10920 5070 10922
rect 5007 10884 5053 10895
rect 5237 11220 5254 11222
rect 5358 11042 5375 11044
rect 5496 11342 5513 11344
rect 5559 11342 5576 11344
rect 5496 11221 5508 11342
rect 5564 11221 5576 11342
rect 5496 11219 5513 11221
rect 5421 11042 5438 11044
rect 5358 10922 5370 11042
rect 5426 10922 5438 11042
rect 5358 10920 5375 10922
rect 5191 10884 5237 10895
rect 5421 10920 5438 10922
rect 5375 10884 5421 10895
rect 4900 10846 4911 10849
rect 4965 10846 4976 10849
rect 5084 10846 5095 10849
rect 5149 10846 5160 10849
rect 5268 10846 5279 10849
rect 5333 10846 5344 10849
rect 4685 10801 4731 10812
rect 4898 10790 4910 10846
rect 4966 10790 4978 10846
rect 4898 10776 4978 10790
rect 5082 10790 5094 10846
rect 5150 10790 5162 10846
rect 5082 10776 5162 10790
rect 5266 10790 5278 10846
rect 5334 10790 5346 10846
rect 5559 11219 5576 11221
rect 5513 10801 5559 10812
rect 5266 10776 5346 10790
rect 4898 10696 4978 10698
rect 4510 10640 4910 10696
rect 4966 10640 4978 10696
rect 4898 10638 4978 10640
rect 4090 10580 4160 10594
rect 5082 10580 5162 10582
rect 4090 10524 4102 10580
rect 4158 10524 5094 10580
rect 5150 10524 5162 10580
rect 4090 10512 4160 10524
rect 5082 10522 5162 10524
rect 5411 10580 5491 10582
rect 5854 10580 5914 10592
rect 5411 10524 5423 10580
rect 5479 10524 5856 10580
rect 5912 10524 5914 10580
rect 5411 10522 5491 10524
rect 5854 10512 5914 10524
rect 3274 10464 3344 10476
rect 5266 10464 5346 10466
rect 3274 10408 3286 10464
rect 3342 10408 5278 10464
rect 5334 10408 5346 10464
rect 3274 10396 3344 10408
rect 5266 10406 5346 10408
rect 4898 10314 4978 10328
rect 4685 10292 4731 10303
rect 4898 10258 4910 10314
rect 4966 10258 4978 10314
rect 5082 10314 5162 10328
rect 5082 10258 5094 10314
rect 5150 10258 5162 10314
rect 5266 10314 5346 10328
rect 5266 10258 5278 10314
rect 5334 10258 5346 10314
rect 5513 10292 5559 10303
rect 4900 10255 4911 10258
rect 4965 10255 4976 10258
rect 5084 10255 5095 10258
rect 5149 10255 5160 10258
rect 5268 10255 5279 10258
rect 5333 10255 5344 10258
rect 4823 10209 4869 10220
rect 4731 10035 4823 10209
rect 4823 10024 4869 10035
rect 5007 10209 5053 10220
rect 5007 10024 5053 10035
rect 5191 10209 5237 10220
rect 5375 10209 5421 10220
rect 5358 10182 5375 10184
rect 5421 10182 5438 10184
rect 5358 10062 5370 10182
rect 5426 10062 5438 10182
rect 5358 10060 5375 10062
rect 5191 10024 5237 10035
rect 5421 10060 5438 10062
rect 5375 10024 5421 10035
rect 4685 9807 4731 9952
rect 4900 9943 4911 9989
rect 4965 9943 4976 9989
rect 4900 9910 4976 9943
rect 5084 9943 5095 9989
rect 5149 9943 5160 9989
rect 5084 9910 5160 9943
rect 5268 9943 5279 9989
rect 5333 9943 5344 9989
rect 5268 9910 5344 9943
rect 5513 9807 5559 9952
rect 4673 9795 4753 9807
rect 4673 9739 4685 9795
rect 4741 9739 4753 9795
rect 4673 9727 4753 9739
rect 5491 9795 5571 9807
rect 5491 9739 5503 9795
rect 5559 9739 5571 9795
rect 5491 9727 5571 9739
rect 3818 9677 3888 9689
rect 4100 9677 4160 9681
rect 5996 9677 6052 12614
rect 6752 12612 6832 12614
rect 8268 12666 8338 12678
rect 9308 12666 9388 12668
rect 10794 12667 10874 12669
rect 8268 12610 8280 12666
rect 8336 12610 9320 12666
rect 9376 12610 9388 12666
rect 8268 12598 8338 12610
rect 6384 12520 6464 12534
rect 6171 12498 6217 12509
rect 6384 12464 6396 12520
rect 6452 12464 6464 12520
rect 6568 12520 6648 12534
rect 6568 12464 6580 12520
rect 6636 12464 6648 12520
rect 6752 12520 6832 12534
rect 6752 12464 6764 12520
rect 6820 12464 6832 12520
rect 6999 12498 7045 12509
rect 6386 12461 6397 12464
rect 6451 12461 6462 12464
rect 6570 12461 6581 12464
rect 6635 12461 6646 12464
rect 6754 12461 6765 12464
rect 6819 12461 6830 12464
rect 6309 12415 6355 12426
rect 6217 12241 6309 12415
rect 6309 12230 6355 12241
rect 6493 12415 6539 12426
rect 6493 12230 6539 12241
rect 6677 12415 6723 12426
rect 6861 12415 6907 12426
rect 6844 12388 6861 12390
rect 6907 12388 6924 12390
rect 6844 12268 6856 12388
rect 6912 12268 6924 12388
rect 6844 12266 6861 12268
rect 6677 12230 6723 12241
rect 6907 12266 6924 12268
rect 6861 12230 6907 12241
rect 6171 12013 6217 12158
rect 6386 12149 6397 12195
rect 6451 12149 6462 12195
rect 6386 12116 6462 12149
rect 6570 12149 6581 12195
rect 6635 12149 6646 12195
rect 6570 12116 6646 12149
rect 6754 12149 6765 12195
rect 6819 12149 6830 12195
rect 6754 12116 6830 12149
rect 6999 12013 7045 12158
rect 6159 12001 6239 12013
rect 6159 11945 6171 12001
rect 6227 11945 6239 12001
rect 6159 11933 6239 11945
rect 6977 12001 7055 12013
rect 6977 11945 6989 12001
rect 7045 11945 7055 12001
rect 6977 11933 7055 11945
rect 8552 11879 8608 12610
rect 9308 12608 9388 12610
rect 10038 12611 10806 12667
rect 10862 12611 10874 12667
rect 8940 12516 9020 12530
rect 8727 12494 8773 12505
rect 8940 12460 8952 12516
rect 9008 12460 9020 12516
rect 9124 12516 9204 12530
rect 9124 12460 9136 12516
rect 9192 12460 9204 12516
rect 9308 12516 9388 12530
rect 9308 12460 9320 12516
rect 9376 12460 9388 12516
rect 9555 12494 9601 12505
rect 8942 12457 8953 12460
rect 9007 12457 9018 12460
rect 9126 12457 9137 12460
rect 9191 12457 9202 12460
rect 9310 12457 9321 12460
rect 9375 12457 9386 12460
rect 8865 12411 8911 12422
rect 8773 12237 8865 12411
rect 8865 12226 8911 12237
rect 9049 12411 9095 12422
rect 9049 12226 9095 12237
rect 9233 12411 9279 12422
rect 9417 12411 9463 12422
rect 9400 12384 9417 12386
rect 9463 12384 9480 12386
rect 9400 12264 9412 12384
rect 9468 12264 9480 12384
rect 9400 12262 9417 12264
rect 9233 12226 9279 12237
rect 9463 12262 9480 12264
rect 9417 12226 9463 12237
rect 8727 12009 8773 12154
rect 8942 12145 8953 12191
rect 9007 12145 9018 12191
rect 8942 12112 9018 12145
rect 9126 12145 9137 12191
rect 9191 12145 9202 12191
rect 9126 12112 9202 12145
rect 9310 12145 9321 12191
rect 9375 12145 9386 12191
rect 9310 12112 9386 12145
rect 9555 12009 9601 12154
rect 8715 11997 8795 12009
rect 8715 11941 8727 11997
rect 8783 11941 8795 11997
rect 8715 11929 8795 11941
rect 9533 11997 9611 12009
rect 9533 11941 9545 11997
rect 9601 11941 9611 11997
rect 9533 11929 9611 11941
rect 9886 11879 9966 11889
rect 8552 11823 9898 11879
rect 9954 11823 9966 11879
rect 9886 11821 9966 11823
rect 9720 11770 9790 11772
rect 8552 11769 9790 11770
rect 8552 11715 9722 11769
rect 9778 11715 9790 11769
rect 8552 11714 9790 11715
rect 8552 10693 8608 11714
rect 9720 11706 9790 11714
rect 9216 11662 9302 11666
rect 9216 11606 9228 11662
rect 9284 11606 9302 11662
rect 9216 11594 9302 11606
rect 8727 11449 8773 11460
rect 8942 11458 9018 11491
rect 8942 11412 8953 11458
rect 9007 11412 9018 11458
rect 9126 11458 9202 11491
rect 9126 11412 9137 11458
rect 9191 11412 9202 11458
rect 9310 11458 9386 11491
rect 9310 11412 9321 11458
rect 9375 11412 9386 11458
rect 9555 11449 9601 11460
rect 8865 11366 8911 11377
rect 8848 11339 8865 11341
rect 9049 11366 9095 11377
rect 8911 11339 8928 11341
rect 8773 11219 8860 11339
rect 8916 11219 8928 11339
rect 8848 11217 8865 11219
rect 8773 10919 8865 11039
rect 8911 11217 8928 11219
rect 9032 11039 9049 11041
rect 9233 11366 9279 11377
rect 9216 11339 9233 11341
rect 9417 11366 9463 11377
rect 9279 11339 9296 11341
rect 9216 11219 9228 11339
rect 9284 11219 9296 11339
rect 9216 11217 9233 11219
rect 9095 11039 9112 11041
rect 9032 10919 9044 11039
rect 9100 10919 9112 11039
rect 9032 10917 9049 10919
rect 8865 10881 8911 10892
rect 9095 10917 9112 10919
rect 9049 10881 9095 10892
rect 9279 11217 9296 11219
rect 9400 11039 9417 11041
rect 9538 11339 9555 11341
rect 9601 11339 9618 11341
rect 9538 11218 9550 11339
rect 9606 11218 9618 11339
rect 9538 11216 9555 11218
rect 9463 11039 9480 11041
rect 9400 10919 9412 11039
rect 9468 10919 9480 11039
rect 9400 10917 9417 10919
rect 9233 10881 9279 10892
rect 9463 10917 9480 10919
rect 9417 10881 9463 10892
rect 8942 10843 8953 10846
rect 9007 10843 9018 10846
rect 9126 10843 9137 10846
rect 9191 10843 9202 10846
rect 9310 10843 9321 10846
rect 9375 10843 9386 10846
rect 8727 10798 8773 10809
rect 8940 10787 8952 10843
rect 9008 10787 9020 10843
rect 8940 10773 9020 10787
rect 9124 10787 9136 10843
rect 9192 10787 9204 10843
rect 9124 10773 9204 10787
rect 9308 10787 9320 10843
rect 9376 10787 9388 10843
rect 9601 11216 9618 11218
rect 9555 10798 9601 10809
rect 9308 10773 9388 10787
rect 8940 10693 9020 10695
rect 8552 10637 8952 10693
rect 9008 10637 9020 10693
rect 8940 10635 9020 10637
rect 8132 10577 8202 10591
rect 9124 10577 9204 10579
rect 8132 10521 8144 10577
rect 8200 10521 9136 10577
rect 9192 10521 9204 10577
rect 8132 10509 8202 10521
rect 9124 10519 9204 10521
rect 9453 10577 9533 10579
rect 9896 10577 9956 10589
rect 9453 10521 9465 10577
rect 9521 10521 9898 10577
rect 9954 10521 9956 10577
rect 9453 10519 9533 10521
rect 9896 10509 9956 10521
rect 7286 10461 7356 10473
rect 9308 10461 9388 10463
rect 7286 10405 7298 10461
rect 7354 10405 9320 10461
rect 9376 10405 9388 10461
rect 7286 10393 7356 10405
rect 9308 10403 9388 10405
rect 8940 10311 9020 10325
rect 8727 10289 8773 10300
rect 8940 10255 8952 10311
rect 9008 10255 9020 10311
rect 9124 10311 9204 10325
rect 9124 10255 9136 10311
rect 9192 10255 9204 10311
rect 9308 10311 9388 10325
rect 9308 10255 9320 10311
rect 9376 10255 9388 10311
rect 9555 10289 9601 10300
rect 8942 10252 8953 10255
rect 9007 10252 9018 10255
rect 9126 10252 9137 10255
rect 9191 10252 9202 10255
rect 9310 10252 9321 10255
rect 9375 10252 9386 10255
rect 8865 10206 8911 10217
rect 8773 10032 8865 10206
rect 8865 10021 8911 10032
rect 9049 10206 9095 10217
rect 9049 10021 9095 10032
rect 9233 10206 9279 10217
rect 9417 10206 9463 10217
rect 9400 10179 9417 10181
rect 9463 10179 9480 10181
rect 9400 10059 9412 10179
rect 9468 10059 9480 10179
rect 9400 10057 9417 10059
rect 9233 10021 9279 10032
rect 9463 10057 9480 10059
rect 9417 10021 9463 10032
rect 8727 9804 8773 9949
rect 8942 9940 8953 9986
rect 9007 9940 9018 9986
rect 8942 9907 9018 9940
rect 9126 9940 9137 9986
rect 9191 9940 9202 9986
rect 9126 9907 9202 9940
rect 9310 9940 9321 9986
rect 9375 9940 9386 9986
rect 9310 9907 9386 9940
rect 9555 9804 9601 9949
rect 8715 9792 8795 9804
rect 8715 9736 8727 9792
rect 8783 9736 8795 9792
rect 8715 9724 8795 9736
rect 9533 9792 9613 9804
rect 9533 9736 9545 9792
rect 9601 9736 9613 9792
rect 9533 9724 9613 9736
rect 3818 9621 3830 9677
rect 3886 9621 4102 9677
rect 4158 9621 6052 9677
rect 7830 9674 7900 9686
rect 8142 9674 8202 9678
rect 10038 9674 10094 12611
rect 10794 12609 10874 12611
rect 12310 12666 12380 12678
rect 13350 12666 13430 12668
rect 14836 12667 14916 12669
rect 12310 12610 12322 12666
rect 12378 12610 13362 12666
rect 13418 12610 13430 12666
rect 12310 12598 12380 12610
rect 10426 12517 10506 12531
rect 10213 12495 10259 12506
rect 10426 12461 10438 12517
rect 10494 12461 10506 12517
rect 10610 12517 10690 12531
rect 10610 12461 10622 12517
rect 10678 12461 10690 12517
rect 10794 12517 10874 12531
rect 10794 12461 10806 12517
rect 10862 12461 10874 12517
rect 11041 12495 11087 12506
rect 10428 12458 10439 12461
rect 10493 12458 10504 12461
rect 10612 12458 10623 12461
rect 10677 12458 10688 12461
rect 10796 12458 10807 12461
rect 10861 12458 10872 12461
rect 10351 12412 10397 12423
rect 10259 12238 10351 12412
rect 10351 12227 10397 12238
rect 10535 12412 10581 12423
rect 10535 12227 10581 12238
rect 10719 12412 10765 12423
rect 10903 12412 10949 12423
rect 10886 12385 10903 12387
rect 10949 12385 10966 12387
rect 10886 12265 10898 12385
rect 10954 12265 10966 12385
rect 10886 12263 10903 12265
rect 10719 12227 10765 12238
rect 10949 12263 10966 12265
rect 10903 12227 10949 12238
rect 10213 12010 10259 12155
rect 10428 12146 10439 12192
rect 10493 12146 10504 12192
rect 10428 12113 10504 12146
rect 10612 12146 10623 12192
rect 10677 12146 10688 12192
rect 10612 12113 10688 12146
rect 10796 12146 10807 12192
rect 10861 12146 10872 12192
rect 10796 12113 10872 12146
rect 11041 12010 11087 12155
rect 10201 11998 10281 12010
rect 10201 11942 10213 11998
rect 10269 11942 10281 11998
rect 10201 11930 10281 11942
rect 11019 11998 11097 12010
rect 11019 11942 11031 11998
rect 11087 11942 11097 11998
rect 11019 11930 11097 11942
rect 12594 11879 12650 12610
rect 13350 12608 13430 12610
rect 14080 12611 14848 12667
rect 14904 12611 14916 12667
rect 12982 12516 13062 12530
rect 12769 12494 12815 12505
rect 12982 12460 12994 12516
rect 13050 12460 13062 12516
rect 13166 12516 13246 12530
rect 13166 12460 13178 12516
rect 13234 12460 13246 12516
rect 13350 12516 13430 12530
rect 13350 12460 13362 12516
rect 13418 12460 13430 12516
rect 13597 12494 13643 12505
rect 12984 12457 12995 12460
rect 13049 12457 13060 12460
rect 13168 12457 13179 12460
rect 13233 12457 13244 12460
rect 13352 12457 13363 12460
rect 13417 12457 13428 12460
rect 12907 12411 12953 12422
rect 12815 12237 12907 12411
rect 12907 12226 12953 12237
rect 13091 12411 13137 12422
rect 13091 12226 13137 12237
rect 13275 12411 13321 12422
rect 13459 12411 13505 12422
rect 13442 12384 13459 12386
rect 13505 12384 13522 12386
rect 13442 12264 13454 12384
rect 13510 12264 13522 12384
rect 13442 12262 13459 12264
rect 13275 12226 13321 12237
rect 13505 12262 13522 12264
rect 13459 12226 13505 12237
rect 12769 12009 12815 12154
rect 12984 12145 12995 12191
rect 13049 12145 13060 12191
rect 12984 12112 13060 12145
rect 13168 12145 13179 12191
rect 13233 12145 13244 12191
rect 13168 12112 13244 12145
rect 13352 12145 13363 12191
rect 13417 12145 13428 12191
rect 13352 12112 13428 12145
rect 13597 12009 13643 12154
rect 12757 11997 12837 12009
rect 12757 11941 12769 11997
rect 12825 11941 12837 11997
rect 12757 11929 12837 11941
rect 13575 11997 13653 12009
rect 13575 11941 13587 11997
rect 13643 11941 13653 11997
rect 13575 11929 13653 11941
rect 13928 11879 14008 11889
rect 12594 11823 13940 11879
rect 13996 11823 14008 11879
rect 13928 11821 14008 11823
rect 13762 11770 13832 11772
rect 12594 11769 13832 11770
rect 12594 11715 13764 11769
rect 13820 11715 13832 11769
rect 12594 11714 13832 11715
rect 12594 10693 12650 11714
rect 13762 11706 13832 11714
rect 13258 11662 13344 11666
rect 13258 11606 13270 11662
rect 13326 11606 13344 11662
rect 13258 11594 13344 11606
rect 12769 11449 12815 11460
rect 12984 11458 13060 11491
rect 12984 11412 12995 11458
rect 13049 11412 13060 11458
rect 13168 11458 13244 11491
rect 13168 11412 13179 11458
rect 13233 11412 13244 11458
rect 13352 11458 13428 11491
rect 13352 11412 13363 11458
rect 13417 11412 13428 11458
rect 13597 11449 13643 11460
rect 12907 11366 12953 11377
rect 12890 11339 12907 11341
rect 13091 11366 13137 11377
rect 12953 11339 12970 11341
rect 12815 11219 12902 11339
rect 12958 11219 12970 11339
rect 12890 11217 12907 11219
rect 12815 10919 12907 11039
rect 12953 11217 12970 11219
rect 13074 11039 13091 11041
rect 13275 11366 13321 11377
rect 13258 11339 13275 11341
rect 13459 11366 13505 11377
rect 13321 11339 13338 11341
rect 13258 11219 13270 11339
rect 13326 11219 13338 11339
rect 13258 11217 13275 11219
rect 13137 11039 13154 11041
rect 13074 10919 13086 11039
rect 13142 10919 13154 11039
rect 13074 10917 13091 10919
rect 12907 10881 12953 10892
rect 13137 10917 13154 10919
rect 13091 10881 13137 10892
rect 13321 11217 13338 11219
rect 13442 11039 13459 11041
rect 13580 11339 13597 11341
rect 13643 11339 13660 11341
rect 13580 11218 13592 11339
rect 13648 11218 13660 11339
rect 13580 11216 13597 11218
rect 13505 11039 13522 11041
rect 13442 10919 13454 11039
rect 13510 10919 13522 11039
rect 13442 10917 13459 10919
rect 13275 10881 13321 10892
rect 13505 10917 13522 10919
rect 13459 10881 13505 10892
rect 12984 10843 12995 10846
rect 13049 10843 13060 10846
rect 13168 10843 13179 10846
rect 13233 10843 13244 10846
rect 13352 10843 13363 10846
rect 13417 10843 13428 10846
rect 12769 10798 12815 10809
rect 12982 10787 12994 10843
rect 13050 10787 13062 10843
rect 12982 10773 13062 10787
rect 13166 10787 13178 10843
rect 13234 10787 13246 10843
rect 13166 10773 13246 10787
rect 13350 10787 13362 10843
rect 13418 10787 13430 10843
rect 13643 11216 13660 11218
rect 13597 10798 13643 10809
rect 13350 10773 13430 10787
rect 12982 10693 13062 10695
rect 12594 10637 12994 10693
rect 13050 10637 13062 10693
rect 12982 10635 13062 10637
rect 12174 10577 12244 10591
rect 13166 10577 13246 10579
rect 12174 10521 12186 10577
rect 12242 10521 13178 10577
rect 13234 10521 13246 10577
rect 12174 10509 12244 10521
rect 13166 10519 13246 10521
rect 13495 10577 13575 10579
rect 13938 10577 13998 10589
rect 13495 10521 13507 10577
rect 13563 10521 13940 10577
rect 13996 10521 13998 10577
rect 13495 10519 13575 10521
rect 13938 10509 13998 10521
rect 11328 10461 11398 10473
rect 13350 10461 13430 10463
rect 11328 10405 11340 10461
rect 11396 10405 13362 10461
rect 13418 10405 13430 10461
rect 11328 10393 11398 10405
rect 13350 10403 13430 10405
rect 12982 10311 13062 10325
rect 12769 10289 12815 10300
rect 12982 10255 12994 10311
rect 13050 10255 13062 10311
rect 13166 10311 13246 10325
rect 13166 10255 13178 10311
rect 13234 10255 13246 10311
rect 13350 10311 13430 10325
rect 13350 10255 13362 10311
rect 13418 10255 13430 10311
rect 13597 10289 13643 10300
rect 12984 10252 12995 10255
rect 13049 10252 13060 10255
rect 13168 10252 13179 10255
rect 13233 10252 13244 10255
rect 13352 10252 13363 10255
rect 13417 10252 13428 10255
rect 12907 10206 12953 10217
rect 12815 10032 12907 10206
rect 12907 10021 12953 10032
rect 13091 10206 13137 10217
rect 13091 10021 13137 10032
rect 13275 10206 13321 10217
rect 13459 10206 13505 10217
rect 13442 10179 13459 10181
rect 13505 10179 13522 10181
rect 13442 10059 13454 10179
rect 13510 10059 13522 10179
rect 13442 10057 13459 10059
rect 13275 10021 13321 10032
rect 13505 10057 13522 10059
rect 13459 10021 13505 10032
rect 12769 9804 12815 9949
rect 12984 9940 12995 9986
rect 13049 9940 13060 9986
rect 12984 9907 13060 9940
rect 13168 9940 13179 9986
rect 13233 9940 13244 9986
rect 13168 9907 13244 9940
rect 13352 9940 13363 9986
rect 13417 9940 13428 9986
rect 13352 9907 13428 9940
rect 13597 9804 13643 9949
rect 12757 9792 12837 9804
rect 12757 9736 12769 9792
rect 12825 9736 12837 9792
rect 12757 9724 12837 9736
rect 13575 9792 13655 9804
rect 13575 9736 13587 9792
rect 13643 9736 13655 9792
rect 13575 9724 13655 9736
rect 3818 9619 3888 9621
rect 4100 9609 4160 9621
rect 7830 9618 7842 9674
rect 7898 9618 8144 9674
rect 8200 9618 10094 9674
rect 11872 9674 11942 9686
rect 12184 9674 12244 9678
rect 14080 9674 14136 12611
rect 14836 12609 14916 12611
rect 16352 12666 16422 12678
rect 17392 12666 17472 12668
rect 18878 12667 18958 12669
rect 16352 12610 16364 12666
rect 16420 12610 17404 12666
rect 17460 12610 17472 12666
rect 16352 12598 16422 12610
rect 14468 12517 14548 12531
rect 14255 12495 14301 12506
rect 14468 12461 14480 12517
rect 14536 12461 14548 12517
rect 14652 12517 14732 12531
rect 14652 12461 14664 12517
rect 14720 12461 14732 12517
rect 14836 12517 14916 12531
rect 14836 12461 14848 12517
rect 14904 12461 14916 12517
rect 15083 12495 15129 12506
rect 14470 12458 14481 12461
rect 14535 12458 14546 12461
rect 14654 12458 14665 12461
rect 14719 12458 14730 12461
rect 14838 12458 14849 12461
rect 14903 12458 14914 12461
rect 14393 12412 14439 12423
rect 14301 12238 14393 12412
rect 14393 12227 14439 12238
rect 14577 12412 14623 12423
rect 14577 12227 14623 12238
rect 14761 12412 14807 12423
rect 14945 12412 14991 12423
rect 14928 12385 14945 12387
rect 14991 12385 15008 12387
rect 14928 12265 14940 12385
rect 14996 12265 15008 12385
rect 14928 12263 14945 12265
rect 14761 12227 14807 12238
rect 14991 12263 15008 12265
rect 14945 12227 14991 12238
rect 14255 12010 14301 12155
rect 14470 12146 14481 12192
rect 14535 12146 14546 12192
rect 14470 12113 14546 12146
rect 14654 12146 14665 12192
rect 14719 12146 14730 12192
rect 14654 12113 14730 12146
rect 14838 12146 14849 12192
rect 14903 12146 14914 12192
rect 14838 12113 14914 12146
rect 15083 12010 15129 12155
rect 14243 11998 14323 12010
rect 14243 11942 14255 11998
rect 14311 11942 14323 11998
rect 14243 11930 14323 11942
rect 15061 11998 15139 12010
rect 15061 11942 15073 11998
rect 15129 11942 15139 11998
rect 15061 11930 15139 11942
rect 16636 11879 16692 12610
rect 17392 12608 17472 12610
rect 18122 12611 18890 12667
rect 18946 12611 18958 12667
rect 17024 12516 17104 12530
rect 16811 12494 16857 12505
rect 17024 12460 17036 12516
rect 17092 12460 17104 12516
rect 17208 12516 17288 12530
rect 17208 12460 17220 12516
rect 17276 12460 17288 12516
rect 17392 12516 17472 12530
rect 17392 12460 17404 12516
rect 17460 12460 17472 12516
rect 17639 12494 17685 12505
rect 17026 12457 17037 12460
rect 17091 12457 17102 12460
rect 17210 12457 17221 12460
rect 17275 12457 17286 12460
rect 17394 12457 17405 12460
rect 17459 12457 17470 12460
rect 16949 12411 16995 12422
rect 16857 12237 16949 12411
rect 16949 12226 16995 12237
rect 17133 12411 17179 12422
rect 17133 12226 17179 12237
rect 17317 12411 17363 12422
rect 17501 12411 17547 12422
rect 17484 12384 17501 12386
rect 17547 12384 17564 12386
rect 17484 12264 17496 12384
rect 17552 12264 17564 12384
rect 17484 12262 17501 12264
rect 17317 12226 17363 12237
rect 17547 12262 17564 12264
rect 17501 12226 17547 12237
rect 16811 12009 16857 12154
rect 17026 12145 17037 12191
rect 17091 12145 17102 12191
rect 17026 12112 17102 12145
rect 17210 12145 17221 12191
rect 17275 12145 17286 12191
rect 17210 12112 17286 12145
rect 17394 12145 17405 12191
rect 17459 12145 17470 12191
rect 17394 12112 17470 12145
rect 17639 12009 17685 12154
rect 16799 11997 16879 12009
rect 16799 11941 16811 11997
rect 16867 11941 16879 11997
rect 16799 11929 16879 11941
rect 17617 11997 17695 12009
rect 17617 11941 17629 11997
rect 17685 11941 17695 11997
rect 17617 11929 17695 11941
rect 17970 11879 18050 11889
rect 16636 11823 17982 11879
rect 18038 11823 18050 11879
rect 17970 11821 18050 11823
rect 17804 11770 17874 11772
rect 16636 11769 17874 11770
rect 16636 11715 17806 11769
rect 17862 11715 17874 11769
rect 16636 11714 17874 11715
rect 16636 10693 16692 11714
rect 17804 11706 17874 11714
rect 17300 11662 17386 11666
rect 17300 11606 17312 11662
rect 17368 11606 17386 11662
rect 17300 11594 17386 11606
rect 16811 11449 16857 11460
rect 17026 11458 17102 11491
rect 17026 11412 17037 11458
rect 17091 11412 17102 11458
rect 17210 11458 17286 11491
rect 17210 11412 17221 11458
rect 17275 11412 17286 11458
rect 17394 11458 17470 11491
rect 17394 11412 17405 11458
rect 17459 11412 17470 11458
rect 17639 11449 17685 11460
rect 16949 11366 16995 11377
rect 16932 11339 16949 11341
rect 17133 11366 17179 11377
rect 16995 11339 17012 11341
rect 16857 11219 16944 11339
rect 17000 11219 17012 11339
rect 16932 11217 16949 11219
rect 16857 10919 16949 11039
rect 16995 11217 17012 11219
rect 17116 11039 17133 11041
rect 17317 11366 17363 11377
rect 17300 11339 17317 11341
rect 17501 11366 17547 11377
rect 17363 11339 17380 11341
rect 17300 11219 17312 11339
rect 17368 11219 17380 11339
rect 17300 11217 17317 11219
rect 17179 11039 17196 11041
rect 17116 10919 17128 11039
rect 17184 10919 17196 11039
rect 17116 10917 17133 10919
rect 16949 10881 16995 10892
rect 17179 10917 17196 10919
rect 17133 10881 17179 10892
rect 17363 11217 17380 11219
rect 17484 11039 17501 11041
rect 17622 11339 17639 11341
rect 17685 11339 17702 11341
rect 17622 11218 17634 11339
rect 17690 11218 17702 11339
rect 17622 11216 17639 11218
rect 17547 11039 17564 11041
rect 17484 10919 17496 11039
rect 17552 10919 17564 11039
rect 17484 10917 17501 10919
rect 17317 10881 17363 10892
rect 17547 10917 17564 10919
rect 17501 10881 17547 10892
rect 17026 10843 17037 10846
rect 17091 10843 17102 10846
rect 17210 10843 17221 10846
rect 17275 10843 17286 10846
rect 17394 10843 17405 10846
rect 17459 10843 17470 10846
rect 16811 10798 16857 10809
rect 17024 10787 17036 10843
rect 17092 10787 17104 10843
rect 17024 10773 17104 10787
rect 17208 10787 17220 10843
rect 17276 10787 17288 10843
rect 17208 10773 17288 10787
rect 17392 10787 17404 10843
rect 17460 10787 17472 10843
rect 17685 11216 17702 11218
rect 17639 10798 17685 10809
rect 17392 10773 17472 10787
rect 17024 10693 17104 10695
rect 16636 10637 17036 10693
rect 17092 10637 17104 10693
rect 17024 10635 17104 10637
rect 16216 10577 16286 10591
rect 17208 10577 17288 10579
rect 16216 10521 16228 10577
rect 16284 10521 17220 10577
rect 17276 10521 17288 10577
rect 16216 10509 16286 10521
rect 17208 10519 17288 10521
rect 17537 10577 17617 10579
rect 17980 10577 18040 10589
rect 17537 10521 17549 10577
rect 17605 10521 17982 10577
rect 18038 10521 18040 10577
rect 17537 10519 17617 10521
rect 17980 10509 18040 10521
rect 15370 10461 15440 10473
rect 17392 10461 17472 10463
rect 15370 10405 15382 10461
rect 15438 10405 17404 10461
rect 17460 10405 17472 10461
rect 15370 10393 15440 10405
rect 17392 10403 17472 10405
rect 17024 10311 17104 10325
rect 16811 10289 16857 10300
rect 17024 10255 17036 10311
rect 17092 10255 17104 10311
rect 17208 10311 17288 10325
rect 17208 10255 17220 10311
rect 17276 10255 17288 10311
rect 17392 10311 17472 10325
rect 17392 10255 17404 10311
rect 17460 10255 17472 10311
rect 17639 10289 17685 10300
rect 17026 10252 17037 10255
rect 17091 10252 17102 10255
rect 17210 10252 17221 10255
rect 17275 10252 17286 10255
rect 17394 10252 17405 10255
rect 17459 10252 17470 10255
rect 16949 10206 16995 10217
rect 16857 10032 16949 10206
rect 16949 10021 16995 10032
rect 17133 10206 17179 10217
rect 17133 10021 17179 10032
rect 17317 10206 17363 10217
rect 17501 10206 17547 10217
rect 17484 10179 17501 10181
rect 17547 10179 17564 10181
rect 17484 10059 17496 10179
rect 17552 10059 17564 10179
rect 17484 10057 17501 10059
rect 17317 10021 17363 10032
rect 17547 10057 17564 10059
rect 17501 10021 17547 10032
rect 16811 9804 16857 9949
rect 17026 9940 17037 9986
rect 17091 9940 17102 9986
rect 17026 9907 17102 9940
rect 17210 9940 17221 9986
rect 17275 9940 17286 9986
rect 17210 9907 17286 9940
rect 17394 9940 17405 9986
rect 17459 9940 17470 9986
rect 17394 9907 17470 9940
rect 17639 9804 17685 9949
rect 16799 9792 16879 9804
rect 16799 9736 16811 9792
rect 16867 9736 16879 9792
rect 16799 9724 16879 9736
rect 17617 9792 17697 9804
rect 17617 9736 17629 9792
rect 17685 9736 17697 9792
rect 17617 9724 17697 9736
rect 11872 9618 11884 9674
rect 11940 9618 12186 9674
rect 12242 9618 14136 9674
rect 15914 9674 15984 9686
rect 16226 9674 16286 9678
rect 18122 9674 18178 12611
rect 18878 12609 18958 12611
rect 20394 12666 20464 12678
rect 21434 12666 21514 12668
rect 22920 12667 23000 12669
rect 20394 12610 20406 12666
rect 20462 12610 21446 12666
rect 21502 12610 21514 12666
rect 20394 12598 20464 12610
rect 18510 12517 18590 12531
rect 18297 12495 18343 12506
rect 18510 12461 18522 12517
rect 18578 12461 18590 12517
rect 18694 12517 18774 12531
rect 18694 12461 18706 12517
rect 18762 12461 18774 12517
rect 18878 12517 18958 12531
rect 18878 12461 18890 12517
rect 18946 12461 18958 12517
rect 19125 12495 19171 12506
rect 18512 12458 18523 12461
rect 18577 12458 18588 12461
rect 18696 12458 18707 12461
rect 18761 12458 18772 12461
rect 18880 12458 18891 12461
rect 18945 12458 18956 12461
rect 18435 12412 18481 12423
rect 18343 12238 18435 12412
rect 18435 12227 18481 12238
rect 18619 12412 18665 12423
rect 18619 12227 18665 12238
rect 18803 12412 18849 12423
rect 18987 12412 19033 12423
rect 18970 12385 18987 12387
rect 19033 12385 19050 12387
rect 18970 12265 18982 12385
rect 19038 12265 19050 12385
rect 18970 12263 18987 12265
rect 18803 12227 18849 12238
rect 19033 12263 19050 12265
rect 18987 12227 19033 12238
rect 18297 12010 18343 12155
rect 18512 12146 18523 12192
rect 18577 12146 18588 12192
rect 18512 12113 18588 12146
rect 18696 12146 18707 12192
rect 18761 12146 18772 12192
rect 18696 12113 18772 12146
rect 18880 12146 18891 12192
rect 18945 12146 18956 12192
rect 18880 12113 18956 12146
rect 19125 12010 19171 12155
rect 18285 11998 18365 12010
rect 18285 11942 18297 11998
rect 18353 11942 18365 11998
rect 18285 11930 18365 11942
rect 19103 11998 19181 12010
rect 19103 11942 19115 11998
rect 19171 11942 19181 11998
rect 19103 11930 19181 11942
rect 20678 11879 20734 12610
rect 21434 12608 21514 12610
rect 22164 12611 22932 12667
rect 22988 12611 23000 12667
rect 21066 12516 21146 12530
rect 20853 12494 20899 12505
rect 21066 12460 21078 12516
rect 21134 12460 21146 12516
rect 21250 12516 21330 12530
rect 21250 12460 21262 12516
rect 21318 12460 21330 12516
rect 21434 12516 21514 12530
rect 21434 12460 21446 12516
rect 21502 12460 21514 12516
rect 21681 12494 21727 12505
rect 21068 12457 21079 12460
rect 21133 12457 21144 12460
rect 21252 12457 21263 12460
rect 21317 12457 21328 12460
rect 21436 12457 21447 12460
rect 21501 12457 21512 12460
rect 20991 12411 21037 12422
rect 20899 12237 20991 12411
rect 20991 12226 21037 12237
rect 21175 12411 21221 12422
rect 21175 12226 21221 12237
rect 21359 12411 21405 12422
rect 21543 12411 21589 12422
rect 21526 12384 21543 12386
rect 21589 12384 21606 12386
rect 21526 12264 21538 12384
rect 21594 12264 21606 12384
rect 21526 12262 21543 12264
rect 21359 12226 21405 12237
rect 21589 12262 21606 12264
rect 21543 12226 21589 12237
rect 20853 12009 20899 12154
rect 21068 12145 21079 12191
rect 21133 12145 21144 12191
rect 21068 12112 21144 12145
rect 21252 12145 21263 12191
rect 21317 12145 21328 12191
rect 21252 12112 21328 12145
rect 21436 12145 21447 12191
rect 21501 12145 21512 12191
rect 21436 12112 21512 12145
rect 21681 12009 21727 12154
rect 20841 11997 20921 12009
rect 20841 11941 20853 11997
rect 20909 11941 20921 11997
rect 20841 11929 20921 11941
rect 21659 11997 21737 12009
rect 21659 11941 21671 11997
rect 21727 11941 21737 11997
rect 21659 11929 21737 11941
rect 22012 11879 22092 11889
rect 20678 11823 22024 11879
rect 22080 11823 22092 11879
rect 22012 11821 22092 11823
rect 21846 11770 21916 11772
rect 20678 11769 21916 11770
rect 20678 11715 21848 11769
rect 21904 11715 21916 11769
rect 20678 11714 21916 11715
rect 20678 10693 20734 11714
rect 21846 11706 21916 11714
rect 21342 11662 21428 11666
rect 21342 11606 21354 11662
rect 21410 11606 21428 11662
rect 21342 11594 21428 11606
rect 20853 11449 20899 11460
rect 21068 11458 21144 11491
rect 21068 11412 21079 11458
rect 21133 11412 21144 11458
rect 21252 11458 21328 11491
rect 21252 11412 21263 11458
rect 21317 11412 21328 11458
rect 21436 11458 21512 11491
rect 21436 11412 21447 11458
rect 21501 11412 21512 11458
rect 21681 11449 21727 11460
rect 20991 11366 21037 11377
rect 20974 11339 20991 11341
rect 21175 11366 21221 11377
rect 21037 11339 21054 11341
rect 20899 11219 20986 11339
rect 21042 11219 21054 11339
rect 20974 11217 20991 11219
rect 20899 10919 20991 11039
rect 21037 11217 21054 11219
rect 21158 11039 21175 11041
rect 21359 11366 21405 11377
rect 21342 11339 21359 11341
rect 21543 11366 21589 11377
rect 21405 11339 21422 11341
rect 21342 11219 21354 11339
rect 21410 11219 21422 11339
rect 21342 11217 21359 11219
rect 21221 11039 21238 11041
rect 21158 10919 21170 11039
rect 21226 10919 21238 11039
rect 21158 10917 21175 10919
rect 20991 10881 21037 10892
rect 21221 10917 21238 10919
rect 21175 10881 21221 10892
rect 21405 11217 21422 11219
rect 21526 11039 21543 11041
rect 21664 11339 21681 11341
rect 21727 11339 21744 11341
rect 21664 11218 21676 11339
rect 21732 11218 21744 11339
rect 21664 11216 21681 11218
rect 21589 11039 21606 11041
rect 21526 10919 21538 11039
rect 21594 10919 21606 11039
rect 21526 10917 21543 10919
rect 21359 10881 21405 10892
rect 21589 10917 21606 10919
rect 21543 10881 21589 10892
rect 21068 10843 21079 10846
rect 21133 10843 21144 10846
rect 21252 10843 21263 10846
rect 21317 10843 21328 10846
rect 21436 10843 21447 10846
rect 21501 10843 21512 10846
rect 20853 10798 20899 10809
rect 21066 10787 21078 10843
rect 21134 10787 21146 10843
rect 21066 10773 21146 10787
rect 21250 10787 21262 10843
rect 21318 10787 21330 10843
rect 21250 10773 21330 10787
rect 21434 10787 21446 10843
rect 21502 10787 21514 10843
rect 21727 11216 21744 11218
rect 21681 10798 21727 10809
rect 21434 10773 21514 10787
rect 21066 10693 21146 10695
rect 20678 10637 21078 10693
rect 21134 10637 21146 10693
rect 21066 10635 21146 10637
rect 20258 10577 20328 10591
rect 21250 10577 21330 10579
rect 20258 10521 20270 10577
rect 20326 10521 21262 10577
rect 21318 10521 21330 10577
rect 20258 10509 20328 10521
rect 21250 10519 21330 10521
rect 21579 10577 21659 10579
rect 22022 10577 22082 10589
rect 21579 10521 21591 10577
rect 21647 10521 22024 10577
rect 22080 10521 22082 10577
rect 21579 10519 21659 10521
rect 22022 10509 22082 10521
rect 19412 10461 19482 10473
rect 21434 10461 21514 10463
rect 19412 10405 19424 10461
rect 19480 10405 21446 10461
rect 21502 10405 21514 10461
rect 19412 10393 19482 10405
rect 21434 10403 21514 10405
rect 21066 10311 21146 10325
rect 20853 10289 20899 10300
rect 21066 10255 21078 10311
rect 21134 10255 21146 10311
rect 21250 10311 21330 10325
rect 21250 10255 21262 10311
rect 21318 10255 21330 10311
rect 21434 10311 21514 10325
rect 21434 10255 21446 10311
rect 21502 10255 21514 10311
rect 21681 10289 21727 10300
rect 21068 10252 21079 10255
rect 21133 10252 21144 10255
rect 21252 10252 21263 10255
rect 21317 10252 21328 10255
rect 21436 10252 21447 10255
rect 21501 10252 21512 10255
rect 20991 10206 21037 10217
rect 20899 10032 20991 10206
rect 20991 10021 21037 10032
rect 21175 10206 21221 10217
rect 21175 10021 21221 10032
rect 21359 10206 21405 10217
rect 21543 10206 21589 10217
rect 21526 10179 21543 10181
rect 21589 10179 21606 10181
rect 21526 10059 21538 10179
rect 21594 10059 21606 10179
rect 21526 10057 21543 10059
rect 21359 10021 21405 10032
rect 21589 10057 21606 10059
rect 21543 10021 21589 10032
rect 20853 9804 20899 9949
rect 21068 9940 21079 9986
rect 21133 9940 21144 9986
rect 21068 9907 21144 9940
rect 21252 9940 21263 9986
rect 21317 9940 21328 9986
rect 21252 9907 21328 9940
rect 21436 9940 21447 9986
rect 21501 9940 21512 9986
rect 21436 9907 21512 9940
rect 21681 9804 21727 9949
rect 20841 9792 20921 9804
rect 20841 9736 20853 9792
rect 20909 9736 20921 9792
rect 20841 9724 20921 9736
rect 21659 9792 21739 9804
rect 21659 9736 21671 9792
rect 21727 9736 21739 9792
rect 21659 9724 21739 9736
rect 15914 9618 15926 9674
rect 15982 9618 16228 9674
rect 16284 9618 18178 9674
rect 19956 9674 20026 9686
rect 20268 9674 20328 9678
rect 22164 9674 22220 12611
rect 22920 12609 23000 12611
rect 24436 12666 24506 12678
rect 25476 12666 25556 12668
rect 26962 12667 27042 12669
rect 24436 12610 24448 12666
rect 24504 12610 25488 12666
rect 25544 12610 25556 12666
rect 24436 12598 24506 12610
rect 22552 12517 22632 12531
rect 22339 12495 22385 12506
rect 22552 12461 22564 12517
rect 22620 12461 22632 12517
rect 22736 12517 22816 12531
rect 22736 12461 22748 12517
rect 22804 12461 22816 12517
rect 22920 12517 23000 12531
rect 22920 12461 22932 12517
rect 22988 12461 23000 12517
rect 23167 12495 23213 12506
rect 22554 12458 22565 12461
rect 22619 12458 22630 12461
rect 22738 12458 22749 12461
rect 22803 12458 22814 12461
rect 22922 12458 22933 12461
rect 22987 12458 22998 12461
rect 22477 12412 22523 12423
rect 22385 12238 22477 12412
rect 22477 12227 22523 12238
rect 22661 12412 22707 12423
rect 22661 12227 22707 12238
rect 22845 12412 22891 12423
rect 23029 12412 23075 12423
rect 23012 12385 23029 12387
rect 23075 12385 23092 12387
rect 23012 12265 23024 12385
rect 23080 12265 23092 12385
rect 23012 12263 23029 12265
rect 22845 12227 22891 12238
rect 23075 12263 23092 12265
rect 23029 12227 23075 12238
rect 22339 12010 22385 12155
rect 22554 12146 22565 12192
rect 22619 12146 22630 12192
rect 22554 12113 22630 12146
rect 22738 12146 22749 12192
rect 22803 12146 22814 12192
rect 22738 12113 22814 12146
rect 22922 12146 22933 12192
rect 22987 12146 22998 12192
rect 22922 12113 22998 12146
rect 23167 12010 23213 12155
rect 22327 11998 22407 12010
rect 22327 11942 22339 11998
rect 22395 11942 22407 11998
rect 22327 11930 22407 11942
rect 23145 11998 23223 12010
rect 23145 11942 23157 11998
rect 23213 11942 23223 11998
rect 23145 11930 23223 11942
rect 24720 11879 24776 12610
rect 25476 12608 25556 12610
rect 26206 12611 26974 12667
rect 27030 12611 27042 12667
rect 25108 12516 25188 12530
rect 24895 12494 24941 12505
rect 25108 12460 25120 12516
rect 25176 12460 25188 12516
rect 25292 12516 25372 12530
rect 25292 12460 25304 12516
rect 25360 12460 25372 12516
rect 25476 12516 25556 12530
rect 25476 12460 25488 12516
rect 25544 12460 25556 12516
rect 25723 12494 25769 12505
rect 25110 12457 25121 12460
rect 25175 12457 25186 12460
rect 25294 12457 25305 12460
rect 25359 12457 25370 12460
rect 25478 12457 25489 12460
rect 25543 12457 25554 12460
rect 25033 12411 25079 12422
rect 24941 12237 25033 12411
rect 25033 12226 25079 12237
rect 25217 12411 25263 12422
rect 25217 12226 25263 12237
rect 25401 12411 25447 12422
rect 25585 12411 25631 12422
rect 25568 12384 25585 12386
rect 25631 12384 25648 12386
rect 25568 12264 25580 12384
rect 25636 12264 25648 12384
rect 25568 12262 25585 12264
rect 25401 12226 25447 12237
rect 25631 12262 25648 12264
rect 25585 12226 25631 12237
rect 24895 12009 24941 12154
rect 25110 12145 25121 12191
rect 25175 12145 25186 12191
rect 25110 12112 25186 12145
rect 25294 12145 25305 12191
rect 25359 12145 25370 12191
rect 25294 12112 25370 12145
rect 25478 12145 25489 12191
rect 25543 12145 25554 12191
rect 25478 12112 25554 12145
rect 25723 12009 25769 12154
rect 24883 11997 24963 12009
rect 24883 11941 24895 11997
rect 24951 11941 24963 11997
rect 24883 11929 24963 11941
rect 25701 11997 25779 12009
rect 25701 11941 25713 11997
rect 25769 11941 25779 11997
rect 25701 11929 25779 11941
rect 26054 11879 26134 11889
rect 24720 11823 26066 11879
rect 26122 11823 26134 11879
rect 26054 11821 26134 11823
rect 25888 11770 25958 11772
rect 24720 11769 25958 11770
rect 24720 11715 25890 11769
rect 25946 11715 25958 11769
rect 24720 11714 25958 11715
rect 24720 10693 24776 11714
rect 25888 11706 25958 11714
rect 25384 11662 25470 11666
rect 25384 11606 25396 11662
rect 25452 11606 25470 11662
rect 25384 11594 25470 11606
rect 24895 11449 24941 11460
rect 25110 11458 25186 11491
rect 25110 11412 25121 11458
rect 25175 11412 25186 11458
rect 25294 11458 25370 11491
rect 25294 11412 25305 11458
rect 25359 11412 25370 11458
rect 25478 11458 25554 11491
rect 25478 11412 25489 11458
rect 25543 11412 25554 11458
rect 25723 11449 25769 11460
rect 25033 11366 25079 11377
rect 25016 11339 25033 11341
rect 25217 11366 25263 11377
rect 25079 11339 25096 11341
rect 24941 11219 25028 11339
rect 25084 11219 25096 11339
rect 25016 11217 25033 11219
rect 24941 10919 25033 11039
rect 25079 11217 25096 11219
rect 25200 11039 25217 11041
rect 25401 11366 25447 11377
rect 25384 11339 25401 11341
rect 25585 11366 25631 11377
rect 25447 11339 25464 11341
rect 25384 11219 25396 11339
rect 25452 11219 25464 11339
rect 25384 11217 25401 11219
rect 25263 11039 25280 11041
rect 25200 10919 25212 11039
rect 25268 10919 25280 11039
rect 25200 10917 25217 10919
rect 25033 10881 25079 10892
rect 25263 10917 25280 10919
rect 25217 10881 25263 10892
rect 25447 11217 25464 11219
rect 25568 11039 25585 11041
rect 25706 11339 25723 11341
rect 25769 11339 25786 11341
rect 25706 11218 25718 11339
rect 25774 11218 25786 11339
rect 25706 11216 25723 11218
rect 25631 11039 25648 11041
rect 25568 10919 25580 11039
rect 25636 10919 25648 11039
rect 25568 10917 25585 10919
rect 25401 10881 25447 10892
rect 25631 10917 25648 10919
rect 25585 10881 25631 10892
rect 25110 10843 25121 10846
rect 25175 10843 25186 10846
rect 25294 10843 25305 10846
rect 25359 10843 25370 10846
rect 25478 10843 25489 10846
rect 25543 10843 25554 10846
rect 24895 10798 24941 10809
rect 25108 10787 25120 10843
rect 25176 10787 25188 10843
rect 25108 10773 25188 10787
rect 25292 10787 25304 10843
rect 25360 10787 25372 10843
rect 25292 10773 25372 10787
rect 25476 10787 25488 10843
rect 25544 10787 25556 10843
rect 25769 11216 25786 11218
rect 25723 10798 25769 10809
rect 25476 10773 25556 10787
rect 25108 10693 25188 10695
rect 24720 10637 25120 10693
rect 25176 10637 25188 10693
rect 25108 10635 25188 10637
rect 24300 10577 24370 10591
rect 25292 10577 25372 10579
rect 24300 10521 24312 10577
rect 24368 10521 25304 10577
rect 25360 10521 25372 10577
rect 24300 10509 24370 10521
rect 25292 10519 25372 10521
rect 25621 10577 25701 10579
rect 26064 10577 26124 10589
rect 25621 10521 25633 10577
rect 25689 10521 26066 10577
rect 26122 10521 26124 10577
rect 25621 10519 25701 10521
rect 26064 10509 26124 10521
rect 23454 10461 23524 10473
rect 25476 10461 25556 10463
rect 23454 10405 23466 10461
rect 23522 10405 25488 10461
rect 25544 10405 25556 10461
rect 23454 10393 23524 10405
rect 25476 10403 25556 10405
rect 25108 10311 25188 10325
rect 24895 10289 24941 10300
rect 25108 10255 25120 10311
rect 25176 10255 25188 10311
rect 25292 10311 25372 10325
rect 25292 10255 25304 10311
rect 25360 10255 25372 10311
rect 25476 10311 25556 10325
rect 25476 10255 25488 10311
rect 25544 10255 25556 10311
rect 25723 10289 25769 10300
rect 25110 10252 25121 10255
rect 25175 10252 25186 10255
rect 25294 10252 25305 10255
rect 25359 10252 25370 10255
rect 25478 10252 25489 10255
rect 25543 10252 25554 10255
rect 25033 10206 25079 10217
rect 24941 10032 25033 10206
rect 25033 10021 25079 10032
rect 25217 10206 25263 10217
rect 25217 10021 25263 10032
rect 25401 10206 25447 10217
rect 25585 10206 25631 10217
rect 25568 10179 25585 10181
rect 25631 10179 25648 10181
rect 25568 10059 25580 10179
rect 25636 10059 25648 10179
rect 25568 10057 25585 10059
rect 25401 10021 25447 10032
rect 25631 10057 25648 10059
rect 25585 10021 25631 10032
rect 24895 9804 24941 9949
rect 25110 9940 25121 9986
rect 25175 9940 25186 9986
rect 25110 9907 25186 9940
rect 25294 9940 25305 9986
rect 25359 9940 25370 9986
rect 25294 9907 25370 9940
rect 25478 9940 25489 9986
rect 25543 9940 25554 9986
rect 25478 9907 25554 9940
rect 25723 9804 25769 9949
rect 24883 9792 24963 9804
rect 24883 9736 24895 9792
rect 24951 9736 24963 9792
rect 24883 9724 24963 9736
rect 25701 9792 25781 9804
rect 25701 9736 25713 9792
rect 25769 9736 25781 9792
rect 25701 9724 25781 9736
rect 19956 9618 19968 9674
rect 20024 9618 20270 9674
rect 20326 9618 22220 9674
rect 23998 9674 24068 9686
rect 24310 9674 24370 9678
rect 26206 9674 26262 12611
rect 26962 12609 27042 12611
rect 28478 12666 28548 12678
rect 29518 12666 29598 12668
rect 31004 12667 31084 12669
rect 28478 12610 28490 12666
rect 28546 12610 29530 12666
rect 29586 12610 29598 12666
rect 28478 12598 28548 12610
rect 26594 12517 26674 12531
rect 26381 12495 26427 12506
rect 26594 12461 26606 12517
rect 26662 12461 26674 12517
rect 26778 12517 26858 12531
rect 26778 12461 26790 12517
rect 26846 12461 26858 12517
rect 26962 12517 27042 12531
rect 26962 12461 26974 12517
rect 27030 12461 27042 12517
rect 27209 12495 27255 12506
rect 26596 12458 26607 12461
rect 26661 12458 26672 12461
rect 26780 12458 26791 12461
rect 26845 12458 26856 12461
rect 26964 12458 26975 12461
rect 27029 12458 27040 12461
rect 26519 12412 26565 12423
rect 26427 12238 26519 12412
rect 26519 12227 26565 12238
rect 26703 12412 26749 12423
rect 26703 12227 26749 12238
rect 26887 12412 26933 12423
rect 27071 12412 27117 12423
rect 27054 12385 27071 12387
rect 27117 12385 27134 12387
rect 27054 12265 27066 12385
rect 27122 12265 27134 12385
rect 27054 12263 27071 12265
rect 26887 12227 26933 12238
rect 27117 12263 27134 12265
rect 27071 12227 27117 12238
rect 26381 12010 26427 12155
rect 26596 12146 26607 12192
rect 26661 12146 26672 12192
rect 26596 12113 26672 12146
rect 26780 12146 26791 12192
rect 26845 12146 26856 12192
rect 26780 12113 26856 12146
rect 26964 12146 26975 12192
rect 27029 12146 27040 12192
rect 26964 12113 27040 12146
rect 27209 12010 27255 12155
rect 26369 11998 26449 12010
rect 26369 11942 26381 11998
rect 26437 11942 26449 11998
rect 26369 11930 26449 11942
rect 27187 11998 27265 12010
rect 27187 11942 27199 11998
rect 27255 11942 27265 11998
rect 27187 11930 27265 11942
rect 28762 11879 28818 12610
rect 29518 12608 29598 12610
rect 30248 12611 31016 12667
rect 31072 12611 31084 12667
rect 29150 12516 29230 12530
rect 28937 12494 28983 12505
rect 29150 12460 29162 12516
rect 29218 12460 29230 12516
rect 29334 12516 29414 12530
rect 29334 12460 29346 12516
rect 29402 12460 29414 12516
rect 29518 12516 29598 12530
rect 29518 12460 29530 12516
rect 29586 12460 29598 12516
rect 29765 12494 29811 12505
rect 29152 12457 29163 12460
rect 29217 12457 29228 12460
rect 29336 12457 29347 12460
rect 29401 12457 29412 12460
rect 29520 12457 29531 12460
rect 29585 12457 29596 12460
rect 29075 12411 29121 12422
rect 28983 12237 29075 12411
rect 29075 12226 29121 12237
rect 29259 12411 29305 12422
rect 29259 12226 29305 12237
rect 29443 12411 29489 12422
rect 29627 12411 29673 12422
rect 29610 12384 29627 12386
rect 29673 12384 29690 12386
rect 29610 12264 29622 12384
rect 29678 12264 29690 12384
rect 29610 12262 29627 12264
rect 29443 12226 29489 12237
rect 29673 12262 29690 12264
rect 29627 12226 29673 12237
rect 28937 12009 28983 12154
rect 29152 12145 29163 12191
rect 29217 12145 29228 12191
rect 29152 12112 29228 12145
rect 29336 12145 29347 12191
rect 29401 12145 29412 12191
rect 29336 12112 29412 12145
rect 29520 12145 29531 12191
rect 29585 12145 29596 12191
rect 29520 12112 29596 12145
rect 29765 12009 29811 12154
rect 28925 11997 29005 12009
rect 28925 11941 28937 11997
rect 28993 11941 29005 11997
rect 28925 11929 29005 11941
rect 29743 11997 29821 12009
rect 29743 11941 29755 11997
rect 29811 11941 29821 11997
rect 29743 11929 29821 11941
rect 30096 11879 30176 11889
rect 28762 11823 30108 11879
rect 30164 11823 30176 11879
rect 30096 11821 30176 11823
rect 29930 11770 30000 11772
rect 28762 11769 30000 11770
rect 28762 11715 29932 11769
rect 29988 11715 30000 11769
rect 28762 11714 30000 11715
rect 28762 10693 28818 11714
rect 29930 11706 30000 11714
rect 29426 11662 29512 11666
rect 29426 11606 29438 11662
rect 29494 11606 29512 11662
rect 29426 11594 29512 11606
rect 28937 11449 28983 11460
rect 29152 11458 29228 11491
rect 29152 11412 29163 11458
rect 29217 11412 29228 11458
rect 29336 11458 29412 11491
rect 29336 11412 29347 11458
rect 29401 11412 29412 11458
rect 29520 11458 29596 11491
rect 29520 11412 29531 11458
rect 29585 11412 29596 11458
rect 29765 11449 29811 11460
rect 29075 11366 29121 11377
rect 29058 11339 29075 11341
rect 29259 11366 29305 11377
rect 29121 11339 29138 11341
rect 28983 11219 29070 11339
rect 29126 11219 29138 11339
rect 29058 11217 29075 11219
rect 28983 10919 29075 11039
rect 29121 11217 29138 11219
rect 29242 11039 29259 11041
rect 29443 11366 29489 11377
rect 29426 11339 29443 11341
rect 29627 11366 29673 11377
rect 29489 11339 29506 11341
rect 29426 11219 29438 11339
rect 29494 11219 29506 11339
rect 29426 11217 29443 11219
rect 29305 11039 29322 11041
rect 29242 10919 29254 11039
rect 29310 10919 29322 11039
rect 29242 10917 29259 10919
rect 29075 10881 29121 10892
rect 29305 10917 29322 10919
rect 29259 10881 29305 10892
rect 29489 11217 29506 11219
rect 29610 11039 29627 11041
rect 29748 11339 29765 11341
rect 29811 11339 29828 11341
rect 29748 11218 29760 11339
rect 29816 11218 29828 11339
rect 29748 11216 29765 11218
rect 29673 11039 29690 11041
rect 29610 10919 29622 11039
rect 29678 10919 29690 11039
rect 29610 10917 29627 10919
rect 29443 10881 29489 10892
rect 29673 10917 29690 10919
rect 29627 10881 29673 10892
rect 29152 10843 29163 10846
rect 29217 10843 29228 10846
rect 29336 10843 29347 10846
rect 29401 10843 29412 10846
rect 29520 10843 29531 10846
rect 29585 10843 29596 10846
rect 28937 10798 28983 10809
rect 29150 10787 29162 10843
rect 29218 10787 29230 10843
rect 29150 10773 29230 10787
rect 29334 10787 29346 10843
rect 29402 10787 29414 10843
rect 29334 10773 29414 10787
rect 29518 10787 29530 10843
rect 29586 10787 29598 10843
rect 29811 11216 29828 11218
rect 29765 10798 29811 10809
rect 29518 10773 29598 10787
rect 29150 10693 29230 10695
rect 28762 10637 29162 10693
rect 29218 10637 29230 10693
rect 29150 10635 29230 10637
rect 28342 10577 28412 10591
rect 29334 10577 29414 10579
rect 28342 10521 28354 10577
rect 28410 10521 29346 10577
rect 29402 10521 29414 10577
rect 28342 10509 28412 10521
rect 29334 10519 29414 10521
rect 29663 10577 29743 10579
rect 30106 10577 30166 10589
rect 29663 10521 29675 10577
rect 29731 10521 30108 10577
rect 30164 10521 30166 10577
rect 29663 10519 29743 10521
rect 30106 10509 30166 10521
rect 28162 10461 28240 10473
rect 29518 10461 29598 10463
rect 28162 10405 28173 10461
rect 28229 10405 29530 10461
rect 29586 10405 29598 10461
rect 28162 10393 28240 10405
rect 29518 10403 29598 10405
rect 29150 10311 29230 10325
rect 28937 10289 28983 10300
rect 29150 10255 29162 10311
rect 29218 10255 29230 10311
rect 29334 10311 29414 10325
rect 29334 10255 29346 10311
rect 29402 10255 29414 10311
rect 29518 10311 29598 10325
rect 29518 10255 29530 10311
rect 29586 10255 29598 10311
rect 29765 10289 29811 10300
rect 29152 10252 29163 10255
rect 29217 10252 29228 10255
rect 29336 10252 29347 10255
rect 29401 10252 29412 10255
rect 29520 10252 29531 10255
rect 29585 10252 29596 10255
rect 29075 10206 29121 10217
rect 28983 10032 29075 10206
rect 29075 10021 29121 10032
rect 29259 10206 29305 10217
rect 29259 10021 29305 10032
rect 29443 10206 29489 10217
rect 29627 10206 29673 10217
rect 29610 10179 29627 10181
rect 29673 10179 29690 10181
rect 29610 10059 29622 10179
rect 29678 10059 29690 10179
rect 29610 10057 29627 10059
rect 29443 10021 29489 10032
rect 29673 10057 29690 10059
rect 29627 10021 29673 10032
rect 28937 9804 28983 9949
rect 29152 9940 29163 9986
rect 29217 9940 29228 9986
rect 29152 9907 29228 9940
rect 29336 9940 29347 9986
rect 29401 9940 29412 9986
rect 29336 9907 29412 9940
rect 29520 9940 29531 9986
rect 29585 9940 29596 9986
rect 29520 9907 29596 9940
rect 29765 9804 29811 9949
rect 28925 9792 29005 9804
rect 28925 9736 28937 9792
rect 28993 9736 29005 9792
rect 28925 9724 29005 9736
rect 29743 9792 29823 9804
rect 29743 9736 29755 9792
rect 29811 9736 29823 9792
rect 29743 9724 29823 9736
rect 23998 9618 24010 9674
rect 24066 9618 24312 9674
rect 24368 9618 26262 9674
rect 28040 9674 28110 9686
rect 28352 9674 28412 9678
rect 30248 9674 30304 12611
rect 31004 12609 31084 12611
rect 30636 12517 30716 12531
rect 30423 12495 30469 12506
rect 30636 12461 30648 12517
rect 30704 12461 30716 12517
rect 30820 12517 30900 12531
rect 30820 12461 30832 12517
rect 30888 12461 30900 12517
rect 31004 12517 31084 12531
rect 31004 12461 31016 12517
rect 31072 12461 31084 12517
rect 31251 12495 31297 12506
rect 30638 12458 30649 12461
rect 30703 12458 30714 12461
rect 30822 12458 30833 12461
rect 30887 12458 30898 12461
rect 31006 12458 31017 12461
rect 31071 12458 31082 12461
rect 30561 12412 30607 12423
rect 30469 12238 30561 12412
rect 30561 12227 30607 12238
rect 30745 12412 30791 12423
rect 30745 12227 30791 12238
rect 30929 12412 30975 12423
rect 31113 12412 31159 12423
rect 31096 12385 31113 12387
rect 31159 12385 31176 12387
rect 31096 12265 31108 12385
rect 31164 12265 31176 12385
rect 31096 12263 31113 12265
rect 30929 12227 30975 12238
rect 31159 12263 31176 12265
rect 31113 12227 31159 12238
rect 30423 12010 30469 12155
rect 30638 12146 30649 12192
rect 30703 12146 30714 12192
rect 30638 12113 30714 12146
rect 30822 12146 30833 12192
rect 30887 12146 30898 12192
rect 30822 12113 30898 12146
rect 31006 12146 31017 12192
rect 31071 12146 31082 12192
rect 31006 12113 31082 12146
rect 31251 12010 31297 12155
rect 30411 11998 30491 12010
rect 30411 11942 30423 11998
rect 30479 11942 30491 11998
rect 30411 11930 30491 11942
rect 31229 11998 31307 12010
rect 31229 11942 31241 11998
rect 31297 11942 31307 11998
rect 31229 11930 31307 11942
rect 28040 9618 28052 9674
rect 28108 9618 28354 9674
rect 28410 9618 30304 9674
rect 7830 9616 7900 9618
rect 8142 9606 8202 9618
rect 11872 9616 11942 9618
rect 12184 9606 12244 9618
rect 15914 9616 15984 9618
rect 16226 9606 16286 9618
rect 19956 9616 20026 9618
rect 20268 9606 20328 9618
rect 23998 9616 24068 9618
rect 24310 9606 24370 9618
rect 28040 9606 28110 9618
rect 28352 9606 28412 9618
rect 493 8753 2040 8809
rect -58 7732 12 7744
rect 493 7732 549 8753
rect 1162 8701 1248 8705
rect 1162 8645 1174 8701
rect 1230 8645 1248 8701
rect 1162 8633 1248 8645
rect 673 8488 719 8499
rect 888 8497 964 8530
rect 888 8451 899 8497
rect 953 8451 964 8497
rect 1072 8497 1148 8530
rect 1072 8451 1083 8497
rect 1137 8451 1148 8497
rect 1256 8497 1332 8530
rect 1256 8451 1267 8497
rect 1321 8451 1332 8497
rect 1501 8488 1547 8499
rect 811 8405 857 8416
rect 794 8378 811 8380
rect 995 8405 1041 8416
rect 857 8378 874 8380
rect 719 8258 806 8378
rect 862 8258 874 8378
rect 794 8256 811 8258
rect 719 7958 811 8078
rect 857 8256 874 8258
rect 978 8078 995 8080
rect 1179 8405 1225 8416
rect 1162 8378 1179 8380
rect 1363 8405 1409 8416
rect 1225 8378 1242 8380
rect 1162 8258 1174 8378
rect 1230 8258 1242 8378
rect 1162 8256 1179 8258
rect 1041 8078 1058 8080
rect 978 7958 990 8078
rect 1046 7958 1058 8078
rect 978 7956 995 7958
rect 811 7920 857 7931
rect 1041 7956 1058 7958
rect 995 7920 1041 7931
rect 1225 8256 1242 8258
rect 1346 8078 1363 8080
rect 1484 8378 1501 8380
rect 1547 8378 1564 8380
rect 1484 8257 1496 8378
rect 1552 8257 1564 8378
rect 1484 8255 1501 8257
rect 1409 8078 1426 8080
rect 1346 7958 1358 8078
rect 1414 7958 1426 8078
rect 1346 7956 1363 7958
rect 1179 7920 1225 7931
rect 1409 7956 1426 7958
rect 1363 7920 1409 7931
rect 888 7882 899 7885
rect 953 7882 964 7885
rect 1072 7882 1083 7885
rect 1137 7882 1148 7885
rect 1256 7882 1267 7885
rect 1321 7882 1332 7885
rect 673 7837 719 7848
rect 886 7826 898 7882
rect 954 7826 966 7882
rect 886 7812 966 7826
rect 1070 7826 1082 7882
rect 1138 7826 1150 7882
rect 1070 7812 1150 7826
rect 1254 7826 1266 7882
rect 1322 7826 1334 7882
rect 1547 8255 1564 8257
rect 1501 7837 1547 7848
rect 1254 7812 1334 7826
rect 886 7732 966 7734
rect -58 7676 -46 7732
rect 10 7676 898 7732
rect 954 7676 966 7732
rect -58 7664 12 7676
rect 886 7674 966 7676
rect 214 7616 284 7628
rect 1070 7616 1150 7618
rect 214 7560 226 7616
rect 282 7560 1082 7616
rect 1138 7560 1150 7616
rect 214 7548 284 7560
rect 1070 7558 1150 7560
rect 1399 7616 1479 7618
rect 1666 7616 1736 7628
rect 1399 7560 1411 7616
rect 1467 7560 1668 7616
rect 1724 7560 1736 7616
rect 1399 7558 1479 7560
rect 1666 7550 1736 7560
rect 1254 7500 1334 7502
rect 498 7444 1266 7500
rect 1322 7444 1334 7500
rect 498 6713 554 7444
rect 1254 7442 1334 7444
rect 886 7350 966 7364
rect 673 7328 719 7339
rect 886 7294 898 7350
rect 954 7294 966 7350
rect 1070 7350 1150 7364
rect 1070 7294 1082 7350
rect 1138 7294 1150 7350
rect 1254 7350 1334 7364
rect 1254 7294 1266 7350
rect 1322 7294 1334 7350
rect 1501 7328 1547 7339
rect 888 7291 899 7294
rect 953 7291 964 7294
rect 1072 7291 1083 7294
rect 1137 7291 1148 7294
rect 1256 7291 1267 7294
rect 1321 7291 1332 7294
rect 811 7245 857 7256
rect 719 7071 811 7245
rect 811 7060 857 7071
rect 995 7245 1041 7256
rect 995 7060 1041 7071
rect 1179 7245 1225 7256
rect 1363 7245 1409 7256
rect 1346 7218 1363 7220
rect 1409 7218 1426 7220
rect 1346 7098 1358 7218
rect 1414 7098 1426 7218
rect 1346 7096 1363 7098
rect 1179 7060 1225 7071
rect 1409 7096 1426 7098
rect 1363 7060 1409 7071
rect 673 6843 719 6988
rect 888 6979 899 7025
rect 953 6979 964 7025
rect 888 6946 964 6979
rect 1072 6979 1083 7025
rect 1137 6979 1148 7025
rect 1072 6946 1148 6979
rect 1256 6979 1267 7025
rect 1321 6979 1332 7025
rect 1256 6946 1332 6979
rect 1501 6843 1547 6988
rect 661 6831 741 6843
rect 661 6775 673 6831
rect 729 6775 741 6831
rect 661 6763 741 6775
rect 1479 6831 1559 6843
rect 1479 6775 1491 6831
rect 1547 6775 1559 6831
rect 1479 6763 1559 6775
rect 1832 6713 1912 6723
rect 498 6657 1844 6713
rect 1900 6657 1912 6713
rect 1832 6655 1912 6657
rect 1666 6604 1736 6606
rect 498 6603 1736 6604
rect 498 6549 1668 6603
rect 1724 6549 1736 6603
rect 498 6548 1736 6549
rect 498 5527 554 6548
rect 1666 6540 1736 6548
rect 1162 6496 1248 6500
rect 1162 6440 1174 6496
rect 1230 6440 1248 6496
rect 1162 6428 1248 6440
rect 673 6283 719 6294
rect 888 6292 964 6325
rect 888 6246 899 6292
rect 953 6246 964 6292
rect 1072 6292 1148 6325
rect 1072 6246 1083 6292
rect 1137 6246 1148 6292
rect 1256 6292 1332 6325
rect 1256 6246 1267 6292
rect 1321 6246 1332 6292
rect 1501 6283 1547 6294
rect 811 6200 857 6211
rect 794 6173 811 6175
rect 995 6200 1041 6211
rect 857 6173 874 6175
rect 719 6053 806 6173
rect 862 6053 874 6173
rect 794 6051 811 6053
rect 719 5753 811 5873
rect 857 6051 874 6053
rect 978 5873 995 5875
rect 1179 6200 1225 6211
rect 1162 6173 1179 6175
rect 1363 6200 1409 6211
rect 1225 6173 1242 6175
rect 1162 6053 1174 6173
rect 1230 6053 1242 6173
rect 1162 6051 1179 6053
rect 1041 5873 1058 5875
rect 978 5753 990 5873
rect 1046 5753 1058 5873
rect 978 5751 995 5753
rect 811 5715 857 5726
rect 1041 5751 1058 5753
rect 995 5715 1041 5726
rect 1225 6051 1242 6053
rect 1346 5873 1363 5875
rect 1484 6173 1501 6175
rect 1547 6173 1564 6175
rect 1484 6052 1496 6173
rect 1552 6052 1564 6173
rect 1484 6050 1501 6052
rect 1409 5873 1426 5875
rect 1346 5753 1358 5873
rect 1414 5753 1426 5873
rect 1346 5751 1363 5753
rect 1179 5715 1225 5726
rect 1409 5751 1426 5753
rect 1363 5715 1409 5726
rect 888 5677 899 5680
rect 953 5677 964 5680
rect 1072 5677 1083 5680
rect 1137 5677 1148 5680
rect 1256 5677 1267 5680
rect 1321 5677 1332 5680
rect 673 5632 719 5643
rect 886 5621 898 5677
rect 954 5621 966 5677
rect 886 5607 966 5621
rect 1070 5621 1082 5677
rect 1138 5621 1150 5677
rect 1070 5607 1150 5621
rect 1254 5621 1266 5677
rect 1322 5621 1334 5677
rect 1547 6050 1564 6052
rect 1501 5632 1547 5643
rect 1254 5607 1334 5621
rect 886 5527 966 5529
rect 498 5471 898 5527
rect 954 5471 966 5527
rect 1984 5527 2040 8753
rect 4505 8753 6052 8809
rect 4010 7732 4096 7744
rect 4505 7732 4561 8753
rect 5174 8701 5260 8705
rect 5174 8645 5186 8701
rect 5242 8645 5260 8701
rect 5174 8633 5260 8645
rect 4685 8488 4731 8499
rect 4900 8497 4976 8530
rect 4900 8451 4911 8497
rect 4965 8451 4976 8497
rect 5084 8497 5160 8530
rect 5084 8451 5095 8497
rect 5149 8451 5160 8497
rect 5268 8497 5344 8530
rect 5268 8451 5279 8497
rect 5333 8451 5344 8497
rect 5513 8488 5559 8499
rect 4823 8405 4869 8416
rect 4806 8378 4823 8380
rect 5007 8405 5053 8416
rect 4869 8378 4886 8380
rect 4731 8258 4818 8378
rect 4874 8258 4886 8378
rect 4806 8256 4823 8258
rect 4731 7958 4823 8078
rect 4869 8256 4886 8258
rect 4990 8078 5007 8080
rect 5191 8405 5237 8416
rect 5174 8378 5191 8380
rect 5375 8405 5421 8416
rect 5237 8378 5254 8380
rect 5174 8258 5186 8378
rect 5242 8258 5254 8378
rect 5174 8256 5191 8258
rect 5053 8078 5070 8080
rect 4990 7958 5002 8078
rect 5058 7958 5070 8078
rect 4990 7956 5007 7958
rect 4823 7920 4869 7931
rect 5053 7956 5070 7958
rect 5007 7920 5053 7931
rect 5237 8256 5254 8258
rect 5358 8078 5375 8080
rect 5496 8378 5513 8380
rect 5559 8378 5576 8380
rect 5496 8257 5508 8378
rect 5564 8257 5576 8378
rect 5496 8255 5513 8257
rect 5421 8078 5438 8080
rect 5358 7958 5370 8078
rect 5426 7958 5438 8078
rect 5358 7956 5375 7958
rect 5191 7920 5237 7931
rect 5421 7956 5438 7958
rect 5375 7920 5421 7931
rect 4900 7882 4911 7885
rect 4965 7882 4976 7885
rect 5084 7882 5095 7885
rect 5149 7882 5160 7885
rect 5268 7882 5279 7885
rect 5333 7882 5344 7885
rect 4685 7837 4731 7848
rect 4898 7826 4910 7882
rect 4966 7826 4978 7882
rect 4898 7812 4978 7826
rect 5082 7826 5094 7882
rect 5150 7826 5162 7882
rect 5082 7812 5162 7826
rect 5266 7826 5278 7882
rect 5334 7826 5346 7882
rect 5559 8255 5576 8257
rect 5513 7837 5559 7848
rect 5266 7812 5346 7826
rect 4898 7732 4978 7734
rect 4010 7676 4022 7732
rect 4078 7676 4910 7732
rect 4966 7676 4978 7732
rect 4010 7664 4096 7676
rect 4898 7674 4978 7676
rect 4226 7616 4296 7628
rect 5082 7616 5162 7618
rect 4226 7560 4238 7616
rect 4294 7560 5094 7616
rect 5150 7560 5162 7616
rect 4226 7548 4296 7560
rect 5082 7558 5162 7560
rect 5411 7616 5491 7618
rect 5678 7616 5748 7628
rect 5411 7560 5423 7616
rect 5479 7560 5680 7616
rect 5736 7560 5748 7616
rect 5411 7558 5491 7560
rect 5678 7550 5748 7560
rect 5266 7500 5346 7502
rect 4510 7444 5278 7500
rect 5334 7444 5346 7500
rect 4510 6713 4566 7444
rect 5266 7442 5346 7444
rect 4898 7350 4978 7364
rect 4685 7328 4731 7339
rect 4898 7294 4910 7350
rect 4966 7294 4978 7350
rect 5082 7350 5162 7364
rect 5082 7294 5094 7350
rect 5150 7294 5162 7350
rect 5266 7350 5346 7364
rect 5266 7294 5278 7350
rect 5334 7294 5346 7350
rect 5513 7328 5559 7339
rect 4900 7291 4911 7294
rect 4965 7291 4976 7294
rect 5084 7291 5095 7294
rect 5149 7291 5160 7294
rect 5268 7291 5279 7294
rect 5333 7291 5344 7294
rect 4823 7245 4869 7256
rect 4731 7071 4823 7245
rect 4823 7060 4869 7071
rect 5007 7245 5053 7256
rect 5007 7060 5053 7071
rect 5191 7245 5237 7256
rect 5375 7245 5421 7256
rect 5358 7218 5375 7220
rect 5421 7218 5438 7220
rect 5358 7098 5370 7218
rect 5426 7098 5438 7218
rect 5358 7096 5375 7098
rect 5191 7060 5237 7071
rect 5421 7096 5438 7098
rect 5375 7060 5421 7071
rect 4685 6843 4731 6988
rect 4900 6979 4911 7025
rect 4965 6979 4976 7025
rect 4900 6946 4976 6979
rect 5084 6979 5095 7025
rect 5149 6979 5160 7025
rect 5084 6946 5160 6979
rect 5268 6979 5279 7025
rect 5333 6979 5344 7025
rect 5268 6946 5344 6979
rect 5513 6843 5559 6988
rect 4673 6831 4753 6843
rect 4673 6775 4685 6831
rect 4741 6775 4753 6831
rect 4673 6763 4753 6775
rect 5491 6831 5571 6843
rect 5491 6775 5503 6831
rect 5559 6775 5571 6831
rect 5491 6763 5571 6775
rect 5844 6713 5924 6723
rect 4510 6657 5856 6713
rect 5912 6657 5924 6713
rect 5844 6655 5924 6657
rect 5678 6604 5748 6606
rect 4510 6603 5748 6604
rect 4510 6549 5680 6603
rect 5736 6549 5748 6603
rect 4510 6548 5748 6549
rect 2648 6496 2734 6500
rect 2648 6440 2660 6496
rect 2716 6440 2734 6496
rect 2648 6428 2734 6440
rect 2159 6283 2205 6294
rect 2374 6292 2450 6325
rect 2374 6246 2385 6292
rect 2439 6246 2450 6292
rect 2558 6292 2634 6325
rect 2558 6246 2569 6292
rect 2623 6246 2634 6292
rect 2742 6292 2818 6325
rect 2742 6246 2753 6292
rect 2807 6246 2818 6292
rect 2987 6283 3033 6294
rect 2297 6200 2343 6211
rect 2280 6173 2297 6175
rect 2481 6200 2527 6211
rect 2343 6173 2360 6175
rect 2205 6053 2292 6173
rect 2348 6053 2360 6173
rect 2280 6051 2297 6053
rect 2205 5753 2297 5873
rect 2343 6051 2360 6053
rect 2464 5873 2481 5875
rect 2665 6200 2711 6211
rect 2648 6173 2665 6175
rect 2849 6200 2895 6211
rect 2711 6173 2728 6175
rect 2648 6053 2660 6173
rect 2716 6053 2728 6173
rect 2648 6051 2665 6053
rect 2527 5873 2544 5875
rect 2464 5753 2476 5873
rect 2532 5753 2544 5873
rect 2464 5751 2481 5753
rect 2297 5715 2343 5726
rect 2527 5751 2544 5753
rect 2481 5715 2527 5726
rect 2711 6051 2728 6053
rect 2832 5873 2849 5875
rect 2970 6173 2987 6175
rect 3033 6173 3050 6175
rect 2970 6052 2982 6173
rect 3038 6052 3050 6173
rect 2970 6050 2987 6052
rect 2895 5873 2912 5875
rect 2832 5753 2844 5873
rect 2900 5753 2912 5873
rect 2832 5751 2849 5753
rect 2665 5715 2711 5726
rect 2895 5751 2912 5753
rect 2849 5715 2895 5726
rect 2374 5677 2385 5680
rect 2439 5677 2450 5680
rect 2558 5677 2569 5680
rect 2623 5677 2634 5680
rect 2742 5677 2753 5680
rect 2807 5677 2818 5680
rect 2159 5632 2205 5643
rect 2372 5621 2384 5677
rect 2440 5621 2452 5677
rect 2372 5607 2452 5621
rect 2556 5621 2568 5677
rect 2624 5621 2636 5677
rect 2556 5607 2636 5621
rect 2740 5621 2752 5677
rect 2808 5621 2820 5677
rect 3033 6050 3050 6052
rect 2987 5632 3033 5643
rect 2740 5607 2820 5621
rect 2372 5527 2452 5529
rect 1984 5471 2384 5527
rect 2440 5471 2452 5527
rect 4510 5527 4566 6548
rect 5678 6540 5748 6548
rect 5174 6496 5260 6500
rect 5174 6440 5186 6496
rect 5242 6440 5260 6496
rect 5174 6428 5260 6440
rect 4685 6283 4731 6294
rect 4900 6292 4976 6325
rect 4900 6246 4911 6292
rect 4965 6246 4976 6292
rect 5084 6292 5160 6325
rect 5084 6246 5095 6292
rect 5149 6246 5160 6292
rect 5268 6292 5344 6325
rect 5268 6246 5279 6292
rect 5333 6246 5344 6292
rect 5513 6283 5559 6294
rect 4823 6200 4869 6211
rect 4806 6173 4823 6175
rect 5007 6200 5053 6211
rect 4869 6173 4886 6175
rect 4731 6053 4818 6173
rect 4874 6053 4886 6173
rect 4806 6051 4823 6053
rect 4731 5753 4823 5873
rect 4869 6051 4886 6053
rect 4990 5873 5007 5875
rect 5191 6200 5237 6211
rect 5174 6173 5191 6175
rect 5375 6200 5421 6211
rect 5237 6173 5254 6175
rect 5174 6053 5186 6173
rect 5242 6053 5254 6173
rect 5174 6051 5191 6053
rect 5053 5873 5070 5875
rect 4990 5753 5002 5873
rect 5058 5753 5070 5873
rect 4990 5751 5007 5753
rect 4823 5715 4869 5726
rect 5053 5751 5070 5753
rect 5007 5715 5053 5726
rect 5237 6051 5254 6053
rect 5358 5873 5375 5875
rect 5496 6173 5513 6175
rect 5559 6173 5576 6175
rect 5496 6052 5508 6173
rect 5564 6052 5576 6173
rect 5496 6050 5513 6052
rect 5421 5873 5438 5875
rect 5358 5753 5370 5873
rect 5426 5753 5438 5873
rect 5358 5751 5375 5753
rect 5191 5715 5237 5726
rect 5421 5751 5438 5753
rect 5375 5715 5421 5726
rect 4900 5677 4911 5680
rect 4965 5677 4976 5680
rect 5084 5677 5095 5680
rect 5149 5677 5160 5680
rect 5268 5677 5279 5680
rect 5333 5677 5344 5680
rect 4685 5632 4731 5643
rect 4898 5621 4910 5677
rect 4966 5621 4978 5677
rect 4898 5607 4978 5621
rect 5082 5621 5094 5677
rect 5150 5621 5162 5677
rect 5082 5607 5162 5621
rect 5266 5621 5278 5677
rect 5334 5621 5346 5677
rect 5559 6050 5576 6052
rect 5513 5632 5559 5643
rect 5266 5607 5346 5621
rect 4898 5527 4978 5529
rect 4510 5471 4910 5527
rect 4966 5471 4978 5527
rect 5996 5527 6052 8753
rect 8547 8753 10094 8809
rect 8052 7732 8138 7744
rect 8547 7732 8603 8753
rect 9216 8701 9302 8705
rect 9216 8645 9228 8701
rect 9284 8645 9302 8701
rect 9216 8633 9302 8645
rect 8727 8488 8773 8499
rect 8942 8497 9018 8530
rect 8942 8451 8953 8497
rect 9007 8451 9018 8497
rect 9126 8497 9202 8530
rect 9126 8451 9137 8497
rect 9191 8451 9202 8497
rect 9310 8497 9386 8530
rect 9310 8451 9321 8497
rect 9375 8451 9386 8497
rect 9555 8488 9601 8499
rect 8865 8405 8911 8416
rect 8848 8378 8865 8380
rect 9049 8405 9095 8416
rect 8911 8378 8928 8380
rect 8773 8258 8860 8378
rect 8916 8258 8928 8378
rect 8848 8256 8865 8258
rect 8773 7958 8865 8078
rect 8911 8256 8928 8258
rect 9032 8078 9049 8080
rect 9233 8405 9279 8416
rect 9216 8378 9233 8380
rect 9417 8405 9463 8416
rect 9279 8378 9296 8380
rect 9216 8258 9228 8378
rect 9284 8258 9296 8378
rect 9216 8256 9233 8258
rect 9095 8078 9112 8080
rect 9032 7958 9044 8078
rect 9100 7958 9112 8078
rect 9032 7956 9049 7958
rect 8865 7920 8911 7931
rect 9095 7956 9112 7958
rect 9049 7920 9095 7931
rect 9279 8256 9296 8258
rect 9400 8078 9417 8080
rect 9538 8378 9555 8380
rect 9601 8378 9618 8380
rect 9538 8257 9550 8378
rect 9606 8257 9618 8378
rect 9538 8255 9555 8257
rect 9463 8078 9480 8080
rect 9400 7958 9412 8078
rect 9468 7958 9480 8078
rect 9400 7956 9417 7958
rect 9233 7920 9279 7931
rect 9463 7956 9480 7958
rect 9417 7920 9463 7931
rect 8942 7882 8953 7885
rect 9007 7882 9018 7885
rect 9126 7882 9137 7885
rect 9191 7882 9202 7885
rect 9310 7882 9321 7885
rect 9375 7882 9386 7885
rect 8727 7837 8773 7848
rect 8940 7826 8952 7882
rect 9008 7826 9020 7882
rect 8940 7812 9020 7826
rect 9124 7826 9136 7882
rect 9192 7826 9204 7882
rect 9124 7812 9204 7826
rect 9308 7826 9320 7882
rect 9376 7826 9388 7882
rect 9601 8255 9618 8257
rect 9555 7837 9601 7848
rect 9308 7812 9388 7826
rect 8940 7732 9020 7734
rect 8052 7676 8064 7732
rect 8120 7676 8952 7732
rect 9008 7676 9020 7732
rect 8052 7664 8138 7676
rect 8940 7674 9020 7676
rect 8268 7616 8338 7628
rect 9124 7616 9204 7618
rect 8268 7560 8280 7616
rect 8336 7560 9136 7616
rect 9192 7560 9204 7616
rect 8268 7548 8338 7560
rect 9124 7558 9204 7560
rect 9453 7616 9533 7618
rect 9720 7616 9790 7628
rect 9453 7560 9465 7616
rect 9521 7560 9722 7616
rect 9778 7560 9790 7616
rect 9453 7558 9533 7560
rect 9720 7550 9790 7560
rect 9308 7500 9388 7502
rect 8552 7444 9320 7500
rect 9376 7444 9388 7500
rect 8552 6713 8608 7444
rect 9308 7442 9388 7444
rect 8940 7350 9020 7364
rect 8727 7328 8773 7339
rect 8940 7294 8952 7350
rect 9008 7294 9020 7350
rect 9124 7350 9204 7364
rect 9124 7294 9136 7350
rect 9192 7294 9204 7350
rect 9308 7350 9388 7364
rect 9308 7294 9320 7350
rect 9376 7294 9388 7350
rect 9555 7328 9601 7339
rect 8942 7291 8953 7294
rect 9007 7291 9018 7294
rect 9126 7291 9137 7294
rect 9191 7291 9202 7294
rect 9310 7291 9321 7294
rect 9375 7291 9386 7294
rect 8865 7245 8911 7256
rect 8773 7071 8865 7245
rect 8865 7060 8911 7071
rect 9049 7245 9095 7256
rect 9049 7060 9095 7071
rect 9233 7245 9279 7256
rect 9417 7245 9463 7256
rect 9400 7218 9417 7220
rect 9463 7218 9480 7220
rect 9400 7098 9412 7218
rect 9468 7098 9480 7218
rect 9400 7096 9417 7098
rect 9233 7060 9279 7071
rect 9463 7096 9480 7098
rect 9417 7060 9463 7071
rect 8727 6843 8773 6988
rect 8942 6979 8953 7025
rect 9007 6979 9018 7025
rect 8942 6946 9018 6979
rect 9126 6979 9137 7025
rect 9191 6979 9202 7025
rect 9126 6946 9202 6979
rect 9310 6979 9321 7025
rect 9375 6979 9386 7025
rect 9310 6946 9386 6979
rect 9555 6843 9601 6988
rect 8715 6831 8795 6843
rect 8715 6775 8727 6831
rect 8783 6775 8795 6831
rect 8715 6763 8795 6775
rect 9533 6831 9613 6843
rect 9533 6775 9545 6831
rect 9601 6775 9613 6831
rect 9533 6763 9613 6775
rect 9886 6713 9966 6723
rect 8552 6657 9898 6713
rect 9954 6657 9966 6713
rect 9886 6655 9966 6657
rect 9720 6604 9790 6606
rect 8552 6603 9790 6604
rect 8552 6549 9722 6603
rect 9778 6549 9790 6603
rect 8552 6548 9790 6549
rect 6660 6496 6746 6500
rect 6660 6440 6672 6496
rect 6728 6440 6746 6496
rect 6660 6428 6746 6440
rect 6171 6283 6217 6294
rect 6386 6292 6462 6325
rect 6386 6246 6397 6292
rect 6451 6246 6462 6292
rect 6570 6292 6646 6325
rect 6570 6246 6581 6292
rect 6635 6246 6646 6292
rect 6754 6292 6830 6325
rect 6754 6246 6765 6292
rect 6819 6246 6830 6292
rect 6999 6283 7045 6294
rect 6309 6200 6355 6211
rect 6292 6173 6309 6175
rect 6493 6200 6539 6211
rect 6355 6173 6372 6175
rect 6217 6053 6304 6173
rect 6360 6053 6372 6173
rect 6292 6051 6309 6053
rect 6217 5753 6309 5873
rect 6355 6051 6372 6053
rect 6476 5873 6493 5875
rect 6677 6200 6723 6211
rect 6660 6173 6677 6175
rect 6861 6200 6907 6211
rect 6723 6173 6740 6175
rect 6660 6053 6672 6173
rect 6728 6053 6740 6173
rect 6660 6051 6677 6053
rect 6539 5873 6556 5875
rect 6476 5753 6488 5873
rect 6544 5753 6556 5873
rect 6476 5751 6493 5753
rect 6309 5715 6355 5726
rect 6539 5751 6556 5753
rect 6493 5715 6539 5726
rect 6723 6051 6740 6053
rect 6844 5873 6861 5875
rect 6982 6173 6999 6175
rect 7045 6173 7062 6175
rect 6982 6052 6994 6173
rect 7050 6052 7062 6173
rect 6982 6050 6999 6052
rect 6907 5873 6924 5875
rect 6844 5753 6856 5873
rect 6912 5753 6924 5873
rect 6844 5751 6861 5753
rect 6677 5715 6723 5726
rect 6907 5751 6924 5753
rect 6861 5715 6907 5726
rect 6386 5677 6397 5680
rect 6451 5677 6462 5680
rect 6570 5677 6581 5680
rect 6635 5677 6646 5680
rect 6754 5677 6765 5680
rect 6819 5677 6830 5680
rect 6171 5632 6217 5643
rect 6384 5621 6396 5677
rect 6452 5621 6464 5677
rect 6384 5607 6464 5621
rect 6568 5621 6580 5677
rect 6636 5621 6648 5677
rect 6568 5607 6648 5621
rect 6752 5621 6764 5677
rect 6820 5621 6832 5677
rect 7045 6050 7062 6052
rect 6999 5632 7045 5643
rect 6752 5607 6832 5621
rect 6384 5527 6464 5529
rect 5996 5471 6396 5527
rect 6452 5471 6464 5527
rect 8552 5527 8608 6548
rect 9720 6540 9790 6548
rect 9216 6496 9302 6500
rect 9216 6440 9228 6496
rect 9284 6440 9302 6496
rect 9216 6428 9302 6440
rect 8727 6283 8773 6294
rect 8942 6292 9018 6325
rect 8942 6246 8953 6292
rect 9007 6246 9018 6292
rect 9126 6292 9202 6325
rect 9126 6246 9137 6292
rect 9191 6246 9202 6292
rect 9310 6292 9386 6325
rect 9310 6246 9321 6292
rect 9375 6246 9386 6292
rect 9555 6283 9601 6294
rect 8865 6200 8911 6211
rect 8848 6173 8865 6175
rect 9049 6200 9095 6211
rect 8911 6173 8928 6175
rect 8773 6053 8860 6173
rect 8916 6053 8928 6173
rect 8848 6051 8865 6053
rect 8773 5753 8865 5873
rect 8911 6051 8928 6053
rect 9032 5873 9049 5875
rect 9233 6200 9279 6211
rect 9216 6173 9233 6175
rect 9417 6200 9463 6211
rect 9279 6173 9296 6175
rect 9216 6053 9228 6173
rect 9284 6053 9296 6173
rect 9216 6051 9233 6053
rect 9095 5873 9112 5875
rect 9032 5753 9044 5873
rect 9100 5753 9112 5873
rect 9032 5751 9049 5753
rect 8865 5715 8911 5726
rect 9095 5751 9112 5753
rect 9049 5715 9095 5726
rect 9279 6051 9296 6053
rect 9400 5873 9417 5875
rect 9538 6173 9555 6175
rect 9601 6173 9618 6175
rect 9538 6052 9550 6173
rect 9606 6052 9618 6173
rect 9538 6050 9555 6052
rect 9463 5873 9480 5875
rect 9400 5753 9412 5873
rect 9468 5753 9480 5873
rect 9400 5751 9417 5753
rect 9233 5715 9279 5726
rect 9463 5751 9480 5753
rect 9417 5715 9463 5726
rect 8942 5677 8953 5680
rect 9007 5677 9018 5680
rect 9126 5677 9137 5680
rect 9191 5677 9202 5680
rect 9310 5677 9321 5680
rect 9375 5677 9386 5680
rect 8727 5632 8773 5643
rect 8940 5621 8952 5677
rect 9008 5621 9020 5677
rect 8940 5607 9020 5621
rect 9124 5621 9136 5677
rect 9192 5621 9204 5677
rect 9124 5607 9204 5621
rect 9308 5621 9320 5677
rect 9376 5621 9388 5677
rect 9601 6050 9618 6052
rect 9555 5632 9601 5643
rect 9308 5607 9388 5621
rect 8940 5527 9020 5529
rect 8552 5471 8952 5527
rect 9008 5471 9020 5527
rect 10038 5527 10094 8753
rect 12589 8753 14136 8809
rect 12094 7732 12180 7744
rect 12589 7732 12645 8753
rect 13258 8701 13344 8705
rect 13258 8645 13270 8701
rect 13326 8645 13344 8701
rect 13258 8633 13344 8645
rect 12769 8488 12815 8499
rect 12984 8497 13060 8530
rect 12984 8451 12995 8497
rect 13049 8451 13060 8497
rect 13168 8497 13244 8530
rect 13168 8451 13179 8497
rect 13233 8451 13244 8497
rect 13352 8497 13428 8530
rect 13352 8451 13363 8497
rect 13417 8451 13428 8497
rect 13597 8488 13643 8499
rect 12907 8405 12953 8416
rect 12890 8378 12907 8380
rect 13091 8405 13137 8416
rect 12953 8378 12970 8380
rect 12815 8258 12902 8378
rect 12958 8258 12970 8378
rect 12890 8256 12907 8258
rect 12815 7958 12907 8078
rect 12953 8256 12970 8258
rect 13074 8078 13091 8080
rect 13275 8405 13321 8416
rect 13258 8378 13275 8380
rect 13459 8405 13505 8416
rect 13321 8378 13338 8380
rect 13258 8258 13270 8378
rect 13326 8258 13338 8378
rect 13258 8256 13275 8258
rect 13137 8078 13154 8080
rect 13074 7958 13086 8078
rect 13142 7958 13154 8078
rect 13074 7956 13091 7958
rect 12907 7920 12953 7931
rect 13137 7956 13154 7958
rect 13091 7920 13137 7931
rect 13321 8256 13338 8258
rect 13442 8078 13459 8080
rect 13580 8378 13597 8380
rect 13643 8378 13660 8380
rect 13580 8257 13592 8378
rect 13648 8257 13660 8378
rect 13580 8255 13597 8257
rect 13505 8078 13522 8080
rect 13442 7958 13454 8078
rect 13510 7958 13522 8078
rect 13442 7956 13459 7958
rect 13275 7920 13321 7931
rect 13505 7956 13522 7958
rect 13459 7920 13505 7931
rect 12984 7882 12995 7885
rect 13049 7882 13060 7885
rect 13168 7882 13179 7885
rect 13233 7882 13244 7885
rect 13352 7882 13363 7885
rect 13417 7882 13428 7885
rect 12769 7837 12815 7848
rect 12982 7826 12994 7882
rect 13050 7826 13062 7882
rect 12982 7812 13062 7826
rect 13166 7826 13178 7882
rect 13234 7826 13246 7882
rect 13166 7812 13246 7826
rect 13350 7826 13362 7882
rect 13418 7826 13430 7882
rect 13643 8255 13660 8257
rect 13597 7837 13643 7848
rect 13350 7812 13430 7826
rect 12982 7732 13062 7734
rect 12094 7676 12106 7732
rect 12162 7676 12994 7732
rect 13050 7676 13062 7732
rect 12094 7664 12180 7676
rect 12982 7674 13062 7676
rect 12310 7616 12380 7628
rect 13166 7616 13246 7618
rect 12310 7560 12322 7616
rect 12378 7560 13178 7616
rect 13234 7560 13246 7616
rect 12310 7548 12380 7560
rect 13166 7558 13246 7560
rect 13495 7616 13575 7618
rect 13762 7616 13832 7628
rect 13495 7560 13507 7616
rect 13563 7560 13764 7616
rect 13820 7560 13832 7616
rect 13495 7558 13575 7560
rect 13762 7550 13832 7560
rect 13350 7500 13430 7502
rect 12594 7444 13362 7500
rect 13418 7444 13430 7500
rect 12594 6713 12650 7444
rect 13350 7442 13430 7444
rect 12982 7350 13062 7364
rect 12769 7328 12815 7339
rect 12982 7294 12994 7350
rect 13050 7294 13062 7350
rect 13166 7350 13246 7364
rect 13166 7294 13178 7350
rect 13234 7294 13246 7350
rect 13350 7350 13430 7364
rect 13350 7294 13362 7350
rect 13418 7294 13430 7350
rect 13597 7328 13643 7339
rect 12984 7291 12995 7294
rect 13049 7291 13060 7294
rect 13168 7291 13179 7294
rect 13233 7291 13244 7294
rect 13352 7291 13363 7294
rect 13417 7291 13428 7294
rect 12907 7245 12953 7256
rect 12815 7071 12907 7245
rect 12907 7060 12953 7071
rect 13091 7245 13137 7256
rect 13091 7060 13137 7071
rect 13275 7245 13321 7256
rect 13459 7245 13505 7256
rect 13442 7218 13459 7220
rect 13505 7218 13522 7220
rect 13442 7098 13454 7218
rect 13510 7098 13522 7218
rect 13442 7096 13459 7098
rect 13275 7060 13321 7071
rect 13505 7096 13522 7098
rect 13459 7060 13505 7071
rect 12769 6843 12815 6988
rect 12984 6979 12995 7025
rect 13049 6979 13060 7025
rect 12984 6946 13060 6979
rect 13168 6979 13179 7025
rect 13233 6979 13244 7025
rect 13168 6946 13244 6979
rect 13352 6979 13363 7025
rect 13417 6979 13428 7025
rect 13352 6946 13428 6979
rect 13597 6843 13643 6988
rect 12757 6831 12837 6843
rect 12757 6775 12769 6831
rect 12825 6775 12837 6831
rect 12757 6763 12837 6775
rect 13575 6831 13655 6843
rect 13575 6775 13587 6831
rect 13643 6775 13655 6831
rect 13575 6763 13655 6775
rect 13928 6713 14008 6723
rect 12594 6657 13940 6713
rect 13996 6657 14008 6713
rect 13928 6655 14008 6657
rect 13762 6604 13832 6606
rect 12594 6603 13832 6604
rect 12594 6549 13764 6603
rect 13820 6549 13832 6603
rect 12594 6548 13832 6549
rect 10702 6496 10788 6500
rect 10702 6440 10714 6496
rect 10770 6440 10788 6496
rect 10702 6428 10788 6440
rect 10213 6283 10259 6294
rect 10428 6292 10504 6325
rect 10428 6246 10439 6292
rect 10493 6246 10504 6292
rect 10612 6292 10688 6325
rect 10612 6246 10623 6292
rect 10677 6246 10688 6292
rect 10796 6292 10872 6325
rect 10796 6246 10807 6292
rect 10861 6246 10872 6292
rect 11041 6283 11087 6294
rect 10351 6200 10397 6211
rect 10334 6173 10351 6175
rect 10535 6200 10581 6211
rect 10397 6173 10414 6175
rect 10259 6053 10346 6173
rect 10402 6053 10414 6173
rect 10334 6051 10351 6053
rect 10259 5753 10351 5873
rect 10397 6051 10414 6053
rect 10518 5873 10535 5875
rect 10719 6200 10765 6211
rect 10702 6173 10719 6175
rect 10903 6200 10949 6211
rect 10765 6173 10782 6175
rect 10702 6053 10714 6173
rect 10770 6053 10782 6173
rect 10702 6051 10719 6053
rect 10581 5873 10598 5875
rect 10518 5753 10530 5873
rect 10586 5753 10598 5873
rect 10518 5751 10535 5753
rect 10351 5715 10397 5726
rect 10581 5751 10598 5753
rect 10535 5715 10581 5726
rect 10765 6051 10782 6053
rect 10886 5873 10903 5875
rect 11024 6173 11041 6175
rect 11087 6173 11104 6175
rect 11024 6052 11036 6173
rect 11092 6052 11104 6173
rect 11024 6050 11041 6052
rect 10949 5873 10966 5875
rect 10886 5753 10898 5873
rect 10954 5753 10966 5873
rect 10886 5751 10903 5753
rect 10719 5715 10765 5726
rect 10949 5751 10966 5753
rect 10903 5715 10949 5726
rect 10428 5677 10439 5680
rect 10493 5677 10504 5680
rect 10612 5677 10623 5680
rect 10677 5677 10688 5680
rect 10796 5677 10807 5680
rect 10861 5677 10872 5680
rect 10213 5632 10259 5643
rect 10426 5621 10438 5677
rect 10494 5621 10506 5677
rect 10426 5607 10506 5621
rect 10610 5621 10622 5677
rect 10678 5621 10690 5677
rect 10610 5607 10690 5621
rect 10794 5621 10806 5677
rect 10862 5621 10874 5677
rect 11087 6050 11104 6052
rect 11041 5632 11087 5643
rect 10794 5607 10874 5621
rect 10426 5527 10506 5529
rect 10038 5471 10438 5527
rect 10494 5471 10506 5527
rect 12594 5527 12650 6548
rect 13762 6540 13832 6548
rect 13258 6496 13344 6500
rect 13258 6440 13270 6496
rect 13326 6440 13344 6496
rect 13258 6428 13344 6440
rect 12769 6283 12815 6294
rect 12984 6292 13060 6325
rect 12984 6246 12995 6292
rect 13049 6246 13060 6292
rect 13168 6292 13244 6325
rect 13168 6246 13179 6292
rect 13233 6246 13244 6292
rect 13352 6292 13428 6325
rect 13352 6246 13363 6292
rect 13417 6246 13428 6292
rect 13597 6283 13643 6294
rect 12907 6200 12953 6211
rect 12890 6173 12907 6175
rect 13091 6200 13137 6211
rect 12953 6173 12970 6175
rect 12815 6053 12902 6173
rect 12958 6053 12970 6173
rect 12890 6051 12907 6053
rect 12815 5753 12907 5873
rect 12953 6051 12970 6053
rect 13074 5873 13091 5875
rect 13275 6200 13321 6211
rect 13258 6173 13275 6175
rect 13459 6200 13505 6211
rect 13321 6173 13338 6175
rect 13258 6053 13270 6173
rect 13326 6053 13338 6173
rect 13258 6051 13275 6053
rect 13137 5873 13154 5875
rect 13074 5753 13086 5873
rect 13142 5753 13154 5873
rect 13074 5751 13091 5753
rect 12907 5715 12953 5726
rect 13137 5751 13154 5753
rect 13091 5715 13137 5726
rect 13321 6051 13338 6053
rect 13442 5873 13459 5875
rect 13580 6173 13597 6175
rect 13643 6173 13660 6175
rect 13580 6052 13592 6173
rect 13648 6052 13660 6173
rect 13580 6050 13597 6052
rect 13505 5873 13522 5875
rect 13442 5753 13454 5873
rect 13510 5753 13522 5873
rect 13442 5751 13459 5753
rect 13275 5715 13321 5726
rect 13505 5751 13522 5753
rect 13459 5715 13505 5726
rect 12984 5677 12995 5680
rect 13049 5677 13060 5680
rect 13168 5677 13179 5680
rect 13233 5677 13244 5680
rect 13352 5677 13363 5680
rect 13417 5677 13428 5680
rect 12769 5632 12815 5643
rect 12982 5621 12994 5677
rect 13050 5621 13062 5677
rect 12982 5607 13062 5621
rect 13166 5621 13178 5677
rect 13234 5621 13246 5677
rect 13166 5607 13246 5621
rect 13350 5621 13362 5677
rect 13418 5621 13430 5677
rect 13643 6050 13660 6052
rect 13597 5632 13643 5643
rect 13350 5607 13430 5621
rect 12982 5527 13062 5529
rect 12594 5471 12994 5527
rect 13050 5471 13062 5527
rect 14080 5527 14136 8753
rect 16631 8753 18178 8809
rect 16136 7732 16222 7744
rect 16631 7732 16687 8753
rect 17300 8701 17386 8705
rect 17300 8645 17312 8701
rect 17368 8645 17386 8701
rect 17300 8633 17386 8645
rect 16811 8488 16857 8499
rect 17026 8497 17102 8530
rect 17026 8451 17037 8497
rect 17091 8451 17102 8497
rect 17210 8497 17286 8530
rect 17210 8451 17221 8497
rect 17275 8451 17286 8497
rect 17394 8497 17470 8530
rect 17394 8451 17405 8497
rect 17459 8451 17470 8497
rect 17639 8488 17685 8499
rect 16949 8405 16995 8416
rect 16932 8378 16949 8380
rect 17133 8405 17179 8416
rect 16995 8378 17012 8380
rect 16857 8258 16944 8378
rect 17000 8258 17012 8378
rect 16932 8256 16949 8258
rect 16857 7958 16949 8078
rect 16995 8256 17012 8258
rect 17116 8078 17133 8080
rect 17317 8405 17363 8416
rect 17300 8378 17317 8380
rect 17501 8405 17547 8416
rect 17363 8378 17380 8380
rect 17300 8258 17312 8378
rect 17368 8258 17380 8378
rect 17300 8256 17317 8258
rect 17179 8078 17196 8080
rect 17116 7958 17128 8078
rect 17184 7958 17196 8078
rect 17116 7956 17133 7958
rect 16949 7920 16995 7931
rect 17179 7956 17196 7958
rect 17133 7920 17179 7931
rect 17363 8256 17380 8258
rect 17484 8078 17501 8080
rect 17622 8378 17639 8380
rect 17685 8378 17702 8380
rect 17622 8257 17634 8378
rect 17690 8257 17702 8378
rect 17622 8255 17639 8257
rect 17547 8078 17564 8080
rect 17484 7958 17496 8078
rect 17552 7958 17564 8078
rect 17484 7956 17501 7958
rect 17317 7920 17363 7931
rect 17547 7956 17564 7958
rect 17501 7920 17547 7931
rect 17026 7882 17037 7885
rect 17091 7882 17102 7885
rect 17210 7882 17221 7885
rect 17275 7882 17286 7885
rect 17394 7882 17405 7885
rect 17459 7882 17470 7885
rect 16811 7837 16857 7848
rect 17024 7826 17036 7882
rect 17092 7826 17104 7882
rect 17024 7812 17104 7826
rect 17208 7826 17220 7882
rect 17276 7826 17288 7882
rect 17208 7812 17288 7826
rect 17392 7826 17404 7882
rect 17460 7826 17472 7882
rect 17685 8255 17702 8257
rect 17639 7837 17685 7848
rect 17392 7812 17472 7826
rect 17024 7732 17104 7734
rect 16136 7676 16148 7732
rect 16204 7676 17036 7732
rect 17092 7676 17104 7732
rect 16136 7664 16222 7676
rect 17024 7674 17104 7676
rect 16352 7616 16422 7628
rect 17208 7616 17288 7618
rect 16352 7560 16364 7616
rect 16420 7560 17220 7616
rect 17276 7560 17288 7616
rect 16352 7548 16422 7560
rect 17208 7558 17288 7560
rect 17537 7616 17617 7618
rect 17804 7616 17874 7628
rect 17537 7560 17549 7616
rect 17605 7560 17806 7616
rect 17862 7560 17874 7616
rect 17537 7558 17617 7560
rect 17804 7550 17874 7560
rect 17392 7500 17472 7502
rect 16636 7444 17404 7500
rect 17460 7444 17472 7500
rect 16636 6713 16692 7444
rect 17392 7442 17472 7444
rect 17024 7350 17104 7364
rect 16811 7328 16857 7339
rect 17024 7294 17036 7350
rect 17092 7294 17104 7350
rect 17208 7350 17288 7364
rect 17208 7294 17220 7350
rect 17276 7294 17288 7350
rect 17392 7350 17472 7364
rect 17392 7294 17404 7350
rect 17460 7294 17472 7350
rect 17639 7328 17685 7339
rect 17026 7291 17037 7294
rect 17091 7291 17102 7294
rect 17210 7291 17221 7294
rect 17275 7291 17286 7294
rect 17394 7291 17405 7294
rect 17459 7291 17470 7294
rect 16949 7245 16995 7256
rect 16857 7071 16949 7245
rect 16949 7060 16995 7071
rect 17133 7245 17179 7256
rect 17133 7060 17179 7071
rect 17317 7245 17363 7256
rect 17501 7245 17547 7256
rect 17484 7218 17501 7220
rect 17547 7218 17564 7220
rect 17484 7098 17496 7218
rect 17552 7098 17564 7218
rect 17484 7096 17501 7098
rect 17317 7060 17363 7071
rect 17547 7096 17564 7098
rect 17501 7060 17547 7071
rect 16811 6843 16857 6988
rect 17026 6979 17037 7025
rect 17091 6979 17102 7025
rect 17026 6946 17102 6979
rect 17210 6979 17221 7025
rect 17275 6979 17286 7025
rect 17210 6946 17286 6979
rect 17394 6979 17405 7025
rect 17459 6979 17470 7025
rect 17394 6946 17470 6979
rect 17639 6843 17685 6988
rect 16799 6831 16879 6843
rect 16799 6775 16811 6831
rect 16867 6775 16879 6831
rect 16799 6763 16879 6775
rect 17617 6831 17697 6843
rect 17617 6775 17629 6831
rect 17685 6775 17697 6831
rect 17617 6763 17697 6775
rect 17970 6713 18050 6723
rect 16636 6657 17982 6713
rect 18038 6657 18050 6713
rect 17970 6655 18050 6657
rect 17804 6604 17874 6606
rect 16636 6603 17874 6604
rect 16636 6549 17806 6603
rect 17862 6549 17874 6603
rect 16636 6548 17874 6549
rect 14744 6496 14830 6500
rect 14744 6440 14756 6496
rect 14812 6440 14830 6496
rect 14744 6428 14830 6440
rect 14255 6283 14301 6294
rect 14470 6292 14546 6325
rect 14470 6246 14481 6292
rect 14535 6246 14546 6292
rect 14654 6292 14730 6325
rect 14654 6246 14665 6292
rect 14719 6246 14730 6292
rect 14838 6292 14914 6325
rect 14838 6246 14849 6292
rect 14903 6246 14914 6292
rect 15083 6283 15129 6294
rect 14393 6200 14439 6211
rect 14376 6173 14393 6175
rect 14577 6200 14623 6211
rect 14439 6173 14456 6175
rect 14301 6053 14388 6173
rect 14444 6053 14456 6173
rect 14376 6051 14393 6053
rect 14301 5753 14393 5873
rect 14439 6051 14456 6053
rect 14560 5873 14577 5875
rect 14761 6200 14807 6211
rect 14744 6173 14761 6175
rect 14945 6200 14991 6211
rect 14807 6173 14824 6175
rect 14744 6053 14756 6173
rect 14812 6053 14824 6173
rect 14744 6051 14761 6053
rect 14623 5873 14640 5875
rect 14560 5753 14572 5873
rect 14628 5753 14640 5873
rect 14560 5751 14577 5753
rect 14393 5715 14439 5726
rect 14623 5751 14640 5753
rect 14577 5715 14623 5726
rect 14807 6051 14824 6053
rect 14928 5873 14945 5875
rect 15066 6173 15083 6175
rect 15129 6173 15146 6175
rect 15066 6052 15078 6173
rect 15134 6052 15146 6173
rect 15066 6050 15083 6052
rect 14991 5873 15008 5875
rect 14928 5753 14940 5873
rect 14996 5753 15008 5873
rect 14928 5751 14945 5753
rect 14761 5715 14807 5726
rect 14991 5751 15008 5753
rect 14945 5715 14991 5726
rect 14470 5677 14481 5680
rect 14535 5677 14546 5680
rect 14654 5677 14665 5680
rect 14719 5677 14730 5680
rect 14838 5677 14849 5680
rect 14903 5677 14914 5680
rect 14255 5632 14301 5643
rect 14468 5621 14480 5677
rect 14536 5621 14548 5677
rect 14468 5607 14548 5621
rect 14652 5621 14664 5677
rect 14720 5621 14732 5677
rect 14652 5607 14732 5621
rect 14836 5621 14848 5677
rect 14904 5621 14916 5677
rect 15129 6050 15146 6052
rect 15083 5632 15129 5643
rect 14836 5607 14916 5621
rect 14468 5527 14548 5529
rect 14080 5471 14480 5527
rect 14536 5471 14548 5527
rect 16636 5527 16692 6548
rect 17804 6540 17874 6548
rect 17300 6496 17386 6500
rect 17300 6440 17312 6496
rect 17368 6440 17386 6496
rect 17300 6428 17386 6440
rect 16811 6283 16857 6294
rect 17026 6292 17102 6325
rect 17026 6246 17037 6292
rect 17091 6246 17102 6292
rect 17210 6292 17286 6325
rect 17210 6246 17221 6292
rect 17275 6246 17286 6292
rect 17394 6292 17470 6325
rect 17394 6246 17405 6292
rect 17459 6246 17470 6292
rect 17639 6283 17685 6294
rect 16949 6200 16995 6211
rect 16932 6173 16949 6175
rect 17133 6200 17179 6211
rect 16995 6173 17012 6175
rect 16857 6053 16944 6173
rect 17000 6053 17012 6173
rect 16932 6051 16949 6053
rect 16857 5753 16949 5873
rect 16995 6051 17012 6053
rect 17116 5873 17133 5875
rect 17317 6200 17363 6211
rect 17300 6173 17317 6175
rect 17501 6200 17547 6211
rect 17363 6173 17380 6175
rect 17300 6053 17312 6173
rect 17368 6053 17380 6173
rect 17300 6051 17317 6053
rect 17179 5873 17196 5875
rect 17116 5753 17128 5873
rect 17184 5753 17196 5873
rect 17116 5751 17133 5753
rect 16949 5715 16995 5726
rect 17179 5751 17196 5753
rect 17133 5715 17179 5726
rect 17363 6051 17380 6053
rect 17484 5873 17501 5875
rect 17622 6173 17639 6175
rect 17685 6173 17702 6175
rect 17622 6052 17634 6173
rect 17690 6052 17702 6173
rect 17622 6050 17639 6052
rect 17547 5873 17564 5875
rect 17484 5753 17496 5873
rect 17552 5753 17564 5873
rect 17484 5751 17501 5753
rect 17317 5715 17363 5726
rect 17547 5751 17564 5753
rect 17501 5715 17547 5726
rect 17026 5677 17037 5680
rect 17091 5677 17102 5680
rect 17210 5677 17221 5680
rect 17275 5677 17286 5680
rect 17394 5677 17405 5680
rect 17459 5677 17470 5680
rect 16811 5632 16857 5643
rect 17024 5621 17036 5677
rect 17092 5621 17104 5677
rect 17024 5607 17104 5621
rect 17208 5621 17220 5677
rect 17276 5621 17288 5677
rect 17208 5607 17288 5621
rect 17392 5621 17404 5677
rect 17460 5621 17472 5677
rect 17685 6050 17702 6052
rect 17639 5632 17685 5643
rect 17392 5607 17472 5621
rect 17024 5527 17104 5529
rect 16636 5471 17036 5527
rect 17092 5471 17104 5527
rect 18122 5527 18178 8753
rect 20673 8753 22220 8809
rect 20178 7732 20264 7744
rect 20673 7732 20729 8753
rect 21342 8701 21428 8705
rect 21342 8645 21354 8701
rect 21410 8645 21428 8701
rect 21342 8633 21428 8645
rect 20853 8488 20899 8499
rect 21068 8497 21144 8530
rect 21068 8451 21079 8497
rect 21133 8451 21144 8497
rect 21252 8497 21328 8530
rect 21252 8451 21263 8497
rect 21317 8451 21328 8497
rect 21436 8497 21512 8530
rect 21436 8451 21447 8497
rect 21501 8451 21512 8497
rect 21681 8488 21727 8499
rect 20991 8405 21037 8416
rect 20974 8378 20991 8380
rect 21175 8405 21221 8416
rect 21037 8378 21054 8380
rect 20899 8258 20986 8378
rect 21042 8258 21054 8378
rect 20974 8256 20991 8258
rect 20899 7958 20991 8078
rect 21037 8256 21054 8258
rect 21158 8078 21175 8080
rect 21359 8405 21405 8416
rect 21342 8378 21359 8380
rect 21543 8405 21589 8416
rect 21405 8378 21422 8380
rect 21342 8258 21354 8378
rect 21410 8258 21422 8378
rect 21342 8256 21359 8258
rect 21221 8078 21238 8080
rect 21158 7958 21170 8078
rect 21226 7958 21238 8078
rect 21158 7956 21175 7958
rect 20991 7920 21037 7931
rect 21221 7956 21238 7958
rect 21175 7920 21221 7931
rect 21405 8256 21422 8258
rect 21526 8078 21543 8080
rect 21664 8378 21681 8380
rect 21727 8378 21744 8380
rect 21664 8257 21676 8378
rect 21732 8257 21744 8378
rect 21664 8255 21681 8257
rect 21589 8078 21606 8080
rect 21526 7958 21538 8078
rect 21594 7958 21606 8078
rect 21526 7956 21543 7958
rect 21359 7920 21405 7931
rect 21589 7956 21606 7958
rect 21543 7920 21589 7931
rect 21068 7882 21079 7885
rect 21133 7882 21144 7885
rect 21252 7882 21263 7885
rect 21317 7882 21328 7885
rect 21436 7882 21447 7885
rect 21501 7882 21512 7885
rect 20853 7837 20899 7848
rect 21066 7826 21078 7882
rect 21134 7826 21146 7882
rect 21066 7812 21146 7826
rect 21250 7826 21262 7882
rect 21318 7826 21330 7882
rect 21250 7812 21330 7826
rect 21434 7826 21446 7882
rect 21502 7826 21514 7882
rect 21727 8255 21744 8257
rect 21681 7837 21727 7848
rect 21434 7812 21514 7826
rect 21066 7732 21146 7734
rect 20178 7676 20190 7732
rect 20246 7676 21078 7732
rect 21134 7676 21146 7732
rect 20178 7664 20264 7676
rect 21066 7674 21146 7676
rect 20394 7616 20464 7628
rect 21250 7616 21330 7618
rect 20394 7560 20406 7616
rect 20462 7560 21262 7616
rect 21318 7560 21330 7616
rect 20394 7548 20464 7560
rect 21250 7558 21330 7560
rect 21579 7616 21659 7618
rect 21846 7616 21916 7628
rect 21579 7560 21591 7616
rect 21647 7560 21848 7616
rect 21904 7560 21916 7616
rect 21579 7558 21659 7560
rect 21846 7550 21916 7560
rect 21434 7500 21514 7502
rect 20678 7444 21446 7500
rect 21502 7444 21514 7500
rect 20678 6713 20734 7444
rect 21434 7442 21514 7444
rect 21066 7350 21146 7364
rect 20853 7328 20899 7339
rect 21066 7294 21078 7350
rect 21134 7294 21146 7350
rect 21250 7350 21330 7364
rect 21250 7294 21262 7350
rect 21318 7294 21330 7350
rect 21434 7350 21514 7364
rect 21434 7294 21446 7350
rect 21502 7294 21514 7350
rect 21681 7328 21727 7339
rect 21068 7291 21079 7294
rect 21133 7291 21144 7294
rect 21252 7291 21263 7294
rect 21317 7291 21328 7294
rect 21436 7291 21447 7294
rect 21501 7291 21512 7294
rect 20991 7245 21037 7256
rect 20899 7071 20991 7245
rect 20991 7060 21037 7071
rect 21175 7245 21221 7256
rect 21175 7060 21221 7071
rect 21359 7245 21405 7256
rect 21543 7245 21589 7256
rect 21526 7218 21543 7220
rect 21589 7218 21606 7220
rect 21526 7098 21538 7218
rect 21594 7098 21606 7218
rect 21526 7096 21543 7098
rect 21359 7060 21405 7071
rect 21589 7096 21606 7098
rect 21543 7060 21589 7071
rect 20853 6843 20899 6988
rect 21068 6979 21079 7025
rect 21133 6979 21144 7025
rect 21068 6946 21144 6979
rect 21252 6979 21263 7025
rect 21317 6979 21328 7025
rect 21252 6946 21328 6979
rect 21436 6979 21447 7025
rect 21501 6979 21512 7025
rect 21436 6946 21512 6979
rect 21681 6843 21727 6988
rect 20841 6831 20921 6843
rect 20841 6775 20853 6831
rect 20909 6775 20921 6831
rect 20841 6763 20921 6775
rect 21659 6831 21739 6843
rect 21659 6775 21671 6831
rect 21727 6775 21739 6831
rect 21659 6763 21739 6775
rect 22012 6713 22092 6723
rect 20678 6657 22024 6713
rect 22080 6657 22092 6713
rect 22012 6655 22092 6657
rect 21846 6604 21916 6606
rect 20678 6603 21916 6604
rect 20678 6549 21848 6603
rect 21904 6549 21916 6603
rect 20678 6548 21916 6549
rect 18786 6496 18872 6500
rect 18786 6440 18798 6496
rect 18854 6440 18872 6496
rect 18786 6428 18872 6440
rect 18297 6283 18343 6294
rect 18512 6292 18588 6325
rect 18512 6246 18523 6292
rect 18577 6246 18588 6292
rect 18696 6292 18772 6325
rect 18696 6246 18707 6292
rect 18761 6246 18772 6292
rect 18880 6292 18956 6325
rect 18880 6246 18891 6292
rect 18945 6246 18956 6292
rect 19125 6283 19171 6294
rect 18435 6200 18481 6211
rect 18418 6173 18435 6175
rect 18619 6200 18665 6211
rect 18481 6173 18498 6175
rect 18343 6053 18430 6173
rect 18486 6053 18498 6173
rect 18418 6051 18435 6053
rect 18343 5753 18435 5873
rect 18481 6051 18498 6053
rect 18602 5873 18619 5875
rect 18803 6200 18849 6211
rect 18786 6173 18803 6175
rect 18987 6200 19033 6211
rect 18849 6173 18866 6175
rect 18786 6053 18798 6173
rect 18854 6053 18866 6173
rect 18786 6051 18803 6053
rect 18665 5873 18682 5875
rect 18602 5753 18614 5873
rect 18670 5753 18682 5873
rect 18602 5751 18619 5753
rect 18435 5715 18481 5726
rect 18665 5751 18682 5753
rect 18619 5715 18665 5726
rect 18849 6051 18866 6053
rect 18970 5873 18987 5875
rect 19108 6173 19125 6175
rect 19171 6173 19188 6175
rect 19108 6052 19120 6173
rect 19176 6052 19188 6173
rect 19108 6050 19125 6052
rect 19033 5873 19050 5875
rect 18970 5753 18982 5873
rect 19038 5753 19050 5873
rect 18970 5751 18987 5753
rect 18803 5715 18849 5726
rect 19033 5751 19050 5753
rect 18987 5715 19033 5726
rect 18512 5677 18523 5680
rect 18577 5677 18588 5680
rect 18696 5677 18707 5680
rect 18761 5677 18772 5680
rect 18880 5677 18891 5680
rect 18945 5677 18956 5680
rect 18297 5632 18343 5643
rect 18510 5621 18522 5677
rect 18578 5621 18590 5677
rect 18510 5607 18590 5621
rect 18694 5621 18706 5677
rect 18762 5621 18774 5677
rect 18694 5607 18774 5621
rect 18878 5621 18890 5677
rect 18946 5621 18958 5677
rect 19171 6050 19188 6052
rect 19125 5632 19171 5643
rect 18878 5607 18958 5621
rect 18510 5527 18590 5529
rect 18122 5471 18522 5527
rect 18578 5471 18590 5527
rect 20678 5527 20734 6548
rect 21846 6540 21916 6548
rect 21342 6496 21428 6500
rect 21342 6440 21354 6496
rect 21410 6440 21428 6496
rect 21342 6428 21428 6440
rect 20853 6283 20899 6294
rect 21068 6292 21144 6325
rect 21068 6246 21079 6292
rect 21133 6246 21144 6292
rect 21252 6292 21328 6325
rect 21252 6246 21263 6292
rect 21317 6246 21328 6292
rect 21436 6292 21512 6325
rect 21436 6246 21447 6292
rect 21501 6246 21512 6292
rect 21681 6283 21727 6294
rect 20991 6200 21037 6211
rect 20974 6173 20991 6175
rect 21175 6200 21221 6211
rect 21037 6173 21054 6175
rect 20899 6053 20986 6173
rect 21042 6053 21054 6173
rect 20974 6051 20991 6053
rect 20899 5753 20991 5873
rect 21037 6051 21054 6053
rect 21158 5873 21175 5875
rect 21359 6200 21405 6211
rect 21342 6173 21359 6175
rect 21543 6200 21589 6211
rect 21405 6173 21422 6175
rect 21342 6053 21354 6173
rect 21410 6053 21422 6173
rect 21342 6051 21359 6053
rect 21221 5873 21238 5875
rect 21158 5753 21170 5873
rect 21226 5753 21238 5873
rect 21158 5751 21175 5753
rect 20991 5715 21037 5726
rect 21221 5751 21238 5753
rect 21175 5715 21221 5726
rect 21405 6051 21422 6053
rect 21526 5873 21543 5875
rect 21664 6173 21681 6175
rect 21727 6173 21744 6175
rect 21664 6052 21676 6173
rect 21732 6052 21744 6173
rect 21664 6050 21681 6052
rect 21589 5873 21606 5875
rect 21526 5753 21538 5873
rect 21594 5753 21606 5873
rect 21526 5751 21543 5753
rect 21359 5715 21405 5726
rect 21589 5751 21606 5753
rect 21543 5715 21589 5726
rect 21068 5677 21079 5680
rect 21133 5677 21144 5680
rect 21252 5677 21263 5680
rect 21317 5677 21328 5680
rect 21436 5677 21447 5680
rect 21501 5677 21512 5680
rect 20853 5632 20899 5643
rect 21066 5621 21078 5677
rect 21134 5621 21146 5677
rect 21066 5607 21146 5621
rect 21250 5621 21262 5677
rect 21318 5621 21330 5677
rect 21250 5607 21330 5621
rect 21434 5621 21446 5677
rect 21502 5621 21514 5677
rect 21727 6050 21744 6052
rect 21681 5632 21727 5643
rect 21434 5607 21514 5621
rect 21066 5527 21146 5529
rect 20678 5471 21078 5527
rect 21134 5471 21146 5527
rect 22164 5527 22220 8753
rect 24715 8753 26262 8809
rect 24220 7732 24306 7744
rect 24715 7732 24771 8753
rect 25384 8701 25470 8705
rect 25384 8645 25396 8701
rect 25452 8645 25470 8701
rect 25384 8633 25470 8645
rect 24895 8488 24941 8499
rect 25110 8497 25186 8530
rect 25110 8451 25121 8497
rect 25175 8451 25186 8497
rect 25294 8497 25370 8530
rect 25294 8451 25305 8497
rect 25359 8451 25370 8497
rect 25478 8497 25554 8530
rect 25478 8451 25489 8497
rect 25543 8451 25554 8497
rect 25723 8488 25769 8499
rect 25033 8405 25079 8416
rect 25016 8378 25033 8380
rect 25217 8405 25263 8416
rect 25079 8378 25096 8380
rect 24941 8258 25028 8378
rect 25084 8258 25096 8378
rect 25016 8256 25033 8258
rect 24941 7958 25033 8078
rect 25079 8256 25096 8258
rect 25200 8078 25217 8080
rect 25401 8405 25447 8416
rect 25384 8378 25401 8380
rect 25585 8405 25631 8416
rect 25447 8378 25464 8380
rect 25384 8258 25396 8378
rect 25452 8258 25464 8378
rect 25384 8256 25401 8258
rect 25263 8078 25280 8080
rect 25200 7958 25212 8078
rect 25268 7958 25280 8078
rect 25200 7956 25217 7958
rect 25033 7920 25079 7931
rect 25263 7956 25280 7958
rect 25217 7920 25263 7931
rect 25447 8256 25464 8258
rect 25568 8078 25585 8080
rect 25706 8378 25723 8380
rect 25769 8378 25786 8380
rect 25706 8257 25718 8378
rect 25774 8257 25786 8378
rect 25706 8255 25723 8257
rect 25631 8078 25648 8080
rect 25568 7958 25580 8078
rect 25636 7958 25648 8078
rect 25568 7956 25585 7958
rect 25401 7920 25447 7931
rect 25631 7956 25648 7958
rect 25585 7920 25631 7931
rect 25110 7882 25121 7885
rect 25175 7882 25186 7885
rect 25294 7882 25305 7885
rect 25359 7882 25370 7885
rect 25478 7882 25489 7885
rect 25543 7882 25554 7885
rect 24895 7837 24941 7848
rect 25108 7826 25120 7882
rect 25176 7826 25188 7882
rect 25108 7812 25188 7826
rect 25292 7826 25304 7882
rect 25360 7826 25372 7882
rect 25292 7812 25372 7826
rect 25476 7826 25488 7882
rect 25544 7826 25556 7882
rect 25769 8255 25786 8257
rect 25723 7837 25769 7848
rect 25476 7812 25556 7826
rect 25108 7732 25188 7734
rect 24220 7676 24232 7732
rect 24288 7676 25120 7732
rect 25176 7676 25188 7732
rect 24220 7664 24306 7676
rect 25108 7674 25188 7676
rect 24436 7616 24506 7628
rect 25292 7616 25372 7618
rect 24436 7560 24448 7616
rect 24504 7560 25304 7616
rect 25360 7560 25372 7616
rect 24436 7548 24506 7560
rect 25292 7558 25372 7560
rect 25621 7616 25701 7618
rect 25888 7616 25958 7628
rect 25621 7560 25633 7616
rect 25689 7560 25890 7616
rect 25946 7560 25958 7616
rect 25621 7558 25701 7560
rect 25888 7550 25958 7560
rect 25476 7500 25556 7502
rect 24720 7444 25488 7500
rect 25544 7444 25556 7500
rect 24720 6713 24776 7444
rect 25476 7442 25556 7444
rect 25108 7350 25188 7364
rect 24895 7328 24941 7339
rect 25108 7294 25120 7350
rect 25176 7294 25188 7350
rect 25292 7350 25372 7364
rect 25292 7294 25304 7350
rect 25360 7294 25372 7350
rect 25476 7350 25556 7364
rect 25476 7294 25488 7350
rect 25544 7294 25556 7350
rect 25723 7328 25769 7339
rect 25110 7291 25121 7294
rect 25175 7291 25186 7294
rect 25294 7291 25305 7294
rect 25359 7291 25370 7294
rect 25478 7291 25489 7294
rect 25543 7291 25554 7294
rect 25033 7245 25079 7256
rect 24941 7071 25033 7245
rect 25033 7060 25079 7071
rect 25217 7245 25263 7256
rect 25217 7060 25263 7071
rect 25401 7245 25447 7256
rect 25585 7245 25631 7256
rect 25568 7218 25585 7220
rect 25631 7218 25648 7220
rect 25568 7098 25580 7218
rect 25636 7098 25648 7218
rect 25568 7096 25585 7098
rect 25401 7060 25447 7071
rect 25631 7096 25648 7098
rect 25585 7060 25631 7071
rect 24895 6843 24941 6988
rect 25110 6979 25121 7025
rect 25175 6979 25186 7025
rect 25110 6946 25186 6979
rect 25294 6979 25305 7025
rect 25359 6979 25370 7025
rect 25294 6946 25370 6979
rect 25478 6979 25489 7025
rect 25543 6979 25554 7025
rect 25478 6946 25554 6979
rect 25723 6843 25769 6988
rect 24883 6831 24963 6843
rect 24883 6775 24895 6831
rect 24951 6775 24963 6831
rect 24883 6763 24963 6775
rect 25701 6831 25781 6843
rect 25701 6775 25713 6831
rect 25769 6775 25781 6831
rect 25701 6763 25781 6775
rect 26054 6713 26134 6723
rect 24720 6657 26066 6713
rect 26122 6657 26134 6713
rect 26054 6655 26134 6657
rect 25888 6604 25958 6606
rect 24720 6603 25958 6604
rect 24720 6549 25890 6603
rect 25946 6549 25958 6603
rect 24720 6548 25958 6549
rect 22828 6496 22914 6500
rect 22828 6440 22840 6496
rect 22896 6440 22914 6496
rect 22828 6428 22914 6440
rect 22339 6283 22385 6294
rect 22554 6292 22630 6325
rect 22554 6246 22565 6292
rect 22619 6246 22630 6292
rect 22738 6292 22814 6325
rect 22738 6246 22749 6292
rect 22803 6246 22814 6292
rect 22922 6292 22998 6325
rect 22922 6246 22933 6292
rect 22987 6246 22998 6292
rect 23167 6283 23213 6294
rect 22477 6200 22523 6211
rect 22460 6173 22477 6175
rect 22661 6200 22707 6211
rect 22523 6173 22540 6175
rect 22385 6053 22472 6173
rect 22528 6053 22540 6173
rect 22460 6051 22477 6053
rect 22385 5753 22477 5873
rect 22523 6051 22540 6053
rect 22644 5873 22661 5875
rect 22845 6200 22891 6211
rect 22828 6173 22845 6175
rect 23029 6200 23075 6211
rect 22891 6173 22908 6175
rect 22828 6053 22840 6173
rect 22896 6053 22908 6173
rect 22828 6051 22845 6053
rect 22707 5873 22724 5875
rect 22644 5753 22656 5873
rect 22712 5753 22724 5873
rect 22644 5751 22661 5753
rect 22477 5715 22523 5726
rect 22707 5751 22724 5753
rect 22661 5715 22707 5726
rect 22891 6051 22908 6053
rect 23012 5873 23029 5875
rect 23150 6173 23167 6175
rect 23213 6173 23230 6175
rect 23150 6052 23162 6173
rect 23218 6052 23230 6173
rect 23150 6050 23167 6052
rect 23075 5873 23092 5875
rect 23012 5753 23024 5873
rect 23080 5753 23092 5873
rect 23012 5751 23029 5753
rect 22845 5715 22891 5726
rect 23075 5751 23092 5753
rect 23029 5715 23075 5726
rect 22554 5677 22565 5680
rect 22619 5677 22630 5680
rect 22738 5677 22749 5680
rect 22803 5677 22814 5680
rect 22922 5677 22933 5680
rect 22987 5677 22998 5680
rect 22339 5632 22385 5643
rect 22552 5621 22564 5677
rect 22620 5621 22632 5677
rect 22552 5607 22632 5621
rect 22736 5621 22748 5677
rect 22804 5621 22816 5677
rect 22736 5607 22816 5621
rect 22920 5621 22932 5677
rect 22988 5621 23000 5677
rect 23213 6050 23230 6052
rect 23167 5632 23213 5643
rect 22920 5607 23000 5621
rect 22552 5527 22632 5529
rect 22164 5471 22564 5527
rect 22620 5471 22632 5527
rect 24720 5527 24776 6548
rect 25888 6540 25958 6548
rect 25384 6496 25470 6500
rect 25384 6440 25396 6496
rect 25452 6440 25470 6496
rect 25384 6428 25470 6440
rect 24895 6283 24941 6294
rect 25110 6292 25186 6325
rect 25110 6246 25121 6292
rect 25175 6246 25186 6292
rect 25294 6292 25370 6325
rect 25294 6246 25305 6292
rect 25359 6246 25370 6292
rect 25478 6292 25554 6325
rect 25478 6246 25489 6292
rect 25543 6246 25554 6292
rect 25723 6283 25769 6294
rect 25033 6200 25079 6211
rect 25016 6173 25033 6175
rect 25217 6200 25263 6211
rect 25079 6173 25096 6175
rect 24941 6053 25028 6173
rect 25084 6053 25096 6173
rect 25016 6051 25033 6053
rect 24941 5753 25033 5873
rect 25079 6051 25096 6053
rect 25200 5873 25217 5875
rect 25401 6200 25447 6211
rect 25384 6173 25401 6175
rect 25585 6200 25631 6211
rect 25447 6173 25464 6175
rect 25384 6053 25396 6173
rect 25452 6053 25464 6173
rect 25384 6051 25401 6053
rect 25263 5873 25280 5875
rect 25200 5753 25212 5873
rect 25268 5753 25280 5873
rect 25200 5751 25217 5753
rect 25033 5715 25079 5726
rect 25263 5751 25280 5753
rect 25217 5715 25263 5726
rect 25447 6051 25464 6053
rect 25568 5873 25585 5875
rect 25706 6173 25723 6175
rect 25769 6173 25786 6175
rect 25706 6052 25718 6173
rect 25774 6052 25786 6173
rect 25706 6050 25723 6052
rect 25631 5873 25648 5875
rect 25568 5753 25580 5873
rect 25636 5753 25648 5873
rect 25568 5751 25585 5753
rect 25401 5715 25447 5726
rect 25631 5751 25648 5753
rect 25585 5715 25631 5726
rect 25110 5677 25121 5680
rect 25175 5677 25186 5680
rect 25294 5677 25305 5680
rect 25359 5677 25370 5680
rect 25478 5677 25489 5680
rect 25543 5677 25554 5680
rect 24895 5632 24941 5643
rect 25108 5621 25120 5677
rect 25176 5621 25188 5677
rect 25108 5607 25188 5621
rect 25292 5621 25304 5677
rect 25360 5621 25372 5677
rect 25292 5607 25372 5621
rect 25476 5621 25488 5677
rect 25544 5621 25556 5677
rect 25769 6050 25786 6052
rect 25723 5632 25769 5643
rect 25476 5607 25556 5621
rect 25108 5527 25188 5529
rect 24720 5471 25120 5527
rect 25176 5471 25188 5527
rect 26206 5527 26262 8753
rect 26870 6496 26956 6500
rect 26870 6440 26882 6496
rect 26938 6440 26956 6496
rect 26870 6428 26956 6440
rect 26381 6283 26427 6294
rect 26596 6292 26672 6325
rect 26596 6246 26607 6292
rect 26661 6246 26672 6292
rect 26780 6292 26856 6325
rect 26780 6246 26791 6292
rect 26845 6246 26856 6292
rect 26964 6292 27040 6325
rect 26964 6246 26975 6292
rect 27029 6246 27040 6292
rect 27209 6283 27255 6294
rect 26519 6200 26565 6211
rect 26502 6173 26519 6175
rect 26703 6200 26749 6211
rect 26565 6173 26582 6175
rect 26427 6053 26514 6173
rect 26570 6053 26582 6173
rect 26502 6051 26519 6053
rect 26427 5753 26519 5873
rect 26565 6051 26582 6053
rect 26686 5873 26703 5875
rect 26887 6200 26933 6211
rect 26870 6173 26887 6175
rect 27071 6200 27117 6211
rect 26933 6173 26950 6175
rect 26870 6053 26882 6173
rect 26938 6053 26950 6173
rect 26870 6051 26887 6053
rect 26749 5873 26766 5875
rect 26686 5753 26698 5873
rect 26754 5753 26766 5873
rect 26686 5751 26703 5753
rect 26519 5715 26565 5726
rect 26749 5751 26766 5753
rect 26703 5715 26749 5726
rect 26933 6051 26950 6053
rect 27054 5873 27071 5875
rect 27192 6173 27209 6175
rect 27255 6173 27272 6175
rect 27192 6052 27204 6173
rect 27260 6052 27272 6173
rect 27192 6050 27209 6052
rect 27117 5873 27134 5875
rect 27054 5753 27066 5873
rect 27122 5753 27134 5873
rect 27054 5751 27071 5753
rect 26887 5715 26933 5726
rect 27117 5751 27134 5753
rect 27071 5715 27117 5726
rect 26596 5677 26607 5680
rect 26661 5677 26672 5680
rect 26780 5677 26791 5680
rect 26845 5677 26856 5680
rect 26964 5677 26975 5680
rect 27029 5677 27040 5680
rect 26381 5632 26427 5643
rect 26594 5621 26606 5677
rect 26662 5621 26674 5677
rect 26594 5607 26674 5621
rect 26778 5621 26790 5677
rect 26846 5621 26858 5677
rect 26778 5607 26858 5621
rect 26962 5621 26974 5677
rect 27030 5621 27042 5677
rect 27255 6050 27272 6052
rect 27209 5632 27255 5643
rect 26962 5607 27042 5621
rect 26594 5527 26674 5529
rect 26206 5471 26606 5527
rect 26662 5471 26674 5527
rect 886 5469 966 5471
rect 2372 5469 2452 5471
rect 4898 5469 4978 5471
rect 6384 5469 6464 5471
rect 8940 5469 9020 5471
rect 10426 5469 10506 5471
rect 12982 5469 13062 5471
rect 14468 5469 14548 5471
rect 17024 5469 17104 5471
rect 18510 5469 18590 5471
rect 21066 5469 21146 5471
rect 22552 5469 22632 5471
rect 25108 5469 25188 5471
rect 26594 5469 26674 5471
rect 78 5411 148 5425
rect 1070 5411 1150 5413
rect 78 5355 90 5411
rect 146 5355 1082 5411
rect 1138 5355 1150 5411
rect 78 5343 148 5355
rect 1070 5353 1150 5355
rect 1399 5411 1479 5413
rect 1842 5411 1902 5421
rect 2556 5411 2636 5413
rect 1399 5355 1411 5411
rect 1467 5355 1844 5411
rect 1900 5355 2568 5411
rect 2624 5355 2636 5411
rect 1399 5353 1479 5355
rect 1842 5343 1902 5355
rect 2556 5353 2636 5355
rect 2885 5411 2965 5413
rect 3152 5411 3222 5423
rect 4090 5411 4160 5425
rect 5082 5411 5162 5413
rect 2885 5355 2897 5411
rect 2953 5355 3154 5411
rect 3210 5355 4022 5411
rect 2885 5353 2965 5355
rect 3152 5345 3222 5355
rect 1254 5295 1334 5297
rect 2740 5295 2820 5297
rect 362 5239 1266 5295
rect 1322 5239 1334 5295
rect -330 4509 -260 4521
rect 362 4509 418 5239
rect 1254 5237 1334 5239
rect 1984 5239 2752 5295
rect 2808 5239 2820 5295
rect 886 5145 966 5159
rect 673 5123 719 5134
rect 886 5089 898 5145
rect 954 5089 966 5145
rect 1070 5145 1150 5159
rect 1070 5089 1082 5145
rect 1138 5089 1150 5145
rect 1254 5145 1334 5159
rect 1254 5089 1266 5145
rect 1322 5089 1334 5145
rect 1501 5123 1547 5134
rect 888 5086 899 5089
rect 953 5086 964 5089
rect 1072 5086 1083 5089
rect 1137 5086 1148 5089
rect 1256 5086 1267 5089
rect 1321 5086 1332 5089
rect 811 5040 857 5051
rect 719 4866 811 5040
rect 811 4855 857 4866
rect 995 5040 1041 5051
rect 995 4855 1041 4866
rect 1179 5040 1225 5051
rect 1363 5040 1409 5051
rect 1346 5013 1363 5015
rect 1409 5013 1426 5015
rect 1346 4893 1358 5013
rect 1414 4893 1426 5013
rect 1346 4891 1363 4893
rect 1179 4855 1225 4866
rect 1409 4891 1426 4893
rect 1363 4855 1409 4866
rect 673 4638 719 4783
rect 888 4774 899 4820
rect 953 4774 964 4820
rect 888 4741 964 4774
rect 1072 4774 1083 4820
rect 1137 4774 1148 4820
rect 1072 4741 1148 4774
rect 1256 4774 1267 4820
rect 1321 4774 1332 4820
rect 1256 4741 1332 4774
rect 1501 4638 1547 4783
rect 661 4626 741 4638
rect 661 4570 673 4626
rect 729 4570 741 4626
rect 661 4558 741 4570
rect 1479 4626 1557 4638
rect 1479 4570 1491 4626
rect 1547 4570 1557 4626
rect 1479 4558 1557 4570
rect -330 4453 -318 4509
rect -262 4453 418 4509
rect 1984 4509 2040 5239
rect 2740 5237 2820 5239
rect 3966 5233 4022 5355
rect 4090 5355 4102 5411
rect 4158 5355 5094 5411
rect 5150 5355 5162 5411
rect 4090 5343 4160 5355
rect 5082 5353 5162 5355
rect 5411 5411 5491 5413
rect 5854 5411 5914 5421
rect 6568 5411 6648 5413
rect 5411 5355 5423 5411
rect 5479 5355 5856 5411
rect 5912 5355 6580 5411
rect 6636 5355 6648 5411
rect 5411 5353 5491 5355
rect 5854 5343 5914 5355
rect 6568 5353 6648 5355
rect 6897 5411 6977 5413
rect 7164 5411 7234 5423
rect 8132 5411 8202 5425
rect 9124 5411 9204 5413
rect 6897 5355 6909 5411
rect 6965 5355 7166 5411
rect 7222 5355 8034 5411
rect 6897 5353 6977 5355
rect 7164 5345 7234 5355
rect 5266 5295 5346 5297
rect 6752 5295 6832 5297
rect 4374 5239 5278 5295
rect 5334 5239 5346 5295
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 2372 5145 2452 5159
rect 2159 5123 2205 5134
rect 2372 5089 2384 5145
rect 2440 5089 2452 5145
rect 2556 5145 2636 5159
rect 2556 5089 2568 5145
rect 2624 5089 2636 5145
rect 2740 5145 2820 5159
rect 2740 5089 2752 5145
rect 2808 5089 2820 5145
rect 2987 5123 3033 5134
rect 2374 5086 2385 5089
rect 2439 5086 2450 5089
rect 2558 5086 2569 5089
rect 2623 5086 2634 5089
rect 2742 5086 2753 5089
rect 2807 5086 2818 5089
rect 2297 5040 2343 5051
rect 2205 4866 2297 5040
rect 2297 4855 2343 4866
rect 2481 5040 2527 5051
rect 2481 4855 2527 4866
rect 2665 5040 2711 5051
rect 2849 5040 2895 5051
rect 2832 5013 2849 5015
rect 2895 5013 2912 5015
rect 2832 4893 2844 5013
rect 2900 4893 2912 5013
rect 2832 4891 2849 4893
rect 2665 4855 2711 4866
rect 2895 4891 2912 4893
rect 2849 4855 2895 4866
rect 2159 4638 2205 4783
rect 2374 4774 2385 4820
rect 2439 4774 2450 4820
rect 2374 4741 2450 4774
rect 2558 4774 2569 4820
rect 2623 4774 2634 4820
rect 2558 4741 2634 4774
rect 2742 4774 2753 4820
rect 2807 4774 2818 4820
rect 2742 4741 2818 4774
rect 2987 4638 3033 4783
rect 2147 4626 2227 4638
rect 2147 4570 2159 4626
rect 2215 4570 2227 4626
rect 2147 4558 2227 4570
rect 2965 4626 3043 4638
rect 2965 4570 2977 4626
rect 3033 4570 3043 4626
rect 2965 4558 3043 4570
rect 3318 4509 3398 4519
rect 1984 4453 3330 4509
rect 3386 4453 3398 4509
rect -330 4441 -260 4453
rect 362 3206 418 4453
rect 3318 4451 3398 4453
rect 3682 4509 3752 4521
rect 4374 4509 4430 5239
rect 5266 5237 5346 5239
rect 5996 5239 6764 5295
rect 6820 5239 6832 5295
rect 4898 5145 4978 5159
rect 4685 5123 4731 5134
rect 4898 5089 4910 5145
rect 4966 5089 4978 5145
rect 5082 5145 5162 5159
rect 5082 5089 5094 5145
rect 5150 5089 5162 5145
rect 5266 5145 5346 5159
rect 5266 5089 5278 5145
rect 5334 5089 5346 5145
rect 5513 5123 5559 5134
rect 4900 5086 4911 5089
rect 4965 5086 4976 5089
rect 5084 5086 5095 5089
rect 5149 5086 5160 5089
rect 5268 5086 5279 5089
rect 5333 5086 5344 5089
rect 4823 5040 4869 5051
rect 4731 4866 4823 5040
rect 4823 4855 4869 4866
rect 5007 5040 5053 5051
rect 5007 4855 5053 4866
rect 5191 5040 5237 5051
rect 5375 5040 5421 5051
rect 5358 5013 5375 5015
rect 5421 5013 5438 5015
rect 5358 4893 5370 5013
rect 5426 4893 5438 5013
rect 5358 4891 5375 4893
rect 5191 4855 5237 4866
rect 5421 4891 5438 4893
rect 5375 4855 5421 4866
rect 4685 4638 4731 4783
rect 4900 4774 4911 4820
rect 4965 4774 4976 4820
rect 4900 4741 4976 4774
rect 5084 4774 5095 4820
rect 5149 4774 5160 4820
rect 5084 4741 5160 4774
rect 5268 4774 5279 4820
rect 5333 4774 5344 4820
rect 5268 4741 5344 4774
rect 5513 4638 5559 4783
rect 4673 4626 4753 4638
rect 4673 4570 4685 4626
rect 4741 4570 4753 4626
rect 4673 4558 4753 4570
rect 5491 4626 5569 4638
rect 5491 4570 5503 4626
rect 5559 4570 5569 4626
rect 5491 4558 5569 4570
rect 3682 4453 3694 4509
rect 3750 4453 4430 4509
rect 5996 4509 6052 5239
rect 6752 5237 6832 5239
rect 7978 5233 8034 5355
rect 8132 5355 8144 5411
rect 8200 5355 9136 5411
rect 9192 5355 9204 5411
rect 8132 5343 8202 5355
rect 9124 5353 9204 5355
rect 9453 5411 9533 5413
rect 9896 5411 9956 5421
rect 10610 5411 10690 5413
rect 9453 5355 9465 5411
rect 9521 5355 9898 5411
rect 9954 5355 10622 5411
rect 10678 5355 10690 5411
rect 9453 5353 9533 5355
rect 9896 5343 9956 5355
rect 10610 5353 10690 5355
rect 10939 5411 11019 5413
rect 11206 5411 11276 5423
rect 12174 5411 12244 5425
rect 13166 5411 13246 5413
rect 10939 5355 10951 5411
rect 11007 5355 11208 5411
rect 11264 5355 12076 5411
rect 10939 5353 11019 5355
rect 11206 5345 11276 5355
rect 9308 5295 9388 5297
rect 10794 5295 10874 5297
rect 8416 5239 9320 5295
rect 9376 5239 9388 5295
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 6384 5145 6464 5159
rect 6171 5123 6217 5134
rect 6384 5089 6396 5145
rect 6452 5089 6464 5145
rect 6568 5145 6648 5159
rect 6568 5089 6580 5145
rect 6636 5089 6648 5145
rect 6752 5145 6832 5159
rect 6752 5089 6764 5145
rect 6820 5089 6832 5145
rect 6999 5123 7045 5134
rect 6386 5086 6397 5089
rect 6451 5086 6462 5089
rect 6570 5086 6581 5089
rect 6635 5086 6646 5089
rect 6754 5086 6765 5089
rect 6819 5086 6830 5089
rect 6309 5040 6355 5051
rect 6217 4866 6309 5040
rect 6309 4855 6355 4866
rect 6493 5040 6539 5051
rect 6493 4855 6539 4866
rect 6677 5040 6723 5051
rect 6861 5040 6907 5051
rect 6844 5013 6861 5015
rect 6907 5013 6924 5015
rect 6844 4893 6856 5013
rect 6912 4893 6924 5013
rect 6844 4891 6861 4893
rect 6677 4855 6723 4866
rect 6907 4891 6924 4893
rect 6861 4855 6907 4866
rect 6171 4638 6217 4783
rect 6386 4774 6397 4820
rect 6451 4774 6462 4820
rect 6386 4741 6462 4774
rect 6570 4774 6581 4820
rect 6635 4774 6646 4820
rect 6570 4741 6646 4774
rect 6754 4774 6765 4820
rect 6819 4774 6830 4820
rect 6754 4741 6830 4774
rect 6999 4638 7045 4783
rect 6159 4626 6239 4638
rect 6159 4570 6171 4626
rect 6227 4570 6239 4626
rect 6159 4558 6239 4570
rect 6977 4626 7055 4638
rect 6977 4570 6989 4626
rect 7045 4570 7055 4626
rect 6977 4558 7055 4570
rect 7330 4509 7410 4519
rect 5996 4453 7342 4509
rect 7398 4453 7410 4509
rect 3682 4441 3752 4453
rect 1842 4398 1912 4400
rect 3142 4399 3222 4401
rect 498 4342 1844 4398
rect 1900 4342 1912 4398
rect 498 3322 554 4342
rect 1842 4330 1912 4342
rect 1984 4343 3154 4399
rect 3210 4343 3222 4399
rect 1162 4291 1248 4295
rect 1162 4235 1174 4291
rect 1230 4235 1248 4291
rect 1162 4223 1248 4235
rect 673 4078 719 4089
rect 888 4087 964 4120
rect 888 4041 899 4087
rect 953 4041 964 4087
rect 1072 4087 1148 4120
rect 1072 4041 1083 4087
rect 1137 4041 1148 4087
rect 1256 4087 1332 4120
rect 1256 4041 1267 4087
rect 1321 4041 1332 4087
rect 1501 4078 1547 4089
rect 811 3995 857 4006
rect 794 3968 811 3970
rect 995 3995 1041 4006
rect 857 3968 874 3970
rect 719 3848 806 3968
rect 862 3848 874 3968
rect 794 3846 811 3848
rect 719 3548 811 3668
rect 857 3846 874 3848
rect 978 3668 995 3670
rect 1179 3995 1225 4006
rect 1162 3968 1179 3970
rect 1363 3995 1409 4006
rect 1225 3968 1242 3970
rect 1162 3848 1174 3968
rect 1230 3848 1242 3968
rect 1162 3846 1179 3848
rect 1041 3668 1058 3670
rect 978 3548 990 3668
rect 1046 3548 1058 3668
rect 978 3546 995 3548
rect 811 3510 857 3521
rect 1041 3546 1058 3548
rect 995 3510 1041 3521
rect 1225 3846 1242 3848
rect 1346 3668 1363 3670
rect 1484 3968 1501 3970
rect 1547 3968 1564 3970
rect 1484 3847 1496 3968
rect 1552 3847 1564 3968
rect 1484 3845 1501 3847
rect 1409 3668 1426 3670
rect 1346 3548 1358 3668
rect 1414 3548 1426 3668
rect 1346 3546 1363 3548
rect 1179 3510 1225 3521
rect 1409 3546 1426 3548
rect 1363 3510 1409 3521
rect 888 3472 899 3475
rect 953 3472 964 3475
rect 1072 3472 1083 3475
rect 1137 3472 1148 3475
rect 1256 3472 1267 3475
rect 1321 3472 1332 3475
rect 673 3427 719 3438
rect 886 3416 898 3472
rect 954 3416 966 3472
rect 886 3402 966 3416
rect 1070 3416 1082 3472
rect 1138 3416 1150 3472
rect 1070 3402 1150 3416
rect 1254 3416 1266 3472
rect 1322 3416 1334 3472
rect 1547 3845 1564 3847
rect 1501 3427 1547 3438
rect 1254 3402 1334 3416
rect 886 3322 966 3324
rect 498 3266 898 3322
rect 954 3266 966 3322
rect 1984 3323 2040 4343
rect 3142 4331 3222 4343
rect 2648 4292 2734 4296
rect 2648 4236 2660 4292
rect 2716 4236 2734 4292
rect 2648 4224 2734 4236
rect 2159 4079 2205 4090
rect 2374 4088 2450 4121
rect 2374 4042 2385 4088
rect 2439 4042 2450 4088
rect 2558 4088 2634 4121
rect 2558 4042 2569 4088
rect 2623 4042 2634 4088
rect 2742 4088 2818 4121
rect 2742 4042 2753 4088
rect 2807 4042 2818 4088
rect 2987 4079 3033 4090
rect 2297 3996 2343 4007
rect 2280 3969 2297 3971
rect 2481 3996 2527 4007
rect 2343 3969 2360 3971
rect 2205 3849 2292 3969
rect 2348 3849 2360 3969
rect 2280 3847 2297 3849
rect 2205 3549 2297 3669
rect 2343 3847 2360 3849
rect 2464 3669 2481 3671
rect 2665 3996 2711 4007
rect 2648 3969 2665 3971
rect 2849 3996 2895 4007
rect 2711 3969 2728 3971
rect 2648 3849 2660 3969
rect 2716 3849 2728 3969
rect 2648 3847 2665 3849
rect 2527 3669 2544 3671
rect 2464 3549 2476 3669
rect 2532 3549 2544 3669
rect 2464 3547 2481 3549
rect 2297 3511 2343 3522
rect 2527 3547 2544 3549
rect 2481 3511 2527 3522
rect 2711 3847 2728 3849
rect 2832 3669 2849 3671
rect 2970 3969 2987 3971
rect 3033 3969 3050 3971
rect 2970 3848 2982 3969
rect 3038 3848 3050 3969
rect 2970 3846 2987 3848
rect 2895 3669 2912 3671
rect 2832 3549 2844 3669
rect 2900 3549 2912 3669
rect 2832 3547 2849 3549
rect 2665 3511 2711 3522
rect 2895 3547 2912 3549
rect 2849 3511 2895 3522
rect 2374 3473 2385 3476
rect 2439 3473 2450 3476
rect 2558 3473 2569 3476
rect 2623 3473 2634 3476
rect 2742 3473 2753 3476
rect 2807 3473 2818 3476
rect 2159 3428 2205 3439
rect 2372 3417 2384 3473
rect 2440 3417 2452 3473
rect 2372 3403 2452 3417
rect 2556 3417 2568 3473
rect 2624 3417 2636 3473
rect 2556 3403 2636 3417
rect 2740 3417 2752 3473
rect 2808 3417 2820 3473
rect 3033 3846 3050 3848
rect 2987 3428 3033 3439
rect 2740 3403 2820 3417
rect 2372 3323 2452 3325
rect 1984 3267 2384 3323
rect 2440 3267 2452 3323
rect 886 3264 966 3266
rect 2372 3265 2452 3267
rect 1070 3206 1150 3208
rect 362 3150 1082 3206
rect 1138 3150 1150 3206
rect 1070 3148 1150 3150
rect 1399 3206 1479 3208
rect 1666 3207 1736 3218
rect 2556 3207 2636 3209
rect 1666 3206 2568 3207
rect 1399 3150 1411 3206
rect 1467 3150 1668 3206
rect 1724 3151 2568 3206
rect 2624 3151 2636 3207
rect 1724 3150 1984 3151
rect 1399 3148 1479 3150
rect 1666 3140 1736 3150
rect 2556 3149 2636 3151
rect 2885 3207 2965 3209
rect 3328 3207 3398 3217
rect 2885 3151 2897 3207
rect 2953 3151 3330 3207
rect 3386 3151 3398 3207
rect 2885 3149 2965 3151
rect 3328 3139 3398 3151
rect 4374 3206 4430 4453
rect 7330 4451 7410 4453
rect 7694 4509 7764 4521
rect 8416 4509 8472 5239
rect 9308 5237 9388 5239
rect 10038 5239 10806 5295
rect 10862 5239 10874 5295
rect 8940 5145 9020 5159
rect 8727 5123 8773 5134
rect 8940 5089 8952 5145
rect 9008 5089 9020 5145
rect 9124 5145 9204 5159
rect 9124 5089 9136 5145
rect 9192 5089 9204 5145
rect 9308 5145 9388 5159
rect 9308 5089 9320 5145
rect 9376 5089 9388 5145
rect 9555 5123 9601 5134
rect 8942 5086 8953 5089
rect 9007 5086 9018 5089
rect 9126 5086 9137 5089
rect 9191 5086 9202 5089
rect 9310 5086 9321 5089
rect 9375 5086 9386 5089
rect 8865 5040 8911 5051
rect 8773 4866 8865 5040
rect 8865 4855 8911 4866
rect 9049 5040 9095 5051
rect 9049 4855 9095 4866
rect 9233 5040 9279 5051
rect 9417 5040 9463 5051
rect 9400 5013 9417 5015
rect 9463 5013 9480 5015
rect 9400 4893 9412 5013
rect 9468 4893 9480 5013
rect 9400 4891 9417 4893
rect 9233 4855 9279 4866
rect 9463 4891 9480 4893
rect 9417 4855 9463 4866
rect 8727 4638 8773 4783
rect 8942 4774 8953 4820
rect 9007 4774 9018 4820
rect 8942 4741 9018 4774
rect 9126 4774 9137 4820
rect 9191 4774 9202 4820
rect 9126 4741 9202 4774
rect 9310 4774 9321 4820
rect 9375 4774 9386 4820
rect 9310 4741 9386 4774
rect 9555 4638 9601 4783
rect 8715 4626 8795 4638
rect 8715 4570 8727 4626
rect 8783 4570 8795 4626
rect 8715 4558 8795 4570
rect 9533 4626 9611 4638
rect 9533 4570 9545 4626
rect 9601 4570 9611 4626
rect 9533 4558 9611 4570
rect 7694 4453 7706 4509
rect 7762 4453 8472 4509
rect 10038 4509 10094 5239
rect 10794 5237 10874 5239
rect 12020 5233 12076 5355
rect 12174 5355 12186 5411
rect 12242 5355 13178 5411
rect 13234 5355 13246 5411
rect 12174 5343 12244 5355
rect 13166 5353 13246 5355
rect 13495 5411 13575 5413
rect 13938 5411 13998 5421
rect 14652 5411 14732 5413
rect 13495 5355 13507 5411
rect 13563 5355 13940 5411
rect 13996 5355 14664 5411
rect 14720 5355 14732 5411
rect 13495 5353 13575 5355
rect 13938 5343 13998 5355
rect 14652 5353 14732 5355
rect 14981 5411 15061 5413
rect 15248 5411 15318 5423
rect 16216 5411 16286 5425
rect 17208 5411 17288 5413
rect 14981 5355 14993 5411
rect 15049 5355 15250 5411
rect 15306 5355 16118 5411
rect 14981 5353 15061 5355
rect 15248 5345 15318 5355
rect 13350 5295 13430 5297
rect 14836 5295 14916 5297
rect 12458 5239 13362 5295
rect 13418 5239 13430 5295
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 10426 5145 10506 5159
rect 10213 5123 10259 5134
rect 10426 5089 10438 5145
rect 10494 5089 10506 5145
rect 10610 5145 10690 5159
rect 10610 5089 10622 5145
rect 10678 5089 10690 5145
rect 10794 5145 10874 5159
rect 10794 5089 10806 5145
rect 10862 5089 10874 5145
rect 11041 5123 11087 5134
rect 10428 5086 10439 5089
rect 10493 5086 10504 5089
rect 10612 5086 10623 5089
rect 10677 5086 10688 5089
rect 10796 5086 10807 5089
rect 10861 5086 10872 5089
rect 10351 5040 10397 5051
rect 10259 4866 10351 5040
rect 10351 4855 10397 4866
rect 10535 5040 10581 5051
rect 10535 4855 10581 4866
rect 10719 5040 10765 5051
rect 10903 5040 10949 5051
rect 10886 5013 10903 5015
rect 10949 5013 10966 5015
rect 10886 4893 10898 5013
rect 10954 4893 10966 5013
rect 10886 4891 10903 4893
rect 10719 4855 10765 4866
rect 10949 4891 10966 4893
rect 10903 4855 10949 4866
rect 10213 4638 10259 4783
rect 10428 4774 10439 4820
rect 10493 4774 10504 4820
rect 10428 4741 10504 4774
rect 10612 4774 10623 4820
rect 10677 4774 10688 4820
rect 10612 4741 10688 4774
rect 10796 4774 10807 4820
rect 10861 4774 10872 4820
rect 10796 4741 10872 4774
rect 11041 4638 11087 4783
rect 10201 4626 10281 4638
rect 10201 4570 10213 4626
rect 10269 4570 10281 4626
rect 10201 4558 10281 4570
rect 11019 4626 11097 4638
rect 11019 4570 11031 4626
rect 11087 4570 11097 4626
rect 11019 4558 11097 4570
rect 11372 4509 11452 4519
rect 10038 4453 11384 4509
rect 11440 4453 11452 4509
rect 7694 4441 7764 4453
rect 5854 4398 5924 4400
rect 7154 4399 7234 4401
rect 4510 4342 5856 4398
rect 5912 4342 5924 4398
rect 4510 3322 4566 4342
rect 5854 4330 5924 4342
rect 5996 4343 7166 4399
rect 7222 4343 7234 4399
rect 5174 4291 5260 4295
rect 5174 4235 5186 4291
rect 5242 4235 5260 4291
rect 5174 4223 5260 4235
rect 4685 4078 4731 4089
rect 4900 4087 4976 4120
rect 4900 4041 4911 4087
rect 4965 4041 4976 4087
rect 5084 4087 5160 4120
rect 5084 4041 5095 4087
rect 5149 4041 5160 4087
rect 5268 4087 5344 4120
rect 5268 4041 5279 4087
rect 5333 4041 5344 4087
rect 5513 4078 5559 4089
rect 4823 3995 4869 4006
rect 4806 3968 4823 3970
rect 5007 3995 5053 4006
rect 4869 3968 4886 3970
rect 4731 3848 4818 3968
rect 4874 3848 4886 3968
rect 4806 3846 4823 3848
rect 4731 3548 4823 3668
rect 4869 3846 4886 3848
rect 4990 3668 5007 3670
rect 5191 3995 5237 4006
rect 5174 3968 5191 3970
rect 5375 3995 5421 4006
rect 5237 3968 5254 3970
rect 5174 3848 5186 3968
rect 5242 3848 5254 3968
rect 5174 3846 5191 3848
rect 5053 3668 5070 3670
rect 4990 3548 5002 3668
rect 5058 3548 5070 3668
rect 4990 3546 5007 3548
rect 4823 3510 4869 3521
rect 5053 3546 5070 3548
rect 5007 3510 5053 3521
rect 5237 3846 5254 3848
rect 5358 3668 5375 3670
rect 5496 3968 5513 3970
rect 5559 3968 5576 3970
rect 5496 3847 5508 3968
rect 5564 3847 5576 3968
rect 5496 3845 5513 3847
rect 5421 3668 5438 3670
rect 5358 3548 5370 3668
rect 5426 3548 5438 3668
rect 5358 3546 5375 3548
rect 5191 3510 5237 3521
rect 5421 3546 5438 3548
rect 5375 3510 5421 3521
rect 4900 3472 4911 3475
rect 4965 3472 4976 3475
rect 5084 3472 5095 3475
rect 5149 3472 5160 3475
rect 5268 3472 5279 3475
rect 5333 3472 5344 3475
rect 4685 3427 4731 3438
rect 4898 3416 4910 3472
rect 4966 3416 4978 3472
rect 4898 3402 4978 3416
rect 5082 3416 5094 3472
rect 5150 3416 5162 3472
rect 5082 3402 5162 3416
rect 5266 3416 5278 3472
rect 5334 3416 5346 3472
rect 5559 3845 5576 3847
rect 5513 3427 5559 3438
rect 5266 3402 5346 3416
rect 4898 3322 4978 3324
rect 4510 3266 4910 3322
rect 4966 3266 4978 3322
rect 5996 3323 6052 4343
rect 7154 4331 7234 4343
rect 6660 4292 6746 4296
rect 6660 4236 6672 4292
rect 6728 4236 6746 4292
rect 6660 4224 6746 4236
rect 6171 4079 6217 4090
rect 6386 4088 6462 4121
rect 6386 4042 6397 4088
rect 6451 4042 6462 4088
rect 6570 4088 6646 4121
rect 6570 4042 6581 4088
rect 6635 4042 6646 4088
rect 6754 4088 6830 4121
rect 6754 4042 6765 4088
rect 6819 4042 6830 4088
rect 6999 4079 7045 4090
rect 6309 3996 6355 4007
rect 6292 3969 6309 3971
rect 6493 3996 6539 4007
rect 6355 3969 6372 3971
rect 6217 3849 6304 3969
rect 6360 3849 6372 3969
rect 6292 3847 6309 3849
rect 6217 3549 6309 3669
rect 6355 3847 6372 3849
rect 6476 3669 6493 3671
rect 6677 3996 6723 4007
rect 6660 3969 6677 3971
rect 6861 3996 6907 4007
rect 6723 3969 6740 3971
rect 6660 3849 6672 3969
rect 6728 3849 6740 3969
rect 6660 3847 6677 3849
rect 6539 3669 6556 3671
rect 6476 3549 6488 3669
rect 6544 3549 6556 3669
rect 6476 3547 6493 3549
rect 6309 3511 6355 3522
rect 6539 3547 6556 3549
rect 6493 3511 6539 3522
rect 6723 3847 6740 3849
rect 6844 3669 6861 3671
rect 6982 3969 6999 3971
rect 7045 3969 7062 3971
rect 6982 3848 6994 3969
rect 7050 3848 7062 3969
rect 6982 3846 6999 3848
rect 6907 3669 6924 3671
rect 6844 3549 6856 3669
rect 6912 3549 6924 3669
rect 6844 3547 6861 3549
rect 6677 3511 6723 3522
rect 6907 3547 6924 3549
rect 6861 3511 6907 3522
rect 6386 3473 6397 3476
rect 6451 3473 6462 3476
rect 6570 3473 6581 3476
rect 6635 3473 6646 3476
rect 6754 3473 6765 3476
rect 6819 3473 6830 3476
rect 6171 3428 6217 3439
rect 6384 3417 6396 3473
rect 6452 3417 6464 3473
rect 6384 3403 6464 3417
rect 6568 3417 6580 3473
rect 6636 3417 6648 3473
rect 6568 3403 6648 3417
rect 6752 3417 6764 3473
rect 6820 3417 6832 3473
rect 7045 3846 7062 3848
rect 6999 3428 7045 3439
rect 6752 3403 6832 3417
rect 6384 3323 6464 3325
rect 5996 3267 6396 3323
rect 6452 3267 6464 3323
rect 4898 3264 4978 3266
rect 6384 3265 6464 3267
rect 5082 3206 5162 3208
rect 4374 3150 5094 3206
rect 5150 3150 5162 3206
rect 5082 3148 5162 3150
rect 5411 3206 5491 3208
rect 5678 3207 5748 3218
rect 6568 3207 6648 3209
rect 5678 3206 6580 3207
rect 5411 3150 5423 3206
rect 5479 3150 5680 3206
rect 5736 3151 6580 3206
rect 6636 3151 6648 3207
rect 5736 3150 5996 3151
rect 5411 3148 5491 3150
rect 5678 3140 5748 3150
rect 6568 3149 6648 3151
rect 6897 3207 6977 3209
rect 7340 3207 7410 3217
rect 6897 3151 6909 3207
rect 6965 3151 7342 3207
rect 7398 3151 7410 3207
rect 6897 3149 6977 3151
rect 7340 3139 7410 3151
rect 8416 3206 8472 4453
rect 11372 4451 11452 4453
rect 11736 4509 11806 4521
rect 12458 4509 12514 5239
rect 13350 5237 13430 5239
rect 14080 5239 14848 5295
rect 14904 5239 14916 5295
rect 12982 5145 13062 5159
rect 12769 5123 12815 5134
rect 12982 5089 12994 5145
rect 13050 5089 13062 5145
rect 13166 5145 13246 5159
rect 13166 5089 13178 5145
rect 13234 5089 13246 5145
rect 13350 5145 13430 5159
rect 13350 5089 13362 5145
rect 13418 5089 13430 5145
rect 13597 5123 13643 5134
rect 12984 5086 12995 5089
rect 13049 5086 13060 5089
rect 13168 5086 13179 5089
rect 13233 5086 13244 5089
rect 13352 5086 13363 5089
rect 13417 5086 13428 5089
rect 12907 5040 12953 5051
rect 12815 4866 12907 5040
rect 12907 4855 12953 4866
rect 13091 5040 13137 5051
rect 13091 4855 13137 4866
rect 13275 5040 13321 5051
rect 13459 5040 13505 5051
rect 13442 5013 13459 5015
rect 13505 5013 13522 5015
rect 13442 4893 13454 5013
rect 13510 4893 13522 5013
rect 13442 4891 13459 4893
rect 13275 4855 13321 4866
rect 13505 4891 13522 4893
rect 13459 4855 13505 4866
rect 12769 4638 12815 4783
rect 12984 4774 12995 4820
rect 13049 4774 13060 4820
rect 12984 4741 13060 4774
rect 13168 4774 13179 4820
rect 13233 4774 13244 4820
rect 13168 4741 13244 4774
rect 13352 4774 13363 4820
rect 13417 4774 13428 4820
rect 13352 4741 13428 4774
rect 13597 4638 13643 4783
rect 12757 4626 12837 4638
rect 12757 4570 12769 4626
rect 12825 4570 12837 4626
rect 12757 4558 12837 4570
rect 13575 4626 13653 4638
rect 13575 4570 13587 4626
rect 13643 4570 13653 4626
rect 13575 4558 13653 4570
rect 11736 4453 11748 4509
rect 11804 4453 12514 4509
rect 14080 4509 14136 5239
rect 14836 5237 14916 5239
rect 16062 5233 16118 5355
rect 16216 5355 16228 5411
rect 16284 5355 17220 5411
rect 17276 5355 17288 5411
rect 16216 5343 16286 5355
rect 17208 5353 17288 5355
rect 17537 5411 17617 5413
rect 17980 5411 18040 5421
rect 18694 5411 18774 5413
rect 17537 5355 17549 5411
rect 17605 5355 17982 5411
rect 18038 5355 18706 5411
rect 18762 5355 18774 5411
rect 17537 5353 17617 5355
rect 17980 5343 18040 5355
rect 18694 5353 18774 5355
rect 19023 5411 19103 5413
rect 19290 5411 19360 5423
rect 20258 5411 20328 5425
rect 21250 5411 21330 5413
rect 19023 5355 19035 5411
rect 19091 5355 19292 5411
rect 19348 5355 20160 5411
rect 19023 5353 19103 5355
rect 19290 5345 19360 5355
rect 17392 5295 17472 5297
rect 18878 5295 18958 5297
rect 16500 5239 17404 5295
rect 17460 5239 17472 5295
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 14468 5145 14548 5159
rect 14255 5123 14301 5134
rect 14468 5089 14480 5145
rect 14536 5089 14548 5145
rect 14652 5145 14732 5159
rect 14652 5089 14664 5145
rect 14720 5089 14732 5145
rect 14836 5145 14916 5159
rect 14836 5089 14848 5145
rect 14904 5089 14916 5145
rect 15083 5123 15129 5134
rect 14470 5086 14481 5089
rect 14535 5086 14546 5089
rect 14654 5086 14665 5089
rect 14719 5086 14730 5089
rect 14838 5086 14849 5089
rect 14903 5086 14914 5089
rect 14393 5040 14439 5051
rect 14301 4866 14393 5040
rect 14393 4855 14439 4866
rect 14577 5040 14623 5051
rect 14577 4855 14623 4866
rect 14761 5040 14807 5051
rect 14945 5040 14991 5051
rect 14928 5013 14945 5015
rect 14991 5013 15008 5015
rect 14928 4893 14940 5013
rect 14996 4893 15008 5013
rect 14928 4891 14945 4893
rect 14761 4855 14807 4866
rect 14991 4891 15008 4893
rect 14945 4855 14991 4866
rect 14255 4638 14301 4783
rect 14470 4774 14481 4820
rect 14535 4774 14546 4820
rect 14470 4741 14546 4774
rect 14654 4774 14665 4820
rect 14719 4774 14730 4820
rect 14654 4741 14730 4774
rect 14838 4774 14849 4820
rect 14903 4774 14914 4820
rect 14838 4741 14914 4774
rect 15083 4638 15129 4783
rect 14243 4626 14323 4638
rect 14243 4570 14255 4626
rect 14311 4570 14323 4626
rect 14243 4558 14323 4570
rect 15061 4626 15139 4638
rect 15061 4570 15073 4626
rect 15129 4570 15139 4626
rect 15061 4558 15139 4570
rect 15414 4509 15494 4519
rect 14080 4453 15426 4509
rect 15482 4453 15494 4509
rect 11736 4441 11806 4453
rect 9896 4398 9966 4400
rect 11196 4399 11276 4401
rect 8552 4342 9898 4398
rect 9954 4342 9966 4398
rect 8552 3322 8608 4342
rect 9896 4330 9966 4342
rect 10038 4343 11208 4399
rect 11264 4343 11276 4399
rect 9216 4291 9302 4295
rect 9216 4235 9228 4291
rect 9284 4235 9302 4291
rect 9216 4223 9302 4235
rect 8727 4078 8773 4089
rect 8942 4087 9018 4120
rect 8942 4041 8953 4087
rect 9007 4041 9018 4087
rect 9126 4087 9202 4120
rect 9126 4041 9137 4087
rect 9191 4041 9202 4087
rect 9310 4087 9386 4120
rect 9310 4041 9321 4087
rect 9375 4041 9386 4087
rect 9555 4078 9601 4089
rect 8865 3995 8911 4006
rect 8848 3968 8865 3970
rect 9049 3995 9095 4006
rect 8911 3968 8928 3970
rect 8773 3848 8860 3968
rect 8916 3848 8928 3968
rect 8848 3846 8865 3848
rect 8773 3548 8865 3668
rect 8911 3846 8928 3848
rect 9032 3668 9049 3670
rect 9233 3995 9279 4006
rect 9216 3968 9233 3970
rect 9417 3995 9463 4006
rect 9279 3968 9296 3970
rect 9216 3848 9228 3968
rect 9284 3848 9296 3968
rect 9216 3846 9233 3848
rect 9095 3668 9112 3670
rect 9032 3548 9044 3668
rect 9100 3548 9112 3668
rect 9032 3546 9049 3548
rect 8865 3510 8911 3521
rect 9095 3546 9112 3548
rect 9049 3510 9095 3521
rect 9279 3846 9296 3848
rect 9400 3668 9417 3670
rect 9538 3968 9555 3970
rect 9601 3968 9618 3970
rect 9538 3847 9550 3968
rect 9606 3847 9618 3968
rect 9538 3845 9555 3847
rect 9463 3668 9480 3670
rect 9400 3548 9412 3668
rect 9468 3548 9480 3668
rect 9400 3546 9417 3548
rect 9233 3510 9279 3521
rect 9463 3546 9480 3548
rect 9417 3510 9463 3521
rect 8942 3472 8953 3475
rect 9007 3472 9018 3475
rect 9126 3472 9137 3475
rect 9191 3472 9202 3475
rect 9310 3472 9321 3475
rect 9375 3472 9386 3475
rect 8727 3427 8773 3438
rect 8940 3416 8952 3472
rect 9008 3416 9020 3472
rect 8940 3402 9020 3416
rect 9124 3416 9136 3472
rect 9192 3416 9204 3472
rect 9124 3402 9204 3416
rect 9308 3416 9320 3472
rect 9376 3416 9388 3472
rect 9601 3845 9618 3847
rect 9555 3427 9601 3438
rect 9308 3402 9388 3416
rect 8940 3322 9020 3324
rect 8552 3266 8952 3322
rect 9008 3266 9020 3322
rect 10038 3323 10094 4343
rect 11196 4331 11276 4343
rect 10702 4292 10788 4296
rect 10702 4236 10714 4292
rect 10770 4236 10788 4292
rect 10702 4224 10788 4236
rect 10213 4079 10259 4090
rect 10428 4088 10504 4121
rect 10428 4042 10439 4088
rect 10493 4042 10504 4088
rect 10612 4088 10688 4121
rect 10612 4042 10623 4088
rect 10677 4042 10688 4088
rect 10796 4088 10872 4121
rect 10796 4042 10807 4088
rect 10861 4042 10872 4088
rect 11041 4079 11087 4090
rect 10351 3996 10397 4007
rect 10334 3969 10351 3971
rect 10535 3996 10581 4007
rect 10397 3969 10414 3971
rect 10259 3849 10346 3969
rect 10402 3849 10414 3969
rect 10334 3847 10351 3849
rect 10259 3549 10351 3669
rect 10397 3847 10414 3849
rect 10518 3669 10535 3671
rect 10719 3996 10765 4007
rect 10702 3969 10719 3971
rect 10903 3996 10949 4007
rect 10765 3969 10782 3971
rect 10702 3849 10714 3969
rect 10770 3849 10782 3969
rect 10702 3847 10719 3849
rect 10581 3669 10598 3671
rect 10518 3549 10530 3669
rect 10586 3549 10598 3669
rect 10518 3547 10535 3549
rect 10351 3511 10397 3522
rect 10581 3547 10598 3549
rect 10535 3511 10581 3522
rect 10765 3847 10782 3849
rect 10886 3669 10903 3671
rect 11024 3969 11041 3971
rect 11087 3969 11104 3971
rect 11024 3848 11036 3969
rect 11092 3848 11104 3969
rect 11024 3846 11041 3848
rect 10949 3669 10966 3671
rect 10886 3549 10898 3669
rect 10954 3549 10966 3669
rect 10886 3547 10903 3549
rect 10719 3511 10765 3522
rect 10949 3547 10966 3549
rect 10903 3511 10949 3522
rect 10428 3473 10439 3476
rect 10493 3473 10504 3476
rect 10612 3473 10623 3476
rect 10677 3473 10688 3476
rect 10796 3473 10807 3476
rect 10861 3473 10872 3476
rect 10213 3428 10259 3439
rect 10426 3417 10438 3473
rect 10494 3417 10506 3473
rect 10426 3403 10506 3417
rect 10610 3417 10622 3473
rect 10678 3417 10690 3473
rect 10610 3403 10690 3417
rect 10794 3417 10806 3473
rect 10862 3417 10874 3473
rect 11087 3846 11104 3848
rect 11041 3428 11087 3439
rect 10794 3403 10874 3417
rect 10426 3323 10506 3325
rect 10038 3267 10438 3323
rect 10494 3267 10506 3323
rect 8940 3264 9020 3266
rect 10426 3265 10506 3267
rect 9124 3206 9204 3208
rect 8416 3150 9136 3206
rect 9192 3150 9204 3206
rect 9124 3148 9204 3150
rect 9453 3206 9533 3208
rect 9720 3207 9790 3218
rect 10610 3207 10690 3209
rect 9720 3206 10622 3207
rect 9453 3150 9465 3206
rect 9521 3150 9722 3206
rect 9778 3151 10622 3206
rect 10678 3151 10690 3207
rect 9778 3150 10038 3151
rect 9453 3148 9533 3150
rect 9720 3140 9790 3150
rect 10610 3149 10690 3151
rect 10939 3207 11019 3209
rect 11382 3207 11452 3217
rect 10939 3151 10951 3207
rect 11007 3151 11384 3207
rect 11440 3151 11452 3207
rect 10939 3149 11019 3151
rect 11382 3139 11452 3151
rect 12458 3206 12514 4453
rect 15414 4451 15494 4453
rect 15778 4509 15848 4521
rect 16500 4509 16556 5239
rect 17392 5237 17472 5239
rect 18122 5239 18890 5295
rect 18946 5239 18958 5295
rect 17024 5145 17104 5159
rect 16811 5123 16857 5134
rect 17024 5089 17036 5145
rect 17092 5089 17104 5145
rect 17208 5145 17288 5159
rect 17208 5089 17220 5145
rect 17276 5089 17288 5145
rect 17392 5145 17472 5159
rect 17392 5089 17404 5145
rect 17460 5089 17472 5145
rect 17639 5123 17685 5134
rect 17026 5086 17037 5089
rect 17091 5086 17102 5089
rect 17210 5086 17221 5089
rect 17275 5086 17286 5089
rect 17394 5086 17405 5089
rect 17459 5086 17470 5089
rect 16949 5040 16995 5051
rect 16857 4866 16949 5040
rect 16949 4855 16995 4866
rect 17133 5040 17179 5051
rect 17133 4855 17179 4866
rect 17317 5040 17363 5051
rect 17501 5040 17547 5051
rect 17484 5013 17501 5015
rect 17547 5013 17564 5015
rect 17484 4893 17496 5013
rect 17552 4893 17564 5013
rect 17484 4891 17501 4893
rect 17317 4855 17363 4866
rect 17547 4891 17564 4893
rect 17501 4855 17547 4866
rect 16811 4638 16857 4783
rect 17026 4774 17037 4820
rect 17091 4774 17102 4820
rect 17026 4741 17102 4774
rect 17210 4774 17221 4820
rect 17275 4774 17286 4820
rect 17210 4741 17286 4774
rect 17394 4774 17405 4820
rect 17459 4774 17470 4820
rect 17394 4741 17470 4774
rect 17639 4638 17685 4783
rect 16799 4626 16879 4638
rect 16799 4570 16811 4626
rect 16867 4570 16879 4626
rect 16799 4558 16879 4570
rect 17617 4626 17695 4638
rect 17617 4570 17629 4626
rect 17685 4570 17695 4626
rect 17617 4558 17695 4570
rect 15778 4453 15790 4509
rect 15846 4453 16556 4509
rect 18122 4509 18178 5239
rect 18878 5237 18958 5239
rect 20104 5233 20160 5355
rect 20258 5355 20270 5411
rect 20326 5355 21262 5411
rect 21318 5355 21330 5411
rect 20258 5343 20328 5355
rect 21250 5353 21330 5355
rect 21579 5411 21659 5413
rect 22022 5411 22082 5421
rect 22736 5411 22816 5413
rect 21579 5355 21591 5411
rect 21647 5355 22024 5411
rect 22080 5355 22748 5411
rect 22804 5355 22816 5411
rect 21579 5353 21659 5355
rect 22022 5343 22082 5355
rect 22736 5353 22816 5355
rect 23065 5411 23145 5413
rect 23332 5411 23402 5423
rect 24300 5411 24370 5425
rect 25292 5411 25372 5413
rect 23065 5355 23077 5411
rect 23133 5355 23334 5411
rect 23390 5355 24202 5411
rect 23065 5353 23145 5355
rect 23332 5345 23402 5355
rect 21434 5295 21514 5297
rect 22920 5295 23000 5297
rect 20542 5239 21446 5295
rect 21502 5239 21514 5295
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 18510 5145 18590 5159
rect 18297 5123 18343 5134
rect 18510 5089 18522 5145
rect 18578 5089 18590 5145
rect 18694 5145 18774 5159
rect 18694 5089 18706 5145
rect 18762 5089 18774 5145
rect 18878 5145 18958 5159
rect 18878 5089 18890 5145
rect 18946 5089 18958 5145
rect 19125 5123 19171 5134
rect 18512 5086 18523 5089
rect 18577 5086 18588 5089
rect 18696 5086 18707 5089
rect 18761 5086 18772 5089
rect 18880 5086 18891 5089
rect 18945 5086 18956 5089
rect 18435 5040 18481 5051
rect 18343 4866 18435 5040
rect 18435 4855 18481 4866
rect 18619 5040 18665 5051
rect 18619 4855 18665 4866
rect 18803 5040 18849 5051
rect 18987 5040 19033 5051
rect 18970 5013 18987 5015
rect 19033 5013 19050 5015
rect 18970 4893 18982 5013
rect 19038 4893 19050 5013
rect 18970 4891 18987 4893
rect 18803 4855 18849 4866
rect 19033 4891 19050 4893
rect 18987 4855 19033 4866
rect 18297 4638 18343 4783
rect 18512 4774 18523 4820
rect 18577 4774 18588 4820
rect 18512 4741 18588 4774
rect 18696 4774 18707 4820
rect 18761 4774 18772 4820
rect 18696 4741 18772 4774
rect 18880 4774 18891 4820
rect 18945 4774 18956 4820
rect 18880 4741 18956 4774
rect 19125 4638 19171 4783
rect 18285 4626 18365 4638
rect 18285 4570 18297 4626
rect 18353 4570 18365 4626
rect 18285 4558 18365 4570
rect 19103 4626 19181 4638
rect 19103 4570 19115 4626
rect 19171 4570 19181 4626
rect 19103 4558 19181 4570
rect 19456 4509 19536 4519
rect 18122 4453 19468 4509
rect 19524 4453 19536 4509
rect 15778 4441 15848 4453
rect 13938 4398 14008 4400
rect 15238 4399 15318 4401
rect 12594 4342 13940 4398
rect 13996 4342 14008 4398
rect 12594 3322 12650 4342
rect 13938 4330 14008 4342
rect 14080 4343 15250 4399
rect 15306 4343 15318 4399
rect 13258 4291 13344 4295
rect 13258 4235 13270 4291
rect 13326 4235 13344 4291
rect 13258 4223 13344 4235
rect 12769 4078 12815 4089
rect 12984 4087 13060 4120
rect 12984 4041 12995 4087
rect 13049 4041 13060 4087
rect 13168 4087 13244 4120
rect 13168 4041 13179 4087
rect 13233 4041 13244 4087
rect 13352 4087 13428 4120
rect 13352 4041 13363 4087
rect 13417 4041 13428 4087
rect 13597 4078 13643 4089
rect 12907 3995 12953 4006
rect 12890 3968 12907 3970
rect 13091 3995 13137 4006
rect 12953 3968 12970 3970
rect 12815 3848 12902 3968
rect 12958 3848 12970 3968
rect 12890 3846 12907 3848
rect 12815 3548 12907 3668
rect 12953 3846 12970 3848
rect 13074 3668 13091 3670
rect 13275 3995 13321 4006
rect 13258 3968 13275 3970
rect 13459 3995 13505 4006
rect 13321 3968 13338 3970
rect 13258 3848 13270 3968
rect 13326 3848 13338 3968
rect 13258 3846 13275 3848
rect 13137 3668 13154 3670
rect 13074 3548 13086 3668
rect 13142 3548 13154 3668
rect 13074 3546 13091 3548
rect 12907 3510 12953 3521
rect 13137 3546 13154 3548
rect 13091 3510 13137 3521
rect 13321 3846 13338 3848
rect 13442 3668 13459 3670
rect 13580 3968 13597 3970
rect 13643 3968 13660 3970
rect 13580 3847 13592 3968
rect 13648 3847 13660 3968
rect 13580 3845 13597 3847
rect 13505 3668 13522 3670
rect 13442 3548 13454 3668
rect 13510 3548 13522 3668
rect 13442 3546 13459 3548
rect 13275 3510 13321 3521
rect 13505 3546 13522 3548
rect 13459 3510 13505 3521
rect 12984 3472 12995 3475
rect 13049 3472 13060 3475
rect 13168 3472 13179 3475
rect 13233 3472 13244 3475
rect 13352 3472 13363 3475
rect 13417 3472 13428 3475
rect 12769 3427 12815 3438
rect 12982 3416 12994 3472
rect 13050 3416 13062 3472
rect 12982 3402 13062 3416
rect 13166 3416 13178 3472
rect 13234 3416 13246 3472
rect 13166 3402 13246 3416
rect 13350 3416 13362 3472
rect 13418 3416 13430 3472
rect 13643 3845 13660 3847
rect 13597 3427 13643 3438
rect 13350 3402 13430 3416
rect 12982 3322 13062 3324
rect 12594 3266 12994 3322
rect 13050 3266 13062 3322
rect 14080 3323 14136 4343
rect 15238 4331 15318 4343
rect 14744 4292 14830 4296
rect 14744 4236 14756 4292
rect 14812 4236 14830 4292
rect 14744 4224 14830 4236
rect 14255 4079 14301 4090
rect 14470 4088 14546 4121
rect 14470 4042 14481 4088
rect 14535 4042 14546 4088
rect 14654 4088 14730 4121
rect 14654 4042 14665 4088
rect 14719 4042 14730 4088
rect 14838 4088 14914 4121
rect 14838 4042 14849 4088
rect 14903 4042 14914 4088
rect 15083 4079 15129 4090
rect 14393 3996 14439 4007
rect 14376 3969 14393 3971
rect 14577 3996 14623 4007
rect 14439 3969 14456 3971
rect 14301 3849 14388 3969
rect 14444 3849 14456 3969
rect 14376 3847 14393 3849
rect 14301 3549 14393 3669
rect 14439 3847 14456 3849
rect 14560 3669 14577 3671
rect 14761 3996 14807 4007
rect 14744 3969 14761 3971
rect 14945 3996 14991 4007
rect 14807 3969 14824 3971
rect 14744 3849 14756 3969
rect 14812 3849 14824 3969
rect 14744 3847 14761 3849
rect 14623 3669 14640 3671
rect 14560 3549 14572 3669
rect 14628 3549 14640 3669
rect 14560 3547 14577 3549
rect 14393 3511 14439 3522
rect 14623 3547 14640 3549
rect 14577 3511 14623 3522
rect 14807 3847 14824 3849
rect 14928 3669 14945 3671
rect 15066 3969 15083 3971
rect 15129 3969 15146 3971
rect 15066 3848 15078 3969
rect 15134 3848 15146 3969
rect 15066 3846 15083 3848
rect 14991 3669 15008 3671
rect 14928 3549 14940 3669
rect 14996 3549 15008 3669
rect 14928 3547 14945 3549
rect 14761 3511 14807 3522
rect 14991 3547 15008 3549
rect 14945 3511 14991 3522
rect 14470 3473 14481 3476
rect 14535 3473 14546 3476
rect 14654 3473 14665 3476
rect 14719 3473 14730 3476
rect 14838 3473 14849 3476
rect 14903 3473 14914 3476
rect 14255 3428 14301 3439
rect 14468 3417 14480 3473
rect 14536 3417 14548 3473
rect 14468 3403 14548 3417
rect 14652 3417 14664 3473
rect 14720 3417 14732 3473
rect 14652 3403 14732 3417
rect 14836 3417 14848 3473
rect 14904 3417 14916 3473
rect 15129 3846 15146 3848
rect 15083 3428 15129 3439
rect 14836 3403 14916 3417
rect 14468 3323 14548 3325
rect 14080 3267 14480 3323
rect 14536 3267 14548 3323
rect 12982 3264 13062 3266
rect 14468 3265 14548 3267
rect 13166 3206 13246 3208
rect 12458 3150 13178 3206
rect 13234 3150 13246 3206
rect 13166 3148 13246 3150
rect 13495 3206 13575 3208
rect 13762 3207 13832 3218
rect 14652 3207 14732 3209
rect 13762 3206 14664 3207
rect 13495 3150 13507 3206
rect 13563 3150 13764 3206
rect 13820 3151 14664 3206
rect 14720 3151 14732 3207
rect 13820 3150 14080 3151
rect 13495 3148 13575 3150
rect 13762 3140 13832 3150
rect 14652 3149 14732 3151
rect 14981 3207 15061 3209
rect 15424 3207 15494 3217
rect 14981 3151 14993 3207
rect 15049 3151 15426 3207
rect 15482 3151 15494 3207
rect 14981 3149 15061 3151
rect 15424 3139 15494 3151
rect 16500 3206 16556 4453
rect 19456 4451 19536 4453
rect 19820 4509 19890 4521
rect 20542 4509 20598 5239
rect 21434 5237 21514 5239
rect 22164 5239 22932 5295
rect 22988 5239 23000 5295
rect 21066 5145 21146 5159
rect 20853 5123 20899 5134
rect 21066 5089 21078 5145
rect 21134 5089 21146 5145
rect 21250 5145 21330 5159
rect 21250 5089 21262 5145
rect 21318 5089 21330 5145
rect 21434 5145 21514 5159
rect 21434 5089 21446 5145
rect 21502 5089 21514 5145
rect 21681 5123 21727 5134
rect 21068 5086 21079 5089
rect 21133 5086 21144 5089
rect 21252 5086 21263 5089
rect 21317 5086 21328 5089
rect 21436 5086 21447 5089
rect 21501 5086 21512 5089
rect 20991 5040 21037 5051
rect 20899 4866 20991 5040
rect 20991 4855 21037 4866
rect 21175 5040 21221 5051
rect 21175 4855 21221 4866
rect 21359 5040 21405 5051
rect 21543 5040 21589 5051
rect 21526 5013 21543 5015
rect 21589 5013 21606 5015
rect 21526 4893 21538 5013
rect 21594 4893 21606 5013
rect 21526 4891 21543 4893
rect 21359 4855 21405 4866
rect 21589 4891 21606 4893
rect 21543 4855 21589 4866
rect 20853 4638 20899 4783
rect 21068 4774 21079 4820
rect 21133 4774 21144 4820
rect 21068 4741 21144 4774
rect 21252 4774 21263 4820
rect 21317 4774 21328 4820
rect 21252 4741 21328 4774
rect 21436 4774 21447 4820
rect 21501 4774 21512 4820
rect 21436 4741 21512 4774
rect 21681 4638 21727 4783
rect 20841 4626 20921 4638
rect 20841 4570 20853 4626
rect 20909 4570 20921 4626
rect 20841 4558 20921 4570
rect 21659 4626 21737 4638
rect 21659 4570 21671 4626
rect 21727 4570 21737 4626
rect 21659 4558 21737 4570
rect 19820 4453 19832 4509
rect 19888 4453 20598 4509
rect 22164 4509 22220 5239
rect 22920 5237 23000 5239
rect 24146 5233 24202 5355
rect 24300 5355 24312 5411
rect 24368 5355 25304 5411
rect 25360 5355 25372 5411
rect 24300 5343 24370 5355
rect 25292 5353 25372 5355
rect 25621 5411 25701 5413
rect 26064 5411 26124 5421
rect 26778 5411 26858 5413
rect 25621 5355 25633 5411
rect 25689 5355 26066 5411
rect 26122 5355 26790 5411
rect 26846 5355 26858 5411
rect 25621 5353 25701 5355
rect 26064 5343 26124 5355
rect 26778 5353 26858 5355
rect 27107 5411 27187 5413
rect 27374 5411 27444 5423
rect 27107 5355 27119 5411
rect 27175 5355 27376 5411
rect 27432 5355 27444 5411
rect 27107 5353 27187 5355
rect 27374 5345 27444 5355
rect 25476 5295 25556 5297
rect 26962 5295 27042 5297
rect 24584 5239 25488 5295
rect 25544 5239 25556 5295
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect 22552 5145 22632 5159
rect 22339 5123 22385 5134
rect 22552 5089 22564 5145
rect 22620 5089 22632 5145
rect 22736 5145 22816 5159
rect 22736 5089 22748 5145
rect 22804 5089 22816 5145
rect 22920 5145 23000 5159
rect 22920 5089 22932 5145
rect 22988 5089 23000 5145
rect 23167 5123 23213 5134
rect 22554 5086 22565 5089
rect 22619 5086 22630 5089
rect 22738 5086 22749 5089
rect 22803 5086 22814 5089
rect 22922 5086 22933 5089
rect 22987 5086 22998 5089
rect 22477 5040 22523 5051
rect 22385 4866 22477 5040
rect 22477 4855 22523 4866
rect 22661 5040 22707 5051
rect 22661 4855 22707 4866
rect 22845 5040 22891 5051
rect 23029 5040 23075 5051
rect 23012 5013 23029 5015
rect 23075 5013 23092 5015
rect 23012 4893 23024 5013
rect 23080 4893 23092 5013
rect 23012 4891 23029 4893
rect 22845 4855 22891 4866
rect 23075 4891 23092 4893
rect 23029 4855 23075 4866
rect 22339 4638 22385 4783
rect 22554 4774 22565 4820
rect 22619 4774 22630 4820
rect 22554 4741 22630 4774
rect 22738 4774 22749 4820
rect 22803 4774 22814 4820
rect 22738 4741 22814 4774
rect 22922 4774 22933 4820
rect 22987 4774 22998 4820
rect 22922 4741 22998 4774
rect 23167 4638 23213 4783
rect 22327 4626 22407 4638
rect 22327 4570 22339 4626
rect 22395 4570 22407 4626
rect 22327 4558 22407 4570
rect 23145 4626 23223 4638
rect 23145 4570 23157 4626
rect 23213 4570 23223 4626
rect 23145 4558 23223 4570
rect 23498 4509 23578 4519
rect 22164 4453 23510 4509
rect 23566 4453 23578 4509
rect 19820 4441 19890 4453
rect 17980 4398 18050 4400
rect 19280 4399 19360 4401
rect 16636 4342 17982 4398
rect 18038 4342 18050 4398
rect 16636 3322 16692 4342
rect 17980 4330 18050 4342
rect 18122 4343 19292 4399
rect 19348 4343 19360 4399
rect 17300 4291 17386 4295
rect 17300 4235 17312 4291
rect 17368 4235 17386 4291
rect 17300 4223 17386 4235
rect 16811 4078 16857 4089
rect 17026 4087 17102 4120
rect 17026 4041 17037 4087
rect 17091 4041 17102 4087
rect 17210 4087 17286 4120
rect 17210 4041 17221 4087
rect 17275 4041 17286 4087
rect 17394 4087 17470 4120
rect 17394 4041 17405 4087
rect 17459 4041 17470 4087
rect 17639 4078 17685 4089
rect 16949 3995 16995 4006
rect 16932 3968 16949 3970
rect 17133 3995 17179 4006
rect 16995 3968 17012 3970
rect 16857 3848 16944 3968
rect 17000 3848 17012 3968
rect 16932 3846 16949 3848
rect 16857 3548 16949 3668
rect 16995 3846 17012 3848
rect 17116 3668 17133 3670
rect 17317 3995 17363 4006
rect 17300 3968 17317 3970
rect 17501 3995 17547 4006
rect 17363 3968 17380 3970
rect 17300 3848 17312 3968
rect 17368 3848 17380 3968
rect 17300 3846 17317 3848
rect 17179 3668 17196 3670
rect 17116 3548 17128 3668
rect 17184 3548 17196 3668
rect 17116 3546 17133 3548
rect 16949 3510 16995 3521
rect 17179 3546 17196 3548
rect 17133 3510 17179 3521
rect 17363 3846 17380 3848
rect 17484 3668 17501 3670
rect 17622 3968 17639 3970
rect 17685 3968 17702 3970
rect 17622 3847 17634 3968
rect 17690 3847 17702 3968
rect 17622 3845 17639 3847
rect 17547 3668 17564 3670
rect 17484 3548 17496 3668
rect 17552 3548 17564 3668
rect 17484 3546 17501 3548
rect 17317 3510 17363 3521
rect 17547 3546 17564 3548
rect 17501 3510 17547 3521
rect 17026 3472 17037 3475
rect 17091 3472 17102 3475
rect 17210 3472 17221 3475
rect 17275 3472 17286 3475
rect 17394 3472 17405 3475
rect 17459 3472 17470 3475
rect 16811 3427 16857 3438
rect 17024 3416 17036 3472
rect 17092 3416 17104 3472
rect 17024 3402 17104 3416
rect 17208 3416 17220 3472
rect 17276 3416 17288 3472
rect 17208 3402 17288 3416
rect 17392 3416 17404 3472
rect 17460 3416 17472 3472
rect 17685 3845 17702 3847
rect 17639 3427 17685 3438
rect 17392 3402 17472 3416
rect 17024 3322 17104 3324
rect 16636 3266 17036 3322
rect 17092 3266 17104 3322
rect 18122 3323 18178 4343
rect 19280 4331 19360 4343
rect 18786 4292 18872 4296
rect 18786 4236 18798 4292
rect 18854 4236 18872 4292
rect 18786 4224 18872 4236
rect 18297 4079 18343 4090
rect 18512 4088 18588 4121
rect 18512 4042 18523 4088
rect 18577 4042 18588 4088
rect 18696 4088 18772 4121
rect 18696 4042 18707 4088
rect 18761 4042 18772 4088
rect 18880 4088 18956 4121
rect 18880 4042 18891 4088
rect 18945 4042 18956 4088
rect 19125 4079 19171 4090
rect 18435 3996 18481 4007
rect 18418 3969 18435 3971
rect 18619 3996 18665 4007
rect 18481 3969 18498 3971
rect 18343 3849 18430 3969
rect 18486 3849 18498 3969
rect 18418 3847 18435 3849
rect 18343 3549 18435 3669
rect 18481 3847 18498 3849
rect 18602 3669 18619 3671
rect 18803 3996 18849 4007
rect 18786 3969 18803 3971
rect 18987 3996 19033 4007
rect 18849 3969 18866 3971
rect 18786 3849 18798 3969
rect 18854 3849 18866 3969
rect 18786 3847 18803 3849
rect 18665 3669 18682 3671
rect 18602 3549 18614 3669
rect 18670 3549 18682 3669
rect 18602 3547 18619 3549
rect 18435 3511 18481 3522
rect 18665 3547 18682 3549
rect 18619 3511 18665 3522
rect 18849 3847 18866 3849
rect 18970 3669 18987 3671
rect 19108 3969 19125 3971
rect 19171 3969 19188 3971
rect 19108 3848 19120 3969
rect 19176 3848 19188 3969
rect 19108 3846 19125 3848
rect 19033 3669 19050 3671
rect 18970 3549 18982 3669
rect 19038 3549 19050 3669
rect 18970 3547 18987 3549
rect 18803 3511 18849 3522
rect 19033 3547 19050 3549
rect 18987 3511 19033 3522
rect 18512 3473 18523 3476
rect 18577 3473 18588 3476
rect 18696 3473 18707 3476
rect 18761 3473 18772 3476
rect 18880 3473 18891 3476
rect 18945 3473 18956 3476
rect 18297 3428 18343 3439
rect 18510 3417 18522 3473
rect 18578 3417 18590 3473
rect 18510 3403 18590 3417
rect 18694 3417 18706 3473
rect 18762 3417 18774 3473
rect 18694 3403 18774 3417
rect 18878 3417 18890 3473
rect 18946 3417 18958 3473
rect 19171 3846 19188 3848
rect 19125 3428 19171 3439
rect 18878 3403 18958 3417
rect 18510 3323 18590 3325
rect 18122 3267 18522 3323
rect 18578 3267 18590 3323
rect 17024 3264 17104 3266
rect 18510 3265 18590 3267
rect 17208 3206 17288 3208
rect 16500 3150 17220 3206
rect 17276 3150 17288 3206
rect 17208 3148 17288 3150
rect 17537 3206 17617 3208
rect 17804 3207 17874 3218
rect 18694 3207 18774 3209
rect 17804 3206 18706 3207
rect 17537 3150 17549 3206
rect 17605 3150 17806 3206
rect 17862 3151 18706 3206
rect 18762 3151 18774 3207
rect 17862 3150 18122 3151
rect 17537 3148 17617 3150
rect 17804 3140 17874 3150
rect 18694 3149 18774 3151
rect 19023 3207 19103 3209
rect 19466 3207 19536 3217
rect 19023 3151 19035 3207
rect 19091 3151 19468 3207
rect 19524 3151 19536 3207
rect 19023 3149 19103 3151
rect 19466 3139 19536 3151
rect 20542 3206 20598 4453
rect 23498 4451 23578 4453
rect 23862 4509 23932 4521
rect 24584 4509 24640 5239
rect 25476 5237 25556 5239
rect 26206 5239 26974 5295
rect 27030 5239 27042 5295
rect 25108 5145 25188 5159
rect 24895 5123 24941 5134
rect 25108 5089 25120 5145
rect 25176 5089 25188 5145
rect 25292 5145 25372 5159
rect 25292 5089 25304 5145
rect 25360 5089 25372 5145
rect 25476 5145 25556 5159
rect 25476 5089 25488 5145
rect 25544 5089 25556 5145
rect 25723 5123 25769 5134
rect 25110 5086 25121 5089
rect 25175 5086 25186 5089
rect 25294 5086 25305 5089
rect 25359 5086 25370 5089
rect 25478 5086 25489 5089
rect 25543 5086 25554 5089
rect 25033 5040 25079 5051
rect 24941 4866 25033 5040
rect 25033 4855 25079 4866
rect 25217 5040 25263 5051
rect 25217 4855 25263 4866
rect 25401 5040 25447 5051
rect 25585 5040 25631 5051
rect 25568 5013 25585 5015
rect 25631 5013 25648 5015
rect 25568 4893 25580 5013
rect 25636 4893 25648 5013
rect 25568 4891 25585 4893
rect 25401 4855 25447 4866
rect 25631 4891 25648 4893
rect 25585 4855 25631 4866
rect 24895 4638 24941 4783
rect 25110 4774 25121 4820
rect 25175 4774 25186 4820
rect 25110 4741 25186 4774
rect 25294 4774 25305 4820
rect 25359 4774 25370 4820
rect 25294 4741 25370 4774
rect 25478 4774 25489 4820
rect 25543 4774 25554 4820
rect 25478 4741 25554 4774
rect 25723 4638 25769 4783
rect 24883 4626 24963 4638
rect 24883 4570 24895 4626
rect 24951 4570 24963 4626
rect 24883 4558 24963 4570
rect 25701 4626 25779 4638
rect 25701 4570 25713 4626
rect 25769 4570 25779 4626
rect 25701 4558 25779 4570
rect 23862 4453 23874 4509
rect 23930 4453 24640 4509
rect 26206 4509 26262 5239
rect 26962 5237 27042 5239
rect 26594 5145 26674 5159
rect 26381 5123 26427 5134
rect 26594 5089 26606 5145
rect 26662 5089 26674 5145
rect 26778 5145 26858 5159
rect 26778 5089 26790 5145
rect 26846 5089 26858 5145
rect 26962 5145 27042 5159
rect 26962 5089 26974 5145
rect 27030 5089 27042 5145
rect 27209 5123 27255 5134
rect 26596 5086 26607 5089
rect 26661 5086 26672 5089
rect 26780 5086 26791 5089
rect 26845 5086 26856 5089
rect 26964 5086 26975 5089
rect 27029 5086 27040 5089
rect 26519 5040 26565 5051
rect 26427 4866 26519 5040
rect 26519 4855 26565 4866
rect 26703 5040 26749 5051
rect 26703 4855 26749 4866
rect 26887 5040 26933 5051
rect 27071 5040 27117 5051
rect 27054 5013 27071 5015
rect 27117 5013 27134 5015
rect 27054 4893 27066 5013
rect 27122 4893 27134 5013
rect 27054 4891 27071 4893
rect 26887 4855 26933 4866
rect 27117 4891 27134 4893
rect 27071 4855 27117 4866
rect 26381 4638 26427 4783
rect 26596 4774 26607 4820
rect 26661 4774 26672 4820
rect 26596 4741 26672 4774
rect 26780 4774 26791 4820
rect 26845 4774 26856 4820
rect 26780 4741 26856 4774
rect 26964 4774 26975 4820
rect 27029 4774 27040 4820
rect 26964 4741 27040 4774
rect 27209 4638 27255 4783
rect 26369 4626 26449 4638
rect 26369 4570 26381 4626
rect 26437 4570 26449 4626
rect 26369 4558 26449 4570
rect 27187 4626 27265 4638
rect 27187 4570 27199 4626
rect 27255 4570 27265 4626
rect 27187 4558 27265 4570
rect 27540 4509 27620 4519
rect 26206 4453 27552 4509
rect 27608 4453 27620 4509
rect 23862 4441 23932 4453
rect 22022 4398 22092 4400
rect 23322 4399 23402 4401
rect 20678 4342 22024 4398
rect 22080 4342 22092 4398
rect 20678 3322 20734 4342
rect 22022 4330 22092 4342
rect 22164 4343 23334 4399
rect 23390 4343 23402 4399
rect 21342 4291 21428 4295
rect 21342 4235 21354 4291
rect 21410 4235 21428 4291
rect 21342 4223 21428 4235
rect 20853 4078 20899 4089
rect 21068 4087 21144 4120
rect 21068 4041 21079 4087
rect 21133 4041 21144 4087
rect 21252 4087 21328 4120
rect 21252 4041 21263 4087
rect 21317 4041 21328 4087
rect 21436 4087 21512 4120
rect 21436 4041 21447 4087
rect 21501 4041 21512 4087
rect 21681 4078 21727 4089
rect 20991 3995 21037 4006
rect 20974 3968 20991 3970
rect 21175 3995 21221 4006
rect 21037 3968 21054 3970
rect 20899 3848 20986 3968
rect 21042 3848 21054 3968
rect 20974 3846 20991 3848
rect 20899 3548 20991 3668
rect 21037 3846 21054 3848
rect 21158 3668 21175 3670
rect 21359 3995 21405 4006
rect 21342 3968 21359 3970
rect 21543 3995 21589 4006
rect 21405 3968 21422 3970
rect 21342 3848 21354 3968
rect 21410 3848 21422 3968
rect 21342 3846 21359 3848
rect 21221 3668 21238 3670
rect 21158 3548 21170 3668
rect 21226 3548 21238 3668
rect 21158 3546 21175 3548
rect 20991 3510 21037 3521
rect 21221 3546 21238 3548
rect 21175 3510 21221 3521
rect 21405 3846 21422 3848
rect 21526 3668 21543 3670
rect 21664 3968 21681 3970
rect 21727 3968 21744 3970
rect 21664 3847 21676 3968
rect 21732 3847 21744 3968
rect 21664 3845 21681 3847
rect 21589 3668 21606 3670
rect 21526 3548 21538 3668
rect 21594 3548 21606 3668
rect 21526 3546 21543 3548
rect 21359 3510 21405 3521
rect 21589 3546 21606 3548
rect 21543 3510 21589 3521
rect 21068 3472 21079 3475
rect 21133 3472 21144 3475
rect 21252 3472 21263 3475
rect 21317 3472 21328 3475
rect 21436 3472 21447 3475
rect 21501 3472 21512 3475
rect 20853 3427 20899 3438
rect 21066 3416 21078 3472
rect 21134 3416 21146 3472
rect 21066 3402 21146 3416
rect 21250 3416 21262 3472
rect 21318 3416 21330 3472
rect 21250 3402 21330 3416
rect 21434 3416 21446 3472
rect 21502 3416 21514 3472
rect 21727 3845 21744 3847
rect 21681 3427 21727 3438
rect 21434 3402 21514 3416
rect 21066 3322 21146 3324
rect 20678 3266 21078 3322
rect 21134 3266 21146 3322
rect 22164 3323 22220 4343
rect 23322 4331 23402 4343
rect 22828 4292 22914 4296
rect 22828 4236 22840 4292
rect 22896 4236 22914 4292
rect 22828 4224 22914 4236
rect 22339 4079 22385 4090
rect 22554 4088 22630 4121
rect 22554 4042 22565 4088
rect 22619 4042 22630 4088
rect 22738 4088 22814 4121
rect 22738 4042 22749 4088
rect 22803 4042 22814 4088
rect 22922 4088 22998 4121
rect 22922 4042 22933 4088
rect 22987 4042 22998 4088
rect 23167 4079 23213 4090
rect 22477 3996 22523 4007
rect 22460 3969 22477 3971
rect 22661 3996 22707 4007
rect 22523 3969 22540 3971
rect 22385 3849 22472 3969
rect 22528 3849 22540 3969
rect 22460 3847 22477 3849
rect 22385 3549 22477 3669
rect 22523 3847 22540 3849
rect 22644 3669 22661 3671
rect 22845 3996 22891 4007
rect 22828 3969 22845 3971
rect 23029 3996 23075 4007
rect 22891 3969 22908 3971
rect 22828 3849 22840 3969
rect 22896 3849 22908 3969
rect 22828 3847 22845 3849
rect 22707 3669 22724 3671
rect 22644 3549 22656 3669
rect 22712 3549 22724 3669
rect 22644 3547 22661 3549
rect 22477 3511 22523 3522
rect 22707 3547 22724 3549
rect 22661 3511 22707 3522
rect 22891 3847 22908 3849
rect 23012 3669 23029 3671
rect 23150 3969 23167 3971
rect 23213 3969 23230 3971
rect 23150 3848 23162 3969
rect 23218 3848 23230 3969
rect 23150 3846 23167 3848
rect 23075 3669 23092 3671
rect 23012 3549 23024 3669
rect 23080 3549 23092 3669
rect 23012 3547 23029 3549
rect 22845 3511 22891 3522
rect 23075 3547 23092 3549
rect 23029 3511 23075 3522
rect 22554 3473 22565 3476
rect 22619 3473 22630 3476
rect 22738 3473 22749 3476
rect 22803 3473 22814 3476
rect 22922 3473 22933 3476
rect 22987 3473 22998 3476
rect 22339 3428 22385 3439
rect 22552 3417 22564 3473
rect 22620 3417 22632 3473
rect 22552 3403 22632 3417
rect 22736 3417 22748 3473
rect 22804 3417 22816 3473
rect 22736 3403 22816 3417
rect 22920 3417 22932 3473
rect 22988 3417 23000 3473
rect 23213 3846 23230 3848
rect 23167 3428 23213 3439
rect 22920 3403 23000 3417
rect 22552 3323 22632 3325
rect 22164 3267 22564 3323
rect 22620 3267 22632 3323
rect 21066 3264 21146 3266
rect 22552 3265 22632 3267
rect 21250 3206 21330 3208
rect 20542 3150 21262 3206
rect 21318 3150 21330 3206
rect 21250 3148 21330 3150
rect 21579 3206 21659 3208
rect 21846 3207 21916 3218
rect 22736 3207 22816 3209
rect 21846 3206 22748 3207
rect 21579 3150 21591 3206
rect 21647 3150 21848 3206
rect 21904 3151 22748 3206
rect 22804 3151 22816 3207
rect 21904 3150 22164 3151
rect 21579 3148 21659 3150
rect 21846 3140 21916 3150
rect 22736 3149 22816 3151
rect 23065 3207 23145 3209
rect 23508 3207 23578 3217
rect 23065 3151 23077 3207
rect 23133 3151 23510 3207
rect 23566 3151 23578 3207
rect 23065 3149 23145 3151
rect 23508 3139 23578 3151
rect 24584 3206 24640 4453
rect 27540 4451 27620 4453
rect 26064 4398 26134 4400
rect 27364 4399 27444 4401
rect 24720 4342 26066 4398
rect 26122 4342 26134 4398
rect 24720 3322 24776 4342
rect 26064 4330 26134 4342
rect 26206 4343 27376 4399
rect 27432 4343 27444 4399
rect 25384 4291 25470 4295
rect 25384 4235 25396 4291
rect 25452 4235 25470 4291
rect 25384 4223 25470 4235
rect 24895 4078 24941 4089
rect 25110 4087 25186 4120
rect 25110 4041 25121 4087
rect 25175 4041 25186 4087
rect 25294 4087 25370 4120
rect 25294 4041 25305 4087
rect 25359 4041 25370 4087
rect 25478 4087 25554 4120
rect 25478 4041 25489 4087
rect 25543 4041 25554 4087
rect 25723 4078 25769 4089
rect 25033 3995 25079 4006
rect 25016 3968 25033 3970
rect 25217 3995 25263 4006
rect 25079 3968 25096 3970
rect 24941 3848 25028 3968
rect 25084 3848 25096 3968
rect 25016 3846 25033 3848
rect 24941 3548 25033 3668
rect 25079 3846 25096 3848
rect 25200 3668 25217 3670
rect 25401 3995 25447 4006
rect 25384 3968 25401 3970
rect 25585 3995 25631 4006
rect 25447 3968 25464 3970
rect 25384 3848 25396 3968
rect 25452 3848 25464 3968
rect 25384 3846 25401 3848
rect 25263 3668 25280 3670
rect 25200 3548 25212 3668
rect 25268 3548 25280 3668
rect 25200 3546 25217 3548
rect 25033 3510 25079 3521
rect 25263 3546 25280 3548
rect 25217 3510 25263 3521
rect 25447 3846 25464 3848
rect 25568 3668 25585 3670
rect 25706 3968 25723 3970
rect 25769 3968 25786 3970
rect 25706 3847 25718 3968
rect 25774 3847 25786 3968
rect 25706 3845 25723 3847
rect 25631 3668 25648 3670
rect 25568 3548 25580 3668
rect 25636 3548 25648 3668
rect 25568 3546 25585 3548
rect 25401 3510 25447 3521
rect 25631 3546 25648 3548
rect 25585 3510 25631 3521
rect 25110 3472 25121 3475
rect 25175 3472 25186 3475
rect 25294 3472 25305 3475
rect 25359 3472 25370 3475
rect 25478 3472 25489 3475
rect 25543 3472 25554 3475
rect 24895 3427 24941 3438
rect 25108 3416 25120 3472
rect 25176 3416 25188 3472
rect 25108 3402 25188 3416
rect 25292 3416 25304 3472
rect 25360 3416 25372 3472
rect 25292 3402 25372 3416
rect 25476 3416 25488 3472
rect 25544 3416 25556 3472
rect 25769 3845 25786 3847
rect 25723 3427 25769 3438
rect 25476 3402 25556 3416
rect 25108 3322 25188 3324
rect 24720 3266 25120 3322
rect 25176 3266 25188 3322
rect 26206 3323 26262 4343
rect 27364 4331 27444 4343
rect 26870 4292 26956 4296
rect 26870 4236 26882 4292
rect 26938 4236 26956 4292
rect 26870 4224 26956 4236
rect 26381 4079 26427 4090
rect 26596 4088 26672 4121
rect 26596 4042 26607 4088
rect 26661 4042 26672 4088
rect 26780 4088 26856 4121
rect 26780 4042 26791 4088
rect 26845 4042 26856 4088
rect 26964 4088 27040 4121
rect 26964 4042 26975 4088
rect 27029 4042 27040 4088
rect 27209 4079 27255 4090
rect 26519 3996 26565 4007
rect 26502 3969 26519 3971
rect 26703 3996 26749 4007
rect 26565 3969 26582 3971
rect 26427 3849 26514 3969
rect 26570 3849 26582 3969
rect 26502 3847 26519 3849
rect 26427 3549 26519 3669
rect 26565 3847 26582 3849
rect 26686 3669 26703 3671
rect 26887 3996 26933 4007
rect 26870 3969 26887 3971
rect 27071 3996 27117 4007
rect 26933 3969 26950 3971
rect 26870 3849 26882 3969
rect 26938 3849 26950 3969
rect 26870 3847 26887 3849
rect 26749 3669 26766 3671
rect 26686 3549 26698 3669
rect 26754 3549 26766 3669
rect 26686 3547 26703 3549
rect 26519 3511 26565 3522
rect 26749 3547 26766 3549
rect 26703 3511 26749 3522
rect 26933 3847 26950 3849
rect 27054 3669 27071 3671
rect 27192 3969 27209 3971
rect 27255 3969 27272 3971
rect 27192 3848 27204 3969
rect 27260 3848 27272 3969
rect 27192 3846 27209 3848
rect 27117 3669 27134 3671
rect 27054 3549 27066 3669
rect 27122 3549 27134 3669
rect 27054 3547 27071 3549
rect 26887 3511 26933 3522
rect 27117 3547 27134 3549
rect 27071 3511 27117 3522
rect 26596 3473 26607 3476
rect 26661 3473 26672 3476
rect 26780 3473 26791 3476
rect 26845 3473 26856 3476
rect 26964 3473 26975 3476
rect 27029 3473 27040 3476
rect 26381 3428 26427 3439
rect 26594 3417 26606 3473
rect 26662 3417 26674 3473
rect 26594 3403 26674 3417
rect 26778 3417 26790 3473
rect 26846 3417 26858 3473
rect 26778 3403 26858 3417
rect 26962 3417 26974 3473
rect 27030 3417 27042 3473
rect 27255 3846 27272 3848
rect 27209 3428 27255 3439
rect 26962 3403 27042 3417
rect 26594 3323 26674 3325
rect 26206 3267 26606 3323
rect 26662 3267 26674 3323
rect 25108 3264 25188 3266
rect 26594 3265 26674 3267
rect 25292 3206 25372 3208
rect 24584 3150 25304 3206
rect 25360 3150 25372 3206
rect 25292 3148 25372 3150
rect 25621 3206 25701 3208
rect 25888 3207 25958 3218
rect 26778 3207 26858 3209
rect 25888 3206 26790 3207
rect 25621 3150 25633 3206
rect 25689 3150 25890 3206
rect 25946 3151 26790 3206
rect 26846 3151 26858 3207
rect 25946 3150 26206 3151
rect 25621 3148 25701 3150
rect 25888 3140 25958 3150
rect 26778 3149 26858 3151
rect 27107 3207 27187 3209
rect 27550 3207 27620 3217
rect 27107 3151 27119 3207
rect 27175 3151 27552 3207
rect 27608 3151 27620 3207
rect 27107 3149 27187 3151
rect 27550 3139 27620 3151
rect 214 3090 284 3102
rect 1254 3090 1334 3092
rect 2740 3091 2820 3093
rect 214 3034 226 3090
rect 282 3034 1266 3090
rect 1322 3034 1334 3090
rect 214 3022 284 3034
rect 498 2303 554 3034
rect 1254 3032 1334 3034
rect 1984 3035 2752 3091
rect 2808 3035 2820 3091
rect 886 2940 966 2954
rect 673 2918 719 2929
rect 886 2884 898 2940
rect 954 2884 966 2940
rect 1070 2940 1150 2954
rect 1070 2884 1082 2940
rect 1138 2884 1150 2940
rect 1254 2940 1334 2954
rect 1254 2884 1266 2940
rect 1322 2884 1334 2940
rect 1501 2918 1547 2929
rect 888 2881 899 2884
rect 953 2881 964 2884
rect 1072 2881 1083 2884
rect 1137 2881 1148 2884
rect 1256 2881 1267 2884
rect 1321 2881 1332 2884
rect 811 2835 857 2846
rect 719 2661 811 2835
rect 811 2650 857 2661
rect 995 2835 1041 2846
rect 995 2650 1041 2661
rect 1179 2835 1225 2846
rect 1363 2835 1409 2846
rect 1346 2808 1363 2810
rect 1409 2808 1426 2810
rect 1346 2688 1358 2808
rect 1414 2688 1426 2808
rect 1346 2686 1363 2688
rect 1179 2650 1225 2661
rect 1409 2686 1426 2688
rect 1363 2650 1409 2661
rect 673 2433 719 2578
rect 888 2569 899 2615
rect 953 2569 964 2615
rect 888 2536 964 2569
rect 1072 2569 1083 2615
rect 1137 2569 1148 2615
rect 1072 2536 1148 2569
rect 1256 2569 1267 2615
rect 1321 2569 1332 2615
rect 1256 2536 1332 2569
rect 1501 2433 1547 2578
rect 661 2421 741 2433
rect 661 2365 673 2421
rect 729 2365 741 2421
rect 661 2353 741 2365
rect 1479 2421 1557 2433
rect 1479 2365 1491 2421
rect 1547 2365 1557 2421
rect 1479 2353 1557 2365
rect 1832 2303 1912 2313
rect 498 2247 1844 2303
rect 1900 2247 1912 2303
rect 1832 2245 1912 2247
rect 1666 2194 1736 2196
rect 498 2193 1736 2194
rect 498 2139 1668 2193
rect 1724 2139 1736 2193
rect 498 2138 1736 2139
rect 498 1117 554 2138
rect 1666 2130 1736 2138
rect 1162 2086 1248 2090
rect 1162 2030 1174 2086
rect 1230 2030 1248 2086
rect 1162 2018 1248 2030
rect 673 1873 719 1884
rect 888 1882 964 1915
rect 888 1836 899 1882
rect 953 1836 964 1882
rect 1072 1882 1148 1915
rect 1072 1836 1083 1882
rect 1137 1836 1148 1882
rect 1256 1882 1332 1915
rect 1256 1836 1267 1882
rect 1321 1836 1332 1882
rect 1501 1873 1547 1884
rect 811 1790 857 1801
rect 794 1763 811 1765
rect 995 1790 1041 1801
rect 857 1763 874 1765
rect 719 1643 806 1763
rect 862 1643 874 1763
rect 794 1641 811 1643
rect 719 1343 811 1463
rect 857 1641 874 1643
rect 978 1463 995 1465
rect 1179 1790 1225 1801
rect 1162 1763 1179 1765
rect 1363 1790 1409 1801
rect 1225 1763 1242 1765
rect 1162 1643 1174 1763
rect 1230 1643 1242 1763
rect 1162 1641 1179 1643
rect 1041 1463 1058 1465
rect 978 1343 990 1463
rect 1046 1343 1058 1463
rect 978 1341 995 1343
rect 811 1305 857 1316
rect 1041 1341 1058 1343
rect 995 1305 1041 1316
rect 1225 1641 1242 1643
rect 1346 1463 1363 1465
rect 1484 1763 1501 1765
rect 1547 1763 1564 1765
rect 1484 1642 1496 1763
rect 1552 1642 1564 1763
rect 1484 1640 1501 1642
rect 1409 1463 1426 1465
rect 1346 1343 1358 1463
rect 1414 1343 1426 1463
rect 1346 1341 1363 1343
rect 1179 1305 1225 1316
rect 1409 1341 1426 1343
rect 1363 1305 1409 1316
rect 888 1267 899 1270
rect 953 1267 964 1270
rect 1072 1267 1083 1270
rect 1137 1267 1148 1270
rect 1256 1267 1267 1270
rect 1321 1267 1332 1270
rect 673 1222 719 1233
rect 886 1211 898 1267
rect 954 1211 966 1267
rect 886 1197 966 1211
rect 1070 1211 1082 1267
rect 1138 1211 1150 1267
rect 1070 1197 1150 1211
rect 1254 1211 1266 1267
rect 1322 1211 1334 1267
rect 1547 1640 1564 1642
rect 1501 1222 1547 1233
rect 1254 1197 1334 1211
rect 886 1117 966 1119
rect 498 1061 898 1117
rect 954 1061 966 1117
rect 886 1059 966 1061
rect 78 1001 148 1015
rect 1070 1001 1150 1003
rect 78 945 90 1001
rect 146 945 1082 1001
rect 1138 945 1150 1001
rect 78 933 148 945
rect 1070 943 1150 945
rect 1399 1001 1479 1003
rect 1842 1001 1902 1013
rect 1399 945 1411 1001
rect 1467 945 1844 1001
rect 1900 945 1902 1001
rect 1399 943 1479 945
rect 1842 933 1902 945
rect -121 885 -41 897
rect 1254 885 1334 887
rect -121 829 -109 885
rect -53 829 1266 885
rect 1322 829 1334 885
rect -121 817 -41 829
rect 1254 827 1334 829
rect 886 735 966 749
rect 673 713 719 724
rect 886 679 898 735
rect 954 679 966 735
rect 1070 735 1150 749
rect 1070 679 1082 735
rect 1138 679 1150 735
rect 1254 735 1334 749
rect 1254 679 1266 735
rect 1322 679 1334 735
rect 1501 713 1547 724
rect 888 676 899 679
rect 953 676 964 679
rect 1072 676 1083 679
rect 1137 676 1148 679
rect 1256 676 1267 679
rect 1321 676 1332 679
rect 811 630 857 641
rect 719 456 811 630
rect 811 445 857 456
rect 995 630 1041 641
rect 995 445 1041 456
rect 1179 630 1225 641
rect 1363 630 1409 641
rect 1346 603 1363 605
rect 1409 603 1426 605
rect 1346 483 1358 603
rect 1414 483 1426 603
rect 1346 481 1363 483
rect 1179 445 1225 456
rect 1409 481 1426 483
rect 1363 445 1409 456
rect 673 228 719 373
rect 888 364 899 410
rect 953 364 964 410
rect 888 331 964 364
rect 1072 364 1083 410
rect 1137 364 1148 410
rect 1072 331 1148 364
rect 1256 364 1267 410
rect 1321 364 1332 410
rect 1256 331 1332 364
rect 1501 228 1547 373
rect 661 216 741 228
rect 661 160 673 216
rect 729 160 741 216
rect 661 148 741 160
rect 1479 216 1559 228
rect 1479 160 1491 216
rect 1547 160 1559 216
rect 1479 148 1559 160
rect -121 98 -35 110
rect 88 98 148 102
rect 1984 98 2040 3035
rect 2740 3033 2820 3035
rect 4226 3090 4296 3102
rect 5266 3090 5346 3092
rect 6752 3091 6832 3093
rect 4226 3034 4238 3090
rect 4294 3034 5278 3090
rect 5334 3034 5346 3090
rect 4226 3022 4296 3034
rect 2372 2941 2452 2955
rect 2159 2919 2205 2930
rect 2372 2885 2384 2941
rect 2440 2885 2452 2941
rect 2556 2941 2636 2955
rect 2556 2885 2568 2941
rect 2624 2885 2636 2941
rect 2740 2941 2820 2955
rect 2740 2885 2752 2941
rect 2808 2885 2820 2941
rect 2987 2919 3033 2930
rect 2374 2882 2385 2885
rect 2439 2882 2450 2885
rect 2558 2882 2569 2885
rect 2623 2882 2634 2885
rect 2742 2882 2753 2885
rect 2807 2882 2818 2885
rect 2297 2836 2343 2847
rect 2205 2662 2297 2836
rect 2297 2651 2343 2662
rect 2481 2836 2527 2847
rect 2481 2651 2527 2662
rect 2665 2836 2711 2847
rect 2849 2836 2895 2847
rect 2832 2809 2849 2811
rect 2895 2809 2912 2811
rect 2832 2689 2844 2809
rect 2900 2689 2912 2809
rect 2832 2687 2849 2689
rect 2665 2651 2711 2662
rect 2895 2687 2912 2689
rect 2849 2651 2895 2662
rect 2159 2434 2205 2579
rect 2374 2570 2385 2616
rect 2439 2570 2450 2616
rect 2374 2537 2450 2570
rect 2558 2570 2569 2616
rect 2623 2570 2634 2616
rect 2558 2537 2634 2570
rect 2742 2570 2753 2616
rect 2807 2570 2818 2616
rect 2742 2537 2818 2570
rect 2987 2434 3033 2579
rect 2147 2422 2227 2434
rect 2147 2366 2159 2422
rect 2215 2366 2227 2422
rect 2147 2354 2227 2366
rect 2965 2422 3043 2434
rect 2965 2366 2977 2422
rect 3033 2366 3043 2422
rect 2965 2354 3043 2366
rect 4510 2303 4566 3034
rect 5266 3032 5346 3034
rect 5996 3035 6764 3091
rect 6820 3035 6832 3091
rect 4898 2940 4978 2954
rect 4685 2918 4731 2929
rect 4898 2884 4910 2940
rect 4966 2884 4978 2940
rect 5082 2940 5162 2954
rect 5082 2884 5094 2940
rect 5150 2884 5162 2940
rect 5266 2940 5346 2954
rect 5266 2884 5278 2940
rect 5334 2884 5346 2940
rect 5513 2918 5559 2929
rect 4900 2881 4911 2884
rect 4965 2881 4976 2884
rect 5084 2881 5095 2884
rect 5149 2881 5160 2884
rect 5268 2881 5279 2884
rect 5333 2881 5344 2884
rect 4823 2835 4869 2846
rect 4731 2661 4823 2835
rect 4823 2650 4869 2661
rect 5007 2835 5053 2846
rect 5007 2650 5053 2661
rect 5191 2835 5237 2846
rect 5375 2835 5421 2846
rect 5358 2808 5375 2810
rect 5421 2808 5438 2810
rect 5358 2688 5370 2808
rect 5426 2688 5438 2808
rect 5358 2686 5375 2688
rect 5191 2650 5237 2661
rect 5421 2686 5438 2688
rect 5375 2650 5421 2661
rect 4685 2433 4731 2578
rect 4900 2569 4911 2615
rect 4965 2569 4976 2615
rect 4900 2536 4976 2569
rect 5084 2569 5095 2615
rect 5149 2569 5160 2615
rect 5084 2536 5160 2569
rect 5268 2569 5279 2615
rect 5333 2569 5344 2615
rect 5268 2536 5344 2569
rect 5513 2433 5559 2578
rect 4673 2421 4753 2433
rect 4673 2365 4685 2421
rect 4741 2365 4753 2421
rect 4673 2353 4753 2365
rect 5491 2421 5569 2433
rect 5491 2365 5503 2421
rect 5559 2365 5569 2421
rect 5491 2353 5569 2365
rect 5844 2303 5924 2313
rect 4510 2247 5856 2303
rect 5912 2247 5924 2303
rect 5844 2245 5924 2247
rect 5678 2194 5748 2196
rect 4510 2193 5748 2194
rect 4510 2139 5680 2193
rect 5736 2139 5748 2193
rect 4510 2138 5748 2139
rect 4510 1117 4566 2138
rect 5678 2130 5748 2138
rect 5174 2086 5260 2090
rect 5174 2030 5186 2086
rect 5242 2030 5260 2086
rect 5174 2018 5260 2030
rect 4685 1873 4731 1884
rect 4900 1882 4976 1915
rect 4900 1836 4911 1882
rect 4965 1836 4976 1882
rect 5084 1882 5160 1915
rect 5084 1836 5095 1882
rect 5149 1836 5160 1882
rect 5268 1882 5344 1915
rect 5268 1836 5279 1882
rect 5333 1836 5344 1882
rect 5513 1873 5559 1884
rect 4823 1790 4869 1801
rect 4806 1763 4823 1765
rect 5007 1790 5053 1801
rect 4869 1763 4886 1765
rect 4731 1643 4818 1763
rect 4874 1643 4886 1763
rect 4806 1641 4823 1643
rect 4731 1343 4823 1463
rect 4869 1641 4886 1643
rect 4990 1463 5007 1465
rect 5191 1790 5237 1801
rect 5174 1763 5191 1765
rect 5375 1790 5421 1801
rect 5237 1763 5254 1765
rect 5174 1643 5186 1763
rect 5242 1643 5254 1763
rect 5174 1641 5191 1643
rect 5053 1463 5070 1465
rect 4990 1343 5002 1463
rect 5058 1343 5070 1463
rect 4990 1341 5007 1343
rect 4823 1305 4869 1316
rect 5053 1341 5070 1343
rect 5007 1305 5053 1316
rect 5237 1641 5254 1643
rect 5358 1463 5375 1465
rect 5496 1763 5513 1765
rect 5559 1763 5576 1765
rect 5496 1642 5508 1763
rect 5564 1642 5576 1763
rect 5496 1640 5513 1642
rect 5421 1463 5438 1465
rect 5358 1343 5370 1463
rect 5426 1343 5438 1463
rect 5358 1341 5375 1343
rect 5191 1305 5237 1316
rect 5421 1341 5438 1343
rect 5375 1305 5421 1316
rect 4900 1267 4911 1270
rect 4965 1267 4976 1270
rect 5084 1267 5095 1270
rect 5149 1267 5160 1270
rect 5268 1267 5279 1270
rect 5333 1267 5344 1270
rect 4685 1222 4731 1233
rect 4898 1211 4910 1267
rect 4966 1211 4978 1267
rect 4898 1197 4978 1211
rect 5082 1211 5094 1267
rect 5150 1211 5162 1267
rect 5082 1197 5162 1211
rect 5266 1211 5278 1267
rect 5334 1211 5346 1267
rect 5559 1640 5576 1642
rect 5513 1222 5559 1233
rect 5266 1197 5346 1211
rect 4898 1117 4978 1119
rect 4510 1061 4910 1117
rect 4966 1061 4978 1117
rect 4898 1059 4978 1061
rect 4090 1001 4160 1015
rect 5082 1001 5162 1003
rect 4090 945 4102 1001
rect 4158 945 5094 1001
rect 5150 945 5162 1001
rect 4090 933 4160 945
rect 5082 943 5162 945
rect 5411 1001 5491 1003
rect 5854 1001 5914 1013
rect 5411 945 5423 1001
rect 5479 945 5856 1001
rect 5912 945 5914 1001
rect 5411 943 5491 945
rect 5854 933 5914 945
rect 3954 885 4024 897
rect 5266 885 5346 887
rect 3954 829 3966 885
rect 4022 829 5278 885
rect 5334 829 5346 885
rect 3954 817 4024 829
rect 5266 827 5346 829
rect 4898 735 4978 749
rect 4685 713 4731 724
rect 4898 679 4910 735
rect 4966 679 4978 735
rect 5082 735 5162 749
rect 5082 679 5094 735
rect 5150 679 5162 735
rect 5266 735 5346 749
rect 5266 679 5278 735
rect 5334 679 5346 735
rect 5513 713 5559 724
rect 4900 676 4911 679
rect 4965 676 4976 679
rect 5084 676 5095 679
rect 5149 676 5160 679
rect 5268 676 5279 679
rect 5333 676 5344 679
rect 4823 630 4869 641
rect 4731 456 4823 630
rect 4823 445 4869 456
rect 5007 630 5053 641
rect 5007 445 5053 456
rect 5191 630 5237 641
rect 5375 630 5421 641
rect 5358 603 5375 605
rect 5421 603 5438 605
rect 5358 483 5370 603
rect 5426 483 5438 603
rect 5358 481 5375 483
rect 5191 445 5237 456
rect 5421 481 5438 483
rect 5375 445 5421 456
rect 4685 228 4731 373
rect 4900 364 4911 410
rect 4965 364 4976 410
rect 4900 331 4976 364
rect 5084 364 5095 410
rect 5149 364 5160 410
rect 5084 331 5160 364
rect 5268 364 5279 410
rect 5333 364 5344 410
rect 5268 331 5344 364
rect 5513 228 5559 373
rect 4673 216 4753 228
rect 4673 160 4685 216
rect 4741 160 4753 216
rect 4673 148 4753 160
rect 5491 216 5571 228
rect 5491 160 5503 216
rect 5559 160 5571 216
rect 5491 148 5571 160
rect -121 42 -109 98
rect -53 42 90 98
rect 146 42 2040 98
rect 3818 98 3888 110
rect 4100 98 4160 102
rect 5996 98 6052 3035
rect 6752 3033 6832 3035
rect 8268 3090 8338 3102
rect 9308 3090 9388 3092
rect 10794 3091 10874 3093
rect 8268 3034 8280 3090
rect 8336 3034 9320 3090
rect 9376 3034 9388 3090
rect 8268 3022 8338 3034
rect 6384 2941 6464 2955
rect 6171 2919 6217 2930
rect 6384 2885 6396 2941
rect 6452 2885 6464 2941
rect 6568 2941 6648 2955
rect 6568 2885 6580 2941
rect 6636 2885 6648 2941
rect 6752 2941 6832 2955
rect 6752 2885 6764 2941
rect 6820 2885 6832 2941
rect 6999 2919 7045 2930
rect 6386 2882 6397 2885
rect 6451 2882 6462 2885
rect 6570 2882 6581 2885
rect 6635 2882 6646 2885
rect 6754 2882 6765 2885
rect 6819 2882 6830 2885
rect 6309 2836 6355 2847
rect 6217 2662 6309 2836
rect 6309 2651 6355 2662
rect 6493 2836 6539 2847
rect 6493 2651 6539 2662
rect 6677 2836 6723 2847
rect 6861 2836 6907 2847
rect 6844 2809 6861 2811
rect 6907 2809 6924 2811
rect 6844 2689 6856 2809
rect 6912 2689 6924 2809
rect 6844 2687 6861 2689
rect 6677 2651 6723 2662
rect 6907 2687 6924 2689
rect 6861 2651 6907 2662
rect 6171 2434 6217 2579
rect 6386 2570 6397 2616
rect 6451 2570 6462 2616
rect 6386 2537 6462 2570
rect 6570 2570 6581 2616
rect 6635 2570 6646 2616
rect 6570 2537 6646 2570
rect 6754 2570 6765 2616
rect 6819 2570 6830 2616
rect 6754 2537 6830 2570
rect 6999 2434 7045 2579
rect 6159 2422 6239 2434
rect 6159 2366 6171 2422
rect 6227 2366 6239 2422
rect 6159 2354 6239 2366
rect 6977 2422 7055 2434
rect 6977 2366 6989 2422
rect 7045 2366 7055 2422
rect 6977 2354 7055 2366
rect 8552 2303 8608 3034
rect 9308 3032 9388 3034
rect 10038 3035 10806 3091
rect 10862 3035 10874 3091
rect 8940 2940 9020 2954
rect 8727 2918 8773 2929
rect 8940 2884 8952 2940
rect 9008 2884 9020 2940
rect 9124 2940 9204 2954
rect 9124 2884 9136 2940
rect 9192 2884 9204 2940
rect 9308 2940 9388 2954
rect 9308 2884 9320 2940
rect 9376 2884 9388 2940
rect 9555 2918 9601 2929
rect 8942 2881 8953 2884
rect 9007 2881 9018 2884
rect 9126 2881 9137 2884
rect 9191 2881 9202 2884
rect 9310 2881 9321 2884
rect 9375 2881 9386 2884
rect 8865 2835 8911 2846
rect 8773 2661 8865 2835
rect 8865 2650 8911 2661
rect 9049 2835 9095 2846
rect 9049 2650 9095 2661
rect 9233 2835 9279 2846
rect 9417 2835 9463 2846
rect 9400 2808 9417 2810
rect 9463 2808 9480 2810
rect 9400 2688 9412 2808
rect 9468 2688 9480 2808
rect 9400 2686 9417 2688
rect 9233 2650 9279 2661
rect 9463 2686 9480 2688
rect 9417 2650 9463 2661
rect 8727 2433 8773 2578
rect 8942 2569 8953 2615
rect 9007 2569 9018 2615
rect 8942 2536 9018 2569
rect 9126 2569 9137 2615
rect 9191 2569 9202 2615
rect 9126 2536 9202 2569
rect 9310 2569 9321 2615
rect 9375 2569 9386 2615
rect 9310 2536 9386 2569
rect 9555 2433 9601 2578
rect 8715 2421 8795 2433
rect 8715 2365 8727 2421
rect 8783 2365 8795 2421
rect 8715 2353 8795 2365
rect 9533 2421 9611 2433
rect 9533 2365 9545 2421
rect 9601 2365 9611 2421
rect 9533 2353 9611 2365
rect 9886 2303 9966 2313
rect 8552 2247 9898 2303
rect 9954 2247 9966 2303
rect 9886 2245 9966 2247
rect 9720 2194 9790 2196
rect 8552 2193 9790 2194
rect 8552 2139 9722 2193
rect 9778 2139 9790 2193
rect 8552 2138 9790 2139
rect 8552 1117 8608 2138
rect 9720 2130 9790 2138
rect 9216 2086 9302 2090
rect 9216 2030 9228 2086
rect 9284 2030 9302 2086
rect 9216 2018 9302 2030
rect 8727 1873 8773 1884
rect 8942 1882 9018 1915
rect 8942 1836 8953 1882
rect 9007 1836 9018 1882
rect 9126 1882 9202 1915
rect 9126 1836 9137 1882
rect 9191 1836 9202 1882
rect 9310 1882 9386 1915
rect 9310 1836 9321 1882
rect 9375 1836 9386 1882
rect 9555 1873 9601 1884
rect 8865 1790 8911 1801
rect 8848 1763 8865 1765
rect 9049 1790 9095 1801
rect 8911 1763 8928 1765
rect 8773 1643 8860 1763
rect 8916 1643 8928 1763
rect 8848 1641 8865 1643
rect 8773 1343 8865 1463
rect 8911 1641 8928 1643
rect 9032 1463 9049 1465
rect 9233 1790 9279 1801
rect 9216 1763 9233 1765
rect 9417 1790 9463 1801
rect 9279 1763 9296 1765
rect 9216 1643 9228 1763
rect 9284 1643 9296 1763
rect 9216 1641 9233 1643
rect 9095 1463 9112 1465
rect 9032 1343 9044 1463
rect 9100 1343 9112 1463
rect 9032 1341 9049 1343
rect 8865 1305 8911 1316
rect 9095 1341 9112 1343
rect 9049 1305 9095 1316
rect 9279 1641 9296 1643
rect 9400 1463 9417 1465
rect 9538 1763 9555 1765
rect 9601 1763 9618 1765
rect 9538 1642 9550 1763
rect 9606 1642 9618 1763
rect 9538 1640 9555 1642
rect 9463 1463 9480 1465
rect 9400 1343 9412 1463
rect 9468 1343 9480 1463
rect 9400 1341 9417 1343
rect 9233 1305 9279 1316
rect 9463 1341 9480 1343
rect 9417 1305 9463 1316
rect 8942 1267 8953 1270
rect 9007 1267 9018 1270
rect 9126 1267 9137 1270
rect 9191 1267 9202 1270
rect 9310 1267 9321 1270
rect 9375 1267 9386 1270
rect 8727 1222 8773 1233
rect 8940 1211 8952 1267
rect 9008 1211 9020 1267
rect 8940 1197 9020 1211
rect 9124 1211 9136 1267
rect 9192 1211 9204 1267
rect 9124 1197 9204 1211
rect 9308 1211 9320 1267
rect 9376 1211 9388 1267
rect 9601 1640 9618 1642
rect 9555 1222 9601 1233
rect 9308 1197 9388 1211
rect 8940 1117 9020 1119
rect 8552 1061 8952 1117
rect 9008 1061 9020 1117
rect 8940 1059 9020 1061
rect 8132 1001 8202 1015
rect 9124 1001 9204 1003
rect 8132 945 8144 1001
rect 8200 945 9136 1001
rect 9192 945 9204 1001
rect 8132 933 8202 945
rect 9124 943 9204 945
rect 9453 1001 9533 1003
rect 9896 1001 9956 1013
rect 9453 945 9465 1001
rect 9521 945 9898 1001
rect 9954 945 9956 1001
rect 9453 943 9533 945
rect 9896 933 9956 945
rect 7966 885 8046 897
rect 9308 885 9388 887
rect 7966 829 7978 885
rect 8034 829 9320 885
rect 9376 829 9388 885
rect 7966 817 8046 829
rect 9308 827 9388 829
rect 8940 735 9020 749
rect 8727 713 8773 724
rect 8940 679 8952 735
rect 9008 679 9020 735
rect 9124 735 9204 749
rect 9124 679 9136 735
rect 9192 679 9204 735
rect 9308 735 9388 749
rect 9308 679 9320 735
rect 9376 679 9388 735
rect 9555 713 9601 724
rect 8942 676 8953 679
rect 9007 676 9018 679
rect 9126 676 9137 679
rect 9191 676 9202 679
rect 9310 676 9321 679
rect 9375 676 9386 679
rect 8865 630 8911 641
rect 8773 456 8865 630
rect 8865 445 8911 456
rect 9049 630 9095 641
rect 9049 445 9095 456
rect 9233 630 9279 641
rect 9417 630 9463 641
rect 9400 603 9417 605
rect 9463 603 9480 605
rect 9400 483 9412 603
rect 9468 483 9480 603
rect 9400 481 9417 483
rect 9233 445 9279 456
rect 9463 481 9480 483
rect 9417 445 9463 456
rect 8727 228 8773 373
rect 8942 364 8953 410
rect 9007 364 9018 410
rect 8942 331 9018 364
rect 9126 364 9137 410
rect 9191 364 9202 410
rect 9126 331 9202 364
rect 9310 364 9321 410
rect 9375 364 9386 410
rect 9310 331 9386 364
rect 9555 228 9601 373
rect 8715 216 8795 228
rect 8715 160 8727 216
rect 8783 160 8795 216
rect 8715 148 8795 160
rect 9533 216 9613 228
rect 9533 160 9545 216
rect 9601 160 9613 216
rect 9533 148 9613 160
rect 3818 42 3830 98
rect 3886 42 4102 98
rect 4158 42 6052 98
rect 7830 98 7900 110
rect 8142 98 8202 102
rect 10038 98 10094 3035
rect 10794 3033 10874 3035
rect 12310 3090 12380 3102
rect 13350 3090 13430 3092
rect 14836 3091 14916 3093
rect 12310 3034 12322 3090
rect 12378 3034 13362 3090
rect 13418 3034 13430 3090
rect 12310 3022 12380 3034
rect 10426 2941 10506 2955
rect 10213 2919 10259 2930
rect 10426 2885 10438 2941
rect 10494 2885 10506 2941
rect 10610 2941 10690 2955
rect 10610 2885 10622 2941
rect 10678 2885 10690 2941
rect 10794 2941 10874 2955
rect 10794 2885 10806 2941
rect 10862 2885 10874 2941
rect 11041 2919 11087 2930
rect 10428 2882 10439 2885
rect 10493 2882 10504 2885
rect 10612 2882 10623 2885
rect 10677 2882 10688 2885
rect 10796 2882 10807 2885
rect 10861 2882 10872 2885
rect 10351 2836 10397 2847
rect 10259 2662 10351 2836
rect 10351 2651 10397 2662
rect 10535 2836 10581 2847
rect 10535 2651 10581 2662
rect 10719 2836 10765 2847
rect 10903 2836 10949 2847
rect 10886 2809 10903 2811
rect 10949 2809 10966 2811
rect 10886 2689 10898 2809
rect 10954 2689 10966 2809
rect 10886 2687 10903 2689
rect 10719 2651 10765 2662
rect 10949 2687 10966 2689
rect 10903 2651 10949 2662
rect 10213 2434 10259 2579
rect 10428 2570 10439 2616
rect 10493 2570 10504 2616
rect 10428 2537 10504 2570
rect 10612 2570 10623 2616
rect 10677 2570 10688 2616
rect 10612 2537 10688 2570
rect 10796 2570 10807 2616
rect 10861 2570 10872 2616
rect 10796 2537 10872 2570
rect 11041 2434 11087 2579
rect 10201 2422 10281 2434
rect 10201 2366 10213 2422
rect 10269 2366 10281 2422
rect 10201 2354 10281 2366
rect 11019 2422 11097 2434
rect 11019 2366 11031 2422
rect 11087 2366 11097 2422
rect 11019 2354 11097 2366
rect 12594 2303 12650 3034
rect 13350 3032 13430 3034
rect 14080 3035 14848 3091
rect 14904 3035 14916 3091
rect 12982 2940 13062 2954
rect 12769 2918 12815 2929
rect 12982 2884 12994 2940
rect 13050 2884 13062 2940
rect 13166 2940 13246 2954
rect 13166 2884 13178 2940
rect 13234 2884 13246 2940
rect 13350 2940 13430 2954
rect 13350 2884 13362 2940
rect 13418 2884 13430 2940
rect 13597 2918 13643 2929
rect 12984 2881 12995 2884
rect 13049 2881 13060 2884
rect 13168 2881 13179 2884
rect 13233 2881 13244 2884
rect 13352 2881 13363 2884
rect 13417 2881 13428 2884
rect 12907 2835 12953 2846
rect 12815 2661 12907 2835
rect 12907 2650 12953 2661
rect 13091 2835 13137 2846
rect 13091 2650 13137 2661
rect 13275 2835 13321 2846
rect 13459 2835 13505 2846
rect 13442 2808 13459 2810
rect 13505 2808 13522 2810
rect 13442 2688 13454 2808
rect 13510 2688 13522 2808
rect 13442 2686 13459 2688
rect 13275 2650 13321 2661
rect 13505 2686 13522 2688
rect 13459 2650 13505 2661
rect 12769 2433 12815 2578
rect 12984 2569 12995 2615
rect 13049 2569 13060 2615
rect 12984 2536 13060 2569
rect 13168 2569 13179 2615
rect 13233 2569 13244 2615
rect 13168 2536 13244 2569
rect 13352 2569 13363 2615
rect 13417 2569 13428 2615
rect 13352 2536 13428 2569
rect 13597 2433 13643 2578
rect 12757 2421 12837 2433
rect 12757 2365 12769 2421
rect 12825 2365 12837 2421
rect 12757 2353 12837 2365
rect 13575 2421 13653 2433
rect 13575 2365 13587 2421
rect 13643 2365 13653 2421
rect 13575 2353 13653 2365
rect 13928 2303 14008 2313
rect 12594 2247 13940 2303
rect 13996 2247 14008 2303
rect 13928 2245 14008 2247
rect 13762 2194 13832 2196
rect 12594 2193 13832 2194
rect 12594 2139 13764 2193
rect 13820 2139 13832 2193
rect 12594 2138 13832 2139
rect 12594 1117 12650 2138
rect 13762 2130 13832 2138
rect 13258 2086 13344 2090
rect 13258 2030 13270 2086
rect 13326 2030 13344 2086
rect 13258 2018 13344 2030
rect 12769 1873 12815 1884
rect 12984 1882 13060 1915
rect 12984 1836 12995 1882
rect 13049 1836 13060 1882
rect 13168 1882 13244 1915
rect 13168 1836 13179 1882
rect 13233 1836 13244 1882
rect 13352 1882 13428 1915
rect 13352 1836 13363 1882
rect 13417 1836 13428 1882
rect 13597 1873 13643 1884
rect 12907 1790 12953 1801
rect 12890 1763 12907 1765
rect 13091 1790 13137 1801
rect 12953 1763 12970 1765
rect 12815 1643 12902 1763
rect 12958 1643 12970 1763
rect 12890 1641 12907 1643
rect 12815 1343 12907 1463
rect 12953 1641 12970 1643
rect 13074 1463 13091 1465
rect 13275 1790 13321 1801
rect 13258 1763 13275 1765
rect 13459 1790 13505 1801
rect 13321 1763 13338 1765
rect 13258 1643 13270 1763
rect 13326 1643 13338 1763
rect 13258 1641 13275 1643
rect 13137 1463 13154 1465
rect 13074 1343 13086 1463
rect 13142 1343 13154 1463
rect 13074 1341 13091 1343
rect 12907 1305 12953 1316
rect 13137 1341 13154 1343
rect 13091 1305 13137 1316
rect 13321 1641 13338 1643
rect 13442 1463 13459 1465
rect 13580 1763 13597 1765
rect 13643 1763 13660 1765
rect 13580 1642 13592 1763
rect 13648 1642 13660 1763
rect 13580 1640 13597 1642
rect 13505 1463 13522 1465
rect 13442 1343 13454 1463
rect 13510 1343 13522 1463
rect 13442 1341 13459 1343
rect 13275 1305 13321 1316
rect 13505 1341 13522 1343
rect 13459 1305 13505 1316
rect 12984 1267 12995 1270
rect 13049 1267 13060 1270
rect 13168 1267 13179 1270
rect 13233 1267 13244 1270
rect 13352 1267 13363 1270
rect 13417 1267 13428 1270
rect 12769 1222 12815 1233
rect 12982 1211 12994 1267
rect 13050 1211 13062 1267
rect 12982 1197 13062 1211
rect 13166 1211 13178 1267
rect 13234 1211 13246 1267
rect 13166 1197 13246 1211
rect 13350 1211 13362 1267
rect 13418 1211 13430 1267
rect 13643 1640 13660 1642
rect 13597 1222 13643 1233
rect 13350 1197 13430 1211
rect 12982 1117 13062 1119
rect 12594 1061 12994 1117
rect 13050 1061 13062 1117
rect 12982 1059 13062 1061
rect 12174 1001 12244 1015
rect 13166 1001 13246 1003
rect 12174 945 12186 1001
rect 12242 945 13178 1001
rect 13234 945 13246 1001
rect 12174 933 12244 945
rect 13166 943 13246 945
rect 13495 1001 13575 1003
rect 13938 1001 13998 1013
rect 13495 945 13507 1001
rect 13563 945 13940 1001
rect 13996 945 13998 1001
rect 13495 943 13575 945
rect 13938 933 13998 945
rect 12008 885 12088 897
rect 13350 885 13430 887
rect 12008 829 12020 885
rect 12076 829 13362 885
rect 13418 829 13430 885
rect 12008 817 12088 829
rect 13350 827 13430 829
rect 12982 735 13062 749
rect 12769 713 12815 724
rect 12982 679 12994 735
rect 13050 679 13062 735
rect 13166 735 13246 749
rect 13166 679 13178 735
rect 13234 679 13246 735
rect 13350 735 13430 749
rect 13350 679 13362 735
rect 13418 679 13430 735
rect 13597 713 13643 724
rect 12984 676 12995 679
rect 13049 676 13060 679
rect 13168 676 13179 679
rect 13233 676 13244 679
rect 13352 676 13363 679
rect 13417 676 13428 679
rect 12907 630 12953 641
rect 12815 456 12907 630
rect 12907 445 12953 456
rect 13091 630 13137 641
rect 13091 445 13137 456
rect 13275 630 13321 641
rect 13459 630 13505 641
rect 13442 603 13459 605
rect 13505 603 13522 605
rect 13442 483 13454 603
rect 13510 483 13522 603
rect 13442 481 13459 483
rect 13275 445 13321 456
rect 13505 481 13522 483
rect 13459 445 13505 456
rect 12769 228 12815 373
rect 12984 364 12995 410
rect 13049 364 13060 410
rect 12984 331 13060 364
rect 13168 364 13179 410
rect 13233 364 13244 410
rect 13168 331 13244 364
rect 13352 364 13363 410
rect 13417 364 13428 410
rect 13352 331 13428 364
rect 13597 228 13643 373
rect 12757 216 12837 228
rect 12757 160 12769 216
rect 12825 160 12837 216
rect 12757 148 12837 160
rect 13575 216 13655 228
rect 13575 160 13587 216
rect 13643 160 13655 216
rect 13575 148 13655 160
rect 7830 42 7842 98
rect 7898 42 8144 98
rect 8200 42 10094 98
rect 11872 98 11942 110
rect 12184 98 12244 102
rect 14080 98 14136 3035
rect 14836 3033 14916 3035
rect 16352 3090 16422 3102
rect 17392 3090 17472 3092
rect 18878 3091 18958 3093
rect 16352 3034 16364 3090
rect 16420 3034 17404 3090
rect 17460 3034 17472 3090
rect 16352 3022 16422 3034
rect 14468 2941 14548 2955
rect 14255 2919 14301 2930
rect 14468 2885 14480 2941
rect 14536 2885 14548 2941
rect 14652 2941 14732 2955
rect 14652 2885 14664 2941
rect 14720 2885 14732 2941
rect 14836 2941 14916 2955
rect 14836 2885 14848 2941
rect 14904 2885 14916 2941
rect 15083 2919 15129 2930
rect 14470 2882 14481 2885
rect 14535 2882 14546 2885
rect 14654 2882 14665 2885
rect 14719 2882 14730 2885
rect 14838 2882 14849 2885
rect 14903 2882 14914 2885
rect 14393 2836 14439 2847
rect 14301 2662 14393 2836
rect 14393 2651 14439 2662
rect 14577 2836 14623 2847
rect 14577 2651 14623 2662
rect 14761 2836 14807 2847
rect 14945 2836 14991 2847
rect 14928 2809 14945 2811
rect 14991 2809 15008 2811
rect 14928 2689 14940 2809
rect 14996 2689 15008 2809
rect 14928 2687 14945 2689
rect 14761 2651 14807 2662
rect 14991 2687 15008 2689
rect 14945 2651 14991 2662
rect 14255 2434 14301 2579
rect 14470 2570 14481 2616
rect 14535 2570 14546 2616
rect 14470 2537 14546 2570
rect 14654 2570 14665 2616
rect 14719 2570 14730 2616
rect 14654 2537 14730 2570
rect 14838 2570 14849 2616
rect 14903 2570 14914 2616
rect 14838 2537 14914 2570
rect 15083 2434 15129 2579
rect 14243 2422 14323 2434
rect 14243 2366 14255 2422
rect 14311 2366 14323 2422
rect 14243 2354 14323 2366
rect 15061 2422 15139 2434
rect 15061 2366 15073 2422
rect 15129 2366 15139 2422
rect 15061 2354 15139 2366
rect 16636 2303 16692 3034
rect 17392 3032 17472 3034
rect 18122 3035 18890 3091
rect 18946 3035 18958 3091
rect 17024 2940 17104 2954
rect 16811 2918 16857 2929
rect 17024 2884 17036 2940
rect 17092 2884 17104 2940
rect 17208 2940 17288 2954
rect 17208 2884 17220 2940
rect 17276 2884 17288 2940
rect 17392 2940 17472 2954
rect 17392 2884 17404 2940
rect 17460 2884 17472 2940
rect 17639 2918 17685 2929
rect 17026 2881 17037 2884
rect 17091 2881 17102 2884
rect 17210 2881 17221 2884
rect 17275 2881 17286 2884
rect 17394 2881 17405 2884
rect 17459 2881 17470 2884
rect 16949 2835 16995 2846
rect 16857 2661 16949 2835
rect 16949 2650 16995 2661
rect 17133 2835 17179 2846
rect 17133 2650 17179 2661
rect 17317 2835 17363 2846
rect 17501 2835 17547 2846
rect 17484 2808 17501 2810
rect 17547 2808 17564 2810
rect 17484 2688 17496 2808
rect 17552 2688 17564 2808
rect 17484 2686 17501 2688
rect 17317 2650 17363 2661
rect 17547 2686 17564 2688
rect 17501 2650 17547 2661
rect 16811 2433 16857 2578
rect 17026 2569 17037 2615
rect 17091 2569 17102 2615
rect 17026 2536 17102 2569
rect 17210 2569 17221 2615
rect 17275 2569 17286 2615
rect 17210 2536 17286 2569
rect 17394 2569 17405 2615
rect 17459 2569 17470 2615
rect 17394 2536 17470 2569
rect 17639 2433 17685 2578
rect 16799 2421 16879 2433
rect 16799 2365 16811 2421
rect 16867 2365 16879 2421
rect 16799 2353 16879 2365
rect 17617 2421 17695 2433
rect 17617 2365 17629 2421
rect 17685 2365 17695 2421
rect 17617 2353 17695 2365
rect 17970 2303 18050 2313
rect 16636 2247 17982 2303
rect 18038 2247 18050 2303
rect 17970 2245 18050 2247
rect 17804 2194 17874 2196
rect 16636 2193 17874 2194
rect 16636 2139 17806 2193
rect 17862 2139 17874 2193
rect 16636 2138 17874 2139
rect 16636 1117 16692 2138
rect 17804 2130 17874 2138
rect 17300 2086 17386 2090
rect 17300 2030 17312 2086
rect 17368 2030 17386 2086
rect 17300 2018 17386 2030
rect 16811 1873 16857 1884
rect 17026 1882 17102 1915
rect 17026 1836 17037 1882
rect 17091 1836 17102 1882
rect 17210 1882 17286 1915
rect 17210 1836 17221 1882
rect 17275 1836 17286 1882
rect 17394 1882 17470 1915
rect 17394 1836 17405 1882
rect 17459 1836 17470 1882
rect 17639 1873 17685 1884
rect 16949 1790 16995 1801
rect 16932 1763 16949 1765
rect 17133 1790 17179 1801
rect 16995 1763 17012 1765
rect 16857 1643 16944 1763
rect 17000 1643 17012 1763
rect 16932 1641 16949 1643
rect 16857 1343 16949 1463
rect 16995 1641 17012 1643
rect 17116 1463 17133 1465
rect 17317 1790 17363 1801
rect 17300 1763 17317 1765
rect 17501 1790 17547 1801
rect 17363 1763 17380 1765
rect 17300 1643 17312 1763
rect 17368 1643 17380 1763
rect 17300 1641 17317 1643
rect 17179 1463 17196 1465
rect 17116 1343 17128 1463
rect 17184 1343 17196 1463
rect 17116 1341 17133 1343
rect 16949 1305 16995 1316
rect 17179 1341 17196 1343
rect 17133 1305 17179 1316
rect 17363 1641 17380 1643
rect 17484 1463 17501 1465
rect 17622 1763 17639 1765
rect 17685 1763 17702 1765
rect 17622 1642 17634 1763
rect 17690 1642 17702 1763
rect 17622 1640 17639 1642
rect 17547 1463 17564 1465
rect 17484 1343 17496 1463
rect 17552 1343 17564 1463
rect 17484 1341 17501 1343
rect 17317 1305 17363 1316
rect 17547 1341 17564 1343
rect 17501 1305 17547 1316
rect 17026 1267 17037 1270
rect 17091 1267 17102 1270
rect 17210 1267 17221 1270
rect 17275 1267 17286 1270
rect 17394 1267 17405 1270
rect 17459 1267 17470 1270
rect 16811 1222 16857 1233
rect 17024 1211 17036 1267
rect 17092 1211 17104 1267
rect 17024 1197 17104 1211
rect 17208 1211 17220 1267
rect 17276 1211 17288 1267
rect 17208 1197 17288 1211
rect 17392 1211 17404 1267
rect 17460 1211 17472 1267
rect 17685 1640 17702 1642
rect 17639 1222 17685 1233
rect 17392 1197 17472 1211
rect 17024 1117 17104 1119
rect 16636 1061 17036 1117
rect 17092 1061 17104 1117
rect 17024 1059 17104 1061
rect 16216 1001 16286 1015
rect 17208 1001 17288 1003
rect 16216 945 16228 1001
rect 16284 945 17220 1001
rect 17276 945 17288 1001
rect 16216 933 16286 945
rect 17208 943 17288 945
rect 17537 1001 17617 1003
rect 17980 1001 18040 1013
rect 17537 945 17549 1001
rect 17605 945 17982 1001
rect 18038 945 18040 1001
rect 17537 943 17617 945
rect 17980 933 18040 945
rect 16050 885 16130 897
rect 17392 885 17472 887
rect 16050 829 16062 885
rect 16118 829 17404 885
rect 17460 829 17472 885
rect 16050 817 16130 829
rect 17392 827 17472 829
rect 17024 735 17104 749
rect 16811 713 16857 724
rect 17024 679 17036 735
rect 17092 679 17104 735
rect 17208 735 17288 749
rect 17208 679 17220 735
rect 17276 679 17288 735
rect 17392 735 17472 749
rect 17392 679 17404 735
rect 17460 679 17472 735
rect 17639 713 17685 724
rect 17026 676 17037 679
rect 17091 676 17102 679
rect 17210 676 17221 679
rect 17275 676 17286 679
rect 17394 676 17405 679
rect 17459 676 17470 679
rect 16949 630 16995 641
rect 16857 456 16949 630
rect 16949 445 16995 456
rect 17133 630 17179 641
rect 17133 445 17179 456
rect 17317 630 17363 641
rect 17501 630 17547 641
rect 17484 603 17501 605
rect 17547 603 17564 605
rect 17484 483 17496 603
rect 17552 483 17564 603
rect 17484 481 17501 483
rect 17317 445 17363 456
rect 17547 481 17564 483
rect 17501 445 17547 456
rect 16811 228 16857 373
rect 17026 364 17037 410
rect 17091 364 17102 410
rect 17026 331 17102 364
rect 17210 364 17221 410
rect 17275 364 17286 410
rect 17210 331 17286 364
rect 17394 364 17405 410
rect 17459 364 17470 410
rect 17394 331 17470 364
rect 17639 228 17685 373
rect 16799 216 16879 228
rect 16799 160 16811 216
rect 16867 160 16879 216
rect 16799 148 16879 160
rect 17617 216 17697 228
rect 17617 160 17629 216
rect 17685 160 17697 216
rect 17617 148 17697 160
rect 11872 42 11884 98
rect 11940 42 12186 98
rect 12242 42 14136 98
rect 15914 98 15984 110
rect 16226 98 16286 102
rect 18122 98 18178 3035
rect 18878 3033 18958 3035
rect 20394 3090 20464 3102
rect 21434 3090 21514 3092
rect 22920 3091 23000 3093
rect 20394 3034 20406 3090
rect 20462 3034 21446 3090
rect 21502 3034 21514 3090
rect 20394 3022 20464 3034
rect 18510 2941 18590 2955
rect 18297 2919 18343 2930
rect 18510 2885 18522 2941
rect 18578 2885 18590 2941
rect 18694 2941 18774 2955
rect 18694 2885 18706 2941
rect 18762 2885 18774 2941
rect 18878 2941 18958 2955
rect 18878 2885 18890 2941
rect 18946 2885 18958 2941
rect 19125 2919 19171 2930
rect 18512 2882 18523 2885
rect 18577 2882 18588 2885
rect 18696 2882 18707 2885
rect 18761 2882 18772 2885
rect 18880 2882 18891 2885
rect 18945 2882 18956 2885
rect 18435 2836 18481 2847
rect 18343 2662 18435 2836
rect 18435 2651 18481 2662
rect 18619 2836 18665 2847
rect 18619 2651 18665 2662
rect 18803 2836 18849 2847
rect 18987 2836 19033 2847
rect 18970 2809 18987 2811
rect 19033 2809 19050 2811
rect 18970 2689 18982 2809
rect 19038 2689 19050 2809
rect 18970 2687 18987 2689
rect 18803 2651 18849 2662
rect 19033 2687 19050 2689
rect 18987 2651 19033 2662
rect 18297 2434 18343 2579
rect 18512 2570 18523 2616
rect 18577 2570 18588 2616
rect 18512 2537 18588 2570
rect 18696 2570 18707 2616
rect 18761 2570 18772 2616
rect 18696 2537 18772 2570
rect 18880 2570 18891 2616
rect 18945 2570 18956 2616
rect 18880 2537 18956 2570
rect 19125 2434 19171 2579
rect 18285 2422 18365 2434
rect 18285 2366 18297 2422
rect 18353 2366 18365 2422
rect 18285 2354 18365 2366
rect 19103 2422 19181 2434
rect 19103 2366 19115 2422
rect 19171 2366 19181 2422
rect 19103 2354 19181 2366
rect 20678 2303 20734 3034
rect 21434 3032 21514 3034
rect 22164 3035 22932 3091
rect 22988 3035 23000 3091
rect 21066 2940 21146 2954
rect 20853 2918 20899 2929
rect 21066 2884 21078 2940
rect 21134 2884 21146 2940
rect 21250 2940 21330 2954
rect 21250 2884 21262 2940
rect 21318 2884 21330 2940
rect 21434 2940 21514 2954
rect 21434 2884 21446 2940
rect 21502 2884 21514 2940
rect 21681 2918 21727 2929
rect 21068 2881 21079 2884
rect 21133 2881 21144 2884
rect 21252 2881 21263 2884
rect 21317 2881 21328 2884
rect 21436 2881 21447 2884
rect 21501 2881 21512 2884
rect 20991 2835 21037 2846
rect 20899 2661 20991 2835
rect 20991 2650 21037 2661
rect 21175 2835 21221 2846
rect 21175 2650 21221 2661
rect 21359 2835 21405 2846
rect 21543 2835 21589 2846
rect 21526 2808 21543 2810
rect 21589 2808 21606 2810
rect 21526 2688 21538 2808
rect 21594 2688 21606 2808
rect 21526 2686 21543 2688
rect 21359 2650 21405 2661
rect 21589 2686 21606 2688
rect 21543 2650 21589 2661
rect 20853 2433 20899 2578
rect 21068 2569 21079 2615
rect 21133 2569 21144 2615
rect 21068 2536 21144 2569
rect 21252 2569 21263 2615
rect 21317 2569 21328 2615
rect 21252 2536 21328 2569
rect 21436 2569 21447 2615
rect 21501 2569 21512 2615
rect 21436 2536 21512 2569
rect 21681 2433 21727 2578
rect 20841 2421 20921 2433
rect 20841 2365 20853 2421
rect 20909 2365 20921 2421
rect 20841 2353 20921 2365
rect 21659 2421 21737 2433
rect 21659 2365 21671 2421
rect 21727 2365 21737 2421
rect 21659 2353 21737 2365
rect 22012 2303 22092 2313
rect 20678 2247 22024 2303
rect 22080 2247 22092 2303
rect 22012 2245 22092 2247
rect 21846 2194 21916 2196
rect 20678 2193 21916 2194
rect 20678 2139 21848 2193
rect 21904 2139 21916 2193
rect 20678 2138 21916 2139
rect 20678 1117 20734 2138
rect 21846 2130 21916 2138
rect 21342 2086 21428 2090
rect 21342 2030 21354 2086
rect 21410 2030 21428 2086
rect 21342 2018 21428 2030
rect 20853 1873 20899 1884
rect 21068 1882 21144 1915
rect 21068 1836 21079 1882
rect 21133 1836 21144 1882
rect 21252 1882 21328 1915
rect 21252 1836 21263 1882
rect 21317 1836 21328 1882
rect 21436 1882 21512 1915
rect 21436 1836 21447 1882
rect 21501 1836 21512 1882
rect 21681 1873 21727 1884
rect 20991 1790 21037 1801
rect 20974 1763 20991 1765
rect 21175 1790 21221 1801
rect 21037 1763 21054 1765
rect 20899 1643 20986 1763
rect 21042 1643 21054 1763
rect 20974 1641 20991 1643
rect 20899 1343 20991 1463
rect 21037 1641 21054 1643
rect 21158 1463 21175 1465
rect 21359 1790 21405 1801
rect 21342 1763 21359 1765
rect 21543 1790 21589 1801
rect 21405 1763 21422 1765
rect 21342 1643 21354 1763
rect 21410 1643 21422 1763
rect 21342 1641 21359 1643
rect 21221 1463 21238 1465
rect 21158 1343 21170 1463
rect 21226 1343 21238 1463
rect 21158 1341 21175 1343
rect 20991 1305 21037 1316
rect 21221 1341 21238 1343
rect 21175 1305 21221 1316
rect 21405 1641 21422 1643
rect 21526 1463 21543 1465
rect 21664 1763 21681 1765
rect 21727 1763 21744 1765
rect 21664 1642 21676 1763
rect 21732 1642 21744 1763
rect 21664 1640 21681 1642
rect 21589 1463 21606 1465
rect 21526 1343 21538 1463
rect 21594 1343 21606 1463
rect 21526 1341 21543 1343
rect 21359 1305 21405 1316
rect 21589 1341 21606 1343
rect 21543 1305 21589 1316
rect 21068 1267 21079 1270
rect 21133 1267 21144 1270
rect 21252 1267 21263 1270
rect 21317 1267 21328 1270
rect 21436 1267 21447 1270
rect 21501 1267 21512 1270
rect 20853 1222 20899 1233
rect 21066 1211 21078 1267
rect 21134 1211 21146 1267
rect 21066 1197 21146 1211
rect 21250 1211 21262 1267
rect 21318 1211 21330 1267
rect 21250 1197 21330 1211
rect 21434 1211 21446 1267
rect 21502 1211 21514 1267
rect 21727 1640 21744 1642
rect 21681 1222 21727 1233
rect 21434 1197 21514 1211
rect 21066 1117 21146 1119
rect 20678 1061 21078 1117
rect 21134 1061 21146 1117
rect 21066 1059 21146 1061
rect 20258 1001 20328 1015
rect 21250 1001 21330 1003
rect 20258 945 20270 1001
rect 20326 945 21262 1001
rect 21318 945 21330 1001
rect 20258 933 20328 945
rect 21250 943 21330 945
rect 21579 1001 21659 1003
rect 22022 1001 22082 1013
rect 21579 945 21591 1001
rect 21647 945 22024 1001
rect 22080 945 22082 1001
rect 21579 943 21659 945
rect 22022 933 22082 945
rect 20092 885 20172 897
rect 21434 885 21514 887
rect 20092 829 20104 885
rect 20160 829 21446 885
rect 21502 829 21514 885
rect 20092 817 20172 829
rect 21434 827 21514 829
rect 21066 735 21146 749
rect 20853 713 20899 724
rect 21066 679 21078 735
rect 21134 679 21146 735
rect 21250 735 21330 749
rect 21250 679 21262 735
rect 21318 679 21330 735
rect 21434 735 21514 749
rect 21434 679 21446 735
rect 21502 679 21514 735
rect 21681 713 21727 724
rect 21068 676 21079 679
rect 21133 676 21144 679
rect 21252 676 21263 679
rect 21317 676 21328 679
rect 21436 676 21447 679
rect 21501 676 21512 679
rect 20991 630 21037 641
rect 20899 456 20991 630
rect 20991 445 21037 456
rect 21175 630 21221 641
rect 21175 445 21221 456
rect 21359 630 21405 641
rect 21543 630 21589 641
rect 21526 603 21543 605
rect 21589 603 21606 605
rect 21526 483 21538 603
rect 21594 483 21606 603
rect 21526 481 21543 483
rect 21359 445 21405 456
rect 21589 481 21606 483
rect 21543 445 21589 456
rect 20853 228 20899 373
rect 21068 364 21079 410
rect 21133 364 21144 410
rect 21068 331 21144 364
rect 21252 364 21263 410
rect 21317 364 21328 410
rect 21252 331 21328 364
rect 21436 364 21447 410
rect 21501 364 21512 410
rect 21436 331 21512 364
rect 21681 228 21727 373
rect 20841 216 20921 228
rect 20841 160 20853 216
rect 20909 160 20921 216
rect 20841 148 20921 160
rect 21659 216 21739 228
rect 21659 160 21671 216
rect 21727 160 21739 216
rect 21659 148 21739 160
rect 15914 42 15926 98
rect 15982 42 16228 98
rect 16284 42 18178 98
rect 19956 98 20026 110
rect 20268 98 20328 102
rect 22164 98 22220 3035
rect 22920 3033 23000 3035
rect 24436 3090 24506 3102
rect 25476 3090 25556 3092
rect 26962 3091 27042 3093
rect 24436 3034 24448 3090
rect 24504 3034 25488 3090
rect 25544 3034 25556 3090
rect 24436 3022 24506 3034
rect 22552 2941 22632 2955
rect 22339 2919 22385 2930
rect 22552 2885 22564 2941
rect 22620 2885 22632 2941
rect 22736 2941 22816 2955
rect 22736 2885 22748 2941
rect 22804 2885 22816 2941
rect 22920 2941 23000 2955
rect 22920 2885 22932 2941
rect 22988 2885 23000 2941
rect 23167 2919 23213 2930
rect 22554 2882 22565 2885
rect 22619 2882 22630 2885
rect 22738 2882 22749 2885
rect 22803 2882 22814 2885
rect 22922 2882 22933 2885
rect 22987 2882 22998 2885
rect 22477 2836 22523 2847
rect 22385 2662 22477 2836
rect 22477 2651 22523 2662
rect 22661 2836 22707 2847
rect 22661 2651 22707 2662
rect 22845 2836 22891 2847
rect 23029 2836 23075 2847
rect 23012 2809 23029 2811
rect 23075 2809 23092 2811
rect 23012 2689 23024 2809
rect 23080 2689 23092 2809
rect 23012 2687 23029 2689
rect 22845 2651 22891 2662
rect 23075 2687 23092 2689
rect 23029 2651 23075 2662
rect 22339 2434 22385 2579
rect 22554 2570 22565 2616
rect 22619 2570 22630 2616
rect 22554 2537 22630 2570
rect 22738 2570 22749 2616
rect 22803 2570 22814 2616
rect 22738 2537 22814 2570
rect 22922 2570 22933 2616
rect 22987 2570 22998 2616
rect 22922 2537 22998 2570
rect 23167 2434 23213 2579
rect 22327 2422 22407 2434
rect 22327 2366 22339 2422
rect 22395 2366 22407 2422
rect 22327 2354 22407 2366
rect 23145 2422 23223 2434
rect 23145 2366 23157 2422
rect 23213 2366 23223 2422
rect 23145 2354 23223 2366
rect 24720 2303 24776 3034
rect 25476 3032 25556 3034
rect 26206 3035 26974 3091
rect 27030 3035 27042 3091
rect 25108 2940 25188 2954
rect 24895 2918 24941 2929
rect 25108 2884 25120 2940
rect 25176 2884 25188 2940
rect 25292 2940 25372 2954
rect 25292 2884 25304 2940
rect 25360 2884 25372 2940
rect 25476 2940 25556 2954
rect 25476 2884 25488 2940
rect 25544 2884 25556 2940
rect 25723 2918 25769 2929
rect 25110 2881 25121 2884
rect 25175 2881 25186 2884
rect 25294 2881 25305 2884
rect 25359 2881 25370 2884
rect 25478 2881 25489 2884
rect 25543 2881 25554 2884
rect 25033 2835 25079 2846
rect 24941 2661 25033 2835
rect 25033 2650 25079 2661
rect 25217 2835 25263 2846
rect 25217 2650 25263 2661
rect 25401 2835 25447 2846
rect 25585 2835 25631 2846
rect 25568 2808 25585 2810
rect 25631 2808 25648 2810
rect 25568 2688 25580 2808
rect 25636 2688 25648 2808
rect 25568 2686 25585 2688
rect 25401 2650 25447 2661
rect 25631 2686 25648 2688
rect 25585 2650 25631 2661
rect 24895 2433 24941 2578
rect 25110 2569 25121 2615
rect 25175 2569 25186 2615
rect 25110 2536 25186 2569
rect 25294 2569 25305 2615
rect 25359 2569 25370 2615
rect 25294 2536 25370 2569
rect 25478 2569 25489 2615
rect 25543 2569 25554 2615
rect 25478 2536 25554 2569
rect 25723 2433 25769 2578
rect 24883 2421 24963 2433
rect 24883 2365 24895 2421
rect 24951 2365 24963 2421
rect 24883 2353 24963 2365
rect 25701 2421 25779 2433
rect 25701 2365 25713 2421
rect 25769 2365 25779 2421
rect 25701 2353 25779 2365
rect 26054 2303 26134 2313
rect 24720 2247 26066 2303
rect 26122 2247 26134 2303
rect 26054 2245 26134 2247
rect 25888 2194 25958 2196
rect 24720 2193 25958 2194
rect 24720 2139 25890 2193
rect 25946 2139 25958 2193
rect 24720 2138 25958 2139
rect 24720 1117 24776 2138
rect 25888 2130 25958 2138
rect 25384 2086 25470 2090
rect 25384 2030 25396 2086
rect 25452 2030 25470 2086
rect 25384 2018 25470 2030
rect 24895 1873 24941 1884
rect 25110 1882 25186 1915
rect 25110 1836 25121 1882
rect 25175 1836 25186 1882
rect 25294 1882 25370 1915
rect 25294 1836 25305 1882
rect 25359 1836 25370 1882
rect 25478 1882 25554 1915
rect 25478 1836 25489 1882
rect 25543 1836 25554 1882
rect 25723 1873 25769 1884
rect 25033 1790 25079 1801
rect 25016 1763 25033 1765
rect 25217 1790 25263 1801
rect 25079 1763 25096 1765
rect 24941 1643 25028 1763
rect 25084 1643 25096 1763
rect 25016 1641 25033 1643
rect 24941 1343 25033 1463
rect 25079 1641 25096 1643
rect 25200 1463 25217 1465
rect 25401 1790 25447 1801
rect 25384 1763 25401 1765
rect 25585 1790 25631 1801
rect 25447 1763 25464 1765
rect 25384 1643 25396 1763
rect 25452 1643 25464 1763
rect 25384 1641 25401 1643
rect 25263 1463 25280 1465
rect 25200 1343 25212 1463
rect 25268 1343 25280 1463
rect 25200 1341 25217 1343
rect 25033 1305 25079 1316
rect 25263 1341 25280 1343
rect 25217 1305 25263 1316
rect 25447 1641 25464 1643
rect 25568 1463 25585 1465
rect 25706 1763 25723 1765
rect 25769 1763 25786 1765
rect 25706 1642 25718 1763
rect 25774 1642 25786 1763
rect 25706 1640 25723 1642
rect 25631 1463 25648 1465
rect 25568 1343 25580 1463
rect 25636 1343 25648 1463
rect 25568 1341 25585 1343
rect 25401 1305 25447 1316
rect 25631 1341 25648 1343
rect 25585 1305 25631 1316
rect 25110 1267 25121 1270
rect 25175 1267 25186 1270
rect 25294 1267 25305 1270
rect 25359 1267 25370 1270
rect 25478 1267 25489 1270
rect 25543 1267 25554 1270
rect 24895 1222 24941 1233
rect 25108 1211 25120 1267
rect 25176 1211 25188 1267
rect 25108 1197 25188 1211
rect 25292 1211 25304 1267
rect 25360 1211 25372 1267
rect 25292 1197 25372 1211
rect 25476 1211 25488 1267
rect 25544 1211 25556 1267
rect 25769 1640 25786 1642
rect 25723 1222 25769 1233
rect 25476 1197 25556 1211
rect 25108 1117 25188 1119
rect 24720 1061 25120 1117
rect 25176 1061 25188 1117
rect 25108 1059 25188 1061
rect 24300 1001 24370 1015
rect 25292 1001 25372 1003
rect 24300 945 24312 1001
rect 24368 945 25304 1001
rect 25360 945 25372 1001
rect 24300 933 24370 945
rect 25292 943 25372 945
rect 25621 1001 25701 1003
rect 26064 1001 26124 1013
rect 25621 945 25633 1001
rect 25689 945 26066 1001
rect 26122 945 26124 1001
rect 25621 943 25701 945
rect 26064 933 26124 945
rect 24134 885 24214 897
rect 25476 885 25556 887
rect 24134 829 24146 885
rect 24202 829 25488 885
rect 25544 829 25556 885
rect 24134 817 24214 829
rect 25476 827 25556 829
rect 25108 735 25188 749
rect 24895 713 24941 724
rect 25108 679 25120 735
rect 25176 679 25188 735
rect 25292 735 25372 749
rect 25292 679 25304 735
rect 25360 679 25372 735
rect 25476 735 25556 749
rect 25476 679 25488 735
rect 25544 679 25556 735
rect 25723 713 25769 724
rect 25110 676 25121 679
rect 25175 676 25186 679
rect 25294 676 25305 679
rect 25359 676 25370 679
rect 25478 676 25489 679
rect 25543 676 25554 679
rect 25033 630 25079 641
rect 24941 456 25033 630
rect 25033 445 25079 456
rect 25217 630 25263 641
rect 25217 445 25263 456
rect 25401 630 25447 641
rect 25585 630 25631 641
rect 25568 603 25585 605
rect 25631 603 25648 605
rect 25568 483 25580 603
rect 25636 483 25648 603
rect 25568 481 25585 483
rect 25401 445 25447 456
rect 25631 481 25648 483
rect 25585 445 25631 456
rect 24895 228 24941 373
rect 25110 364 25121 410
rect 25175 364 25186 410
rect 25110 331 25186 364
rect 25294 364 25305 410
rect 25359 364 25370 410
rect 25294 331 25370 364
rect 25478 364 25489 410
rect 25543 364 25554 410
rect 25478 331 25554 364
rect 25723 228 25769 373
rect 24883 216 24963 228
rect 24883 160 24895 216
rect 24951 160 24963 216
rect 24883 148 24963 160
rect 25701 216 25781 228
rect 25701 160 25713 216
rect 25769 160 25781 216
rect 25701 148 25781 160
rect 19956 42 19968 98
rect 20024 42 20270 98
rect 20326 42 22220 98
rect 23998 98 24068 110
rect 24310 98 24370 102
rect 26206 98 26262 3035
rect 26962 3033 27042 3035
rect 26594 2941 26674 2955
rect 26381 2919 26427 2930
rect 26594 2885 26606 2941
rect 26662 2885 26674 2941
rect 26778 2941 26858 2955
rect 26778 2885 26790 2941
rect 26846 2885 26858 2941
rect 26962 2941 27042 2955
rect 26962 2885 26974 2941
rect 27030 2885 27042 2941
rect 27209 2919 27255 2930
rect 26596 2882 26607 2885
rect 26661 2882 26672 2885
rect 26780 2882 26791 2885
rect 26845 2882 26856 2885
rect 26964 2882 26975 2885
rect 27029 2882 27040 2885
rect 26519 2836 26565 2847
rect 26427 2662 26519 2836
rect 26519 2651 26565 2662
rect 26703 2836 26749 2847
rect 26703 2651 26749 2662
rect 26887 2836 26933 2847
rect 27071 2836 27117 2847
rect 27054 2809 27071 2811
rect 27117 2809 27134 2811
rect 27054 2689 27066 2809
rect 27122 2689 27134 2809
rect 27054 2687 27071 2689
rect 26887 2651 26933 2662
rect 27117 2687 27134 2689
rect 27071 2651 27117 2662
rect 26381 2434 26427 2579
rect 26596 2570 26607 2616
rect 26661 2570 26672 2616
rect 26596 2537 26672 2570
rect 26780 2570 26791 2616
rect 26845 2570 26856 2616
rect 26780 2537 26856 2570
rect 26964 2570 26975 2616
rect 27029 2570 27040 2616
rect 26964 2537 27040 2570
rect 27209 2434 27255 2579
rect 26369 2422 26449 2434
rect 26369 2366 26381 2422
rect 26437 2366 26449 2422
rect 26369 2354 26449 2366
rect 27187 2422 27265 2434
rect 27187 2366 27199 2422
rect 27255 2366 27265 2422
rect 27187 2354 27265 2366
rect 23998 42 24010 98
rect 24066 42 24312 98
rect 24368 42 26262 98
rect -121 30 -35 42
rect 88 30 148 42
rect 3818 30 3888 42
rect 4100 30 4160 42
rect 7830 30 7900 42
rect 8142 30 8202 42
rect 11872 30 11942 42
rect 12184 30 12244 42
rect 15914 30 15984 42
rect 16226 30 16286 42
rect 19956 30 20026 42
rect 20268 30 20328 42
rect 23998 30 24068 42
rect 24310 30 24370 42
<< via1 >>
rect 12050 19033 12106 19089
rect 19898 19033 19954 19089
rect 16092 18857 16148 18913
rect 23940 18857 23996 18913
rect 3912 18681 3968 18737
rect 11760 18681 11816 18737
rect 20134 18681 20190 18737
rect 27982 18681 28038 18737
rect 8008 18505 8064 18561
rect 15856 18505 15912 18561
rect 24176 18505 24232 18561
rect 32024 18505 32080 18561
rect 5186 18224 5242 18280
rect 4818 17837 4823 17957
rect 4823 17837 4869 17957
rect 4869 17837 4874 17957
rect 5186 17837 5191 17957
rect 5191 17837 5237 17957
rect 5237 17837 5242 17957
rect 5002 17537 5007 17657
rect 5007 17537 5053 17657
rect 5053 17537 5058 17657
rect 5508 17836 5513 17957
rect 5513 17836 5559 17957
rect 5559 17836 5564 17957
rect 5370 17537 5375 17657
rect 5375 17537 5421 17657
rect 5421 17537 5426 17657
rect 4910 17418 4911 17461
rect 4911 17418 4965 17461
rect 4965 17418 4966 17461
rect 4910 17405 4966 17418
rect 5094 17418 5095 17461
rect 5095 17418 5149 17461
rect 5149 17418 5150 17461
rect 5094 17405 5150 17418
rect 5278 17418 5279 17461
rect 5279 17418 5333 17461
rect 5333 17418 5334 17461
rect 5278 17405 5334 17418
rect 3558 17255 3614 17311
rect 4910 17255 4966 17311
rect 4238 17139 4294 17195
rect 5094 17139 5150 17195
rect 5423 17139 5479 17195
rect 5680 17139 5736 17195
rect 5278 17023 5334 17079
rect 4910 16916 4966 16929
rect 4910 16873 4911 16916
rect 4911 16873 4965 16916
rect 4965 16873 4966 16916
rect 5094 16916 5150 16929
rect 5094 16873 5095 16916
rect 5095 16873 5149 16916
rect 5149 16873 5150 16916
rect 5278 16916 5334 16929
rect 5278 16873 5279 16916
rect 5279 16873 5333 16916
rect 5333 16873 5334 16916
rect 5370 16677 5375 16797
rect 5375 16677 5421 16797
rect 5421 16677 5426 16797
rect 4685 16354 4741 16410
rect 5503 16354 5559 16410
rect 5856 16236 5912 16292
rect 5680 16128 5736 16182
rect 5186 16019 5242 16075
rect 4818 15632 4823 15752
rect 4823 15632 4869 15752
rect 4869 15632 4874 15752
rect 5186 15632 5191 15752
rect 5191 15632 5237 15752
rect 5237 15632 5242 15752
rect 5002 15332 5007 15452
rect 5007 15332 5053 15452
rect 5053 15332 5058 15452
rect 5508 15631 5513 15752
rect 5513 15631 5559 15752
rect 5559 15631 5564 15752
rect 5370 15332 5375 15452
rect 5375 15332 5421 15452
rect 5421 15332 5426 15452
rect 4910 15213 4911 15256
rect 4911 15213 4965 15256
rect 4965 15213 4966 15256
rect 4910 15200 4966 15213
rect 5094 15213 5095 15256
rect 5095 15213 5149 15256
rect 5149 15213 5150 15256
rect 5094 15200 5150 15213
rect 5278 15213 5279 15256
rect 5279 15213 5333 15256
rect 5333 15213 5334 15256
rect 5278 15200 5334 15213
rect 4910 15050 4966 15106
rect 9228 18221 9284 18277
rect 8860 17834 8865 17954
rect 8865 17834 8911 17954
rect 8911 17834 8916 17954
rect 9228 17834 9233 17954
rect 9233 17834 9279 17954
rect 9279 17834 9284 17954
rect 9044 17534 9049 17654
rect 9049 17534 9095 17654
rect 9095 17534 9100 17654
rect 9550 17833 9555 17954
rect 9555 17833 9601 17954
rect 9601 17833 9606 17954
rect 9412 17534 9417 17654
rect 9417 17534 9463 17654
rect 9463 17534 9468 17654
rect 8952 17415 8953 17458
rect 8953 17415 9007 17458
rect 9007 17415 9008 17458
rect 8952 17402 9008 17415
rect 9136 17415 9137 17458
rect 9137 17415 9191 17458
rect 9191 17415 9192 17458
rect 9136 17402 9192 17415
rect 9320 17415 9321 17458
rect 9321 17415 9375 17458
rect 9375 17415 9376 17458
rect 9320 17402 9376 17415
rect 7570 17252 7626 17308
rect 8952 17252 9008 17308
rect 8280 17136 8336 17192
rect 9136 17136 9192 17192
rect 9465 17136 9521 17192
rect 9722 17136 9778 17192
rect 9320 17020 9376 17076
rect 8952 16913 9008 16926
rect 8952 16870 8953 16913
rect 8953 16870 9007 16913
rect 9007 16870 9008 16913
rect 9136 16913 9192 16926
rect 9136 16870 9137 16913
rect 9137 16870 9191 16913
rect 9191 16870 9192 16913
rect 9320 16913 9376 16926
rect 9320 16870 9321 16913
rect 9321 16870 9375 16913
rect 9375 16870 9376 16913
rect 9412 16674 9417 16794
rect 9417 16674 9463 16794
rect 9463 16674 9468 16794
rect 8727 16351 8783 16407
rect 9545 16351 9601 16407
rect 9898 16233 9954 16289
rect 9722 16125 9778 16179
rect 6672 16019 6728 16075
rect 6304 15632 6309 15752
rect 6309 15632 6355 15752
rect 6355 15632 6360 15752
rect 6672 15632 6677 15752
rect 6677 15632 6723 15752
rect 6723 15632 6728 15752
rect 6488 15332 6493 15452
rect 6493 15332 6539 15452
rect 6539 15332 6544 15452
rect 6994 15631 6999 15752
rect 6999 15631 7045 15752
rect 7045 15631 7050 15752
rect 6856 15332 6861 15452
rect 6861 15332 6907 15452
rect 6907 15332 6912 15452
rect 6396 15213 6397 15256
rect 6397 15213 6451 15256
rect 6451 15213 6452 15256
rect 6396 15200 6452 15213
rect 6580 15213 6581 15256
rect 6581 15213 6635 15256
rect 6635 15213 6636 15256
rect 6580 15200 6636 15213
rect 6764 15213 6765 15256
rect 6765 15213 6819 15256
rect 6819 15213 6820 15256
rect 6764 15200 6820 15213
rect 6396 15050 6452 15106
rect 9228 16016 9284 16072
rect 8860 15629 8865 15749
rect 8865 15629 8911 15749
rect 8911 15629 8916 15749
rect 9228 15629 9233 15749
rect 9233 15629 9279 15749
rect 9279 15629 9284 15749
rect 9044 15329 9049 15449
rect 9049 15329 9095 15449
rect 9095 15329 9100 15449
rect 9550 15628 9555 15749
rect 9555 15628 9601 15749
rect 9601 15628 9606 15749
rect 9412 15329 9417 15449
rect 9417 15329 9463 15449
rect 9463 15329 9468 15449
rect 8952 15210 8953 15253
rect 8953 15210 9007 15253
rect 9007 15210 9008 15253
rect 8952 15197 9008 15210
rect 9136 15210 9137 15253
rect 9137 15210 9191 15253
rect 9191 15210 9192 15253
rect 9136 15197 9192 15210
rect 9320 15210 9321 15253
rect 9321 15210 9375 15253
rect 9375 15210 9376 15253
rect 9320 15197 9376 15210
rect 8952 15047 9008 15103
rect 13270 18221 13326 18277
rect 12902 17834 12907 17954
rect 12907 17834 12953 17954
rect 12953 17834 12958 17954
rect 13270 17834 13275 17954
rect 13275 17834 13321 17954
rect 13321 17834 13326 17954
rect 13086 17534 13091 17654
rect 13091 17534 13137 17654
rect 13137 17534 13142 17654
rect 13592 17833 13597 17954
rect 13597 17833 13643 17954
rect 13643 17833 13648 17954
rect 13454 17534 13459 17654
rect 13459 17534 13505 17654
rect 13505 17534 13510 17654
rect 12994 17415 12995 17458
rect 12995 17415 13049 17458
rect 13049 17415 13050 17458
rect 12994 17402 13050 17415
rect 13178 17415 13179 17458
rect 13179 17415 13233 17458
rect 13233 17415 13234 17458
rect 13178 17402 13234 17415
rect 13362 17415 13363 17458
rect 13363 17415 13417 17458
rect 13417 17415 13418 17458
rect 13362 17402 13418 17415
rect 11612 17252 11668 17308
rect 12994 17252 13050 17308
rect 12322 17136 12378 17192
rect 13178 17136 13234 17192
rect 13507 17136 13563 17192
rect 13764 17136 13820 17192
rect 13362 17020 13418 17076
rect 12994 16913 13050 16926
rect 12994 16870 12995 16913
rect 12995 16870 13049 16913
rect 13049 16870 13050 16913
rect 13178 16913 13234 16926
rect 13178 16870 13179 16913
rect 13179 16870 13233 16913
rect 13233 16870 13234 16913
rect 13362 16913 13418 16926
rect 13362 16870 13363 16913
rect 13363 16870 13417 16913
rect 13417 16870 13418 16913
rect 13454 16674 13459 16794
rect 13459 16674 13505 16794
rect 13505 16674 13510 16794
rect 12769 16351 12825 16407
rect 13587 16351 13643 16407
rect 13940 16233 13996 16289
rect 13764 16125 13820 16179
rect 10714 16016 10770 16072
rect 10346 15629 10351 15749
rect 10351 15629 10397 15749
rect 10397 15629 10402 15749
rect 10714 15629 10719 15749
rect 10719 15629 10765 15749
rect 10765 15629 10770 15749
rect 10530 15329 10535 15449
rect 10535 15329 10581 15449
rect 10581 15329 10586 15449
rect 11036 15628 11041 15749
rect 11041 15628 11087 15749
rect 11087 15628 11092 15749
rect 10898 15329 10903 15449
rect 10903 15329 10949 15449
rect 10949 15329 10954 15449
rect 10438 15210 10439 15253
rect 10439 15210 10493 15253
rect 10493 15210 10494 15253
rect 10438 15197 10494 15210
rect 10622 15210 10623 15253
rect 10623 15210 10677 15253
rect 10677 15210 10678 15253
rect 10622 15197 10678 15210
rect 10806 15210 10807 15253
rect 10807 15210 10861 15253
rect 10861 15210 10862 15253
rect 10806 15197 10862 15210
rect 10438 15047 10494 15103
rect 13270 16016 13326 16072
rect 12902 15629 12907 15749
rect 12907 15629 12953 15749
rect 12953 15629 12958 15749
rect 13270 15629 13275 15749
rect 13275 15629 13321 15749
rect 13321 15629 13326 15749
rect 13086 15329 13091 15449
rect 13091 15329 13137 15449
rect 13137 15329 13142 15449
rect 13592 15628 13597 15749
rect 13597 15628 13643 15749
rect 13643 15628 13648 15749
rect 13454 15329 13459 15449
rect 13459 15329 13505 15449
rect 13505 15329 13510 15449
rect 12994 15210 12995 15253
rect 12995 15210 13049 15253
rect 13049 15210 13050 15253
rect 12994 15197 13050 15210
rect 13178 15210 13179 15253
rect 13179 15210 13233 15253
rect 13233 15210 13234 15253
rect 13178 15197 13234 15210
rect 13362 15210 13363 15253
rect 13363 15210 13417 15253
rect 13417 15210 13418 15253
rect 13362 15197 13418 15210
rect 12994 15047 13050 15103
rect 17312 18221 17368 18277
rect 16944 17834 16949 17954
rect 16949 17834 16995 17954
rect 16995 17834 17000 17954
rect 17312 17834 17317 17954
rect 17317 17834 17363 17954
rect 17363 17834 17368 17954
rect 17128 17534 17133 17654
rect 17133 17534 17179 17654
rect 17179 17534 17184 17654
rect 17634 17833 17639 17954
rect 17639 17833 17685 17954
rect 17685 17833 17690 17954
rect 17496 17534 17501 17654
rect 17501 17534 17547 17654
rect 17547 17534 17552 17654
rect 17036 17415 17037 17458
rect 17037 17415 17091 17458
rect 17091 17415 17092 17458
rect 17036 17402 17092 17415
rect 17220 17415 17221 17458
rect 17221 17415 17275 17458
rect 17275 17415 17276 17458
rect 17220 17402 17276 17415
rect 17404 17415 17405 17458
rect 17405 17415 17459 17458
rect 17459 17415 17460 17458
rect 17404 17402 17460 17415
rect 15654 17252 15710 17308
rect 17036 17252 17092 17308
rect 16364 17136 16420 17192
rect 17220 17136 17276 17192
rect 17549 17136 17605 17192
rect 17806 17136 17862 17192
rect 17404 17020 17460 17076
rect 17036 16913 17092 16926
rect 17036 16870 17037 16913
rect 17037 16870 17091 16913
rect 17091 16870 17092 16913
rect 17220 16913 17276 16926
rect 17220 16870 17221 16913
rect 17221 16870 17275 16913
rect 17275 16870 17276 16913
rect 17404 16913 17460 16926
rect 17404 16870 17405 16913
rect 17405 16870 17459 16913
rect 17459 16870 17460 16913
rect 17496 16674 17501 16794
rect 17501 16674 17547 16794
rect 17547 16674 17552 16794
rect 16811 16351 16867 16407
rect 17629 16351 17685 16407
rect 17982 16233 18038 16289
rect 17806 16125 17862 16179
rect 14756 16016 14812 16072
rect 14388 15629 14393 15749
rect 14393 15629 14439 15749
rect 14439 15629 14444 15749
rect 14756 15629 14761 15749
rect 14761 15629 14807 15749
rect 14807 15629 14812 15749
rect 14572 15329 14577 15449
rect 14577 15329 14623 15449
rect 14623 15329 14628 15449
rect 15078 15628 15083 15749
rect 15083 15628 15129 15749
rect 15129 15628 15134 15749
rect 14940 15329 14945 15449
rect 14945 15329 14991 15449
rect 14991 15329 14996 15449
rect 14480 15210 14481 15253
rect 14481 15210 14535 15253
rect 14535 15210 14536 15253
rect 14480 15197 14536 15210
rect 14664 15210 14665 15253
rect 14665 15210 14719 15253
rect 14719 15210 14720 15253
rect 14664 15197 14720 15210
rect 14848 15210 14849 15253
rect 14849 15210 14903 15253
rect 14903 15210 14904 15253
rect 14848 15197 14904 15210
rect 14480 15047 14536 15103
rect 17312 16016 17368 16072
rect 16944 15629 16949 15749
rect 16949 15629 16995 15749
rect 16995 15629 17000 15749
rect 17312 15629 17317 15749
rect 17317 15629 17363 15749
rect 17363 15629 17368 15749
rect 17128 15329 17133 15449
rect 17133 15329 17179 15449
rect 17179 15329 17184 15449
rect 17634 15628 17639 15749
rect 17639 15628 17685 15749
rect 17685 15628 17690 15749
rect 17496 15329 17501 15449
rect 17501 15329 17547 15449
rect 17547 15329 17552 15449
rect 17036 15210 17037 15253
rect 17037 15210 17091 15253
rect 17091 15210 17092 15253
rect 17036 15197 17092 15210
rect 17220 15210 17221 15253
rect 17221 15210 17275 15253
rect 17275 15210 17276 15253
rect 17220 15197 17276 15210
rect 17404 15210 17405 15253
rect 17405 15210 17459 15253
rect 17459 15210 17460 15253
rect 17404 15197 17460 15210
rect 17036 15047 17092 15103
rect 21354 18221 21410 18277
rect 20986 17834 20991 17954
rect 20991 17834 21037 17954
rect 21037 17834 21042 17954
rect 21354 17834 21359 17954
rect 21359 17834 21405 17954
rect 21405 17834 21410 17954
rect 21170 17534 21175 17654
rect 21175 17534 21221 17654
rect 21221 17534 21226 17654
rect 21676 17833 21681 17954
rect 21681 17833 21727 17954
rect 21727 17833 21732 17954
rect 21538 17534 21543 17654
rect 21543 17534 21589 17654
rect 21589 17534 21594 17654
rect 21078 17415 21079 17458
rect 21079 17415 21133 17458
rect 21133 17415 21134 17458
rect 21078 17402 21134 17415
rect 21262 17415 21263 17458
rect 21263 17415 21317 17458
rect 21317 17415 21318 17458
rect 21262 17402 21318 17415
rect 21446 17415 21447 17458
rect 21447 17415 21501 17458
rect 21501 17415 21502 17458
rect 21446 17402 21502 17415
rect 19696 17252 19752 17308
rect 21078 17252 21134 17308
rect 20406 17136 20462 17192
rect 21262 17136 21318 17192
rect 21591 17136 21647 17192
rect 21848 17136 21904 17192
rect 21446 17020 21502 17076
rect 21078 16913 21134 16926
rect 21078 16870 21079 16913
rect 21079 16870 21133 16913
rect 21133 16870 21134 16913
rect 21262 16913 21318 16926
rect 21262 16870 21263 16913
rect 21263 16870 21317 16913
rect 21317 16870 21318 16913
rect 21446 16913 21502 16926
rect 21446 16870 21447 16913
rect 21447 16870 21501 16913
rect 21501 16870 21502 16913
rect 21538 16674 21543 16794
rect 21543 16674 21589 16794
rect 21589 16674 21594 16794
rect 20853 16351 20909 16407
rect 21671 16351 21727 16407
rect 22024 16233 22080 16289
rect 21848 16125 21904 16179
rect 18798 16016 18854 16072
rect 18430 15629 18435 15749
rect 18435 15629 18481 15749
rect 18481 15629 18486 15749
rect 18798 15629 18803 15749
rect 18803 15629 18849 15749
rect 18849 15629 18854 15749
rect 18614 15329 18619 15449
rect 18619 15329 18665 15449
rect 18665 15329 18670 15449
rect 19120 15628 19125 15749
rect 19125 15628 19171 15749
rect 19171 15628 19176 15749
rect 18982 15329 18987 15449
rect 18987 15329 19033 15449
rect 19033 15329 19038 15449
rect 18522 15210 18523 15253
rect 18523 15210 18577 15253
rect 18577 15210 18578 15253
rect 18522 15197 18578 15210
rect 18706 15210 18707 15253
rect 18707 15210 18761 15253
rect 18761 15210 18762 15253
rect 18706 15197 18762 15210
rect 18890 15210 18891 15253
rect 18891 15210 18945 15253
rect 18945 15210 18946 15253
rect 18890 15197 18946 15210
rect 18522 15047 18578 15103
rect 21354 16016 21410 16072
rect 20986 15629 20991 15749
rect 20991 15629 21037 15749
rect 21037 15629 21042 15749
rect 21354 15629 21359 15749
rect 21359 15629 21405 15749
rect 21405 15629 21410 15749
rect 21170 15329 21175 15449
rect 21175 15329 21221 15449
rect 21221 15329 21226 15449
rect 21676 15628 21681 15749
rect 21681 15628 21727 15749
rect 21727 15628 21732 15749
rect 21538 15329 21543 15449
rect 21543 15329 21589 15449
rect 21589 15329 21594 15449
rect 21078 15210 21079 15253
rect 21079 15210 21133 15253
rect 21133 15210 21134 15253
rect 21078 15197 21134 15210
rect 21262 15210 21263 15253
rect 21263 15210 21317 15253
rect 21317 15210 21318 15253
rect 21262 15197 21318 15210
rect 21446 15210 21447 15253
rect 21447 15210 21501 15253
rect 21501 15210 21502 15253
rect 21446 15197 21502 15210
rect 21078 15047 21134 15103
rect 25396 18221 25452 18277
rect 25028 17834 25033 17954
rect 25033 17834 25079 17954
rect 25079 17834 25084 17954
rect 25396 17834 25401 17954
rect 25401 17834 25447 17954
rect 25447 17834 25452 17954
rect 25212 17534 25217 17654
rect 25217 17534 25263 17654
rect 25263 17534 25268 17654
rect 25718 17833 25723 17954
rect 25723 17833 25769 17954
rect 25769 17833 25774 17954
rect 25580 17534 25585 17654
rect 25585 17534 25631 17654
rect 25631 17534 25636 17654
rect 25120 17415 25121 17458
rect 25121 17415 25175 17458
rect 25175 17415 25176 17458
rect 25120 17402 25176 17415
rect 25304 17415 25305 17458
rect 25305 17415 25359 17458
rect 25359 17415 25360 17458
rect 25304 17402 25360 17415
rect 25488 17415 25489 17458
rect 25489 17415 25543 17458
rect 25543 17415 25544 17458
rect 25488 17402 25544 17415
rect 23738 17252 23794 17308
rect 25120 17252 25176 17308
rect 24448 17136 24504 17192
rect 25304 17136 25360 17192
rect 25633 17136 25689 17192
rect 25890 17136 25946 17192
rect 25488 17020 25544 17076
rect 25120 16913 25176 16926
rect 25120 16870 25121 16913
rect 25121 16870 25175 16913
rect 25175 16870 25176 16913
rect 25304 16913 25360 16926
rect 25304 16870 25305 16913
rect 25305 16870 25359 16913
rect 25359 16870 25360 16913
rect 25488 16913 25544 16926
rect 25488 16870 25489 16913
rect 25489 16870 25543 16913
rect 25543 16870 25544 16913
rect 25580 16674 25585 16794
rect 25585 16674 25631 16794
rect 25631 16674 25636 16794
rect 24895 16351 24951 16407
rect 25713 16351 25769 16407
rect 26066 16233 26122 16289
rect 25890 16125 25946 16179
rect 22840 16016 22896 16072
rect 22472 15629 22477 15749
rect 22477 15629 22523 15749
rect 22523 15629 22528 15749
rect 22840 15629 22845 15749
rect 22845 15629 22891 15749
rect 22891 15629 22896 15749
rect 22656 15329 22661 15449
rect 22661 15329 22707 15449
rect 22707 15329 22712 15449
rect 23162 15628 23167 15749
rect 23167 15628 23213 15749
rect 23213 15628 23218 15749
rect 23024 15329 23029 15449
rect 23029 15329 23075 15449
rect 23075 15329 23080 15449
rect 22564 15210 22565 15253
rect 22565 15210 22619 15253
rect 22619 15210 22620 15253
rect 22564 15197 22620 15210
rect 22748 15210 22749 15253
rect 22749 15210 22803 15253
rect 22803 15210 22804 15253
rect 22748 15197 22804 15210
rect 22932 15210 22933 15253
rect 22933 15210 22987 15253
rect 22987 15210 22988 15253
rect 22932 15197 22988 15210
rect 22564 15047 22620 15103
rect 25396 16016 25452 16072
rect 25028 15629 25033 15749
rect 25033 15629 25079 15749
rect 25079 15629 25084 15749
rect 25396 15629 25401 15749
rect 25401 15629 25447 15749
rect 25447 15629 25452 15749
rect 25212 15329 25217 15449
rect 25217 15329 25263 15449
rect 25263 15329 25268 15449
rect 25718 15628 25723 15749
rect 25723 15628 25769 15749
rect 25769 15628 25774 15749
rect 25580 15329 25585 15449
rect 25585 15329 25631 15449
rect 25631 15329 25636 15449
rect 25120 15210 25121 15253
rect 25121 15210 25175 15253
rect 25175 15210 25176 15253
rect 25120 15197 25176 15210
rect 25304 15210 25305 15253
rect 25305 15210 25359 15253
rect 25359 15210 25360 15253
rect 25304 15197 25360 15210
rect 25488 15210 25489 15253
rect 25489 15210 25543 15253
rect 25543 15210 25544 15253
rect 25488 15197 25544 15210
rect 25120 15047 25176 15103
rect 29438 18221 29494 18277
rect 29070 17834 29075 17954
rect 29075 17834 29121 17954
rect 29121 17834 29126 17954
rect 29438 17834 29443 17954
rect 29443 17834 29489 17954
rect 29489 17834 29494 17954
rect 29254 17534 29259 17654
rect 29259 17534 29305 17654
rect 29305 17534 29310 17654
rect 29760 17833 29765 17954
rect 29765 17833 29811 17954
rect 29811 17833 29816 17954
rect 29622 17534 29627 17654
rect 29627 17534 29673 17654
rect 29673 17534 29678 17654
rect 29162 17415 29163 17458
rect 29163 17415 29217 17458
rect 29217 17415 29218 17458
rect 29162 17402 29218 17415
rect 29346 17415 29347 17458
rect 29347 17415 29401 17458
rect 29401 17415 29402 17458
rect 29346 17402 29402 17415
rect 29530 17415 29531 17458
rect 29531 17415 29585 17458
rect 29585 17415 29586 17458
rect 29530 17402 29586 17415
rect 27780 17252 27836 17308
rect 29162 17252 29218 17308
rect 28490 17136 28546 17192
rect 29346 17136 29402 17192
rect 29675 17136 29731 17192
rect 29932 17136 29988 17192
rect 29530 17020 29586 17076
rect 29162 16913 29218 16926
rect 29162 16870 29163 16913
rect 29163 16870 29217 16913
rect 29217 16870 29218 16913
rect 29346 16913 29402 16926
rect 29346 16870 29347 16913
rect 29347 16870 29401 16913
rect 29401 16870 29402 16913
rect 29530 16913 29586 16926
rect 29530 16870 29531 16913
rect 29531 16870 29585 16913
rect 29585 16870 29586 16913
rect 29622 16674 29627 16794
rect 29627 16674 29673 16794
rect 29673 16674 29678 16794
rect 28937 16351 28993 16407
rect 29755 16351 29811 16407
rect 30108 16233 30164 16289
rect 29932 16125 29988 16179
rect 26882 16016 26938 16072
rect 26514 15629 26519 15749
rect 26519 15629 26565 15749
rect 26565 15629 26570 15749
rect 26882 15629 26887 15749
rect 26887 15629 26933 15749
rect 26933 15629 26938 15749
rect 26698 15329 26703 15449
rect 26703 15329 26749 15449
rect 26749 15329 26754 15449
rect 27204 15628 27209 15749
rect 27209 15628 27255 15749
rect 27255 15628 27260 15749
rect 27066 15329 27071 15449
rect 27071 15329 27117 15449
rect 27117 15329 27122 15449
rect 26606 15210 26607 15253
rect 26607 15210 26661 15253
rect 26661 15210 26662 15253
rect 26606 15197 26662 15210
rect 26790 15210 26791 15253
rect 26791 15210 26845 15253
rect 26845 15210 26846 15253
rect 26790 15197 26846 15210
rect 26974 15210 26975 15253
rect 26975 15210 27029 15253
rect 27029 15210 27030 15253
rect 26974 15197 27030 15210
rect 26606 15047 26662 15103
rect 29438 16016 29494 16072
rect 29070 15629 29075 15749
rect 29075 15629 29121 15749
rect 29121 15629 29126 15749
rect 29438 15629 29443 15749
rect 29443 15629 29489 15749
rect 29489 15629 29494 15749
rect 29254 15329 29259 15449
rect 29259 15329 29305 15449
rect 29305 15329 29310 15449
rect 29760 15628 29765 15749
rect 29765 15628 29811 15749
rect 29811 15628 29816 15749
rect 29622 15329 29627 15449
rect 29627 15329 29673 15449
rect 29673 15329 29678 15449
rect 29162 15210 29163 15253
rect 29163 15210 29217 15253
rect 29217 15210 29218 15253
rect 29162 15197 29218 15210
rect 29346 15210 29347 15253
rect 29347 15210 29401 15253
rect 29401 15210 29402 15253
rect 29346 15197 29402 15210
rect 29530 15210 29531 15253
rect 29531 15210 29585 15253
rect 29585 15210 29586 15253
rect 29530 15197 29586 15210
rect 29162 15047 29218 15103
rect 30924 16016 30980 16072
rect 30556 15629 30561 15749
rect 30561 15629 30607 15749
rect 30607 15629 30612 15749
rect 30924 15629 30929 15749
rect 30929 15629 30975 15749
rect 30975 15629 30980 15749
rect 30740 15329 30745 15449
rect 30745 15329 30791 15449
rect 30791 15329 30796 15449
rect 31246 15628 31251 15749
rect 31251 15628 31297 15749
rect 31297 15628 31302 15749
rect 31108 15329 31113 15449
rect 31113 15329 31159 15449
rect 31159 15329 31164 15449
rect 30648 15210 30649 15253
rect 30649 15210 30703 15253
rect 30703 15210 30704 15253
rect 30648 15197 30704 15210
rect 30832 15210 30833 15253
rect 30833 15210 30887 15253
rect 30887 15210 30888 15253
rect 30832 15197 30888 15210
rect 31016 15210 31017 15253
rect 31017 15210 31071 15253
rect 31071 15210 31072 15253
rect 31016 15197 31072 15210
rect 30648 15047 30704 15103
rect 4102 14934 4158 14990
rect 5094 14934 5150 14990
rect 5423 14934 5479 14990
rect 5856 14934 5912 14990
rect 6580 14934 6636 14990
rect 6909 14934 6965 14990
rect 7166 14934 7222 14990
rect 7706 14934 7762 14990
rect 8144 14931 8200 14987
rect 9136 14931 9192 14987
rect 9465 14931 9521 14987
rect 9898 14931 9954 14987
rect 10622 14931 10678 14987
rect 10951 14931 11007 14987
rect 11208 14931 11264 14987
rect 11760 14931 11816 14987
rect 12186 14931 12242 14987
rect 13178 14931 13234 14987
rect 13507 14931 13563 14987
rect 13940 14931 13996 14987
rect 14664 14931 14720 14987
rect 14993 14931 15049 14987
rect 15250 14931 15306 14987
rect 15856 14931 15912 14987
rect 16228 14931 16284 14987
rect 17220 14931 17276 14987
rect 17549 14931 17605 14987
rect 17982 14931 18038 14987
rect 18706 14931 18762 14987
rect 19035 14931 19091 14987
rect 19292 14931 19348 14987
rect 19898 14931 19954 14987
rect 20270 14931 20326 14987
rect 21262 14931 21318 14987
rect 21591 14931 21647 14987
rect 22024 14931 22080 14987
rect 22748 14931 22804 14987
rect 23077 14931 23133 14987
rect 23334 14931 23390 14987
rect 23940 14931 23996 14987
rect 24312 14931 24368 14987
rect 25304 14931 25360 14987
rect 25633 14931 25689 14987
rect 26066 14931 26122 14987
rect 26790 14931 26846 14987
rect 27119 14931 27175 14987
rect 27376 14931 27432 14987
rect 27982 14931 28038 14987
rect 28354 14931 28410 14987
rect 29346 14931 29402 14987
rect 29675 14931 29731 14987
rect 30108 14931 30164 14987
rect 30832 14931 30888 14987
rect 31161 14931 31217 14987
rect 31418 14931 31474 14987
rect 32024 14931 32080 14987
rect 5278 14818 5334 14874
rect 6764 14818 6820 14874
rect 4910 14711 4966 14724
rect 4910 14668 4911 14711
rect 4911 14668 4965 14711
rect 4965 14668 4966 14711
rect 5094 14711 5150 14724
rect 5094 14668 5095 14711
rect 5095 14668 5149 14711
rect 5149 14668 5150 14711
rect 5278 14711 5334 14724
rect 5278 14668 5279 14711
rect 5279 14668 5333 14711
rect 5333 14668 5334 14711
rect 5370 14472 5375 14592
rect 5375 14472 5421 14592
rect 5421 14472 5426 14592
rect 4685 14149 4741 14205
rect 5503 14149 5559 14205
rect 3912 14032 3968 14088
rect 9320 14815 9376 14871
rect 6396 14711 6452 14724
rect 6396 14668 6397 14711
rect 6397 14668 6451 14711
rect 6451 14668 6452 14711
rect 6580 14711 6636 14724
rect 6580 14668 6581 14711
rect 6581 14668 6635 14711
rect 6635 14668 6636 14711
rect 6764 14711 6820 14724
rect 6764 14668 6765 14711
rect 6765 14668 6819 14711
rect 6819 14668 6820 14711
rect 6856 14472 6861 14592
rect 6861 14472 6907 14592
rect 6907 14472 6912 14592
rect 6171 14149 6227 14205
rect 6989 14149 7045 14205
rect 7342 14032 7398 14088
rect 10806 14815 10862 14871
rect 8952 14708 9008 14721
rect 8952 14665 8953 14708
rect 8953 14665 9007 14708
rect 9007 14665 9008 14708
rect 9136 14708 9192 14721
rect 9136 14665 9137 14708
rect 9137 14665 9191 14708
rect 9191 14665 9192 14708
rect 9320 14708 9376 14721
rect 9320 14665 9321 14708
rect 9321 14665 9375 14708
rect 9375 14665 9376 14708
rect 9412 14469 9417 14589
rect 9417 14469 9463 14589
rect 9463 14469 9468 14589
rect 8727 14146 8783 14202
rect 9545 14146 9601 14202
rect 8008 14029 8064 14085
rect 13362 14815 13418 14871
rect 10438 14708 10494 14721
rect 10438 14665 10439 14708
rect 10439 14665 10493 14708
rect 10493 14665 10494 14708
rect 10622 14708 10678 14721
rect 10622 14665 10623 14708
rect 10623 14665 10677 14708
rect 10677 14665 10678 14708
rect 10806 14708 10862 14721
rect 10806 14665 10807 14708
rect 10807 14665 10861 14708
rect 10861 14665 10862 14708
rect 10898 14469 10903 14589
rect 10903 14469 10949 14589
rect 10949 14469 10954 14589
rect 10213 14146 10269 14202
rect 11031 14146 11087 14202
rect 11384 14029 11440 14085
rect 5856 13921 5912 13977
rect 7166 13922 7222 13978
rect 5186 13814 5242 13870
rect 4818 13427 4823 13547
rect 4823 13427 4869 13547
rect 4869 13427 4874 13547
rect 5186 13427 5191 13547
rect 5191 13427 5237 13547
rect 5237 13427 5242 13547
rect 5002 13127 5007 13247
rect 5007 13127 5053 13247
rect 5053 13127 5058 13247
rect 5508 13426 5513 13547
rect 5513 13426 5559 13547
rect 5559 13426 5564 13547
rect 5370 13127 5375 13247
rect 5375 13127 5421 13247
rect 5421 13127 5426 13247
rect 4910 13008 4911 13051
rect 4911 13008 4965 13051
rect 4965 13008 4966 13051
rect 4910 12995 4966 13008
rect 5094 13008 5095 13051
rect 5095 13008 5149 13051
rect 5149 13008 5150 13051
rect 5094 12995 5150 13008
rect 5278 13008 5279 13051
rect 5279 13008 5333 13051
rect 5333 13008 5334 13051
rect 5278 12995 5334 13008
rect 4910 12845 4966 12901
rect 6672 13815 6728 13871
rect 6304 13428 6309 13548
rect 6309 13428 6355 13548
rect 6355 13428 6360 13548
rect 6672 13428 6677 13548
rect 6677 13428 6723 13548
rect 6723 13428 6728 13548
rect 6488 13128 6493 13248
rect 6493 13128 6539 13248
rect 6539 13128 6544 13248
rect 6994 13427 6999 13548
rect 6999 13427 7045 13548
rect 7045 13427 7050 13548
rect 6856 13128 6861 13248
rect 6861 13128 6907 13248
rect 6907 13128 6912 13248
rect 6396 13009 6397 13052
rect 6397 13009 6451 13052
rect 6451 13009 6452 13052
rect 6396 12996 6452 13009
rect 6580 13009 6581 13052
rect 6581 13009 6635 13052
rect 6635 13009 6636 13052
rect 6580 12996 6636 13009
rect 6764 13009 6765 13052
rect 6765 13009 6819 13052
rect 6819 13009 6820 13052
rect 6764 12996 6820 13009
rect 6396 12846 6452 12902
rect 5094 12729 5150 12785
rect 5423 12729 5479 12785
rect 5680 12729 5736 12785
rect 6580 12730 6636 12786
rect 6909 12730 6965 12786
rect 7342 12730 7398 12786
rect 14848 14815 14904 14871
rect 12994 14708 13050 14721
rect 12994 14665 12995 14708
rect 12995 14665 13049 14708
rect 13049 14665 13050 14708
rect 13178 14708 13234 14721
rect 13178 14665 13179 14708
rect 13179 14665 13233 14708
rect 13233 14665 13234 14708
rect 13362 14708 13418 14721
rect 13362 14665 13363 14708
rect 13363 14665 13417 14708
rect 13417 14665 13418 14708
rect 13454 14469 13459 14589
rect 13459 14469 13505 14589
rect 13505 14469 13510 14589
rect 12769 14146 12825 14202
rect 13587 14146 13643 14202
rect 12050 14029 12106 14085
rect 17404 14815 17460 14871
rect 14480 14708 14536 14721
rect 14480 14665 14481 14708
rect 14481 14665 14535 14708
rect 14535 14665 14536 14708
rect 14664 14708 14720 14721
rect 14664 14665 14665 14708
rect 14665 14665 14719 14708
rect 14719 14665 14720 14708
rect 14848 14708 14904 14721
rect 14848 14665 14849 14708
rect 14849 14665 14903 14708
rect 14903 14665 14904 14708
rect 14940 14469 14945 14589
rect 14945 14469 14991 14589
rect 14991 14469 14996 14589
rect 14255 14146 14311 14202
rect 15073 14146 15129 14202
rect 15426 14029 15482 14085
rect 9898 13918 9954 13974
rect 11208 13919 11264 13975
rect 9228 13811 9284 13867
rect 8860 13424 8865 13544
rect 8865 13424 8911 13544
rect 8911 13424 8916 13544
rect 9228 13424 9233 13544
rect 9233 13424 9279 13544
rect 9279 13424 9284 13544
rect 9044 13124 9049 13244
rect 9049 13124 9095 13244
rect 9095 13124 9100 13244
rect 9550 13423 9555 13544
rect 9555 13423 9601 13544
rect 9601 13423 9606 13544
rect 9412 13124 9417 13244
rect 9417 13124 9463 13244
rect 9463 13124 9468 13244
rect 8952 13005 8953 13048
rect 8953 13005 9007 13048
rect 9007 13005 9008 13048
rect 8952 12992 9008 13005
rect 9136 13005 9137 13048
rect 9137 13005 9191 13048
rect 9191 13005 9192 13048
rect 9136 12992 9192 13005
rect 9320 13005 9321 13048
rect 9321 13005 9375 13048
rect 9375 13005 9376 13048
rect 9320 12992 9376 13005
rect 8952 12842 9008 12898
rect 10714 13812 10770 13868
rect 10346 13425 10351 13545
rect 10351 13425 10397 13545
rect 10397 13425 10402 13545
rect 10714 13425 10719 13545
rect 10719 13425 10765 13545
rect 10765 13425 10770 13545
rect 10530 13125 10535 13245
rect 10535 13125 10581 13245
rect 10581 13125 10586 13245
rect 11036 13424 11041 13545
rect 11041 13424 11087 13545
rect 11087 13424 11092 13545
rect 10898 13125 10903 13245
rect 10903 13125 10949 13245
rect 10949 13125 10954 13245
rect 10438 13006 10439 13049
rect 10439 13006 10493 13049
rect 10493 13006 10494 13049
rect 10438 12993 10494 13006
rect 10622 13006 10623 13049
rect 10623 13006 10677 13049
rect 10677 13006 10678 13049
rect 10622 12993 10678 13006
rect 10806 13006 10807 13049
rect 10807 13006 10861 13049
rect 10861 13006 10862 13049
rect 10806 12993 10862 13006
rect 10438 12843 10494 12899
rect 9136 12726 9192 12782
rect 9465 12726 9521 12782
rect 9722 12726 9778 12782
rect 10622 12727 10678 12783
rect 10951 12727 11007 12783
rect 11384 12727 11440 12783
rect 18890 14815 18946 14871
rect 17036 14708 17092 14721
rect 17036 14665 17037 14708
rect 17037 14665 17091 14708
rect 17091 14665 17092 14708
rect 17220 14708 17276 14721
rect 17220 14665 17221 14708
rect 17221 14665 17275 14708
rect 17275 14665 17276 14708
rect 17404 14708 17460 14721
rect 17404 14665 17405 14708
rect 17405 14665 17459 14708
rect 17459 14665 17460 14708
rect 17496 14469 17501 14589
rect 17501 14469 17547 14589
rect 17547 14469 17552 14589
rect 16811 14146 16867 14202
rect 17629 14146 17685 14202
rect 16092 14029 16148 14085
rect 21446 14815 21502 14871
rect 18522 14708 18578 14721
rect 18522 14665 18523 14708
rect 18523 14665 18577 14708
rect 18577 14665 18578 14708
rect 18706 14708 18762 14721
rect 18706 14665 18707 14708
rect 18707 14665 18761 14708
rect 18761 14665 18762 14708
rect 18890 14708 18946 14721
rect 18890 14665 18891 14708
rect 18891 14665 18945 14708
rect 18945 14665 18946 14708
rect 18982 14469 18987 14589
rect 18987 14469 19033 14589
rect 19033 14469 19038 14589
rect 18297 14146 18353 14202
rect 19115 14146 19171 14202
rect 19468 14029 19524 14085
rect 13940 13918 13996 13974
rect 15250 13919 15306 13975
rect 13270 13811 13326 13867
rect 12902 13424 12907 13544
rect 12907 13424 12953 13544
rect 12953 13424 12958 13544
rect 13270 13424 13275 13544
rect 13275 13424 13321 13544
rect 13321 13424 13326 13544
rect 13086 13124 13091 13244
rect 13091 13124 13137 13244
rect 13137 13124 13142 13244
rect 13592 13423 13597 13544
rect 13597 13423 13643 13544
rect 13643 13423 13648 13544
rect 13454 13124 13459 13244
rect 13459 13124 13505 13244
rect 13505 13124 13510 13244
rect 12994 13005 12995 13048
rect 12995 13005 13049 13048
rect 13049 13005 13050 13048
rect 12994 12992 13050 13005
rect 13178 13005 13179 13048
rect 13179 13005 13233 13048
rect 13233 13005 13234 13048
rect 13178 12992 13234 13005
rect 13362 13005 13363 13048
rect 13363 13005 13417 13048
rect 13417 13005 13418 13048
rect 13362 12992 13418 13005
rect 12994 12842 13050 12898
rect 14756 13812 14812 13868
rect 14388 13425 14393 13545
rect 14393 13425 14439 13545
rect 14439 13425 14444 13545
rect 14756 13425 14761 13545
rect 14761 13425 14807 13545
rect 14807 13425 14812 13545
rect 14572 13125 14577 13245
rect 14577 13125 14623 13245
rect 14623 13125 14628 13245
rect 15078 13424 15083 13545
rect 15083 13424 15129 13545
rect 15129 13424 15134 13545
rect 14940 13125 14945 13245
rect 14945 13125 14991 13245
rect 14991 13125 14996 13245
rect 14480 13006 14481 13049
rect 14481 13006 14535 13049
rect 14535 13006 14536 13049
rect 14480 12993 14536 13006
rect 14664 13006 14665 13049
rect 14665 13006 14719 13049
rect 14719 13006 14720 13049
rect 14664 12993 14720 13006
rect 14848 13006 14849 13049
rect 14849 13006 14903 13049
rect 14903 13006 14904 13049
rect 14848 12993 14904 13006
rect 14480 12843 14536 12899
rect 13178 12726 13234 12782
rect 13507 12726 13563 12782
rect 13764 12726 13820 12782
rect 14664 12727 14720 12783
rect 14993 12727 15049 12783
rect 15426 12727 15482 12783
rect 22932 14815 22988 14871
rect 21078 14708 21134 14721
rect 21078 14665 21079 14708
rect 21079 14665 21133 14708
rect 21133 14665 21134 14708
rect 21262 14708 21318 14721
rect 21262 14665 21263 14708
rect 21263 14665 21317 14708
rect 21317 14665 21318 14708
rect 21446 14708 21502 14721
rect 21446 14665 21447 14708
rect 21447 14665 21501 14708
rect 21501 14665 21502 14708
rect 21538 14469 21543 14589
rect 21543 14469 21589 14589
rect 21589 14469 21594 14589
rect 20853 14146 20909 14202
rect 21671 14146 21727 14202
rect 20134 14029 20190 14085
rect 25488 14815 25544 14871
rect 22564 14708 22620 14721
rect 22564 14665 22565 14708
rect 22565 14665 22619 14708
rect 22619 14665 22620 14708
rect 22748 14708 22804 14721
rect 22748 14665 22749 14708
rect 22749 14665 22803 14708
rect 22803 14665 22804 14708
rect 22932 14708 22988 14721
rect 22932 14665 22933 14708
rect 22933 14665 22987 14708
rect 22987 14665 22988 14708
rect 23024 14469 23029 14589
rect 23029 14469 23075 14589
rect 23075 14469 23080 14589
rect 22339 14146 22395 14202
rect 23157 14146 23213 14202
rect 23510 14029 23566 14085
rect 17982 13918 18038 13974
rect 19292 13919 19348 13975
rect 17312 13811 17368 13867
rect 16944 13424 16949 13544
rect 16949 13424 16995 13544
rect 16995 13424 17000 13544
rect 17312 13424 17317 13544
rect 17317 13424 17363 13544
rect 17363 13424 17368 13544
rect 17128 13124 17133 13244
rect 17133 13124 17179 13244
rect 17179 13124 17184 13244
rect 17634 13423 17639 13544
rect 17639 13423 17685 13544
rect 17685 13423 17690 13544
rect 17496 13124 17501 13244
rect 17501 13124 17547 13244
rect 17547 13124 17552 13244
rect 17036 13005 17037 13048
rect 17037 13005 17091 13048
rect 17091 13005 17092 13048
rect 17036 12992 17092 13005
rect 17220 13005 17221 13048
rect 17221 13005 17275 13048
rect 17275 13005 17276 13048
rect 17220 12992 17276 13005
rect 17404 13005 17405 13048
rect 17405 13005 17459 13048
rect 17459 13005 17460 13048
rect 17404 12992 17460 13005
rect 17036 12842 17092 12898
rect 18798 13812 18854 13868
rect 18430 13425 18435 13545
rect 18435 13425 18481 13545
rect 18481 13425 18486 13545
rect 18798 13425 18803 13545
rect 18803 13425 18849 13545
rect 18849 13425 18854 13545
rect 18614 13125 18619 13245
rect 18619 13125 18665 13245
rect 18665 13125 18670 13245
rect 19120 13424 19125 13545
rect 19125 13424 19171 13545
rect 19171 13424 19176 13545
rect 18982 13125 18987 13245
rect 18987 13125 19033 13245
rect 19033 13125 19038 13245
rect 18522 13006 18523 13049
rect 18523 13006 18577 13049
rect 18577 13006 18578 13049
rect 18522 12993 18578 13006
rect 18706 13006 18707 13049
rect 18707 13006 18761 13049
rect 18761 13006 18762 13049
rect 18706 12993 18762 13006
rect 18890 13006 18891 13049
rect 18891 13006 18945 13049
rect 18945 13006 18946 13049
rect 18890 12993 18946 13006
rect 18522 12843 18578 12899
rect 17220 12726 17276 12782
rect 17549 12726 17605 12782
rect 17806 12726 17862 12782
rect 18706 12727 18762 12783
rect 19035 12727 19091 12783
rect 19468 12727 19524 12783
rect 26974 14815 27030 14871
rect 25120 14708 25176 14721
rect 25120 14665 25121 14708
rect 25121 14665 25175 14708
rect 25175 14665 25176 14708
rect 25304 14708 25360 14721
rect 25304 14665 25305 14708
rect 25305 14665 25359 14708
rect 25359 14665 25360 14708
rect 25488 14708 25544 14721
rect 25488 14665 25489 14708
rect 25489 14665 25543 14708
rect 25543 14665 25544 14708
rect 25580 14469 25585 14589
rect 25585 14469 25631 14589
rect 25631 14469 25636 14589
rect 24895 14146 24951 14202
rect 25713 14146 25769 14202
rect 24176 14029 24232 14085
rect 29530 14815 29586 14871
rect 26606 14708 26662 14721
rect 26606 14665 26607 14708
rect 26607 14665 26661 14708
rect 26661 14665 26662 14708
rect 26790 14708 26846 14721
rect 26790 14665 26791 14708
rect 26791 14665 26845 14708
rect 26845 14665 26846 14708
rect 26974 14708 27030 14721
rect 26974 14665 26975 14708
rect 26975 14665 27029 14708
rect 27029 14665 27030 14708
rect 27066 14469 27071 14589
rect 27071 14469 27117 14589
rect 27117 14469 27122 14589
rect 26381 14146 26437 14202
rect 27199 14146 27255 14202
rect 27552 14029 27608 14085
rect 22024 13918 22080 13974
rect 23334 13919 23390 13975
rect 21354 13811 21410 13867
rect 20986 13424 20991 13544
rect 20991 13424 21037 13544
rect 21037 13424 21042 13544
rect 21354 13424 21359 13544
rect 21359 13424 21405 13544
rect 21405 13424 21410 13544
rect 21170 13124 21175 13244
rect 21175 13124 21221 13244
rect 21221 13124 21226 13244
rect 21676 13423 21681 13544
rect 21681 13423 21727 13544
rect 21727 13423 21732 13544
rect 21538 13124 21543 13244
rect 21543 13124 21589 13244
rect 21589 13124 21594 13244
rect 21078 13005 21079 13048
rect 21079 13005 21133 13048
rect 21133 13005 21134 13048
rect 21078 12992 21134 13005
rect 21262 13005 21263 13048
rect 21263 13005 21317 13048
rect 21317 13005 21318 13048
rect 21262 12992 21318 13005
rect 21446 13005 21447 13048
rect 21447 13005 21501 13048
rect 21501 13005 21502 13048
rect 21446 12992 21502 13005
rect 21078 12842 21134 12898
rect 22840 13812 22896 13868
rect 22472 13425 22477 13545
rect 22477 13425 22523 13545
rect 22523 13425 22528 13545
rect 22840 13425 22845 13545
rect 22845 13425 22891 13545
rect 22891 13425 22896 13545
rect 22656 13125 22661 13245
rect 22661 13125 22707 13245
rect 22707 13125 22712 13245
rect 23162 13424 23167 13545
rect 23167 13424 23213 13545
rect 23213 13424 23218 13545
rect 23024 13125 23029 13245
rect 23029 13125 23075 13245
rect 23075 13125 23080 13245
rect 22564 13006 22565 13049
rect 22565 13006 22619 13049
rect 22619 13006 22620 13049
rect 22564 12993 22620 13006
rect 22748 13006 22749 13049
rect 22749 13006 22803 13049
rect 22803 13006 22804 13049
rect 22748 12993 22804 13006
rect 22932 13006 22933 13049
rect 22933 13006 22987 13049
rect 22987 13006 22988 13049
rect 22932 12993 22988 13006
rect 22564 12843 22620 12899
rect 21262 12726 21318 12782
rect 21591 12726 21647 12782
rect 21848 12726 21904 12782
rect 22748 12727 22804 12783
rect 23077 12727 23133 12783
rect 23510 12727 23566 12783
rect 31016 14815 31072 14871
rect 29162 14708 29218 14721
rect 29162 14665 29163 14708
rect 29163 14665 29217 14708
rect 29217 14665 29218 14708
rect 29346 14708 29402 14721
rect 29346 14665 29347 14708
rect 29347 14665 29401 14708
rect 29401 14665 29402 14708
rect 29530 14708 29586 14721
rect 29530 14665 29531 14708
rect 29531 14665 29585 14708
rect 29585 14665 29586 14708
rect 29622 14469 29627 14589
rect 29627 14469 29673 14589
rect 29673 14469 29678 14589
rect 28937 14146 28993 14202
rect 29755 14146 29811 14202
rect 28173 14029 28229 14085
rect 30648 14708 30704 14721
rect 30648 14665 30649 14708
rect 30649 14665 30703 14708
rect 30703 14665 30704 14708
rect 30832 14708 30888 14721
rect 30832 14665 30833 14708
rect 30833 14665 30887 14708
rect 30887 14665 30888 14708
rect 31016 14708 31072 14721
rect 31016 14665 31017 14708
rect 31017 14665 31071 14708
rect 31071 14665 31072 14708
rect 31108 14469 31113 14589
rect 31113 14469 31159 14589
rect 31159 14469 31164 14589
rect 30423 14146 30479 14202
rect 31241 14146 31297 14202
rect 31594 14029 31650 14085
rect 26066 13918 26122 13974
rect 27376 13919 27432 13975
rect 25396 13811 25452 13867
rect 25028 13424 25033 13544
rect 25033 13424 25079 13544
rect 25079 13424 25084 13544
rect 25396 13424 25401 13544
rect 25401 13424 25447 13544
rect 25447 13424 25452 13544
rect 25212 13124 25217 13244
rect 25217 13124 25263 13244
rect 25263 13124 25268 13244
rect 25718 13423 25723 13544
rect 25723 13423 25769 13544
rect 25769 13423 25774 13544
rect 25580 13124 25585 13244
rect 25585 13124 25631 13244
rect 25631 13124 25636 13244
rect 25120 13005 25121 13048
rect 25121 13005 25175 13048
rect 25175 13005 25176 13048
rect 25120 12992 25176 13005
rect 25304 13005 25305 13048
rect 25305 13005 25359 13048
rect 25359 13005 25360 13048
rect 25304 12992 25360 13005
rect 25488 13005 25489 13048
rect 25489 13005 25543 13048
rect 25543 13005 25544 13048
rect 25488 12992 25544 13005
rect 25120 12842 25176 12898
rect 26882 13812 26938 13868
rect 26514 13425 26519 13545
rect 26519 13425 26565 13545
rect 26565 13425 26570 13545
rect 26882 13425 26887 13545
rect 26887 13425 26933 13545
rect 26933 13425 26938 13545
rect 26698 13125 26703 13245
rect 26703 13125 26749 13245
rect 26749 13125 26754 13245
rect 27204 13424 27209 13545
rect 27209 13424 27255 13545
rect 27255 13424 27260 13545
rect 27066 13125 27071 13245
rect 27071 13125 27117 13245
rect 27117 13125 27122 13245
rect 26606 13006 26607 13049
rect 26607 13006 26661 13049
rect 26661 13006 26662 13049
rect 26606 12993 26662 13006
rect 26790 13006 26791 13049
rect 26791 13006 26845 13049
rect 26845 13006 26846 13049
rect 26790 12993 26846 13006
rect 26974 13006 26975 13049
rect 26975 13006 27029 13049
rect 27029 13006 27030 13049
rect 26974 12993 27030 13006
rect 26606 12843 26662 12899
rect 25304 12726 25360 12782
rect 25633 12726 25689 12782
rect 25890 12726 25946 12782
rect 26790 12727 26846 12783
rect 27119 12727 27175 12783
rect 27552 12727 27608 12783
rect 30108 13918 30164 13974
rect 31418 13919 31474 13975
rect 29438 13811 29494 13867
rect 29070 13424 29075 13544
rect 29075 13424 29121 13544
rect 29121 13424 29126 13544
rect 29438 13424 29443 13544
rect 29443 13424 29489 13544
rect 29489 13424 29494 13544
rect 29254 13124 29259 13244
rect 29259 13124 29305 13244
rect 29305 13124 29310 13244
rect 29760 13423 29765 13544
rect 29765 13423 29811 13544
rect 29811 13423 29816 13544
rect 29622 13124 29627 13244
rect 29627 13124 29673 13244
rect 29673 13124 29678 13244
rect 29162 13005 29163 13048
rect 29163 13005 29217 13048
rect 29217 13005 29218 13048
rect 29162 12992 29218 13005
rect 29346 13005 29347 13048
rect 29347 13005 29401 13048
rect 29401 13005 29402 13048
rect 29346 12992 29402 13005
rect 29530 13005 29531 13048
rect 29531 13005 29585 13048
rect 29585 13005 29586 13048
rect 29530 12992 29586 13005
rect 29162 12842 29218 12898
rect 30924 13812 30980 13868
rect 30556 13425 30561 13545
rect 30561 13425 30607 13545
rect 30607 13425 30612 13545
rect 30924 13425 30929 13545
rect 30929 13425 30975 13545
rect 30975 13425 30980 13545
rect 30740 13125 30745 13245
rect 30745 13125 30791 13245
rect 30791 13125 30796 13245
rect 31246 13424 31251 13545
rect 31251 13424 31297 13545
rect 31297 13424 31302 13545
rect 31108 13125 31113 13245
rect 31113 13125 31159 13245
rect 31159 13125 31164 13245
rect 30648 13006 30649 13049
rect 30649 13006 30703 13049
rect 30703 13006 30704 13049
rect 30648 12993 30704 13006
rect 30832 13006 30833 13049
rect 30833 13006 30887 13049
rect 30887 13006 30888 13049
rect 30832 12993 30888 13006
rect 31016 13006 31017 13049
rect 31017 13006 31071 13049
rect 31071 13006 31072 13049
rect 31016 12993 31072 13006
rect 30648 12843 30704 12899
rect 29346 12726 29402 12782
rect 29675 12726 29731 12782
rect 29932 12726 29988 12782
rect 30832 12727 30888 12783
rect 31161 12727 31217 12783
rect 31594 12727 31650 12783
rect 4238 12613 4294 12669
rect 5278 12613 5334 12669
rect 6764 12614 6820 12670
rect 4910 12506 4966 12519
rect 4910 12463 4911 12506
rect 4911 12463 4965 12506
rect 4965 12463 4966 12506
rect 5094 12506 5150 12519
rect 5094 12463 5095 12506
rect 5095 12463 5149 12506
rect 5149 12463 5150 12506
rect 5278 12506 5334 12519
rect 5278 12463 5279 12506
rect 5279 12463 5333 12506
rect 5333 12463 5334 12506
rect 5370 12267 5375 12387
rect 5375 12267 5421 12387
rect 5421 12267 5426 12387
rect 4685 11944 4741 12000
rect 5503 11944 5559 12000
rect 5856 11826 5912 11882
rect 5680 11718 5736 11772
rect 5186 11609 5242 11665
rect 4818 11222 4823 11342
rect 4823 11222 4869 11342
rect 4869 11222 4874 11342
rect 5186 11222 5191 11342
rect 5191 11222 5237 11342
rect 5237 11222 5242 11342
rect 5002 10922 5007 11042
rect 5007 10922 5053 11042
rect 5053 10922 5058 11042
rect 5508 11221 5513 11342
rect 5513 11221 5559 11342
rect 5559 11221 5564 11342
rect 5370 10922 5375 11042
rect 5375 10922 5421 11042
rect 5421 10922 5426 11042
rect 4910 10803 4911 10846
rect 4911 10803 4965 10846
rect 4965 10803 4966 10846
rect 4910 10790 4966 10803
rect 5094 10803 5095 10846
rect 5095 10803 5149 10846
rect 5149 10803 5150 10846
rect 5094 10790 5150 10803
rect 5278 10803 5279 10846
rect 5279 10803 5333 10846
rect 5333 10803 5334 10846
rect 5278 10790 5334 10803
rect 4910 10640 4966 10696
rect 4102 10524 4158 10580
rect 5094 10524 5150 10580
rect 5423 10524 5479 10580
rect 5856 10524 5912 10580
rect 3286 10408 3342 10464
rect 5278 10408 5334 10464
rect 4910 10301 4966 10314
rect 4910 10258 4911 10301
rect 4911 10258 4965 10301
rect 4965 10258 4966 10301
rect 5094 10301 5150 10314
rect 5094 10258 5095 10301
rect 5095 10258 5149 10301
rect 5149 10258 5150 10301
rect 5278 10301 5334 10314
rect 5278 10258 5279 10301
rect 5279 10258 5333 10301
rect 5333 10258 5334 10301
rect 5370 10062 5375 10182
rect 5375 10062 5421 10182
rect 5421 10062 5426 10182
rect 4685 9739 4741 9795
rect 5503 9739 5559 9795
rect 8280 12610 8336 12666
rect 9320 12610 9376 12666
rect 6396 12507 6452 12520
rect 6396 12464 6397 12507
rect 6397 12464 6451 12507
rect 6451 12464 6452 12507
rect 6580 12507 6636 12520
rect 6580 12464 6581 12507
rect 6581 12464 6635 12507
rect 6635 12464 6636 12507
rect 6764 12507 6820 12520
rect 6764 12464 6765 12507
rect 6765 12464 6819 12507
rect 6819 12464 6820 12507
rect 6856 12268 6861 12388
rect 6861 12268 6907 12388
rect 6907 12268 6912 12388
rect 6171 11945 6227 12001
rect 6989 11945 7045 12001
rect 10806 12611 10862 12667
rect 8952 12503 9008 12516
rect 8952 12460 8953 12503
rect 8953 12460 9007 12503
rect 9007 12460 9008 12503
rect 9136 12503 9192 12516
rect 9136 12460 9137 12503
rect 9137 12460 9191 12503
rect 9191 12460 9192 12503
rect 9320 12503 9376 12516
rect 9320 12460 9321 12503
rect 9321 12460 9375 12503
rect 9375 12460 9376 12503
rect 9412 12264 9417 12384
rect 9417 12264 9463 12384
rect 9463 12264 9468 12384
rect 8727 11941 8783 11997
rect 9545 11941 9601 11997
rect 9898 11823 9954 11879
rect 9722 11715 9778 11769
rect 9228 11606 9284 11662
rect 8860 11219 8865 11339
rect 8865 11219 8911 11339
rect 8911 11219 8916 11339
rect 9228 11219 9233 11339
rect 9233 11219 9279 11339
rect 9279 11219 9284 11339
rect 9044 10919 9049 11039
rect 9049 10919 9095 11039
rect 9095 10919 9100 11039
rect 9550 11218 9555 11339
rect 9555 11218 9601 11339
rect 9601 11218 9606 11339
rect 9412 10919 9417 11039
rect 9417 10919 9463 11039
rect 9463 10919 9468 11039
rect 8952 10800 8953 10843
rect 8953 10800 9007 10843
rect 9007 10800 9008 10843
rect 8952 10787 9008 10800
rect 9136 10800 9137 10843
rect 9137 10800 9191 10843
rect 9191 10800 9192 10843
rect 9136 10787 9192 10800
rect 9320 10800 9321 10843
rect 9321 10800 9375 10843
rect 9375 10800 9376 10843
rect 9320 10787 9376 10800
rect 8952 10637 9008 10693
rect 8144 10521 8200 10577
rect 9136 10521 9192 10577
rect 9465 10521 9521 10577
rect 9898 10521 9954 10577
rect 7298 10405 7354 10461
rect 9320 10405 9376 10461
rect 8952 10298 9008 10311
rect 8952 10255 8953 10298
rect 8953 10255 9007 10298
rect 9007 10255 9008 10298
rect 9136 10298 9192 10311
rect 9136 10255 9137 10298
rect 9137 10255 9191 10298
rect 9191 10255 9192 10298
rect 9320 10298 9376 10311
rect 9320 10255 9321 10298
rect 9321 10255 9375 10298
rect 9375 10255 9376 10298
rect 9412 10059 9417 10179
rect 9417 10059 9463 10179
rect 9463 10059 9468 10179
rect 8727 9736 8783 9792
rect 9545 9736 9601 9792
rect 3830 9621 3886 9677
rect 4102 9621 4158 9677
rect 12322 12610 12378 12666
rect 13362 12610 13418 12666
rect 10438 12504 10494 12517
rect 10438 12461 10439 12504
rect 10439 12461 10493 12504
rect 10493 12461 10494 12504
rect 10622 12504 10678 12517
rect 10622 12461 10623 12504
rect 10623 12461 10677 12504
rect 10677 12461 10678 12504
rect 10806 12504 10862 12517
rect 10806 12461 10807 12504
rect 10807 12461 10861 12504
rect 10861 12461 10862 12504
rect 10898 12265 10903 12385
rect 10903 12265 10949 12385
rect 10949 12265 10954 12385
rect 10213 11942 10269 11998
rect 11031 11942 11087 11998
rect 14848 12611 14904 12667
rect 12994 12503 13050 12516
rect 12994 12460 12995 12503
rect 12995 12460 13049 12503
rect 13049 12460 13050 12503
rect 13178 12503 13234 12516
rect 13178 12460 13179 12503
rect 13179 12460 13233 12503
rect 13233 12460 13234 12503
rect 13362 12503 13418 12516
rect 13362 12460 13363 12503
rect 13363 12460 13417 12503
rect 13417 12460 13418 12503
rect 13454 12264 13459 12384
rect 13459 12264 13505 12384
rect 13505 12264 13510 12384
rect 12769 11941 12825 11997
rect 13587 11941 13643 11997
rect 13940 11823 13996 11879
rect 13764 11715 13820 11769
rect 13270 11606 13326 11662
rect 12902 11219 12907 11339
rect 12907 11219 12953 11339
rect 12953 11219 12958 11339
rect 13270 11219 13275 11339
rect 13275 11219 13321 11339
rect 13321 11219 13326 11339
rect 13086 10919 13091 11039
rect 13091 10919 13137 11039
rect 13137 10919 13142 11039
rect 13592 11218 13597 11339
rect 13597 11218 13643 11339
rect 13643 11218 13648 11339
rect 13454 10919 13459 11039
rect 13459 10919 13505 11039
rect 13505 10919 13510 11039
rect 12994 10800 12995 10843
rect 12995 10800 13049 10843
rect 13049 10800 13050 10843
rect 12994 10787 13050 10800
rect 13178 10800 13179 10843
rect 13179 10800 13233 10843
rect 13233 10800 13234 10843
rect 13178 10787 13234 10800
rect 13362 10800 13363 10843
rect 13363 10800 13417 10843
rect 13417 10800 13418 10843
rect 13362 10787 13418 10800
rect 12994 10637 13050 10693
rect 12186 10521 12242 10577
rect 13178 10521 13234 10577
rect 13507 10521 13563 10577
rect 13940 10521 13996 10577
rect 11340 10405 11396 10461
rect 13362 10405 13418 10461
rect 12994 10298 13050 10311
rect 12994 10255 12995 10298
rect 12995 10255 13049 10298
rect 13049 10255 13050 10298
rect 13178 10298 13234 10311
rect 13178 10255 13179 10298
rect 13179 10255 13233 10298
rect 13233 10255 13234 10298
rect 13362 10298 13418 10311
rect 13362 10255 13363 10298
rect 13363 10255 13417 10298
rect 13417 10255 13418 10298
rect 13454 10059 13459 10179
rect 13459 10059 13505 10179
rect 13505 10059 13510 10179
rect 12769 9736 12825 9792
rect 13587 9736 13643 9792
rect 7842 9618 7898 9674
rect 8144 9618 8200 9674
rect 16364 12610 16420 12666
rect 17404 12610 17460 12666
rect 14480 12504 14536 12517
rect 14480 12461 14481 12504
rect 14481 12461 14535 12504
rect 14535 12461 14536 12504
rect 14664 12504 14720 12517
rect 14664 12461 14665 12504
rect 14665 12461 14719 12504
rect 14719 12461 14720 12504
rect 14848 12504 14904 12517
rect 14848 12461 14849 12504
rect 14849 12461 14903 12504
rect 14903 12461 14904 12504
rect 14940 12265 14945 12385
rect 14945 12265 14991 12385
rect 14991 12265 14996 12385
rect 14255 11942 14311 11998
rect 15073 11942 15129 11998
rect 18890 12611 18946 12667
rect 17036 12503 17092 12516
rect 17036 12460 17037 12503
rect 17037 12460 17091 12503
rect 17091 12460 17092 12503
rect 17220 12503 17276 12516
rect 17220 12460 17221 12503
rect 17221 12460 17275 12503
rect 17275 12460 17276 12503
rect 17404 12503 17460 12516
rect 17404 12460 17405 12503
rect 17405 12460 17459 12503
rect 17459 12460 17460 12503
rect 17496 12264 17501 12384
rect 17501 12264 17547 12384
rect 17547 12264 17552 12384
rect 16811 11941 16867 11997
rect 17629 11941 17685 11997
rect 17982 11823 18038 11879
rect 17806 11715 17862 11769
rect 17312 11606 17368 11662
rect 16944 11219 16949 11339
rect 16949 11219 16995 11339
rect 16995 11219 17000 11339
rect 17312 11219 17317 11339
rect 17317 11219 17363 11339
rect 17363 11219 17368 11339
rect 17128 10919 17133 11039
rect 17133 10919 17179 11039
rect 17179 10919 17184 11039
rect 17634 11218 17639 11339
rect 17639 11218 17685 11339
rect 17685 11218 17690 11339
rect 17496 10919 17501 11039
rect 17501 10919 17547 11039
rect 17547 10919 17552 11039
rect 17036 10800 17037 10843
rect 17037 10800 17091 10843
rect 17091 10800 17092 10843
rect 17036 10787 17092 10800
rect 17220 10800 17221 10843
rect 17221 10800 17275 10843
rect 17275 10800 17276 10843
rect 17220 10787 17276 10800
rect 17404 10800 17405 10843
rect 17405 10800 17459 10843
rect 17459 10800 17460 10843
rect 17404 10787 17460 10800
rect 17036 10637 17092 10693
rect 16228 10521 16284 10577
rect 17220 10521 17276 10577
rect 17549 10521 17605 10577
rect 17982 10521 18038 10577
rect 15382 10405 15438 10461
rect 17404 10405 17460 10461
rect 17036 10298 17092 10311
rect 17036 10255 17037 10298
rect 17037 10255 17091 10298
rect 17091 10255 17092 10298
rect 17220 10298 17276 10311
rect 17220 10255 17221 10298
rect 17221 10255 17275 10298
rect 17275 10255 17276 10298
rect 17404 10298 17460 10311
rect 17404 10255 17405 10298
rect 17405 10255 17459 10298
rect 17459 10255 17460 10298
rect 17496 10059 17501 10179
rect 17501 10059 17547 10179
rect 17547 10059 17552 10179
rect 16811 9736 16867 9792
rect 17629 9736 17685 9792
rect 11884 9618 11940 9674
rect 12186 9618 12242 9674
rect 20406 12610 20462 12666
rect 21446 12610 21502 12666
rect 18522 12504 18578 12517
rect 18522 12461 18523 12504
rect 18523 12461 18577 12504
rect 18577 12461 18578 12504
rect 18706 12504 18762 12517
rect 18706 12461 18707 12504
rect 18707 12461 18761 12504
rect 18761 12461 18762 12504
rect 18890 12504 18946 12517
rect 18890 12461 18891 12504
rect 18891 12461 18945 12504
rect 18945 12461 18946 12504
rect 18982 12265 18987 12385
rect 18987 12265 19033 12385
rect 19033 12265 19038 12385
rect 18297 11942 18353 11998
rect 19115 11942 19171 11998
rect 22932 12611 22988 12667
rect 21078 12503 21134 12516
rect 21078 12460 21079 12503
rect 21079 12460 21133 12503
rect 21133 12460 21134 12503
rect 21262 12503 21318 12516
rect 21262 12460 21263 12503
rect 21263 12460 21317 12503
rect 21317 12460 21318 12503
rect 21446 12503 21502 12516
rect 21446 12460 21447 12503
rect 21447 12460 21501 12503
rect 21501 12460 21502 12503
rect 21538 12264 21543 12384
rect 21543 12264 21589 12384
rect 21589 12264 21594 12384
rect 20853 11941 20909 11997
rect 21671 11941 21727 11997
rect 22024 11823 22080 11879
rect 21848 11715 21904 11769
rect 21354 11606 21410 11662
rect 20986 11219 20991 11339
rect 20991 11219 21037 11339
rect 21037 11219 21042 11339
rect 21354 11219 21359 11339
rect 21359 11219 21405 11339
rect 21405 11219 21410 11339
rect 21170 10919 21175 11039
rect 21175 10919 21221 11039
rect 21221 10919 21226 11039
rect 21676 11218 21681 11339
rect 21681 11218 21727 11339
rect 21727 11218 21732 11339
rect 21538 10919 21543 11039
rect 21543 10919 21589 11039
rect 21589 10919 21594 11039
rect 21078 10800 21079 10843
rect 21079 10800 21133 10843
rect 21133 10800 21134 10843
rect 21078 10787 21134 10800
rect 21262 10800 21263 10843
rect 21263 10800 21317 10843
rect 21317 10800 21318 10843
rect 21262 10787 21318 10800
rect 21446 10800 21447 10843
rect 21447 10800 21501 10843
rect 21501 10800 21502 10843
rect 21446 10787 21502 10800
rect 21078 10637 21134 10693
rect 20270 10521 20326 10577
rect 21262 10521 21318 10577
rect 21591 10521 21647 10577
rect 22024 10521 22080 10577
rect 19424 10405 19480 10461
rect 21446 10405 21502 10461
rect 21078 10298 21134 10311
rect 21078 10255 21079 10298
rect 21079 10255 21133 10298
rect 21133 10255 21134 10298
rect 21262 10298 21318 10311
rect 21262 10255 21263 10298
rect 21263 10255 21317 10298
rect 21317 10255 21318 10298
rect 21446 10298 21502 10311
rect 21446 10255 21447 10298
rect 21447 10255 21501 10298
rect 21501 10255 21502 10298
rect 21538 10059 21543 10179
rect 21543 10059 21589 10179
rect 21589 10059 21594 10179
rect 20853 9736 20909 9792
rect 21671 9736 21727 9792
rect 15926 9618 15982 9674
rect 16228 9618 16284 9674
rect 24448 12610 24504 12666
rect 25488 12610 25544 12666
rect 22564 12504 22620 12517
rect 22564 12461 22565 12504
rect 22565 12461 22619 12504
rect 22619 12461 22620 12504
rect 22748 12504 22804 12517
rect 22748 12461 22749 12504
rect 22749 12461 22803 12504
rect 22803 12461 22804 12504
rect 22932 12504 22988 12517
rect 22932 12461 22933 12504
rect 22933 12461 22987 12504
rect 22987 12461 22988 12504
rect 23024 12265 23029 12385
rect 23029 12265 23075 12385
rect 23075 12265 23080 12385
rect 22339 11942 22395 11998
rect 23157 11942 23213 11998
rect 26974 12611 27030 12667
rect 25120 12503 25176 12516
rect 25120 12460 25121 12503
rect 25121 12460 25175 12503
rect 25175 12460 25176 12503
rect 25304 12503 25360 12516
rect 25304 12460 25305 12503
rect 25305 12460 25359 12503
rect 25359 12460 25360 12503
rect 25488 12503 25544 12516
rect 25488 12460 25489 12503
rect 25489 12460 25543 12503
rect 25543 12460 25544 12503
rect 25580 12264 25585 12384
rect 25585 12264 25631 12384
rect 25631 12264 25636 12384
rect 24895 11941 24951 11997
rect 25713 11941 25769 11997
rect 26066 11823 26122 11879
rect 25890 11715 25946 11769
rect 25396 11606 25452 11662
rect 25028 11219 25033 11339
rect 25033 11219 25079 11339
rect 25079 11219 25084 11339
rect 25396 11219 25401 11339
rect 25401 11219 25447 11339
rect 25447 11219 25452 11339
rect 25212 10919 25217 11039
rect 25217 10919 25263 11039
rect 25263 10919 25268 11039
rect 25718 11218 25723 11339
rect 25723 11218 25769 11339
rect 25769 11218 25774 11339
rect 25580 10919 25585 11039
rect 25585 10919 25631 11039
rect 25631 10919 25636 11039
rect 25120 10800 25121 10843
rect 25121 10800 25175 10843
rect 25175 10800 25176 10843
rect 25120 10787 25176 10800
rect 25304 10800 25305 10843
rect 25305 10800 25359 10843
rect 25359 10800 25360 10843
rect 25304 10787 25360 10800
rect 25488 10800 25489 10843
rect 25489 10800 25543 10843
rect 25543 10800 25544 10843
rect 25488 10787 25544 10800
rect 25120 10637 25176 10693
rect 24312 10521 24368 10577
rect 25304 10521 25360 10577
rect 25633 10521 25689 10577
rect 26066 10521 26122 10577
rect 23466 10405 23522 10461
rect 25488 10405 25544 10461
rect 25120 10298 25176 10311
rect 25120 10255 25121 10298
rect 25121 10255 25175 10298
rect 25175 10255 25176 10298
rect 25304 10298 25360 10311
rect 25304 10255 25305 10298
rect 25305 10255 25359 10298
rect 25359 10255 25360 10298
rect 25488 10298 25544 10311
rect 25488 10255 25489 10298
rect 25489 10255 25543 10298
rect 25543 10255 25544 10298
rect 25580 10059 25585 10179
rect 25585 10059 25631 10179
rect 25631 10059 25636 10179
rect 24895 9736 24951 9792
rect 25713 9736 25769 9792
rect 19968 9618 20024 9674
rect 20270 9618 20326 9674
rect 28490 12610 28546 12666
rect 29530 12610 29586 12666
rect 26606 12504 26662 12517
rect 26606 12461 26607 12504
rect 26607 12461 26661 12504
rect 26661 12461 26662 12504
rect 26790 12504 26846 12517
rect 26790 12461 26791 12504
rect 26791 12461 26845 12504
rect 26845 12461 26846 12504
rect 26974 12504 27030 12517
rect 26974 12461 26975 12504
rect 26975 12461 27029 12504
rect 27029 12461 27030 12504
rect 27066 12265 27071 12385
rect 27071 12265 27117 12385
rect 27117 12265 27122 12385
rect 26381 11942 26437 11998
rect 27199 11942 27255 11998
rect 31016 12611 31072 12667
rect 29162 12503 29218 12516
rect 29162 12460 29163 12503
rect 29163 12460 29217 12503
rect 29217 12460 29218 12503
rect 29346 12503 29402 12516
rect 29346 12460 29347 12503
rect 29347 12460 29401 12503
rect 29401 12460 29402 12503
rect 29530 12503 29586 12516
rect 29530 12460 29531 12503
rect 29531 12460 29585 12503
rect 29585 12460 29586 12503
rect 29622 12264 29627 12384
rect 29627 12264 29673 12384
rect 29673 12264 29678 12384
rect 28937 11941 28993 11997
rect 29755 11941 29811 11997
rect 30108 11823 30164 11879
rect 29932 11715 29988 11769
rect 29438 11606 29494 11662
rect 29070 11219 29075 11339
rect 29075 11219 29121 11339
rect 29121 11219 29126 11339
rect 29438 11219 29443 11339
rect 29443 11219 29489 11339
rect 29489 11219 29494 11339
rect 29254 10919 29259 11039
rect 29259 10919 29305 11039
rect 29305 10919 29310 11039
rect 29760 11218 29765 11339
rect 29765 11218 29811 11339
rect 29811 11218 29816 11339
rect 29622 10919 29627 11039
rect 29627 10919 29673 11039
rect 29673 10919 29678 11039
rect 29162 10800 29163 10843
rect 29163 10800 29217 10843
rect 29217 10800 29218 10843
rect 29162 10787 29218 10800
rect 29346 10800 29347 10843
rect 29347 10800 29401 10843
rect 29401 10800 29402 10843
rect 29346 10787 29402 10800
rect 29530 10800 29531 10843
rect 29531 10800 29585 10843
rect 29585 10800 29586 10843
rect 29530 10787 29586 10800
rect 29162 10637 29218 10693
rect 28354 10521 28410 10577
rect 29346 10521 29402 10577
rect 29675 10521 29731 10577
rect 30108 10521 30164 10577
rect 28173 10405 28229 10461
rect 29530 10405 29586 10461
rect 29162 10298 29218 10311
rect 29162 10255 29163 10298
rect 29163 10255 29217 10298
rect 29217 10255 29218 10298
rect 29346 10298 29402 10311
rect 29346 10255 29347 10298
rect 29347 10255 29401 10298
rect 29401 10255 29402 10298
rect 29530 10298 29586 10311
rect 29530 10255 29531 10298
rect 29531 10255 29585 10298
rect 29585 10255 29586 10298
rect 29622 10059 29627 10179
rect 29627 10059 29673 10179
rect 29673 10059 29678 10179
rect 28937 9736 28993 9792
rect 29755 9736 29811 9792
rect 24010 9618 24066 9674
rect 24312 9618 24368 9674
rect 30648 12504 30704 12517
rect 30648 12461 30649 12504
rect 30649 12461 30703 12504
rect 30703 12461 30704 12504
rect 30832 12504 30888 12517
rect 30832 12461 30833 12504
rect 30833 12461 30887 12504
rect 30887 12461 30888 12504
rect 31016 12504 31072 12517
rect 31016 12461 31017 12504
rect 31017 12461 31071 12504
rect 31071 12461 31072 12504
rect 31108 12265 31113 12385
rect 31113 12265 31159 12385
rect 31159 12265 31164 12385
rect 30423 11942 30479 11998
rect 31241 11942 31297 11998
rect 28052 9618 28108 9674
rect 28354 9618 28410 9674
rect 1174 8645 1230 8701
rect 806 8258 811 8378
rect 811 8258 857 8378
rect 857 8258 862 8378
rect 1174 8258 1179 8378
rect 1179 8258 1225 8378
rect 1225 8258 1230 8378
rect 990 7958 995 8078
rect 995 7958 1041 8078
rect 1041 7958 1046 8078
rect 1496 8257 1501 8378
rect 1501 8257 1547 8378
rect 1547 8257 1552 8378
rect 1358 7958 1363 8078
rect 1363 7958 1409 8078
rect 1409 7958 1414 8078
rect 898 7839 899 7882
rect 899 7839 953 7882
rect 953 7839 954 7882
rect 898 7826 954 7839
rect 1082 7839 1083 7882
rect 1083 7839 1137 7882
rect 1137 7839 1138 7882
rect 1082 7826 1138 7839
rect 1266 7839 1267 7882
rect 1267 7839 1321 7882
rect 1321 7839 1322 7882
rect 1266 7826 1322 7839
rect -46 7676 10 7732
rect 898 7676 954 7732
rect 226 7560 282 7616
rect 1082 7560 1138 7616
rect 1411 7560 1467 7616
rect 1668 7560 1724 7616
rect 1266 7444 1322 7500
rect 898 7337 954 7350
rect 898 7294 899 7337
rect 899 7294 953 7337
rect 953 7294 954 7337
rect 1082 7337 1138 7350
rect 1082 7294 1083 7337
rect 1083 7294 1137 7337
rect 1137 7294 1138 7337
rect 1266 7337 1322 7350
rect 1266 7294 1267 7337
rect 1267 7294 1321 7337
rect 1321 7294 1322 7337
rect 1358 7098 1363 7218
rect 1363 7098 1409 7218
rect 1409 7098 1414 7218
rect 673 6775 729 6831
rect 1491 6775 1547 6831
rect 1844 6657 1900 6713
rect 1668 6549 1724 6603
rect 1174 6440 1230 6496
rect 806 6053 811 6173
rect 811 6053 857 6173
rect 857 6053 862 6173
rect 1174 6053 1179 6173
rect 1179 6053 1225 6173
rect 1225 6053 1230 6173
rect 990 5753 995 5873
rect 995 5753 1041 5873
rect 1041 5753 1046 5873
rect 1496 6052 1501 6173
rect 1501 6052 1547 6173
rect 1547 6052 1552 6173
rect 1358 5753 1363 5873
rect 1363 5753 1409 5873
rect 1409 5753 1414 5873
rect 898 5634 899 5677
rect 899 5634 953 5677
rect 953 5634 954 5677
rect 898 5621 954 5634
rect 1082 5634 1083 5677
rect 1083 5634 1137 5677
rect 1137 5634 1138 5677
rect 1082 5621 1138 5634
rect 1266 5634 1267 5677
rect 1267 5634 1321 5677
rect 1321 5634 1322 5677
rect 1266 5621 1322 5634
rect 898 5471 954 5527
rect 5186 8645 5242 8701
rect 4818 8258 4823 8378
rect 4823 8258 4869 8378
rect 4869 8258 4874 8378
rect 5186 8258 5191 8378
rect 5191 8258 5237 8378
rect 5237 8258 5242 8378
rect 5002 7958 5007 8078
rect 5007 7958 5053 8078
rect 5053 7958 5058 8078
rect 5508 8257 5513 8378
rect 5513 8257 5559 8378
rect 5559 8257 5564 8378
rect 5370 7958 5375 8078
rect 5375 7958 5421 8078
rect 5421 7958 5426 8078
rect 4910 7839 4911 7882
rect 4911 7839 4965 7882
rect 4965 7839 4966 7882
rect 4910 7826 4966 7839
rect 5094 7839 5095 7882
rect 5095 7839 5149 7882
rect 5149 7839 5150 7882
rect 5094 7826 5150 7839
rect 5278 7839 5279 7882
rect 5279 7839 5333 7882
rect 5333 7839 5334 7882
rect 5278 7826 5334 7839
rect 4022 7676 4078 7732
rect 4910 7676 4966 7732
rect 4238 7560 4294 7616
rect 5094 7560 5150 7616
rect 5423 7560 5479 7616
rect 5680 7560 5736 7616
rect 5278 7444 5334 7500
rect 4910 7337 4966 7350
rect 4910 7294 4911 7337
rect 4911 7294 4965 7337
rect 4965 7294 4966 7337
rect 5094 7337 5150 7350
rect 5094 7294 5095 7337
rect 5095 7294 5149 7337
rect 5149 7294 5150 7337
rect 5278 7337 5334 7350
rect 5278 7294 5279 7337
rect 5279 7294 5333 7337
rect 5333 7294 5334 7337
rect 5370 7098 5375 7218
rect 5375 7098 5421 7218
rect 5421 7098 5426 7218
rect 4685 6775 4741 6831
rect 5503 6775 5559 6831
rect 5856 6657 5912 6713
rect 5680 6549 5736 6603
rect 2660 6440 2716 6496
rect 2292 6053 2297 6173
rect 2297 6053 2343 6173
rect 2343 6053 2348 6173
rect 2660 6053 2665 6173
rect 2665 6053 2711 6173
rect 2711 6053 2716 6173
rect 2476 5753 2481 5873
rect 2481 5753 2527 5873
rect 2527 5753 2532 5873
rect 2982 6052 2987 6173
rect 2987 6052 3033 6173
rect 3033 6052 3038 6173
rect 2844 5753 2849 5873
rect 2849 5753 2895 5873
rect 2895 5753 2900 5873
rect 2384 5634 2385 5677
rect 2385 5634 2439 5677
rect 2439 5634 2440 5677
rect 2384 5621 2440 5634
rect 2568 5634 2569 5677
rect 2569 5634 2623 5677
rect 2623 5634 2624 5677
rect 2568 5621 2624 5634
rect 2752 5634 2753 5677
rect 2753 5634 2807 5677
rect 2807 5634 2808 5677
rect 2752 5621 2808 5634
rect 2384 5471 2440 5527
rect 5186 6440 5242 6496
rect 4818 6053 4823 6173
rect 4823 6053 4869 6173
rect 4869 6053 4874 6173
rect 5186 6053 5191 6173
rect 5191 6053 5237 6173
rect 5237 6053 5242 6173
rect 5002 5753 5007 5873
rect 5007 5753 5053 5873
rect 5053 5753 5058 5873
rect 5508 6052 5513 6173
rect 5513 6052 5559 6173
rect 5559 6052 5564 6173
rect 5370 5753 5375 5873
rect 5375 5753 5421 5873
rect 5421 5753 5426 5873
rect 4910 5634 4911 5677
rect 4911 5634 4965 5677
rect 4965 5634 4966 5677
rect 4910 5621 4966 5634
rect 5094 5634 5095 5677
rect 5095 5634 5149 5677
rect 5149 5634 5150 5677
rect 5094 5621 5150 5634
rect 5278 5634 5279 5677
rect 5279 5634 5333 5677
rect 5333 5634 5334 5677
rect 5278 5621 5334 5634
rect 4910 5471 4966 5527
rect 9228 8645 9284 8701
rect 8860 8258 8865 8378
rect 8865 8258 8911 8378
rect 8911 8258 8916 8378
rect 9228 8258 9233 8378
rect 9233 8258 9279 8378
rect 9279 8258 9284 8378
rect 9044 7958 9049 8078
rect 9049 7958 9095 8078
rect 9095 7958 9100 8078
rect 9550 8257 9555 8378
rect 9555 8257 9601 8378
rect 9601 8257 9606 8378
rect 9412 7958 9417 8078
rect 9417 7958 9463 8078
rect 9463 7958 9468 8078
rect 8952 7839 8953 7882
rect 8953 7839 9007 7882
rect 9007 7839 9008 7882
rect 8952 7826 9008 7839
rect 9136 7839 9137 7882
rect 9137 7839 9191 7882
rect 9191 7839 9192 7882
rect 9136 7826 9192 7839
rect 9320 7839 9321 7882
rect 9321 7839 9375 7882
rect 9375 7839 9376 7882
rect 9320 7826 9376 7839
rect 8064 7676 8120 7732
rect 8952 7676 9008 7732
rect 8280 7560 8336 7616
rect 9136 7560 9192 7616
rect 9465 7560 9521 7616
rect 9722 7560 9778 7616
rect 9320 7444 9376 7500
rect 8952 7337 9008 7350
rect 8952 7294 8953 7337
rect 8953 7294 9007 7337
rect 9007 7294 9008 7337
rect 9136 7337 9192 7350
rect 9136 7294 9137 7337
rect 9137 7294 9191 7337
rect 9191 7294 9192 7337
rect 9320 7337 9376 7350
rect 9320 7294 9321 7337
rect 9321 7294 9375 7337
rect 9375 7294 9376 7337
rect 9412 7098 9417 7218
rect 9417 7098 9463 7218
rect 9463 7098 9468 7218
rect 8727 6775 8783 6831
rect 9545 6775 9601 6831
rect 9898 6657 9954 6713
rect 9722 6549 9778 6603
rect 6672 6440 6728 6496
rect 6304 6053 6309 6173
rect 6309 6053 6355 6173
rect 6355 6053 6360 6173
rect 6672 6053 6677 6173
rect 6677 6053 6723 6173
rect 6723 6053 6728 6173
rect 6488 5753 6493 5873
rect 6493 5753 6539 5873
rect 6539 5753 6544 5873
rect 6994 6052 6999 6173
rect 6999 6052 7045 6173
rect 7045 6052 7050 6173
rect 6856 5753 6861 5873
rect 6861 5753 6907 5873
rect 6907 5753 6912 5873
rect 6396 5634 6397 5677
rect 6397 5634 6451 5677
rect 6451 5634 6452 5677
rect 6396 5621 6452 5634
rect 6580 5634 6581 5677
rect 6581 5634 6635 5677
rect 6635 5634 6636 5677
rect 6580 5621 6636 5634
rect 6764 5634 6765 5677
rect 6765 5634 6819 5677
rect 6819 5634 6820 5677
rect 6764 5621 6820 5634
rect 6396 5471 6452 5527
rect 9228 6440 9284 6496
rect 8860 6053 8865 6173
rect 8865 6053 8911 6173
rect 8911 6053 8916 6173
rect 9228 6053 9233 6173
rect 9233 6053 9279 6173
rect 9279 6053 9284 6173
rect 9044 5753 9049 5873
rect 9049 5753 9095 5873
rect 9095 5753 9100 5873
rect 9550 6052 9555 6173
rect 9555 6052 9601 6173
rect 9601 6052 9606 6173
rect 9412 5753 9417 5873
rect 9417 5753 9463 5873
rect 9463 5753 9468 5873
rect 8952 5634 8953 5677
rect 8953 5634 9007 5677
rect 9007 5634 9008 5677
rect 8952 5621 9008 5634
rect 9136 5634 9137 5677
rect 9137 5634 9191 5677
rect 9191 5634 9192 5677
rect 9136 5621 9192 5634
rect 9320 5634 9321 5677
rect 9321 5634 9375 5677
rect 9375 5634 9376 5677
rect 9320 5621 9376 5634
rect 8952 5471 9008 5527
rect 13270 8645 13326 8701
rect 12902 8258 12907 8378
rect 12907 8258 12953 8378
rect 12953 8258 12958 8378
rect 13270 8258 13275 8378
rect 13275 8258 13321 8378
rect 13321 8258 13326 8378
rect 13086 7958 13091 8078
rect 13091 7958 13137 8078
rect 13137 7958 13142 8078
rect 13592 8257 13597 8378
rect 13597 8257 13643 8378
rect 13643 8257 13648 8378
rect 13454 7958 13459 8078
rect 13459 7958 13505 8078
rect 13505 7958 13510 8078
rect 12994 7839 12995 7882
rect 12995 7839 13049 7882
rect 13049 7839 13050 7882
rect 12994 7826 13050 7839
rect 13178 7839 13179 7882
rect 13179 7839 13233 7882
rect 13233 7839 13234 7882
rect 13178 7826 13234 7839
rect 13362 7839 13363 7882
rect 13363 7839 13417 7882
rect 13417 7839 13418 7882
rect 13362 7826 13418 7839
rect 12106 7676 12162 7732
rect 12994 7676 13050 7732
rect 12322 7560 12378 7616
rect 13178 7560 13234 7616
rect 13507 7560 13563 7616
rect 13764 7560 13820 7616
rect 13362 7444 13418 7500
rect 12994 7337 13050 7350
rect 12994 7294 12995 7337
rect 12995 7294 13049 7337
rect 13049 7294 13050 7337
rect 13178 7337 13234 7350
rect 13178 7294 13179 7337
rect 13179 7294 13233 7337
rect 13233 7294 13234 7337
rect 13362 7337 13418 7350
rect 13362 7294 13363 7337
rect 13363 7294 13417 7337
rect 13417 7294 13418 7337
rect 13454 7098 13459 7218
rect 13459 7098 13505 7218
rect 13505 7098 13510 7218
rect 12769 6775 12825 6831
rect 13587 6775 13643 6831
rect 13940 6657 13996 6713
rect 13764 6549 13820 6603
rect 10714 6440 10770 6496
rect 10346 6053 10351 6173
rect 10351 6053 10397 6173
rect 10397 6053 10402 6173
rect 10714 6053 10719 6173
rect 10719 6053 10765 6173
rect 10765 6053 10770 6173
rect 10530 5753 10535 5873
rect 10535 5753 10581 5873
rect 10581 5753 10586 5873
rect 11036 6052 11041 6173
rect 11041 6052 11087 6173
rect 11087 6052 11092 6173
rect 10898 5753 10903 5873
rect 10903 5753 10949 5873
rect 10949 5753 10954 5873
rect 10438 5634 10439 5677
rect 10439 5634 10493 5677
rect 10493 5634 10494 5677
rect 10438 5621 10494 5634
rect 10622 5634 10623 5677
rect 10623 5634 10677 5677
rect 10677 5634 10678 5677
rect 10622 5621 10678 5634
rect 10806 5634 10807 5677
rect 10807 5634 10861 5677
rect 10861 5634 10862 5677
rect 10806 5621 10862 5634
rect 10438 5471 10494 5527
rect 13270 6440 13326 6496
rect 12902 6053 12907 6173
rect 12907 6053 12953 6173
rect 12953 6053 12958 6173
rect 13270 6053 13275 6173
rect 13275 6053 13321 6173
rect 13321 6053 13326 6173
rect 13086 5753 13091 5873
rect 13091 5753 13137 5873
rect 13137 5753 13142 5873
rect 13592 6052 13597 6173
rect 13597 6052 13643 6173
rect 13643 6052 13648 6173
rect 13454 5753 13459 5873
rect 13459 5753 13505 5873
rect 13505 5753 13510 5873
rect 12994 5634 12995 5677
rect 12995 5634 13049 5677
rect 13049 5634 13050 5677
rect 12994 5621 13050 5634
rect 13178 5634 13179 5677
rect 13179 5634 13233 5677
rect 13233 5634 13234 5677
rect 13178 5621 13234 5634
rect 13362 5634 13363 5677
rect 13363 5634 13417 5677
rect 13417 5634 13418 5677
rect 13362 5621 13418 5634
rect 12994 5471 13050 5527
rect 17312 8645 17368 8701
rect 16944 8258 16949 8378
rect 16949 8258 16995 8378
rect 16995 8258 17000 8378
rect 17312 8258 17317 8378
rect 17317 8258 17363 8378
rect 17363 8258 17368 8378
rect 17128 7958 17133 8078
rect 17133 7958 17179 8078
rect 17179 7958 17184 8078
rect 17634 8257 17639 8378
rect 17639 8257 17685 8378
rect 17685 8257 17690 8378
rect 17496 7958 17501 8078
rect 17501 7958 17547 8078
rect 17547 7958 17552 8078
rect 17036 7839 17037 7882
rect 17037 7839 17091 7882
rect 17091 7839 17092 7882
rect 17036 7826 17092 7839
rect 17220 7839 17221 7882
rect 17221 7839 17275 7882
rect 17275 7839 17276 7882
rect 17220 7826 17276 7839
rect 17404 7839 17405 7882
rect 17405 7839 17459 7882
rect 17459 7839 17460 7882
rect 17404 7826 17460 7839
rect 16148 7676 16204 7732
rect 17036 7676 17092 7732
rect 16364 7560 16420 7616
rect 17220 7560 17276 7616
rect 17549 7560 17605 7616
rect 17806 7560 17862 7616
rect 17404 7444 17460 7500
rect 17036 7337 17092 7350
rect 17036 7294 17037 7337
rect 17037 7294 17091 7337
rect 17091 7294 17092 7337
rect 17220 7337 17276 7350
rect 17220 7294 17221 7337
rect 17221 7294 17275 7337
rect 17275 7294 17276 7337
rect 17404 7337 17460 7350
rect 17404 7294 17405 7337
rect 17405 7294 17459 7337
rect 17459 7294 17460 7337
rect 17496 7098 17501 7218
rect 17501 7098 17547 7218
rect 17547 7098 17552 7218
rect 16811 6775 16867 6831
rect 17629 6775 17685 6831
rect 17982 6657 18038 6713
rect 17806 6549 17862 6603
rect 14756 6440 14812 6496
rect 14388 6053 14393 6173
rect 14393 6053 14439 6173
rect 14439 6053 14444 6173
rect 14756 6053 14761 6173
rect 14761 6053 14807 6173
rect 14807 6053 14812 6173
rect 14572 5753 14577 5873
rect 14577 5753 14623 5873
rect 14623 5753 14628 5873
rect 15078 6052 15083 6173
rect 15083 6052 15129 6173
rect 15129 6052 15134 6173
rect 14940 5753 14945 5873
rect 14945 5753 14991 5873
rect 14991 5753 14996 5873
rect 14480 5634 14481 5677
rect 14481 5634 14535 5677
rect 14535 5634 14536 5677
rect 14480 5621 14536 5634
rect 14664 5634 14665 5677
rect 14665 5634 14719 5677
rect 14719 5634 14720 5677
rect 14664 5621 14720 5634
rect 14848 5634 14849 5677
rect 14849 5634 14903 5677
rect 14903 5634 14904 5677
rect 14848 5621 14904 5634
rect 14480 5471 14536 5527
rect 17312 6440 17368 6496
rect 16944 6053 16949 6173
rect 16949 6053 16995 6173
rect 16995 6053 17000 6173
rect 17312 6053 17317 6173
rect 17317 6053 17363 6173
rect 17363 6053 17368 6173
rect 17128 5753 17133 5873
rect 17133 5753 17179 5873
rect 17179 5753 17184 5873
rect 17634 6052 17639 6173
rect 17639 6052 17685 6173
rect 17685 6052 17690 6173
rect 17496 5753 17501 5873
rect 17501 5753 17547 5873
rect 17547 5753 17552 5873
rect 17036 5634 17037 5677
rect 17037 5634 17091 5677
rect 17091 5634 17092 5677
rect 17036 5621 17092 5634
rect 17220 5634 17221 5677
rect 17221 5634 17275 5677
rect 17275 5634 17276 5677
rect 17220 5621 17276 5634
rect 17404 5634 17405 5677
rect 17405 5634 17459 5677
rect 17459 5634 17460 5677
rect 17404 5621 17460 5634
rect 17036 5471 17092 5527
rect 21354 8645 21410 8701
rect 20986 8258 20991 8378
rect 20991 8258 21037 8378
rect 21037 8258 21042 8378
rect 21354 8258 21359 8378
rect 21359 8258 21405 8378
rect 21405 8258 21410 8378
rect 21170 7958 21175 8078
rect 21175 7958 21221 8078
rect 21221 7958 21226 8078
rect 21676 8257 21681 8378
rect 21681 8257 21727 8378
rect 21727 8257 21732 8378
rect 21538 7958 21543 8078
rect 21543 7958 21589 8078
rect 21589 7958 21594 8078
rect 21078 7839 21079 7882
rect 21079 7839 21133 7882
rect 21133 7839 21134 7882
rect 21078 7826 21134 7839
rect 21262 7839 21263 7882
rect 21263 7839 21317 7882
rect 21317 7839 21318 7882
rect 21262 7826 21318 7839
rect 21446 7839 21447 7882
rect 21447 7839 21501 7882
rect 21501 7839 21502 7882
rect 21446 7826 21502 7839
rect 20190 7676 20246 7732
rect 21078 7676 21134 7732
rect 20406 7560 20462 7616
rect 21262 7560 21318 7616
rect 21591 7560 21647 7616
rect 21848 7560 21904 7616
rect 21446 7444 21502 7500
rect 21078 7337 21134 7350
rect 21078 7294 21079 7337
rect 21079 7294 21133 7337
rect 21133 7294 21134 7337
rect 21262 7337 21318 7350
rect 21262 7294 21263 7337
rect 21263 7294 21317 7337
rect 21317 7294 21318 7337
rect 21446 7337 21502 7350
rect 21446 7294 21447 7337
rect 21447 7294 21501 7337
rect 21501 7294 21502 7337
rect 21538 7098 21543 7218
rect 21543 7098 21589 7218
rect 21589 7098 21594 7218
rect 20853 6775 20909 6831
rect 21671 6775 21727 6831
rect 22024 6657 22080 6713
rect 21848 6549 21904 6603
rect 18798 6440 18854 6496
rect 18430 6053 18435 6173
rect 18435 6053 18481 6173
rect 18481 6053 18486 6173
rect 18798 6053 18803 6173
rect 18803 6053 18849 6173
rect 18849 6053 18854 6173
rect 18614 5753 18619 5873
rect 18619 5753 18665 5873
rect 18665 5753 18670 5873
rect 19120 6052 19125 6173
rect 19125 6052 19171 6173
rect 19171 6052 19176 6173
rect 18982 5753 18987 5873
rect 18987 5753 19033 5873
rect 19033 5753 19038 5873
rect 18522 5634 18523 5677
rect 18523 5634 18577 5677
rect 18577 5634 18578 5677
rect 18522 5621 18578 5634
rect 18706 5634 18707 5677
rect 18707 5634 18761 5677
rect 18761 5634 18762 5677
rect 18706 5621 18762 5634
rect 18890 5634 18891 5677
rect 18891 5634 18945 5677
rect 18945 5634 18946 5677
rect 18890 5621 18946 5634
rect 18522 5471 18578 5527
rect 21354 6440 21410 6496
rect 20986 6053 20991 6173
rect 20991 6053 21037 6173
rect 21037 6053 21042 6173
rect 21354 6053 21359 6173
rect 21359 6053 21405 6173
rect 21405 6053 21410 6173
rect 21170 5753 21175 5873
rect 21175 5753 21221 5873
rect 21221 5753 21226 5873
rect 21676 6052 21681 6173
rect 21681 6052 21727 6173
rect 21727 6052 21732 6173
rect 21538 5753 21543 5873
rect 21543 5753 21589 5873
rect 21589 5753 21594 5873
rect 21078 5634 21079 5677
rect 21079 5634 21133 5677
rect 21133 5634 21134 5677
rect 21078 5621 21134 5634
rect 21262 5634 21263 5677
rect 21263 5634 21317 5677
rect 21317 5634 21318 5677
rect 21262 5621 21318 5634
rect 21446 5634 21447 5677
rect 21447 5634 21501 5677
rect 21501 5634 21502 5677
rect 21446 5621 21502 5634
rect 21078 5471 21134 5527
rect 25396 8645 25452 8701
rect 25028 8258 25033 8378
rect 25033 8258 25079 8378
rect 25079 8258 25084 8378
rect 25396 8258 25401 8378
rect 25401 8258 25447 8378
rect 25447 8258 25452 8378
rect 25212 7958 25217 8078
rect 25217 7958 25263 8078
rect 25263 7958 25268 8078
rect 25718 8257 25723 8378
rect 25723 8257 25769 8378
rect 25769 8257 25774 8378
rect 25580 7958 25585 8078
rect 25585 7958 25631 8078
rect 25631 7958 25636 8078
rect 25120 7839 25121 7882
rect 25121 7839 25175 7882
rect 25175 7839 25176 7882
rect 25120 7826 25176 7839
rect 25304 7839 25305 7882
rect 25305 7839 25359 7882
rect 25359 7839 25360 7882
rect 25304 7826 25360 7839
rect 25488 7839 25489 7882
rect 25489 7839 25543 7882
rect 25543 7839 25544 7882
rect 25488 7826 25544 7839
rect 24232 7676 24288 7732
rect 25120 7676 25176 7732
rect 24448 7560 24504 7616
rect 25304 7560 25360 7616
rect 25633 7560 25689 7616
rect 25890 7560 25946 7616
rect 25488 7444 25544 7500
rect 25120 7337 25176 7350
rect 25120 7294 25121 7337
rect 25121 7294 25175 7337
rect 25175 7294 25176 7337
rect 25304 7337 25360 7350
rect 25304 7294 25305 7337
rect 25305 7294 25359 7337
rect 25359 7294 25360 7337
rect 25488 7337 25544 7350
rect 25488 7294 25489 7337
rect 25489 7294 25543 7337
rect 25543 7294 25544 7337
rect 25580 7098 25585 7218
rect 25585 7098 25631 7218
rect 25631 7098 25636 7218
rect 24895 6775 24951 6831
rect 25713 6775 25769 6831
rect 26066 6657 26122 6713
rect 25890 6549 25946 6603
rect 22840 6440 22896 6496
rect 22472 6053 22477 6173
rect 22477 6053 22523 6173
rect 22523 6053 22528 6173
rect 22840 6053 22845 6173
rect 22845 6053 22891 6173
rect 22891 6053 22896 6173
rect 22656 5753 22661 5873
rect 22661 5753 22707 5873
rect 22707 5753 22712 5873
rect 23162 6052 23167 6173
rect 23167 6052 23213 6173
rect 23213 6052 23218 6173
rect 23024 5753 23029 5873
rect 23029 5753 23075 5873
rect 23075 5753 23080 5873
rect 22564 5634 22565 5677
rect 22565 5634 22619 5677
rect 22619 5634 22620 5677
rect 22564 5621 22620 5634
rect 22748 5634 22749 5677
rect 22749 5634 22803 5677
rect 22803 5634 22804 5677
rect 22748 5621 22804 5634
rect 22932 5634 22933 5677
rect 22933 5634 22987 5677
rect 22987 5634 22988 5677
rect 22932 5621 22988 5634
rect 22564 5471 22620 5527
rect 25396 6440 25452 6496
rect 25028 6053 25033 6173
rect 25033 6053 25079 6173
rect 25079 6053 25084 6173
rect 25396 6053 25401 6173
rect 25401 6053 25447 6173
rect 25447 6053 25452 6173
rect 25212 5753 25217 5873
rect 25217 5753 25263 5873
rect 25263 5753 25268 5873
rect 25718 6052 25723 6173
rect 25723 6052 25769 6173
rect 25769 6052 25774 6173
rect 25580 5753 25585 5873
rect 25585 5753 25631 5873
rect 25631 5753 25636 5873
rect 25120 5634 25121 5677
rect 25121 5634 25175 5677
rect 25175 5634 25176 5677
rect 25120 5621 25176 5634
rect 25304 5634 25305 5677
rect 25305 5634 25359 5677
rect 25359 5634 25360 5677
rect 25304 5621 25360 5634
rect 25488 5634 25489 5677
rect 25489 5634 25543 5677
rect 25543 5634 25544 5677
rect 25488 5621 25544 5634
rect 25120 5471 25176 5527
rect 26882 6440 26938 6496
rect 26514 6053 26519 6173
rect 26519 6053 26565 6173
rect 26565 6053 26570 6173
rect 26882 6053 26887 6173
rect 26887 6053 26933 6173
rect 26933 6053 26938 6173
rect 26698 5753 26703 5873
rect 26703 5753 26749 5873
rect 26749 5753 26754 5873
rect 27204 6052 27209 6173
rect 27209 6052 27255 6173
rect 27255 6052 27260 6173
rect 27066 5753 27071 5873
rect 27071 5753 27117 5873
rect 27117 5753 27122 5873
rect 26606 5634 26607 5677
rect 26607 5634 26661 5677
rect 26661 5634 26662 5677
rect 26606 5621 26662 5634
rect 26790 5634 26791 5677
rect 26791 5634 26845 5677
rect 26845 5634 26846 5677
rect 26790 5621 26846 5634
rect 26974 5634 26975 5677
rect 26975 5634 27029 5677
rect 27029 5634 27030 5677
rect 26974 5621 27030 5634
rect 26606 5471 26662 5527
rect 90 5355 146 5411
rect 1082 5355 1138 5411
rect 1411 5355 1467 5411
rect 1844 5355 1900 5411
rect 2568 5355 2624 5411
rect 2897 5355 2953 5411
rect 3154 5355 3210 5411
rect 1266 5239 1322 5295
rect 2752 5239 2808 5295
rect 898 5132 954 5145
rect 898 5089 899 5132
rect 899 5089 953 5132
rect 953 5089 954 5132
rect 1082 5132 1138 5145
rect 1082 5089 1083 5132
rect 1083 5089 1137 5132
rect 1137 5089 1138 5132
rect 1266 5132 1322 5145
rect 1266 5089 1267 5132
rect 1267 5089 1321 5132
rect 1321 5089 1322 5132
rect 1358 4893 1363 5013
rect 1363 4893 1409 5013
rect 1409 4893 1414 5013
rect 673 4570 729 4626
rect 1491 4570 1547 4626
rect -318 4453 -262 4509
rect 4102 5355 4158 5411
rect 5094 5355 5150 5411
rect 5423 5355 5479 5411
rect 5856 5355 5912 5411
rect 6580 5355 6636 5411
rect 6909 5355 6965 5411
rect 7166 5355 7222 5411
rect 5278 5239 5334 5295
rect 3966 5167 4022 5223
rect 2384 5132 2440 5145
rect 2384 5089 2385 5132
rect 2385 5089 2439 5132
rect 2439 5089 2440 5132
rect 2568 5132 2624 5145
rect 2568 5089 2569 5132
rect 2569 5089 2623 5132
rect 2623 5089 2624 5132
rect 2752 5132 2808 5145
rect 2752 5089 2753 5132
rect 2753 5089 2807 5132
rect 2807 5089 2808 5132
rect 2844 4893 2849 5013
rect 2849 4893 2895 5013
rect 2895 4893 2900 5013
rect 2159 4570 2215 4626
rect 2977 4570 3033 4626
rect 3330 4453 3386 4509
rect 6764 5239 6820 5295
rect 4910 5132 4966 5145
rect 4910 5089 4911 5132
rect 4911 5089 4965 5132
rect 4965 5089 4966 5132
rect 5094 5132 5150 5145
rect 5094 5089 5095 5132
rect 5095 5089 5149 5132
rect 5149 5089 5150 5132
rect 5278 5132 5334 5145
rect 5278 5089 5279 5132
rect 5279 5089 5333 5132
rect 5333 5089 5334 5132
rect 5370 4893 5375 5013
rect 5375 4893 5421 5013
rect 5421 4893 5426 5013
rect 4685 4570 4741 4626
rect 5503 4570 5559 4626
rect 3694 4453 3750 4509
rect 8144 5355 8200 5411
rect 9136 5355 9192 5411
rect 9465 5355 9521 5411
rect 9898 5355 9954 5411
rect 10622 5355 10678 5411
rect 10951 5355 11007 5411
rect 11208 5355 11264 5411
rect 9320 5239 9376 5295
rect 7978 5167 8034 5223
rect 6396 5132 6452 5145
rect 6396 5089 6397 5132
rect 6397 5089 6451 5132
rect 6451 5089 6452 5132
rect 6580 5132 6636 5145
rect 6580 5089 6581 5132
rect 6581 5089 6635 5132
rect 6635 5089 6636 5132
rect 6764 5132 6820 5145
rect 6764 5089 6765 5132
rect 6765 5089 6819 5132
rect 6819 5089 6820 5132
rect 6856 4893 6861 5013
rect 6861 4893 6907 5013
rect 6907 4893 6912 5013
rect 6171 4570 6227 4626
rect 6989 4570 7045 4626
rect 7342 4453 7398 4509
rect 1844 4342 1900 4398
rect 3154 4343 3210 4399
rect 1174 4235 1230 4291
rect 806 3848 811 3968
rect 811 3848 857 3968
rect 857 3848 862 3968
rect 1174 3848 1179 3968
rect 1179 3848 1225 3968
rect 1225 3848 1230 3968
rect 990 3548 995 3668
rect 995 3548 1041 3668
rect 1041 3548 1046 3668
rect 1496 3847 1501 3968
rect 1501 3847 1547 3968
rect 1547 3847 1552 3968
rect 1358 3548 1363 3668
rect 1363 3548 1409 3668
rect 1409 3548 1414 3668
rect 898 3429 899 3472
rect 899 3429 953 3472
rect 953 3429 954 3472
rect 898 3416 954 3429
rect 1082 3429 1083 3472
rect 1083 3429 1137 3472
rect 1137 3429 1138 3472
rect 1082 3416 1138 3429
rect 1266 3429 1267 3472
rect 1267 3429 1321 3472
rect 1321 3429 1322 3472
rect 1266 3416 1322 3429
rect 898 3266 954 3322
rect 2660 4236 2716 4292
rect 2292 3849 2297 3969
rect 2297 3849 2343 3969
rect 2343 3849 2348 3969
rect 2660 3849 2665 3969
rect 2665 3849 2711 3969
rect 2711 3849 2716 3969
rect 2476 3549 2481 3669
rect 2481 3549 2527 3669
rect 2527 3549 2532 3669
rect 2982 3848 2987 3969
rect 2987 3848 3033 3969
rect 3033 3848 3038 3969
rect 2844 3549 2849 3669
rect 2849 3549 2895 3669
rect 2895 3549 2900 3669
rect 2384 3430 2385 3473
rect 2385 3430 2439 3473
rect 2439 3430 2440 3473
rect 2384 3417 2440 3430
rect 2568 3430 2569 3473
rect 2569 3430 2623 3473
rect 2623 3430 2624 3473
rect 2568 3417 2624 3430
rect 2752 3430 2753 3473
rect 2753 3430 2807 3473
rect 2807 3430 2808 3473
rect 2752 3417 2808 3430
rect 2384 3267 2440 3323
rect 1082 3150 1138 3206
rect 1411 3150 1467 3206
rect 1668 3150 1724 3206
rect 2568 3151 2624 3207
rect 2897 3151 2953 3207
rect 3330 3151 3386 3207
rect 10806 5239 10862 5295
rect 8952 5132 9008 5145
rect 8952 5089 8953 5132
rect 8953 5089 9007 5132
rect 9007 5089 9008 5132
rect 9136 5132 9192 5145
rect 9136 5089 9137 5132
rect 9137 5089 9191 5132
rect 9191 5089 9192 5132
rect 9320 5132 9376 5145
rect 9320 5089 9321 5132
rect 9321 5089 9375 5132
rect 9375 5089 9376 5132
rect 9412 4893 9417 5013
rect 9417 4893 9463 5013
rect 9463 4893 9468 5013
rect 8727 4570 8783 4626
rect 9545 4570 9601 4626
rect 7706 4453 7762 4509
rect 12186 5355 12242 5411
rect 13178 5355 13234 5411
rect 13507 5355 13563 5411
rect 13940 5355 13996 5411
rect 14664 5355 14720 5411
rect 14993 5355 15049 5411
rect 15250 5355 15306 5411
rect 13362 5239 13418 5295
rect 12020 5167 12076 5223
rect 10438 5132 10494 5145
rect 10438 5089 10439 5132
rect 10439 5089 10493 5132
rect 10493 5089 10494 5132
rect 10622 5132 10678 5145
rect 10622 5089 10623 5132
rect 10623 5089 10677 5132
rect 10677 5089 10678 5132
rect 10806 5132 10862 5145
rect 10806 5089 10807 5132
rect 10807 5089 10861 5132
rect 10861 5089 10862 5132
rect 10898 4893 10903 5013
rect 10903 4893 10949 5013
rect 10949 4893 10954 5013
rect 10213 4570 10269 4626
rect 11031 4570 11087 4626
rect 11384 4453 11440 4509
rect 5856 4342 5912 4398
rect 7166 4343 7222 4399
rect 5186 4235 5242 4291
rect 4818 3848 4823 3968
rect 4823 3848 4869 3968
rect 4869 3848 4874 3968
rect 5186 3848 5191 3968
rect 5191 3848 5237 3968
rect 5237 3848 5242 3968
rect 5002 3548 5007 3668
rect 5007 3548 5053 3668
rect 5053 3548 5058 3668
rect 5508 3847 5513 3968
rect 5513 3847 5559 3968
rect 5559 3847 5564 3968
rect 5370 3548 5375 3668
rect 5375 3548 5421 3668
rect 5421 3548 5426 3668
rect 4910 3429 4911 3472
rect 4911 3429 4965 3472
rect 4965 3429 4966 3472
rect 4910 3416 4966 3429
rect 5094 3429 5095 3472
rect 5095 3429 5149 3472
rect 5149 3429 5150 3472
rect 5094 3416 5150 3429
rect 5278 3429 5279 3472
rect 5279 3429 5333 3472
rect 5333 3429 5334 3472
rect 5278 3416 5334 3429
rect 4910 3266 4966 3322
rect 6672 4236 6728 4292
rect 6304 3849 6309 3969
rect 6309 3849 6355 3969
rect 6355 3849 6360 3969
rect 6672 3849 6677 3969
rect 6677 3849 6723 3969
rect 6723 3849 6728 3969
rect 6488 3549 6493 3669
rect 6493 3549 6539 3669
rect 6539 3549 6544 3669
rect 6994 3848 6999 3969
rect 6999 3848 7045 3969
rect 7045 3848 7050 3969
rect 6856 3549 6861 3669
rect 6861 3549 6907 3669
rect 6907 3549 6912 3669
rect 6396 3430 6397 3473
rect 6397 3430 6451 3473
rect 6451 3430 6452 3473
rect 6396 3417 6452 3430
rect 6580 3430 6581 3473
rect 6581 3430 6635 3473
rect 6635 3430 6636 3473
rect 6580 3417 6636 3430
rect 6764 3430 6765 3473
rect 6765 3430 6819 3473
rect 6819 3430 6820 3473
rect 6764 3417 6820 3430
rect 6396 3267 6452 3323
rect 5094 3150 5150 3206
rect 5423 3150 5479 3206
rect 5680 3150 5736 3206
rect 6580 3151 6636 3207
rect 6909 3151 6965 3207
rect 7342 3151 7398 3207
rect 14848 5239 14904 5295
rect 12994 5132 13050 5145
rect 12994 5089 12995 5132
rect 12995 5089 13049 5132
rect 13049 5089 13050 5132
rect 13178 5132 13234 5145
rect 13178 5089 13179 5132
rect 13179 5089 13233 5132
rect 13233 5089 13234 5132
rect 13362 5132 13418 5145
rect 13362 5089 13363 5132
rect 13363 5089 13417 5132
rect 13417 5089 13418 5132
rect 13454 4893 13459 5013
rect 13459 4893 13505 5013
rect 13505 4893 13510 5013
rect 12769 4570 12825 4626
rect 13587 4570 13643 4626
rect 11748 4453 11804 4509
rect 16228 5355 16284 5411
rect 17220 5355 17276 5411
rect 17549 5355 17605 5411
rect 17982 5355 18038 5411
rect 18706 5355 18762 5411
rect 19035 5355 19091 5411
rect 19292 5355 19348 5411
rect 17404 5239 17460 5295
rect 16062 5167 16118 5223
rect 14480 5132 14536 5145
rect 14480 5089 14481 5132
rect 14481 5089 14535 5132
rect 14535 5089 14536 5132
rect 14664 5132 14720 5145
rect 14664 5089 14665 5132
rect 14665 5089 14719 5132
rect 14719 5089 14720 5132
rect 14848 5132 14904 5145
rect 14848 5089 14849 5132
rect 14849 5089 14903 5132
rect 14903 5089 14904 5132
rect 14940 4893 14945 5013
rect 14945 4893 14991 5013
rect 14991 4893 14996 5013
rect 14255 4570 14311 4626
rect 15073 4570 15129 4626
rect 15426 4453 15482 4509
rect 9898 4342 9954 4398
rect 11208 4343 11264 4399
rect 9228 4235 9284 4291
rect 8860 3848 8865 3968
rect 8865 3848 8911 3968
rect 8911 3848 8916 3968
rect 9228 3848 9233 3968
rect 9233 3848 9279 3968
rect 9279 3848 9284 3968
rect 9044 3548 9049 3668
rect 9049 3548 9095 3668
rect 9095 3548 9100 3668
rect 9550 3847 9555 3968
rect 9555 3847 9601 3968
rect 9601 3847 9606 3968
rect 9412 3548 9417 3668
rect 9417 3548 9463 3668
rect 9463 3548 9468 3668
rect 8952 3429 8953 3472
rect 8953 3429 9007 3472
rect 9007 3429 9008 3472
rect 8952 3416 9008 3429
rect 9136 3429 9137 3472
rect 9137 3429 9191 3472
rect 9191 3429 9192 3472
rect 9136 3416 9192 3429
rect 9320 3429 9321 3472
rect 9321 3429 9375 3472
rect 9375 3429 9376 3472
rect 9320 3416 9376 3429
rect 8952 3266 9008 3322
rect 10714 4236 10770 4292
rect 10346 3849 10351 3969
rect 10351 3849 10397 3969
rect 10397 3849 10402 3969
rect 10714 3849 10719 3969
rect 10719 3849 10765 3969
rect 10765 3849 10770 3969
rect 10530 3549 10535 3669
rect 10535 3549 10581 3669
rect 10581 3549 10586 3669
rect 11036 3848 11041 3969
rect 11041 3848 11087 3969
rect 11087 3848 11092 3969
rect 10898 3549 10903 3669
rect 10903 3549 10949 3669
rect 10949 3549 10954 3669
rect 10438 3430 10439 3473
rect 10439 3430 10493 3473
rect 10493 3430 10494 3473
rect 10438 3417 10494 3430
rect 10622 3430 10623 3473
rect 10623 3430 10677 3473
rect 10677 3430 10678 3473
rect 10622 3417 10678 3430
rect 10806 3430 10807 3473
rect 10807 3430 10861 3473
rect 10861 3430 10862 3473
rect 10806 3417 10862 3430
rect 10438 3267 10494 3323
rect 9136 3150 9192 3206
rect 9465 3150 9521 3206
rect 9722 3150 9778 3206
rect 10622 3151 10678 3207
rect 10951 3151 11007 3207
rect 11384 3151 11440 3207
rect 18890 5239 18946 5295
rect 17036 5132 17092 5145
rect 17036 5089 17037 5132
rect 17037 5089 17091 5132
rect 17091 5089 17092 5132
rect 17220 5132 17276 5145
rect 17220 5089 17221 5132
rect 17221 5089 17275 5132
rect 17275 5089 17276 5132
rect 17404 5132 17460 5145
rect 17404 5089 17405 5132
rect 17405 5089 17459 5132
rect 17459 5089 17460 5132
rect 17496 4893 17501 5013
rect 17501 4893 17547 5013
rect 17547 4893 17552 5013
rect 16811 4570 16867 4626
rect 17629 4570 17685 4626
rect 15790 4453 15846 4509
rect 20270 5355 20326 5411
rect 21262 5355 21318 5411
rect 21591 5355 21647 5411
rect 22024 5355 22080 5411
rect 22748 5355 22804 5411
rect 23077 5355 23133 5411
rect 23334 5355 23390 5411
rect 21446 5239 21502 5295
rect 20104 5167 20160 5223
rect 18522 5132 18578 5145
rect 18522 5089 18523 5132
rect 18523 5089 18577 5132
rect 18577 5089 18578 5132
rect 18706 5132 18762 5145
rect 18706 5089 18707 5132
rect 18707 5089 18761 5132
rect 18761 5089 18762 5132
rect 18890 5132 18946 5145
rect 18890 5089 18891 5132
rect 18891 5089 18945 5132
rect 18945 5089 18946 5132
rect 18982 4893 18987 5013
rect 18987 4893 19033 5013
rect 19033 4893 19038 5013
rect 18297 4570 18353 4626
rect 19115 4570 19171 4626
rect 19468 4453 19524 4509
rect 13940 4342 13996 4398
rect 15250 4343 15306 4399
rect 13270 4235 13326 4291
rect 12902 3848 12907 3968
rect 12907 3848 12953 3968
rect 12953 3848 12958 3968
rect 13270 3848 13275 3968
rect 13275 3848 13321 3968
rect 13321 3848 13326 3968
rect 13086 3548 13091 3668
rect 13091 3548 13137 3668
rect 13137 3548 13142 3668
rect 13592 3847 13597 3968
rect 13597 3847 13643 3968
rect 13643 3847 13648 3968
rect 13454 3548 13459 3668
rect 13459 3548 13505 3668
rect 13505 3548 13510 3668
rect 12994 3429 12995 3472
rect 12995 3429 13049 3472
rect 13049 3429 13050 3472
rect 12994 3416 13050 3429
rect 13178 3429 13179 3472
rect 13179 3429 13233 3472
rect 13233 3429 13234 3472
rect 13178 3416 13234 3429
rect 13362 3429 13363 3472
rect 13363 3429 13417 3472
rect 13417 3429 13418 3472
rect 13362 3416 13418 3429
rect 12994 3266 13050 3322
rect 14756 4236 14812 4292
rect 14388 3849 14393 3969
rect 14393 3849 14439 3969
rect 14439 3849 14444 3969
rect 14756 3849 14761 3969
rect 14761 3849 14807 3969
rect 14807 3849 14812 3969
rect 14572 3549 14577 3669
rect 14577 3549 14623 3669
rect 14623 3549 14628 3669
rect 15078 3848 15083 3969
rect 15083 3848 15129 3969
rect 15129 3848 15134 3969
rect 14940 3549 14945 3669
rect 14945 3549 14991 3669
rect 14991 3549 14996 3669
rect 14480 3430 14481 3473
rect 14481 3430 14535 3473
rect 14535 3430 14536 3473
rect 14480 3417 14536 3430
rect 14664 3430 14665 3473
rect 14665 3430 14719 3473
rect 14719 3430 14720 3473
rect 14664 3417 14720 3430
rect 14848 3430 14849 3473
rect 14849 3430 14903 3473
rect 14903 3430 14904 3473
rect 14848 3417 14904 3430
rect 14480 3267 14536 3323
rect 13178 3150 13234 3206
rect 13507 3150 13563 3206
rect 13764 3150 13820 3206
rect 14664 3151 14720 3207
rect 14993 3151 15049 3207
rect 15426 3151 15482 3207
rect 22932 5239 22988 5295
rect 21078 5132 21134 5145
rect 21078 5089 21079 5132
rect 21079 5089 21133 5132
rect 21133 5089 21134 5132
rect 21262 5132 21318 5145
rect 21262 5089 21263 5132
rect 21263 5089 21317 5132
rect 21317 5089 21318 5132
rect 21446 5132 21502 5145
rect 21446 5089 21447 5132
rect 21447 5089 21501 5132
rect 21501 5089 21502 5132
rect 21538 4893 21543 5013
rect 21543 4893 21589 5013
rect 21589 4893 21594 5013
rect 20853 4570 20909 4626
rect 21671 4570 21727 4626
rect 19832 4453 19888 4509
rect 24312 5355 24368 5411
rect 25304 5355 25360 5411
rect 25633 5355 25689 5411
rect 26066 5355 26122 5411
rect 26790 5355 26846 5411
rect 27119 5355 27175 5411
rect 27376 5355 27432 5411
rect 25488 5239 25544 5295
rect 24146 5167 24202 5223
rect 22564 5132 22620 5145
rect 22564 5089 22565 5132
rect 22565 5089 22619 5132
rect 22619 5089 22620 5132
rect 22748 5132 22804 5145
rect 22748 5089 22749 5132
rect 22749 5089 22803 5132
rect 22803 5089 22804 5132
rect 22932 5132 22988 5145
rect 22932 5089 22933 5132
rect 22933 5089 22987 5132
rect 22987 5089 22988 5132
rect 23024 4893 23029 5013
rect 23029 4893 23075 5013
rect 23075 4893 23080 5013
rect 22339 4570 22395 4626
rect 23157 4570 23213 4626
rect 23510 4453 23566 4509
rect 17982 4342 18038 4398
rect 19292 4343 19348 4399
rect 17312 4235 17368 4291
rect 16944 3848 16949 3968
rect 16949 3848 16995 3968
rect 16995 3848 17000 3968
rect 17312 3848 17317 3968
rect 17317 3848 17363 3968
rect 17363 3848 17368 3968
rect 17128 3548 17133 3668
rect 17133 3548 17179 3668
rect 17179 3548 17184 3668
rect 17634 3847 17639 3968
rect 17639 3847 17685 3968
rect 17685 3847 17690 3968
rect 17496 3548 17501 3668
rect 17501 3548 17547 3668
rect 17547 3548 17552 3668
rect 17036 3429 17037 3472
rect 17037 3429 17091 3472
rect 17091 3429 17092 3472
rect 17036 3416 17092 3429
rect 17220 3429 17221 3472
rect 17221 3429 17275 3472
rect 17275 3429 17276 3472
rect 17220 3416 17276 3429
rect 17404 3429 17405 3472
rect 17405 3429 17459 3472
rect 17459 3429 17460 3472
rect 17404 3416 17460 3429
rect 17036 3266 17092 3322
rect 18798 4236 18854 4292
rect 18430 3849 18435 3969
rect 18435 3849 18481 3969
rect 18481 3849 18486 3969
rect 18798 3849 18803 3969
rect 18803 3849 18849 3969
rect 18849 3849 18854 3969
rect 18614 3549 18619 3669
rect 18619 3549 18665 3669
rect 18665 3549 18670 3669
rect 19120 3848 19125 3969
rect 19125 3848 19171 3969
rect 19171 3848 19176 3969
rect 18982 3549 18987 3669
rect 18987 3549 19033 3669
rect 19033 3549 19038 3669
rect 18522 3430 18523 3473
rect 18523 3430 18577 3473
rect 18577 3430 18578 3473
rect 18522 3417 18578 3430
rect 18706 3430 18707 3473
rect 18707 3430 18761 3473
rect 18761 3430 18762 3473
rect 18706 3417 18762 3430
rect 18890 3430 18891 3473
rect 18891 3430 18945 3473
rect 18945 3430 18946 3473
rect 18890 3417 18946 3430
rect 18522 3267 18578 3323
rect 17220 3150 17276 3206
rect 17549 3150 17605 3206
rect 17806 3150 17862 3206
rect 18706 3151 18762 3207
rect 19035 3151 19091 3207
rect 19468 3151 19524 3207
rect 26974 5239 27030 5295
rect 25120 5132 25176 5145
rect 25120 5089 25121 5132
rect 25121 5089 25175 5132
rect 25175 5089 25176 5132
rect 25304 5132 25360 5145
rect 25304 5089 25305 5132
rect 25305 5089 25359 5132
rect 25359 5089 25360 5132
rect 25488 5132 25544 5145
rect 25488 5089 25489 5132
rect 25489 5089 25543 5132
rect 25543 5089 25544 5132
rect 25580 4893 25585 5013
rect 25585 4893 25631 5013
rect 25631 4893 25636 5013
rect 24895 4570 24951 4626
rect 25713 4570 25769 4626
rect 23874 4453 23930 4509
rect 26606 5132 26662 5145
rect 26606 5089 26607 5132
rect 26607 5089 26661 5132
rect 26661 5089 26662 5132
rect 26790 5132 26846 5145
rect 26790 5089 26791 5132
rect 26791 5089 26845 5132
rect 26845 5089 26846 5132
rect 26974 5132 27030 5145
rect 26974 5089 26975 5132
rect 26975 5089 27029 5132
rect 27029 5089 27030 5132
rect 27066 4893 27071 5013
rect 27071 4893 27117 5013
rect 27117 4893 27122 5013
rect 26381 4570 26437 4626
rect 27199 4570 27255 4626
rect 27552 4453 27608 4509
rect 22024 4342 22080 4398
rect 23334 4343 23390 4399
rect 21354 4235 21410 4291
rect 20986 3848 20991 3968
rect 20991 3848 21037 3968
rect 21037 3848 21042 3968
rect 21354 3848 21359 3968
rect 21359 3848 21405 3968
rect 21405 3848 21410 3968
rect 21170 3548 21175 3668
rect 21175 3548 21221 3668
rect 21221 3548 21226 3668
rect 21676 3847 21681 3968
rect 21681 3847 21727 3968
rect 21727 3847 21732 3968
rect 21538 3548 21543 3668
rect 21543 3548 21589 3668
rect 21589 3548 21594 3668
rect 21078 3429 21079 3472
rect 21079 3429 21133 3472
rect 21133 3429 21134 3472
rect 21078 3416 21134 3429
rect 21262 3429 21263 3472
rect 21263 3429 21317 3472
rect 21317 3429 21318 3472
rect 21262 3416 21318 3429
rect 21446 3429 21447 3472
rect 21447 3429 21501 3472
rect 21501 3429 21502 3472
rect 21446 3416 21502 3429
rect 21078 3266 21134 3322
rect 22840 4236 22896 4292
rect 22472 3849 22477 3969
rect 22477 3849 22523 3969
rect 22523 3849 22528 3969
rect 22840 3849 22845 3969
rect 22845 3849 22891 3969
rect 22891 3849 22896 3969
rect 22656 3549 22661 3669
rect 22661 3549 22707 3669
rect 22707 3549 22712 3669
rect 23162 3848 23167 3969
rect 23167 3848 23213 3969
rect 23213 3848 23218 3969
rect 23024 3549 23029 3669
rect 23029 3549 23075 3669
rect 23075 3549 23080 3669
rect 22564 3430 22565 3473
rect 22565 3430 22619 3473
rect 22619 3430 22620 3473
rect 22564 3417 22620 3430
rect 22748 3430 22749 3473
rect 22749 3430 22803 3473
rect 22803 3430 22804 3473
rect 22748 3417 22804 3430
rect 22932 3430 22933 3473
rect 22933 3430 22987 3473
rect 22987 3430 22988 3473
rect 22932 3417 22988 3430
rect 22564 3267 22620 3323
rect 21262 3150 21318 3206
rect 21591 3150 21647 3206
rect 21848 3150 21904 3206
rect 22748 3151 22804 3207
rect 23077 3151 23133 3207
rect 23510 3151 23566 3207
rect 26066 4342 26122 4398
rect 27376 4343 27432 4399
rect 25396 4235 25452 4291
rect 25028 3848 25033 3968
rect 25033 3848 25079 3968
rect 25079 3848 25084 3968
rect 25396 3848 25401 3968
rect 25401 3848 25447 3968
rect 25447 3848 25452 3968
rect 25212 3548 25217 3668
rect 25217 3548 25263 3668
rect 25263 3548 25268 3668
rect 25718 3847 25723 3968
rect 25723 3847 25769 3968
rect 25769 3847 25774 3968
rect 25580 3548 25585 3668
rect 25585 3548 25631 3668
rect 25631 3548 25636 3668
rect 25120 3429 25121 3472
rect 25121 3429 25175 3472
rect 25175 3429 25176 3472
rect 25120 3416 25176 3429
rect 25304 3429 25305 3472
rect 25305 3429 25359 3472
rect 25359 3429 25360 3472
rect 25304 3416 25360 3429
rect 25488 3429 25489 3472
rect 25489 3429 25543 3472
rect 25543 3429 25544 3472
rect 25488 3416 25544 3429
rect 25120 3266 25176 3322
rect 26882 4236 26938 4292
rect 26514 3849 26519 3969
rect 26519 3849 26565 3969
rect 26565 3849 26570 3969
rect 26882 3849 26887 3969
rect 26887 3849 26933 3969
rect 26933 3849 26938 3969
rect 26698 3549 26703 3669
rect 26703 3549 26749 3669
rect 26749 3549 26754 3669
rect 27204 3848 27209 3969
rect 27209 3848 27255 3969
rect 27255 3848 27260 3969
rect 27066 3549 27071 3669
rect 27071 3549 27117 3669
rect 27117 3549 27122 3669
rect 26606 3430 26607 3473
rect 26607 3430 26661 3473
rect 26661 3430 26662 3473
rect 26606 3417 26662 3430
rect 26790 3430 26791 3473
rect 26791 3430 26845 3473
rect 26845 3430 26846 3473
rect 26790 3417 26846 3430
rect 26974 3430 26975 3473
rect 26975 3430 27029 3473
rect 27029 3430 27030 3473
rect 26974 3417 27030 3430
rect 26606 3267 26662 3323
rect 25304 3150 25360 3206
rect 25633 3150 25689 3206
rect 25890 3150 25946 3206
rect 26790 3151 26846 3207
rect 27119 3151 27175 3207
rect 27552 3151 27608 3207
rect 226 3034 282 3090
rect 1266 3034 1322 3090
rect 2752 3035 2808 3091
rect 898 2927 954 2940
rect 898 2884 899 2927
rect 899 2884 953 2927
rect 953 2884 954 2927
rect 1082 2927 1138 2940
rect 1082 2884 1083 2927
rect 1083 2884 1137 2927
rect 1137 2884 1138 2927
rect 1266 2927 1322 2940
rect 1266 2884 1267 2927
rect 1267 2884 1321 2927
rect 1321 2884 1322 2927
rect 1358 2688 1363 2808
rect 1363 2688 1409 2808
rect 1409 2688 1414 2808
rect 673 2365 729 2421
rect 1491 2365 1547 2421
rect 1844 2247 1900 2303
rect 1668 2139 1724 2193
rect 1174 2030 1230 2086
rect 806 1643 811 1763
rect 811 1643 857 1763
rect 857 1643 862 1763
rect 1174 1643 1179 1763
rect 1179 1643 1225 1763
rect 1225 1643 1230 1763
rect 990 1343 995 1463
rect 995 1343 1041 1463
rect 1041 1343 1046 1463
rect 1496 1642 1501 1763
rect 1501 1642 1547 1763
rect 1547 1642 1552 1763
rect 1358 1343 1363 1463
rect 1363 1343 1409 1463
rect 1409 1343 1414 1463
rect 898 1224 899 1267
rect 899 1224 953 1267
rect 953 1224 954 1267
rect 898 1211 954 1224
rect 1082 1224 1083 1267
rect 1083 1224 1137 1267
rect 1137 1224 1138 1267
rect 1082 1211 1138 1224
rect 1266 1224 1267 1267
rect 1267 1224 1321 1267
rect 1321 1224 1322 1267
rect 1266 1211 1322 1224
rect 898 1061 954 1117
rect 90 945 146 1001
rect 1082 945 1138 1001
rect 1411 945 1467 1001
rect 1844 945 1900 1001
rect -109 829 -53 885
rect 1266 829 1322 885
rect 898 722 954 735
rect 898 679 899 722
rect 899 679 953 722
rect 953 679 954 722
rect 1082 722 1138 735
rect 1082 679 1083 722
rect 1083 679 1137 722
rect 1137 679 1138 722
rect 1266 722 1322 735
rect 1266 679 1267 722
rect 1267 679 1321 722
rect 1321 679 1322 722
rect 1358 483 1363 603
rect 1363 483 1409 603
rect 1409 483 1414 603
rect 673 160 729 216
rect 1491 160 1547 216
rect 4238 3034 4294 3090
rect 5278 3034 5334 3090
rect 2384 2928 2440 2941
rect 2384 2885 2385 2928
rect 2385 2885 2439 2928
rect 2439 2885 2440 2928
rect 2568 2928 2624 2941
rect 2568 2885 2569 2928
rect 2569 2885 2623 2928
rect 2623 2885 2624 2928
rect 2752 2928 2808 2941
rect 2752 2885 2753 2928
rect 2753 2885 2807 2928
rect 2807 2885 2808 2928
rect 2844 2689 2849 2809
rect 2849 2689 2895 2809
rect 2895 2689 2900 2809
rect 2159 2366 2215 2422
rect 2977 2366 3033 2422
rect 6764 3035 6820 3091
rect 4910 2927 4966 2940
rect 4910 2884 4911 2927
rect 4911 2884 4965 2927
rect 4965 2884 4966 2927
rect 5094 2927 5150 2940
rect 5094 2884 5095 2927
rect 5095 2884 5149 2927
rect 5149 2884 5150 2927
rect 5278 2927 5334 2940
rect 5278 2884 5279 2927
rect 5279 2884 5333 2927
rect 5333 2884 5334 2927
rect 5370 2688 5375 2808
rect 5375 2688 5421 2808
rect 5421 2688 5426 2808
rect 4685 2365 4741 2421
rect 5503 2365 5559 2421
rect 5856 2247 5912 2303
rect 5680 2139 5736 2193
rect 5186 2030 5242 2086
rect 4818 1643 4823 1763
rect 4823 1643 4869 1763
rect 4869 1643 4874 1763
rect 5186 1643 5191 1763
rect 5191 1643 5237 1763
rect 5237 1643 5242 1763
rect 5002 1343 5007 1463
rect 5007 1343 5053 1463
rect 5053 1343 5058 1463
rect 5508 1642 5513 1763
rect 5513 1642 5559 1763
rect 5559 1642 5564 1763
rect 5370 1343 5375 1463
rect 5375 1343 5421 1463
rect 5421 1343 5426 1463
rect 4910 1224 4911 1267
rect 4911 1224 4965 1267
rect 4965 1224 4966 1267
rect 4910 1211 4966 1224
rect 5094 1224 5095 1267
rect 5095 1224 5149 1267
rect 5149 1224 5150 1267
rect 5094 1211 5150 1224
rect 5278 1224 5279 1267
rect 5279 1224 5333 1267
rect 5333 1224 5334 1267
rect 5278 1211 5334 1224
rect 4910 1061 4966 1117
rect 4102 945 4158 1001
rect 5094 945 5150 1001
rect 5423 945 5479 1001
rect 5856 945 5912 1001
rect 3966 829 4022 885
rect 5278 829 5334 885
rect 4910 722 4966 735
rect 4910 679 4911 722
rect 4911 679 4965 722
rect 4965 679 4966 722
rect 5094 722 5150 735
rect 5094 679 5095 722
rect 5095 679 5149 722
rect 5149 679 5150 722
rect 5278 722 5334 735
rect 5278 679 5279 722
rect 5279 679 5333 722
rect 5333 679 5334 722
rect 5370 483 5375 603
rect 5375 483 5421 603
rect 5421 483 5426 603
rect 4685 160 4741 216
rect 5503 160 5559 216
rect -109 42 -53 98
rect 90 42 146 98
rect 8280 3034 8336 3090
rect 9320 3034 9376 3090
rect 6396 2928 6452 2941
rect 6396 2885 6397 2928
rect 6397 2885 6451 2928
rect 6451 2885 6452 2928
rect 6580 2928 6636 2941
rect 6580 2885 6581 2928
rect 6581 2885 6635 2928
rect 6635 2885 6636 2928
rect 6764 2928 6820 2941
rect 6764 2885 6765 2928
rect 6765 2885 6819 2928
rect 6819 2885 6820 2928
rect 6856 2689 6861 2809
rect 6861 2689 6907 2809
rect 6907 2689 6912 2809
rect 6171 2366 6227 2422
rect 6989 2366 7045 2422
rect 10806 3035 10862 3091
rect 8952 2927 9008 2940
rect 8952 2884 8953 2927
rect 8953 2884 9007 2927
rect 9007 2884 9008 2927
rect 9136 2927 9192 2940
rect 9136 2884 9137 2927
rect 9137 2884 9191 2927
rect 9191 2884 9192 2927
rect 9320 2927 9376 2940
rect 9320 2884 9321 2927
rect 9321 2884 9375 2927
rect 9375 2884 9376 2927
rect 9412 2688 9417 2808
rect 9417 2688 9463 2808
rect 9463 2688 9468 2808
rect 8727 2365 8783 2421
rect 9545 2365 9601 2421
rect 9898 2247 9954 2303
rect 9722 2139 9778 2193
rect 9228 2030 9284 2086
rect 8860 1643 8865 1763
rect 8865 1643 8911 1763
rect 8911 1643 8916 1763
rect 9228 1643 9233 1763
rect 9233 1643 9279 1763
rect 9279 1643 9284 1763
rect 9044 1343 9049 1463
rect 9049 1343 9095 1463
rect 9095 1343 9100 1463
rect 9550 1642 9555 1763
rect 9555 1642 9601 1763
rect 9601 1642 9606 1763
rect 9412 1343 9417 1463
rect 9417 1343 9463 1463
rect 9463 1343 9468 1463
rect 8952 1224 8953 1267
rect 8953 1224 9007 1267
rect 9007 1224 9008 1267
rect 8952 1211 9008 1224
rect 9136 1224 9137 1267
rect 9137 1224 9191 1267
rect 9191 1224 9192 1267
rect 9136 1211 9192 1224
rect 9320 1224 9321 1267
rect 9321 1224 9375 1267
rect 9375 1224 9376 1267
rect 9320 1211 9376 1224
rect 8952 1061 9008 1117
rect 8144 945 8200 1001
rect 9136 945 9192 1001
rect 9465 945 9521 1001
rect 9898 945 9954 1001
rect 7978 829 8034 885
rect 9320 829 9376 885
rect 8952 722 9008 735
rect 8952 679 8953 722
rect 8953 679 9007 722
rect 9007 679 9008 722
rect 9136 722 9192 735
rect 9136 679 9137 722
rect 9137 679 9191 722
rect 9191 679 9192 722
rect 9320 722 9376 735
rect 9320 679 9321 722
rect 9321 679 9375 722
rect 9375 679 9376 722
rect 9412 483 9417 603
rect 9417 483 9463 603
rect 9463 483 9468 603
rect 8727 160 8783 216
rect 9545 160 9601 216
rect 3830 42 3886 98
rect 4102 42 4158 98
rect 12322 3034 12378 3090
rect 13362 3034 13418 3090
rect 10438 2928 10494 2941
rect 10438 2885 10439 2928
rect 10439 2885 10493 2928
rect 10493 2885 10494 2928
rect 10622 2928 10678 2941
rect 10622 2885 10623 2928
rect 10623 2885 10677 2928
rect 10677 2885 10678 2928
rect 10806 2928 10862 2941
rect 10806 2885 10807 2928
rect 10807 2885 10861 2928
rect 10861 2885 10862 2928
rect 10898 2689 10903 2809
rect 10903 2689 10949 2809
rect 10949 2689 10954 2809
rect 10213 2366 10269 2422
rect 11031 2366 11087 2422
rect 14848 3035 14904 3091
rect 12994 2927 13050 2940
rect 12994 2884 12995 2927
rect 12995 2884 13049 2927
rect 13049 2884 13050 2927
rect 13178 2927 13234 2940
rect 13178 2884 13179 2927
rect 13179 2884 13233 2927
rect 13233 2884 13234 2927
rect 13362 2927 13418 2940
rect 13362 2884 13363 2927
rect 13363 2884 13417 2927
rect 13417 2884 13418 2927
rect 13454 2688 13459 2808
rect 13459 2688 13505 2808
rect 13505 2688 13510 2808
rect 12769 2365 12825 2421
rect 13587 2365 13643 2421
rect 13940 2247 13996 2303
rect 13764 2139 13820 2193
rect 13270 2030 13326 2086
rect 12902 1643 12907 1763
rect 12907 1643 12953 1763
rect 12953 1643 12958 1763
rect 13270 1643 13275 1763
rect 13275 1643 13321 1763
rect 13321 1643 13326 1763
rect 13086 1343 13091 1463
rect 13091 1343 13137 1463
rect 13137 1343 13142 1463
rect 13592 1642 13597 1763
rect 13597 1642 13643 1763
rect 13643 1642 13648 1763
rect 13454 1343 13459 1463
rect 13459 1343 13505 1463
rect 13505 1343 13510 1463
rect 12994 1224 12995 1267
rect 12995 1224 13049 1267
rect 13049 1224 13050 1267
rect 12994 1211 13050 1224
rect 13178 1224 13179 1267
rect 13179 1224 13233 1267
rect 13233 1224 13234 1267
rect 13178 1211 13234 1224
rect 13362 1224 13363 1267
rect 13363 1224 13417 1267
rect 13417 1224 13418 1267
rect 13362 1211 13418 1224
rect 12994 1061 13050 1117
rect 12186 945 12242 1001
rect 13178 945 13234 1001
rect 13507 945 13563 1001
rect 13940 945 13996 1001
rect 12020 829 12076 885
rect 13362 829 13418 885
rect 12994 722 13050 735
rect 12994 679 12995 722
rect 12995 679 13049 722
rect 13049 679 13050 722
rect 13178 722 13234 735
rect 13178 679 13179 722
rect 13179 679 13233 722
rect 13233 679 13234 722
rect 13362 722 13418 735
rect 13362 679 13363 722
rect 13363 679 13417 722
rect 13417 679 13418 722
rect 13454 483 13459 603
rect 13459 483 13505 603
rect 13505 483 13510 603
rect 12769 160 12825 216
rect 13587 160 13643 216
rect 7842 42 7898 98
rect 8144 42 8200 98
rect 16364 3034 16420 3090
rect 17404 3034 17460 3090
rect 14480 2928 14536 2941
rect 14480 2885 14481 2928
rect 14481 2885 14535 2928
rect 14535 2885 14536 2928
rect 14664 2928 14720 2941
rect 14664 2885 14665 2928
rect 14665 2885 14719 2928
rect 14719 2885 14720 2928
rect 14848 2928 14904 2941
rect 14848 2885 14849 2928
rect 14849 2885 14903 2928
rect 14903 2885 14904 2928
rect 14940 2689 14945 2809
rect 14945 2689 14991 2809
rect 14991 2689 14996 2809
rect 14255 2366 14311 2422
rect 15073 2366 15129 2422
rect 18890 3035 18946 3091
rect 17036 2927 17092 2940
rect 17036 2884 17037 2927
rect 17037 2884 17091 2927
rect 17091 2884 17092 2927
rect 17220 2927 17276 2940
rect 17220 2884 17221 2927
rect 17221 2884 17275 2927
rect 17275 2884 17276 2927
rect 17404 2927 17460 2940
rect 17404 2884 17405 2927
rect 17405 2884 17459 2927
rect 17459 2884 17460 2927
rect 17496 2688 17501 2808
rect 17501 2688 17547 2808
rect 17547 2688 17552 2808
rect 16811 2365 16867 2421
rect 17629 2365 17685 2421
rect 17982 2247 18038 2303
rect 17806 2139 17862 2193
rect 17312 2030 17368 2086
rect 16944 1643 16949 1763
rect 16949 1643 16995 1763
rect 16995 1643 17000 1763
rect 17312 1643 17317 1763
rect 17317 1643 17363 1763
rect 17363 1643 17368 1763
rect 17128 1343 17133 1463
rect 17133 1343 17179 1463
rect 17179 1343 17184 1463
rect 17634 1642 17639 1763
rect 17639 1642 17685 1763
rect 17685 1642 17690 1763
rect 17496 1343 17501 1463
rect 17501 1343 17547 1463
rect 17547 1343 17552 1463
rect 17036 1224 17037 1267
rect 17037 1224 17091 1267
rect 17091 1224 17092 1267
rect 17036 1211 17092 1224
rect 17220 1224 17221 1267
rect 17221 1224 17275 1267
rect 17275 1224 17276 1267
rect 17220 1211 17276 1224
rect 17404 1224 17405 1267
rect 17405 1224 17459 1267
rect 17459 1224 17460 1267
rect 17404 1211 17460 1224
rect 17036 1061 17092 1117
rect 16228 945 16284 1001
rect 17220 945 17276 1001
rect 17549 945 17605 1001
rect 17982 945 18038 1001
rect 16062 829 16118 885
rect 17404 829 17460 885
rect 17036 722 17092 735
rect 17036 679 17037 722
rect 17037 679 17091 722
rect 17091 679 17092 722
rect 17220 722 17276 735
rect 17220 679 17221 722
rect 17221 679 17275 722
rect 17275 679 17276 722
rect 17404 722 17460 735
rect 17404 679 17405 722
rect 17405 679 17459 722
rect 17459 679 17460 722
rect 17496 483 17501 603
rect 17501 483 17547 603
rect 17547 483 17552 603
rect 16811 160 16867 216
rect 17629 160 17685 216
rect 11884 42 11940 98
rect 12186 42 12242 98
rect 20406 3034 20462 3090
rect 21446 3034 21502 3090
rect 18522 2928 18578 2941
rect 18522 2885 18523 2928
rect 18523 2885 18577 2928
rect 18577 2885 18578 2928
rect 18706 2928 18762 2941
rect 18706 2885 18707 2928
rect 18707 2885 18761 2928
rect 18761 2885 18762 2928
rect 18890 2928 18946 2941
rect 18890 2885 18891 2928
rect 18891 2885 18945 2928
rect 18945 2885 18946 2928
rect 18982 2689 18987 2809
rect 18987 2689 19033 2809
rect 19033 2689 19038 2809
rect 18297 2366 18353 2422
rect 19115 2366 19171 2422
rect 22932 3035 22988 3091
rect 21078 2927 21134 2940
rect 21078 2884 21079 2927
rect 21079 2884 21133 2927
rect 21133 2884 21134 2927
rect 21262 2927 21318 2940
rect 21262 2884 21263 2927
rect 21263 2884 21317 2927
rect 21317 2884 21318 2927
rect 21446 2927 21502 2940
rect 21446 2884 21447 2927
rect 21447 2884 21501 2927
rect 21501 2884 21502 2927
rect 21538 2688 21543 2808
rect 21543 2688 21589 2808
rect 21589 2688 21594 2808
rect 20853 2365 20909 2421
rect 21671 2365 21727 2421
rect 22024 2247 22080 2303
rect 21848 2139 21904 2193
rect 21354 2030 21410 2086
rect 20986 1643 20991 1763
rect 20991 1643 21037 1763
rect 21037 1643 21042 1763
rect 21354 1643 21359 1763
rect 21359 1643 21405 1763
rect 21405 1643 21410 1763
rect 21170 1343 21175 1463
rect 21175 1343 21221 1463
rect 21221 1343 21226 1463
rect 21676 1642 21681 1763
rect 21681 1642 21727 1763
rect 21727 1642 21732 1763
rect 21538 1343 21543 1463
rect 21543 1343 21589 1463
rect 21589 1343 21594 1463
rect 21078 1224 21079 1267
rect 21079 1224 21133 1267
rect 21133 1224 21134 1267
rect 21078 1211 21134 1224
rect 21262 1224 21263 1267
rect 21263 1224 21317 1267
rect 21317 1224 21318 1267
rect 21262 1211 21318 1224
rect 21446 1224 21447 1267
rect 21447 1224 21501 1267
rect 21501 1224 21502 1267
rect 21446 1211 21502 1224
rect 21078 1061 21134 1117
rect 20270 945 20326 1001
rect 21262 945 21318 1001
rect 21591 945 21647 1001
rect 22024 945 22080 1001
rect 20104 829 20160 885
rect 21446 829 21502 885
rect 21078 722 21134 735
rect 21078 679 21079 722
rect 21079 679 21133 722
rect 21133 679 21134 722
rect 21262 722 21318 735
rect 21262 679 21263 722
rect 21263 679 21317 722
rect 21317 679 21318 722
rect 21446 722 21502 735
rect 21446 679 21447 722
rect 21447 679 21501 722
rect 21501 679 21502 722
rect 21538 483 21543 603
rect 21543 483 21589 603
rect 21589 483 21594 603
rect 20853 160 20909 216
rect 21671 160 21727 216
rect 15926 42 15982 98
rect 16228 42 16284 98
rect 24448 3034 24504 3090
rect 25488 3034 25544 3090
rect 22564 2928 22620 2941
rect 22564 2885 22565 2928
rect 22565 2885 22619 2928
rect 22619 2885 22620 2928
rect 22748 2928 22804 2941
rect 22748 2885 22749 2928
rect 22749 2885 22803 2928
rect 22803 2885 22804 2928
rect 22932 2928 22988 2941
rect 22932 2885 22933 2928
rect 22933 2885 22987 2928
rect 22987 2885 22988 2928
rect 23024 2689 23029 2809
rect 23029 2689 23075 2809
rect 23075 2689 23080 2809
rect 22339 2366 22395 2422
rect 23157 2366 23213 2422
rect 26974 3035 27030 3091
rect 25120 2927 25176 2940
rect 25120 2884 25121 2927
rect 25121 2884 25175 2927
rect 25175 2884 25176 2927
rect 25304 2927 25360 2940
rect 25304 2884 25305 2927
rect 25305 2884 25359 2927
rect 25359 2884 25360 2927
rect 25488 2927 25544 2940
rect 25488 2884 25489 2927
rect 25489 2884 25543 2927
rect 25543 2884 25544 2927
rect 25580 2688 25585 2808
rect 25585 2688 25631 2808
rect 25631 2688 25636 2808
rect 24895 2365 24951 2421
rect 25713 2365 25769 2421
rect 26066 2247 26122 2303
rect 25890 2139 25946 2193
rect 25396 2030 25452 2086
rect 25028 1643 25033 1763
rect 25033 1643 25079 1763
rect 25079 1643 25084 1763
rect 25396 1643 25401 1763
rect 25401 1643 25447 1763
rect 25447 1643 25452 1763
rect 25212 1343 25217 1463
rect 25217 1343 25263 1463
rect 25263 1343 25268 1463
rect 25718 1642 25723 1763
rect 25723 1642 25769 1763
rect 25769 1642 25774 1763
rect 25580 1343 25585 1463
rect 25585 1343 25631 1463
rect 25631 1343 25636 1463
rect 25120 1224 25121 1267
rect 25121 1224 25175 1267
rect 25175 1224 25176 1267
rect 25120 1211 25176 1224
rect 25304 1224 25305 1267
rect 25305 1224 25359 1267
rect 25359 1224 25360 1267
rect 25304 1211 25360 1224
rect 25488 1224 25489 1267
rect 25489 1224 25543 1267
rect 25543 1224 25544 1267
rect 25488 1211 25544 1224
rect 25120 1061 25176 1117
rect 24312 945 24368 1001
rect 25304 945 25360 1001
rect 25633 945 25689 1001
rect 26066 945 26122 1001
rect 24146 829 24202 885
rect 25488 829 25544 885
rect 25120 722 25176 735
rect 25120 679 25121 722
rect 25121 679 25175 722
rect 25175 679 25176 722
rect 25304 722 25360 735
rect 25304 679 25305 722
rect 25305 679 25359 722
rect 25359 679 25360 722
rect 25488 722 25544 735
rect 25488 679 25489 722
rect 25489 679 25543 722
rect 25543 679 25544 722
rect 25580 483 25585 603
rect 25585 483 25631 603
rect 25631 483 25636 603
rect 24895 160 24951 216
rect 25713 160 25769 216
rect 19968 42 20024 98
rect 20270 42 20326 98
rect 26606 2928 26662 2941
rect 26606 2885 26607 2928
rect 26607 2885 26661 2928
rect 26661 2885 26662 2928
rect 26790 2928 26846 2941
rect 26790 2885 26791 2928
rect 26791 2885 26845 2928
rect 26845 2885 26846 2928
rect 26974 2928 27030 2941
rect 26974 2885 26975 2928
rect 26975 2885 27029 2928
rect 27029 2885 27030 2928
rect 27066 2689 27071 2809
rect 27071 2689 27117 2809
rect 27117 2689 27122 2809
rect 26381 2366 26437 2422
rect 27199 2366 27255 2422
rect 24010 42 24066 98
rect 24312 42 24368 98
<< metal2 >>
rect 3900 18737 3970 18749
rect 3900 18681 3912 18737
rect 3968 18681 3970 18737
rect 3900 18679 3970 18681
rect 3546 17311 3616 17323
rect 3546 17255 3558 17311
rect 3614 17255 3616 17311
rect 3546 17253 3616 17255
rect 3274 10464 3344 10476
rect 3274 10408 3286 10464
rect 3342 10408 3344 10464
rect 3274 10396 3344 10408
rect -201 9514 10 9524
rect -201 9414 -46 9514
rect -201 9404 10 9414
rect 3286 9514 3342 10396
rect 3286 9404 3342 9414
rect -201 9004 10 9014
rect -201 8904 -46 9004
rect -201 8894 10 8904
rect -46 7744 10 8894
rect 806 8701 1552 8713
rect 806 8645 1174 8701
rect 1230 8645 1552 8701
rect 806 8633 1552 8645
rect 806 8380 862 8633
rect 1174 8380 1230 8633
rect 1496 8380 1552 8633
rect 794 8378 874 8380
rect 794 8258 806 8378
rect 862 8258 874 8378
rect 794 8256 874 8258
rect 1162 8378 1242 8380
rect 1162 8258 1174 8378
rect 1230 8258 1242 8378
rect 1162 8256 1242 8258
rect 1484 8378 1564 8380
rect 1484 8257 1496 8378
rect 1552 8257 1564 8378
rect 806 8248 862 8256
rect 1174 8248 1230 8256
rect 1484 8255 1564 8257
rect 1496 8247 1552 8255
rect 990 8080 1046 8088
rect 1358 8080 1414 8088
rect 978 8078 1467 8080
rect 978 7958 990 8078
rect 1046 7958 1358 8078
rect 1414 7958 1467 8078
rect 978 7956 1467 7958
rect 990 7948 1046 7956
rect 1358 7948 1467 7956
rect 886 7882 966 7892
rect 886 7826 898 7882
rect 954 7826 966 7882
rect 886 7816 966 7826
rect 1070 7882 1150 7892
rect 1070 7826 1082 7882
rect 1138 7826 1150 7882
rect 1070 7816 1150 7826
rect 1254 7882 1334 7892
rect 1254 7826 1266 7882
rect 1322 7826 1334 7882
rect 1254 7816 1334 7826
rect -58 7732 12 7744
rect 898 7734 954 7816
rect -58 7676 -46 7732
rect 10 7676 12 7732
rect -58 7664 12 7676
rect 886 7732 966 7734
rect 886 7676 898 7732
rect 954 7676 966 7732
rect 886 7674 966 7676
rect 214 7616 284 7628
rect 214 7560 226 7616
rect 282 7560 284 7616
rect 214 7548 284 7560
rect 78 5411 148 5425
rect 78 5355 90 5411
rect 146 5355 148 5411
rect 78 5343 148 5355
rect -330 4509 -260 4521
rect -330 4453 -318 4509
rect -262 4453 -260 4509
rect -330 4441 -260 4453
rect -318 -55 -262 4441
rect 90 1015 146 5343
rect 226 3102 282 7548
rect 898 7360 954 7674
rect 1082 7618 1138 7816
rect 1070 7616 1150 7618
rect 1070 7560 1082 7616
rect 1138 7560 1150 7616
rect 1070 7558 1150 7560
rect 1082 7360 1138 7558
rect 1266 7502 1322 7816
rect 1399 7618 1467 7948
rect 1399 7616 1479 7618
rect 1399 7560 1411 7616
rect 1467 7560 1479 7616
rect 1399 7558 1479 7560
rect 1666 7616 1736 7628
rect 1666 7560 1668 7616
rect 1724 7560 1736 7616
rect 1254 7500 1334 7502
rect 1254 7444 1266 7500
rect 1322 7444 1334 7500
rect 1254 7442 1334 7444
rect 1266 7360 1322 7442
rect 886 7350 966 7360
rect 886 7294 898 7350
rect 954 7294 966 7350
rect 886 7284 966 7294
rect 1070 7350 1150 7360
rect 1070 7294 1082 7350
rect 1138 7294 1150 7350
rect 1070 7284 1150 7294
rect 1254 7350 1334 7360
rect 1254 7294 1266 7350
rect 1322 7294 1334 7350
rect 1254 7284 1334 7294
rect 1399 7228 1467 7558
rect 1666 7550 1736 7560
rect 1358 7220 1467 7228
rect 1346 7218 1467 7220
rect 1346 7098 1358 7218
rect 1414 7098 1467 7218
rect 1346 7096 1467 7098
rect 1358 7088 1414 7096
rect 661 6831 1559 6843
rect 661 6775 673 6831
rect 729 6775 1491 6831
rect 1547 6775 1559 6831
rect 661 6763 1559 6775
rect 1668 6606 1724 7550
rect 1832 6713 1912 6723
rect 1832 6657 1844 6713
rect 1900 6657 1912 6713
rect 1832 6655 1912 6657
rect 1666 6603 1736 6606
rect 1666 6549 1668 6603
rect 1724 6549 1736 6603
rect 1666 6537 1736 6549
rect 806 6496 1552 6508
rect 806 6440 1174 6496
rect 1230 6440 1552 6496
rect 806 6428 1552 6440
rect 806 6175 862 6428
rect 1174 6175 1230 6428
rect 1496 6175 1552 6428
rect 794 6173 874 6175
rect 794 6053 806 6173
rect 862 6053 874 6173
rect 794 6051 874 6053
rect 1162 6173 1242 6175
rect 1162 6053 1174 6173
rect 1230 6053 1242 6173
rect 1162 6051 1242 6053
rect 1484 6173 1564 6175
rect 1484 6052 1496 6173
rect 1552 6052 1564 6173
rect 806 6043 862 6051
rect 1174 6043 1230 6051
rect 1484 6050 1564 6052
rect 1496 6042 1552 6050
rect 990 5875 1046 5883
rect 1358 5875 1414 5883
rect 978 5873 1467 5875
rect 978 5753 990 5873
rect 1046 5753 1358 5873
rect 1414 5753 1467 5873
rect 978 5751 1467 5753
rect 990 5743 1046 5751
rect 1358 5743 1467 5751
rect 886 5677 966 5687
rect 886 5621 898 5677
rect 954 5621 966 5677
rect 886 5611 966 5621
rect 1070 5677 1150 5687
rect 1070 5621 1082 5677
rect 1138 5621 1150 5677
rect 1070 5611 1150 5621
rect 1254 5677 1334 5687
rect 1254 5621 1266 5677
rect 1322 5621 1334 5677
rect 1254 5611 1334 5621
rect 898 5529 954 5611
rect 886 5527 966 5529
rect 886 5471 898 5527
rect 954 5471 966 5527
rect 886 5469 966 5471
rect 898 5155 954 5469
rect 1082 5413 1138 5611
rect 1070 5411 1150 5413
rect 1070 5355 1082 5411
rect 1138 5355 1150 5411
rect 1070 5353 1150 5355
rect 1082 5155 1138 5353
rect 1266 5297 1322 5611
rect 1399 5413 1467 5743
rect 1844 5421 1900 6655
rect 2292 6496 3038 6508
rect 2292 6440 2660 6496
rect 2716 6440 3038 6496
rect 2292 6428 3038 6440
rect 2292 6175 2348 6428
rect 2660 6175 2716 6428
rect 2982 6175 3038 6428
rect 2280 6173 2360 6175
rect 2280 6053 2292 6173
rect 2348 6053 2360 6173
rect 2280 6051 2360 6053
rect 2648 6173 2728 6175
rect 2648 6053 2660 6173
rect 2716 6053 2728 6173
rect 2648 6051 2728 6053
rect 2970 6173 3050 6175
rect 2970 6052 2982 6173
rect 3038 6052 3050 6173
rect 2292 6043 2348 6051
rect 2660 6043 2716 6051
rect 2970 6050 3050 6052
rect 2982 6042 3038 6050
rect 2476 5875 2532 5883
rect 2844 5875 2900 5883
rect 2464 5873 2953 5875
rect 2464 5753 2476 5873
rect 2532 5753 2844 5873
rect 2900 5753 2953 5873
rect 2464 5751 2953 5753
rect 2476 5743 2532 5751
rect 2844 5743 2953 5751
rect 2372 5677 2452 5687
rect 2372 5621 2384 5677
rect 2440 5621 2452 5677
rect 2372 5611 2452 5621
rect 2556 5677 2636 5687
rect 2556 5621 2568 5677
rect 2624 5621 2636 5677
rect 2556 5611 2636 5621
rect 2740 5677 2820 5687
rect 2740 5621 2752 5677
rect 2808 5621 2820 5677
rect 2740 5611 2820 5621
rect 2384 5529 2440 5611
rect 2372 5527 2452 5529
rect 2372 5471 2384 5527
rect 2440 5471 2452 5527
rect 2372 5469 2452 5471
rect 1399 5411 1479 5413
rect 1399 5355 1411 5411
rect 1467 5355 1479 5411
rect 1399 5353 1479 5355
rect 1842 5411 1902 5421
rect 1842 5355 1844 5411
rect 1900 5355 1902 5411
rect 1254 5295 1334 5297
rect 1254 5239 1266 5295
rect 1322 5239 1334 5295
rect 1254 5237 1334 5239
rect 1266 5155 1322 5237
rect 886 5145 966 5155
rect 886 5089 898 5145
rect 954 5089 966 5145
rect 886 5079 966 5089
rect 1070 5145 1150 5155
rect 1070 5089 1082 5145
rect 1138 5089 1150 5145
rect 1070 5079 1150 5089
rect 1254 5145 1334 5155
rect 1254 5089 1266 5145
rect 1322 5089 1334 5145
rect 1254 5079 1334 5089
rect 1399 5023 1467 5353
rect 1842 5343 1902 5355
rect 1358 5015 1467 5023
rect 1346 5013 1467 5015
rect 1346 4893 1358 5013
rect 1414 4893 1467 5013
rect 1346 4891 1467 4893
rect 1358 4883 1414 4891
rect 661 4626 1557 4638
rect 661 4570 673 4626
rect 729 4570 1491 4626
rect 1547 4570 1557 4626
rect 661 4558 1557 4570
rect 1844 4400 1900 5343
rect 2384 5155 2440 5469
rect 2568 5413 2624 5611
rect 2556 5411 2636 5413
rect 2556 5355 2568 5411
rect 2624 5355 2636 5411
rect 2556 5353 2636 5355
rect 2568 5155 2624 5353
rect 2752 5297 2808 5611
rect 2885 5413 2953 5743
rect 2885 5411 2965 5413
rect 2885 5355 2897 5411
rect 2953 5355 2965 5411
rect 2885 5353 2965 5355
rect 3152 5411 3222 5423
rect 3152 5355 3154 5411
rect 3210 5355 3478 5411
rect 2740 5295 2820 5297
rect 2740 5239 2752 5295
rect 2808 5239 2820 5295
rect 2740 5237 2820 5239
rect 2752 5155 2808 5237
rect 2372 5145 2452 5155
rect 2372 5089 2384 5145
rect 2440 5089 2452 5145
rect 2372 5079 2452 5089
rect 2556 5145 2636 5155
rect 2556 5089 2568 5145
rect 2624 5089 2636 5145
rect 2556 5079 2636 5089
rect 2740 5145 2820 5155
rect 2740 5089 2752 5145
rect 2808 5089 2820 5145
rect 2740 5079 2820 5089
rect 2885 5023 2953 5353
rect 3152 5345 3222 5355
rect 2844 5015 2953 5023
rect 2832 5013 2953 5015
rect 2832 4893 2844 5013
rect 2900 4893 2953 5013
rect 2832 4891 2953 4893
rect 2844 4883 2900 4891
rect 2147 4626 3043 4638
rect 2147 4570 2159 4626
rect 2215 4570 2977 4626
rect 3033 4570 3043 4626
rect 2147 4558 3043 4570
rect 3154 4401 3210 5345
rect 3318 4509 3398 4519
rect 3318 4453 3330 4509
rect 3386 4453 3398 4509
rect 3318 4451 3398 4453
rect 1842 4398 1912 4400
rect 1842 4342 1844 4398
rect 1900 4342 1912 4398
rect 1842 4330 1912 4342
rect 3142 4399 3222 4401
rect 3142 4343 3154 4399
rect 3210 4343 3222 4399
rect 3142 4331 3222 4343
rect 806 4291 1552 4303
rect 806 4235 1174 4291
rect 1230 4235 1552 4291
rect 806 4223 1552 4235
rect 806 3970 862 4223
rect 1174 3970 1230 4223
rect 1496 3970 1552 4223
rect 2292 4292 3038 4304
rect 2292 4236 2660 4292
rect 2716 4236 3038 4292
rect 2292 4224 3038 4236
rect 2292 3971 2348 4224
rect 2660 3971 2716 4224
rect 2982 3971 3038 4224
rect 794 3968 874 3970
rect 794 3848 806 3968
rect 862 3848 874 3968
rect 794 3846 874 3848
rect 1162 3968 1242 3970
rect 1162 3848 1174 3968
rect 1230 3848 1242 3968
rect 1162 3846 1242 3848
rect 1484 3968 1564 3970
rect 1484 3847 1496 3968
rect 1552 3847 1564 3968
rect 2280 3969 2360 3971
rect 2280 3849 2292 3969
rect 2348 3849 2360 3969
rect 2280 3847 2360 3849
rect 2648 3969 2728 3971
rect 2648 3849 2660 3969
rect 2716 3849 2728 3969
rect 2648 3847 2728 3849
rect 2970 3969 3050 3971
rect 2970 3848 2982 3969
rect 3038 3848 3050 3969
rect 806 3838 862 3846
rect 1174 3838 1230 3846
rect 1484 3845 1564 3847
rect 1496 3837 1552 3845
rect 2292 3839 2348 3847
rect 2660 3839 2716 3847
rect 2970 3846 3050 3848
rect 2982 3838 3038 3846
rect 990 3670 1046 3678
rect 1358 3670 1414 3678
rect 2476 3671 2532 3679
rect 2844 3671 2900 3679
rect 978 3668 1467 3670
rect 978 3548 990 3668
rect 1046 3548 1358 3668
rect 1414 3548 1467 3668
rect 978 3546 1467 3548
rect 2464 3669 2953 3671
rect 2464 3549 2476 3669
rect 2532 3549 2844 3669
rect 2900 3549 2953 3669
rect 2464 3547 2953 3549
rect 990 3538 1046 3546
rect 1358 3538 1467 3546
rect 2476 3539 2532 3547
rect 2844 3539 2953 3547
rect 886 3472 966 3482
rect 886 3416 898 3472
rect 954 3416 966 3472
rect 886 3406 966 3416
rect 1070 3472 1150 3482
rect 1070 3416 1082 3472
rect 1138 3416 1150 3472
rect 1070 3406 1150 3416
rect 1254 3472 1334 3482
rect 1254 3416 1266 3472
rect 1322 3416 1334 3472
rect 1254 3406 1334 3416
rect 898 3324 954 3406
rect 886 3322 966 3324
rect 886 3266 898 3322
rect 954 3266 966 3322
rect 886 3264 966 3266
rect 214 3090 284 3102
rect 214 3034 226 3090
rect 282 3034 284 3090
rect 214 3022 284 3034
rect 898 2950 954 3264
rect 1082 3208 1138 3406
rect 1070 3206 1150 3208
rect 1070 3150 1082 3206
rect 1138 3150 1150 3206
rect 1070 3148 1150 3150
rect 1082 2950 1138 3148
rect 1266 3092 1322 3406
rect 1399 3208 1467 3538
rect 2372 3473 2452 3483
rect 2372 3417 2384 3473
rect 2440 3417 2452 3473
rect 2372 3407 2452 3417
rect 2556 3473 2636 3483
rect 2556 3417 2568 3473
rect 2624 3417 2636 3473
rect 2556 3407 2636 3417
rect 2740 3473 2820 3483
rect 2740 3417 2752 3473
rect 2808 3417 2820 3473
rect 2740 3407 2820 3417
rect 2384 3325 2440 3407
rect 2372 3323 2452 3325
rect 2372 3267 2384 3323
rect 2440 3267 2452 3323
rect 2372 3265 2452 3267
rect 1399 3206 1479 3208
rect 1399 3150 1411 3206
rect 1467 3150 1479 3206
rect 1399 3148 1479 3150
rect 1666 3206 1736 3218
rect 1666 3150 1668 3206
rect 1724 3150 1736 3206
rect 1254 3090 1334 3092
rect 1254 3034 1266 3090
rect 1322 3034 1334 3090
rect 1254 3032 1334 3034
rect 1266 2950 1322 3032
rect 886 2940 966 2950
rect 886 2884 898 2940
rect 954 2884 966 2940
rect 886 2874 966 2884
rect 1070 2940 1150 2950
rect 1070 2884 1082 2940
rect 1138 2884 1150 2940
rect 1070 2874 1150 2884
rect 1254 2940 1334 2950
rect 1254 2884 1266 2940
rect 1322 2884 1334 2940
rect 1254 2874 1334 2884
rect 1399 2818 1467 3148
rect 1666 3140 1736 3150
rect 1358 2810 1467 2818
rect 1346 2808 1467 2810
rect 1346 2688 1358 2808
rect 1414 2688 1467 2808
rect 1346 2686 1467 2688
rect 1358 2678 1414 2686
rect 661 2421 1557 2433
rect 661 2365 673 2421
rect 729 2365 1491 2421
rect 1547 2365 1557 2421
rect 661 2353 1557 2365
rect 1668 2196 1724 3140
rect 2384 2951 2440 3265
rect 2568 3209 2624 3407
rect 2556 3207 2636 3209
rect 2556 3151 2568 3207
rect 2624 3151 2636 3207
rect 2556 3149 2636 3151
rect 2568 2951 2624 3149
rect 2752 3093 2808 3407
rect 2885 3209 2953 3539
rect 3330 3217 3386 4451
rect 2885 3207 2965 3209
rect 2885 3151 2897 3207
rect 2953 3151 2965 3207
rect 2885 3149 2965 3151
rect 3328 3207 3398 3217
rect 3558 3207 3614 17253
rect 3912 14090 3968 18679
rect 4818 18280 5564 18292
rect 4818 18224 5186 18280
rect 5242 18224 5564 18280
rect 4818 18212 5564 18224
rect 4818 17959 4874 18212
rect 5186 17959 5242 18212
rect 5508 17959 5564 18212
rect 4806 17957 4886 17959
rect 4806 17837 4818 17957
rect 4874 17837 4886 17957
rect 4806 17835 4886 17837
rect 5174 17957 5254 17959
rect 5174 17837 5186 17957
rect 5242 17837 5254 17957
rect 5174 17835 5254 17837
rect 5496 17957 5576 17959
rect 5496 17836 5508 17957
rect 5564 17836 5576 17957
rect 4818 17827 4874 17835
rect 5186 17827 5242 17835
rect 5496 17834 5576 17836
rect 5508 17826 5564 17834
rect 5002 17659 5058 17667
rect 5370 17659 5426 17667
rect 4990 17657 5479 17659
rect 4990 17537 5002 17657
rect 5058 17537 5370 17657
rect 5426 17537 5479 17657
rect 4990 17535 5479 17537
rect 5002 17527 5058 17535
rect 5370 17527 5479 17535
rect 4898 17461 4978 17471
rect 4898 17405 4910 17461
rect 4966 17405 4978 17461
rect 4898 17395 4978 17405
rect 5082 17461 5162 17471
rect 5082 17405 5094 17461
rect 5150 17405 5162 17461
rect 5082 17395 5162 17405
rect 5266 17461 5346 17471
rect 5266 17405 5278 17461
rect 5334 17405 5346 17461
rect 5266 17395 5346 17405
rect 4910 17313 4966 17395
rect 4898 17311 4978 17313
rect 4898 17255 4910 17311
rect 4966 17255 4978 17311
rect 4898 17253 4978 17255
rect 4226 17195 4296 17207
rect 4226 17139 4238 17195
rect 4294 17139 4296 17195
rect 4226 17127 4296 17139
rect 4090 14990 4160 15004
rect 4090 14934 4102 14990
rect 4158 14934 4160 14990
rect 4090 14922 4160 14934
rect 3900 14088 3970 14090
rect 3900 14032 3912 14088
rect 3968 14032 3970 14088
rect 3900 14020 3970 14032
rect 4102 10594 4158 14922
rect 4238 12681 4294 17127
rect 4910 16939 4966 17253
rect 5094 17197 5150 17395
rect 5082 17195 5162 17197
rect 5082 17139 5094 17195
rect 5150 17139 5162 17195
rect 5082 17137 5162 17139
rect 5094 16939 5150 17137
rect 5278 17081 5334 17395
rect 5411 17197 5479 17527
rect 7558 17308 7628 17320
rect 7558 17252 7570 17308
rect 7626 17252 7628 17308
rect 7558 17250 7628 17252
rect 5411 17195 5491 17197
rect 5411 17139 5423 17195
rect 5479 17139 5491 17195
rect 5411 17137 5491 17139
rect 5678 17195 5748 17207
rect 5678 17139 5680 17195
rect 5736 17139 5748 17195
rect 5266 17079 5346 17081
rect 5266 17023 5278 17079
rect 5334 17023 5346 17079
rect 5266 17021 5346 17023
rect 5278 16939 5334 17021
rect 4898 16929 4978 16939
rect 4898 16873 4910 16929
rect 4966 16873 4978 16929
rect 4898 16863 4978 16873
rect 5082 16929 5162 16939
rect 5082 16873 5094 16929
rect 5150 16873 5162 16929
rect 5082 16863 5162 16873
rect 5266 16929 5346 16939
rect 5266 16873 5278 16929
rect 5334 16873 5346 16929
rect 5266 16863 5346 16873
rect 5411 16807 5479 17137
rect 5678 17129 5748 17139
rect 5370 16799 5479 16807
rect 5358 16797 5479 16799
rect 5358 16677 5370 16797
rect 5426 16677 5479 16797
rect 5358 16675 5479 16677
rect 5370 16667 5426 16675
rect 4673 16410 5571 16422
rect 4673 16354 4685 16410
rect 4741 16354 5503 16410
rect 5559 16354 5571 16410
rect 4673 16342 5571 16354
rect 5680 16185 5736 17129
rect 5844 16292 5924 16302
rect 5844 16236 5856 16292
rect 5912 16236 5924 16292
rect 5844 16234 5924 16236
rect 5678 16182 5748 16185
rect 5678 16128 5680 16182
rect 5736 16128 5748 16182
rect 5678 16116 5748 16128
rect 4818 16075 5564 16087
rect 4818 16019 5186 16075
rect 5242 16019 5564 16075
rect 4818 16007 5564 16019
rect 4818 15754 4874 16007
rect 5186 15754 5242 16007
rect 5508 15754 5564 16007
rect 4806 15752 4886 15754
rect 4806 15632 4818 15752
rect 4874 15632 4886 15752
rect 4806 15630 4886 15632
rect 5174 15752 5254 15754
rect 5174 15632 5186 15752
rect 5242 15632 5254 15752
rect 5174 15630 5254 15632
rect 5496 15752 5576 15754
rect 5496 15631 5508 15752
rect 5564 15631 5576 15752
rect 4818 15622 4874 15630
rect 5186 15622 5242 15630
rect 5496 15629 5576 15631
rect 5508 15621 5564 15629
rect 5002 15454 5058 15462
rect 5370 15454 5426 15462
rect 4990 15452 5479 15454
rect 4990 15332 5002 15452
rect 5058 15332 5370 15452
rect 5426 15332 5479 15452
rect 4990 15330 5479 15332
rect 5002 15322 5058 15330
rect 5370 15322 5479 15330
rect 4898 15256 4978 15266
rect 4898 15200 4910 15256
rect 4966 15200 4978 15256
rect 4898 15190 4978 15200
rect 5082 15256 5162 15266
rect 5082 15200 5094 15256
rect 5150 15200 5162 15256
rect 5082 15190 5162 15200
rect 5266 15256 5346 15266
rect 5266 15200 5278 15256
rect 5334 15200 5346 15256
rect 5266 15190 5346 15200
rect 4910 15108 4966 15190
rect 4898 15106 4978 15108
rect 4898 15050 4910 15106
rect 4966 15050 4978 15106
rect 4898 15048 4978 15050
rect 4910 14734 4966 15048
rect 5094 14992 5150 15190
rect 5082 14990 5162 14992
rect 5082 14934 5094 14990
rect 5150 14934 5162 14990
rect 5082 14932 5162 14934
rect 5094 14734 5150 14932
rect 5278 14876 5334 15190
rect 5411 14992 5479 15322
rect 5856 15000 5912 16234
rect 6304 16075 7050 16087
rect 6304 16019 6672 16075
rect 6728 16019 7050 16075
rect 6304 16007 7050 16019
rect 6304 15754 6360 16007
rect 6672 15754 6728 16007
rect 6994 15754 7050 16007
rect 6292 15752 6372 15754
rect 6292 15632 6304 15752
rect 6360 15632 6372 15752
rect 6292 15630 6372 15632
rect 6660 15752 6740 15754
rect 6660 15632 6672 15752
rect 6728 15632 6740 15752
rect 6660 15630 6740 15632
rect 6982 15752 7062 15754
rect 6982 15631 6994 15752
rect 7050 15631 7062 15752
rect 6304 15622 6360 15630
rect 6672 15622 6728 15630
rect 6982 15629 7062 15631
rect 6994 15621 7050 15629
rect 6488 15454 6544 15462
rect 6856 15454 6912 15462
rect 6476 15452 6965 15454
rect 6476 15332 6488 15452
rect 6544 15332 6856 15452
rect 6912 15332 6965 15452
rect 6476 15330 6965 15332
rect 6488 15322 6544 15330
rect 6856 15322 6965 15330
rect 6384 15256 6464 15266
rect 6384 15200 6396 15256
rect 6452 15200 6464 15256
rect 6384 15190 6464 15200
rect 6568 15256 6648 15266
rect 6568 15200 6580 15256
rect 6636 15200 6648 15256
rect 6568 15190 6648 15200
rect 6752 15256 6832 15266
rect 6752 15200 6764 15256
rect 6820 15200 6832 15256
rect 6752 15190 6832 15200
rect 6396 15108 6452 15190
rect 6384 15106 6464 15108
rect 6384 15050 6396 15106
rect 6452 15050 6464 15106
rect 6384 15048 6464 15050
rect 5411 14990 5491 14992
rect 5411 14934 5423 14990
rect 5479 14934 5491 14990
rect 5411 14932 5491 14934
rect 5854 14990 5914 15000
rect 5854 14934 5856 14990
rect 5912 14934 5914 14990
rect 5266 14874 5346 14876
rect 5266 14818 5278 14874
rect 5334 14818 5346 14874
rect 5266 14816 5346 14818
rect 5278 14734 5334 14816
rect 4898 14724 4978 14734
rect 4898 14668 4910 14724
rect 4966 14668 4978 14724
rect 4898 14658 4978 14668
rect 5082 14724 5162 14734
rect 5082 14668 5094 14724
rect 5150 14668 5162 14724
rect 5082 14658 5162 14668
rect 5266 14724 5346 14734
rect 5266 14668 5278 14724
rect 5334 14668 5346 14724
rect 5266 14658 5346 14668
rect 5411 14602 5479 14932
rect 5854 14922 5914 14934
rect 5370 14594 5479 14602
rect 5358 14592 5479 14594
rect 5358 14472 5370 14592
rect 5426 14472 5479 14592
rect 5358 14470 5479 14472
rect 5370 14462 5426 14470
rect 4673 14205 5569 14217
rect 4673 14149 4685 14205
rect 4741 14149 5503 14205
rect 5559 14149 5569 14205
rect 4673 14137 5569 14149
rect 5856 13979 5912 14922
rect 6396 14734 6452 15048
rect 6580 14992 6636 15190
rect 6568 14990 6648 14992
rect 6568 14934 6580 14990
rect 6636 14934 6648 14990
rect 6568 14932 6648 14934
rect 6580 14734 6636 14932
rect 6764 14876 6820 15190
rect 6897 14992 6965 15322
rect 6897 14990 6977 14992
rect 6897 14934 6909 14990
rect 6965 14934 6977 14990
rect 6897 14932 6977 14934
rect 7164 14990 7234 15002
rect 7164 14934 7166 14990
rect 7222 14934 7490 14990
rect 6752 14874 6832 14876
rect 6752 14818 6764 14874
rect 6820 14818 6832 14874
rect 6752 14816 6832 14818
rect 6764 14734 6820 14816
rect 6384 14724 6464 14734
rect 6384 14668 6396 14724
rect 6452 14668 6464 14724
rect 6384 14658 6464 14668
rect 6568 14724 6648 14734
rect 6568 14668 6580 14724
rect 6636 14668 6648 14724
rect 6568 14658 6648 14668
rect 6752 14724 6832 14734
rect 6752 14668 6764 14724
rect 6820 14668 6832 14724
rect 6752 14658 6832 14668
rect 6897 14602 6965 14932
rect 7164 14924 7234 14934
rect 6856 14594 6965 14602
rect 6844 14592 6965 14594
rect 6844 14472 6856 14592
rect 6912 14472 6965 14592
rect 6844 14470 6965 14472
rect 6856 14462 6912 14470
rect 6159 14205 7055 14217
rect 6159 14149 6171 14205
rect 6227 14149 6989 14205
rect 7045 14149 7055 14205
rect 6159 14137 7055 14149
rect 7166 13980 7222 14924
rect 7330 14088 7410 14098
rect 7330 14032 7342 14088
rect 7398 14032 7410 14088
rect 7330 14030 7410 14032
rect 5854 13977 5924 13979
rect 5854 13921 5856 13977
rect 5912 13921 5924 13977
rect 5854 13909 5924 13921
rect 7154 13978 7234 13980
rect 7154 13922 7166 13978
rect 7222 13922 7234 13978
rect 7154 13910 7234 13922
rect 4818 13870 5564 13882
rect 4818 13814 5186 13870
rect 5242 13814 5564 13870
rect 4818 13802 5564 13814
rect 4818 13549 4874 13802
rect 5186 13549 5242 13802
rect 5508 13549 5564 13802
rect 6304 13871 7050 13883
rect 6304 13815 6672 13871
rect 6728 13815 7050 13871
rect 6304 13803 7050 13815
rect 6304 13550 6360 13803
rect 6672 13550 6728 13803
rect 6994 13550 7050 13803
rect 4806 13547 4886 13549
rect 4806 13427 4818 13547
rect 4874 13427 4886 13547
rect 4806 13425 4886 13427
rect 5174 13547 5254 13549
rect 5174 13427 5186 13547
rect 5242 13427 5254 13547
rect 5174 13425 5254 13427
rect 5496 13547 5576 13549
rect 5496 13426 5508 13547
rect 5564 13426 5576 13547
rect 6292 13548 6372 13550
rect 6292 13428 6304 13548
rect 6360 13428 6372 13548
rect 6292 13426 6372 13428
rect 6660 13548 6740 13550
rect 6660 13428 6672 13548
rect 6728 13428 6740 13548
rect 6660 13426 6740 13428
rect 6982 13548 7062 13550
rect 6982 13427 6994 13548
rect 7050 13427 7062 13548
rect 4818 13417 4874 13425
rect 5186 13417 5242 13425
rect 5496 13424 5576 13426
rect 5508 13416 5564 13424
rect 6304 13418 6360 13426
rect 6672 13418 6728 13426
rect 6982 13425 7062 13427
rect 6994 13417 7050 13425
rect 5002 13249 5058 13257
rect 5370 13249 5426 13257
rect 6488 13250 6544 13258
rect 6856 13250 6912 13258
rect 4990 13247 5479 13249
rect 4990 13127 5002 13247
rect 5058 13127 5370 13247
rect 5426 13127 5479 13247
rect 4990 13125 5479 13127
rect 6476 13248 6965 13250
rect 6476 13128 6488 13248
rect 6544 13128 6856 13248
rect 6912 13128 6965 13248
rect 6476 13126 6965 13128
rect 5002 13117 5058 13125
rect 5370 13117 5479 13125
rect 6488 13118 6544 13126
rect 6856 13118 6965 13126
rect 4898 13051 4978 13061
rect 4898 12995 4910 13051
rect 4966 12995 4978 13051
rect 4898 12985 4978 12995
rect 5082 13051 5162 13061
rect 5082 12995 5094 13051
rect 5150 12995 5162 13051
rect 5082 12985 5162 12995
rect 5266 13051 5346 13061
rect 5266 12995 5278 13051
rect 5334 12995 5346 13051
rect 5266 12985 5346 12995
rect 4910 12903 4966 12985
rect 4898 12901 4978 12903
rect 4898 12845 4910 12901
rect 4966 12845 4978 12901
rect 4898 12843 4978 12845
rect 4226 12669 4296 12681
rect 4226 12613 4238 12669
rect 4294 12613 4296 12669
rect 4226 12601 4296 12613
rect 4910 12529 4966 12843
rect 5094 12787 5150 12985
rect 5082 12785 5162 12787
rect 5082 12729 5094 12785
rect 5150 12729 5162 12785
rect 5082 12727 5162 12729
rect 5094 12529 5150 12727
rect 5278 12671 5334 12985
rect 5411 12787 5479 13117
rect 6384 13052 6464 13062
rect 6384 12996 6396 13052
rect 6452 12996 6464 13052
rect 6384 12986 6464 12996
rect 6568 13052 6648 13062
rect 6568 12996 6580 13052
rect 6636 12996 6648 13052
rect 6568 12986 6648 12996
rect 6752 13052 6832 13062
rect 6752 12996 6764 13052
rect 6820 12996 6832 13052
rect 6752 12986 6832 12996
rect 6396 12904 6452 12986
rect 6384 12902 6464 12904
rect 6384 12846 6396 12902
rect 6452 12846 6464 12902
rect 6384 12844 6464 12846
rect 5411 12785 5491 12787
rect 5411 12729 5423 12785
rect 5479 12729 5491 12785
rect 5411 12727 5491 12729
rect 5678 12785 5748 12797
rect 5678 12729 5680 12785
rect 5736 12729 5748 12785
rect 5266 12669 5346 12671
rect 5266 12613 5278 12669
rect 5334 12613 5346 12669
rect 5266 12611 5346 12613
rect 5278 12529 5334 12611
rect 4898 12519 4978 12529
rect 4898 12463 4910 12519
rect 4966 12463 4978 12519
rect 4898 12453 4978 12463
rect 5082 12519 5162 12529
rect 5082 12463 5094 12519
rect 5150 12463 5162 12519
rect 5082 12453 5162 12463
rect 5266 12519 5346 12529
rect 5266 12463 5278 12519
rect 5334 12463 5346 12519
rect 5266 12453 5346 12463
rect 5411 12397 5479 12727
rect 5678 12719 5748 12729
rect 5370 12389 5479 12397
rect 5358 12387 5479 12389
rect 5358 12267 5370 12387
rect 5426 12267 5479 12387
rect 5358 12265 5479 12267
rect 5370 12257 5426 12265
rect 4673 12000 5569 12012
rect 4673 11944 4685 12000
rect 4741 11944 5503 12000
rect 5559 11944 5569 12000
rect 4673 11932 5569 11944
rect 5680 11775 5736 12719
rect 6396 12530 6452 12844
rect 6580 12788 6636 12986
rect 6568 12786 6648 12788
rect 6568 12730 6580 12786
rect 6636 12730 6648 12786
rect 6568 12728 6648 12730
rect 6580 12530 6636 12728
rect 6764 12672 6820 12986
rect 6897 12788 6965 13118
rect 7342 12796 7398 14030
rect 6897 12786 6977 12788
rect 6897 12730 6909 12786
rect 6965 12730 6977 12786
rect 6897 12728 6977 12730
rect 7340 12786 7410 12796
rect 7340 12730 7342 12786
rect 7398 12730 7490 12786
rect 6752 12670 6832 12672
rect 6752 12614 6764 12670
rect 6820 12614 6832 12670
rect 6752 12612 6832 12614
rect 6764 12530 6820 12612
rect 6384 12520 6464 12530
rect 6384 12464 6396 12520
rect 6452 12464 6464 12520
rect 6384 12454 6464 12464
rect 6568 12520 6648 12530
rect 6568 12464 6580 12520
rect 6636 12464 6648 12520
rect 6568 12454 6648 12464
rect 6752 12520 6832 12530
rect 6752 12464 6764 12520
rect 6820 12464 6832 12520
rect 6752 12454 6832 12464
rect 6897 12398 6965 12728
rect 7340 12718 7410 12730
rect 6856 12390 6965 12398
rect 6844 12388 6965 12390
rect 6844 12268 6856 12388
rect 6912 12268 6965 12388
rect 6844 12266 6965 12268
rect 6856 12258 6912 12266
rect 6159 12001 7055 12013
rect 6159 11945 6171 12001
rect 6227 11945 6989 12001
rect 7045 11945 7055 12001
rect 6159 11933 7055 11945
rect 5844 11882 5924 11892
rect 5844 11826 5856 11882
rect 5912 11826 5924 11882
rect 5844 11824 5924 11826
rect 5678 11772 5748 11775
rect 5678 11718 5680 11772
rect 5736 11718 5748 11772
rect 5678 11706 5748 11718
rect 4818 11665 5564 11677
rect 4818 11609 5186 11665
rect 5242 11609 5564 11665
rect 4818 11597 5564 11609
rect 4818 11344 4874 11597
rect 5186 11344 5242 11597
rect 5508 11344 5564 11597
rect 4806 11342 4886 11344
rect 4806 11222 4818 11342
rect 4874 11222 4886 11342
rect 4806 11220 4886 11222
rect 5174 11342 5254 11344
rect 5174 11222 5186 11342
rect 5242 11222 5254 11342
rect 5174 11220 5254 11222
rect 5496 11342 5576 11344
rect 5496 11221 5508 11342
rect 5564 11221 5576 11342
rect 4818 11212 4874 11220
rect 5186 11212 5242 11220
rect 5496 11219 5576 11221
rect 5508 11211 5564 11219
rect 5002 11044 5058 11052
rect 5370 11044 5426 11052
rect 4990 11042 5479 11044
rect 4990 10922 5002 11042
rect 5058 10922 5370 11042
rect 5426 10922 5479 11042
rect 4990 10920 5479 10922
rect 5002 10912 5058 10920
rect 5370 10912 5479 10920
rect 4898 10846 4978 10856
rect 4898 10790 4910 10846
rect 4966 10790 4978 10846
rect 4898 10780 4978 10790
rect 5082 10846 5162 10856
rect 5082 10790 5094 10846
rect 5150 10790 5162 10846
rect 5082 10780 5162 10790
rect 5266 10846 5346 10856
rect 5266 10790 5278 10846
rect 5334 10790 5346 10846
rect 5266 10780 5346 10790
rect 4910 10698 4966 10780
rect 4898 10696 4978 10698
rect 4898 10640 4910 10696
rect 4966 10640 4978 10696
rect 4898 10638 4978 10640
rect 4090 10580 4160 10594
rect 4090 10524 4102 10580
rect 4158 10524 4160 10580
rect 4090 10512 4160 10524
rect 3818 9677 3888 9689
rect 4102 9681 4158 10512
rect 4910 10324 4966 10638
rect 5094 10582 5150 10780
rect 5082 10580 5162 10582
rect 5082 10524 5094 10580
rect 5150 10524 5162 10580
rect 5082 10522 5162 10524
rect 5094 10324 5150 10522
rect 5278 10466 5334 10780
rect 5411 10582 5479 10912
rect 5856 10592 5912 11824
rect 5411 10580 5491 10582
rect 5411 10524 5423 10580
rect 5479 10524 5491 10580
rect 5411 10522 5491 10524
rect 5854 10580 5914 10592
rect 5854 10524 5856 10580
rect 5912 10524 5914 10580
rect 5266 10464 5346 10466
rect 5266 10408 5278 10464
rect 5334 10408 5346 10464
rect 5266 10406 5346 10408
rect 5278 10324 5334 10406
rect 4898 10314 4978 10324
rect 4898 10258 4910 10314
rect 4966 10258 4978 10314
rect 4898 10248 4978 10258
rect 5082 10314 5162 10324
rect 5082 10258 5094 10314
rect 5150 10258 5162 10314
rect 5082 10248 5162 10258
rect 5266 10314 5346 10324
rect 5266 10258 5278 10314
rect 5334 10258 5346 10314
rect 5266 10248 5346 10258
rect 5411 10192 5479 10522
rect 5854 10512 5914 10524
rect 7286 10461 7356 10473
rect 7286 10405 7298 10461
rect 7354 10405 7356 10461
rect 7286 10393 7356 10405
rect 5370 10184 5479 10192
rect 5358 10182 5479 10184
rect 5358 10062 5370 10182
rect 5426 10062 5479 10182
rect 5358 10060 5479 10062
rect 5370 10052 5426 10060
rect 4673 9795 5571 9807
rect 4673 9739 4685 9795
rect 4741 9739 5503 9795
rect 5559 9739 5571 9795
rect 4673 9727 5571 9739
rect 3818 9621 3830 9677
rect 3886 9621 3888 9677
rect 3818 9619 3888 9621
rect 4100 9677 4160 9681
rect 4100 9621 4102 9677
rect 4158 9621 4160 9677
rect 3830 9007 3886 9619
rect 4100 9609 4160 9621
rect 7298 9514 7354 10393
rect 7298 9404 7354 9414
rect 3682 4509 3752 4521
rect 3682 4453 3694 4509
rect 3750 4453 3752 4509
rect 3682 4441 3752 4453
rect 3328 3151 3330 3207
rect 3386 3151 3614 3207
rect 2740 3091 2820 3093
rect 2740 3035 2752 3091
rect 2808 3035 2820 3091
rect 2740 3033 2820 3035
rect 2752 2951 2808 3033
rect 2372 2941 2452 2951
rect 2372 2885 2384 2941
rect 2440 2885 2452 2941
rect 2372 2875 2452 2885
rect 2556 2941 2636 2951
rect 2556 2885 2568 2941
rect 2624 2885 2636 2941
rect 2556 2875 2636 2885
rect 2740 2941 2820 2951
rect 2740 2885 2752 2941
rect 2808 2885 2820 2941
rect 2740 2875 2820 2885
rect 2885 2819 2953 3149
rect 3328 3139 3398 3151
rect 2844 2811 2953 2819
rect 2832 2809 2953 2811
rect 2832 2689 2844 2809
rect 2900 2689 2953 2809
rect 2832 2687 2953 2689
rect 2844 2679 2900 2687
rect 2147 2422 3043 2434
rect 2147 2366 2159 2422
rect 2215 2366 2977 2422
rect 3033 2366 3043 2422
rect 2147 2354 3043 2366
rect 1832 2303 1912 2313
rect 1832 2247 1844 2303
rect 1900 2247 1912 2303
rect 1832 2245 1912 2247
rect 1666 2193 1736 2196
rect 1666 2139 1668 2193
rect 1724 2139 1736 2193
rect 1666 2127 1736 2139
rect 806 2086 1552 2098
rect 806 2030 1174 2086
rect 1230 2030 1552 2086
rect 806 2018 1552 2030
rect 806 1765 862 2018
rect 1174 1765 1230 2018
rect 1496 1765 1552 2018
rect 794 1763 874 1765
rect 794 1643 806 1763
rect 862 1643 874 1763
rect 794 1641 874 1643
rect 1162 1763 1242 1765
rect 1162 1643 1174 1763
rect 1230 1643 1242 1763
rect 1162 1641 1242 1643
rect 1484 1763 1564 1765
rect 1484 1642 1496 1763
rect 1552 1642 1564 1763
rect 806 1633 862 1641
rect 1174 1633 1230 1641
rect 1484 1640 1564 1642
rect 1496 1632 1552 1640
rect 990 1465 1046 1473
rect 1358 1465 1414 1473
rect 978 1463 1467 1465
rect 978 1343 990 1463
rect 1046 1343 1358 1463
rect 1414 1343 1467 1463
rect 978 1341 1467 1343
rect 990 1333 1046 1341
rect 1358 1333 1467 1341
rect 886 1267 966 1277
rect 886 1211 898 1267
rect 954 1211 966 1267
rect 886 1201 966 1211
rect 1070 1267 1150 1277
rect 1070 1211 1082 1267
rect 1138 1211 1150 1267
rect 1070 1201 1150 1211
rect 1254 1267 1334 1277
rect 1254 1211 1266 1267
rect 1322 1211 1334 1267
rect 1254 1201 1334 1211
rect 898 1119 954 1201
rect 886 1117 966 1119
rect 886 1061 898 1117
rect 954 1061 966 1117
rect 886 1059 966 1061
rect 78 1001 148 1015
rect 78 945 90 1001
rect 146 945 148 1001
rect 78 933 148 945
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect -121 98 -35 110
rect 90 102 146 933
rect 898 745 954 1059
rect 1082 1003 1138 1201
rect 1070 1001 1150 1003
rect 1070 945 1082 1001
rect 1138 945 1150 1001
rect 1070 943 1150 945
rect 1082 745 1138 943
rect 1266 887 1322 1201
rect 1399 1003 1467 1333
rect 1844 1013 1900 2245
rect 1399 1001 1479 1003
rect 1399 945 1411 1001
rect 1467 945 1479 1001
rect 1399 943 1479 945
rect 1842 1001 1902 1013
rect 1842 945 1844 1001
rect 1900 945 1902 1001
rect 1254 885 1334 887
rect 1254 829 1266 885
rect 1322 829 1334 885
rect 1254 827 1334 829
rect 1266 745 1322 827
rect 886 735 966 745
rect 886 679 898 735
rect 954 679 966 735
rect 886 669 966 679
rect 1070 735 1150 745
rect 1070 679 1082 735
rect 1138 679 1150 735
rect 1070 669 1150 679
rect 1254 735 1334 745
rect 1254 679 1266 735
rect 1322 679 1334 735
rect 1254 669 1334 679
rect 1399 613 1467 943
rect 1842 933 1902 945
rect 1358 605 1467 613
rect 1346 603 1467 605
rect 1346 483 1358 603
rect 1414 483 1467 603
rect 1346 481 1467 483
rect 1358 473 1414 481
rect 661 216 1559 228
rect 661 160 673 216
rect 729 160 1491 216
rect 1547 160 1559 216
rect 661 148 1559 160
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect 88 98 148 102
rect 88 42 90 98
rect 146 42 148 98
rect 88 30 148 42
rect -473 -65 -262 -55
rect -473 -165 -318 -65
rect -473 -175 -262 -165
rect 3694 -65 3750 4441
rect 3830 110 3886 8907
rect 4818 8701 5564 8713
rect 4818 8645 5186 8701
rect 5242 8645 5564 8701
rect 4818 8633 5564 8645
rect 4818 8380 4874 8633
rect 5186 8380 5242 8633
rect 5508 8380 5564 8633
rect 4806 8378 4886 8380
rect 4806 8258 4818 8378
rect 4874 8258 4886 8378
rect 4806 8256 4886 8258
rect 5174 8378 5254 8380
rect 5174 8258 5186 8378
rect 5242 8258 5254 8378
rect 5174 8256 5254 8258
rect 5496 8378 5576 8380
rect 5496 8257 5508 8378
rect 5564 8257 5576 8378
rect 4818 8248 4874 8256
rect 5186 8248 5242 8256
rect 5496 8255 5576 8257
rect 5508 8247 5564 8255
rect 5002 8080 5058 8088
rect 5370 8080 5426 8088
rect 4990 8078 5479 8080
rect 4990 7958 5002 8078
rect 5058 7958 5370 8078
rect 5426 7958 5479 8078
rect 4990 7956 5479 7958
rect 5002 7948 5058 7956
rect 5370 7948 5479 7956
rect 4898 7882 4978 7892
rect 4898 7826 4910 7882
rect 4966 7826 4978 7882
rect 4898 7816 4978 7826
rect 5082 7882 5162 7892
rect 5082 7826 5094 7882
rect 5150 7826 5162 7882
rect 5082 7816 5162 7826
rect 5266 7882 5346 7892
rect 5266 7826 5278 7882
rect 5334 7826 5346 7882
rect 5266 7816 5346 7826
rect 4010 7732 4096 7744
rect 4910 7734 4966 7816
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 4898 7732 4978 7734
rect 4898 7676 4910 7732
rect 4966 7676 4978 7732
rect 4898 7674 4978 7676
rect 4226 7616 4296 7628
rect 4226 7560 4238 7616
rect 4294 7560 4296 7616
rect 4226 7548 4296 7560
rect 4090 5411 4160 5425
rect 4090 5355 4102 5411
rect 4158 5355 4160 5411
rect 4090 5343 4160 5355
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 3966 897 4022 5165
rect 4102 1015 4158 5343
rect 4238 3102 4294 7548
rect 4910 7360 4966 7674
rect 5094 7618 5150 7816
rect 5082 7616 5162 7618
rect 5082 7560 5094 7616
rect 5150 7560 5162 7616
rect 5082 7558 5162 7560
rect 5094 7360 5150 7558
rect 5278 7502 5334 7816
rect 5411 7618 5479 7948
rect 5411 7616 5491 7618
rect 5411 7560 5423 7616
rect 5479 7560 5491 7616
rect 5411 7558 5491 7560
rect 5678 7616 5748 7628
rect 5678 7560 5680 7616
rect 5736 7560 5748 7616
rect 5266 7500 5346 7502
rect 5266 7444 5278 7500
rect 5334 7444 5346 7500
rect 5266 7442 5346 7444
rect 5278 7360 5334 7442
rect 4898 7350 4978 7360
rect 4898 7294 4910 7350
rect 4966 7294 4978 7350
rect 4898 7284 4978 7294
rect 5082 7350 5162 7360
rect 5082 7294 5094 7350
rect 5150 7294 5162 7350
rect 5082 7284 5162 7294
rect 5266 7350 5346 7360
rect 5266 7294 5278 7350
rect 5334 7294 5346 7350
rect 5266 7284 5346 7294
rect 5411 7228 5479 7558
rect 5678 7550 5748 7560
rect 5370 7220 5479 7228
rect 5358 7218 5479 7220
rect 5358 7098 5370 7218
rect 5426 7098 5479 7218
rect 5358 7096 5479 7098
rect 5370 7088 5426 7096
rect 4673 6831 5571 6843
rect 4673 6775 4685 6831
rect 4741 6775 5503 6831
rect 5559 6775 5571 6831
rect 4673 6763 5571 6775
rect 5680 6606 5736 7550
rect 5844 6713 5924 6723
rect 5844 6657 5856 6713
rect 5912 6657 5924 6713
rect 5844 6655 5924 6657
rect 5678 6603 5748 6606
rect 5678 6549 5680 6603
rect 5736 6549 5748 6603
rect 5678 6537 5748 6549
rect 4818 6496 5564 6508
rect 4818 6440 5186 6496
rect 5242 6440 5564 6496
rect 4818 6428 5564 6440
rect 4818 6175 4874 6428
rect 5186 6175 5242 6428
rect 5508 6175 5564 6428
rect 4806 6173 4886 6175
rect 4806 6053 4818 6173
rect 4874 6053 4886 6173
rect 4806 6051 4886 6053
rect 5174 6173 5254 6175
rect 5174 6053 5186 6173
rect 5242 6053 5254 6173
rect 5174 6051 5254 6053
rect 5496 6173 5576 6175
rect 5496 6052 5508 6173
rect 5564 6052 5576 6173
rect 4818 6043 4874 6051
rect 5186 6043 5242 6051
rect 5496 6050 5576 6052
rect 5508 6042 5564 6050
rect 5002 5875 5058 5883
rect 5370 5875 5426 5883
rect 4990 5873 5479 5875
rect 4990 5753 5002 5873
rect 5058 5753 5370 5873
rect 5426 5753 5479 5873
rect 4990 5751 5479 5753
rect 5002 5743 5058 5751
rect 5370 5743 5479 5751
rect 4898 5677 4978 5687
rect 4898 5621 4910 5677
rect 4966 5621 4978 5677
rect 4898 5611 4978 5621
rect 5082 5677 5162 5687
rect 5082 5621 5094 5677
rect 5150 5621 5162 5677
rect 5082 5611 5162 5621
rect 5266 5677 5346 5687
rect 5266 5621 5278 5677
rect 5334 5621 5346 5677
rect 5266 5611 5346 5621
rect 4910 5529 4966 5611
rect 4898 5527 4978 5529
rect 4898 5471 4910 5527
rect 4966 5471 4978 5527
rect 4898 5469 4978 5471
rect 4910 5155 4966 5469
rect 5094 5413 5150 5611
rect 5082 5411 5162 5413
rect 5082 5355 5094 5411
rect 5150 5355 5162 5411
rect 5082 5353 5162 5355
rect 5094 5155 5150 5353
rect 5278 5297 5334 5611
rect 5411 5413 5479 5743
rect 5856 5421 5912 6655
rect 6304 6496 7050 6508
rect 6304 6440 6672 6496
rect 6728 6440 7050 6496
rect 6304 6428 7050 6440
rect 6304 6175 6360 6428
rect 6672 6175 6728 6428
rect 6994 6175 7050 6428
rect 6292 6173 6372 6175
rect 6292 6053 6304 6173
rect 6360 6053 6372 6173
rect 6292 6051 6372 6053
rect 6660 6173 6740 6175
rect 6660 6053 6672 6173
rect 6728 6053 6740 6173
rect 6660 6051 6740 6053
rect 6982 6173 7062 6175
rect 6982 6052 6994 6173
rect 7050 6052 7062 6173
rect 6304 6043 6360 6051
rect 6672 6043 6728 6051
rect 6982 6050 7062 6052
rect 6994 6042 7050 6050
rect 6488 5875 6544 5883
rect 6856 5875 6912 5883
rect 6476 5873 6965 5875
rect 6476 5753 6488 5873
rect 6544 5753 6856 5873
rect 6912 5753 6965 5873
rect 6476 5751 6965 5753
rect 6488 5743 6544 5751
rect 6856 5743 6965 5751
rect 6384 5677 6464 5687
rect 6384 5621 6396 5677
rect 6452 5621 6464 5677
rect 6384 5611 6464 5621
rect 6568 5677 6648 5687
rect 6568 5621 6580 5677
rect 6636 5621 6648 5677
rect 6568 5611 6648 5621
rect 6752 5677 6832 5687
rect 6752 5621 6764 5677
rect 6820 5621 6832 5677
rect 6752 5611 6832 5621
rect 6396 5529 6452 5611
rect 6384 5527 6464 5529
rect 6384 5471 6396 5527
rect 6452 5471 6464 5527
rect 6384 5469 6464 5471
rect 5411 5411 5491 5413
rect 5411 5355 5423 5411
rect 5479 5355 5491 5411
rect 5411 5353 5491 5355
rect 5854 5411 5914 5421
rect 5854 5355 5856 5411
rect 5912 5355 5914 5411
rect 5266 5295 5346 5297
rect 5266 5239 5278 5295
rect 5334 5239 5346 5295
rect 5266 5237 5346 5239
rect 5278 5155 5334 5237
rect 4898 5145 4978 5155
rect 4898 5089 4910 5145
rect 4966 5089 4978 5145
rect 4898 5079 4978 5089
rect 5082 5145 5162 5155
rect 5082 5089 5094 5145
rect 5150 5089 5162 5145
rect 5082 5079 5162 5089
rect 5266 5145 5346 5155
rect 5266 5089 5278 5145
rect 5334 5089 5346 5145
rect 5266 5079 5346 5089
rect 5411 5023 5479 5353
rect 5854 5343 5914 5355
rect 5370 5015 5479 5023
rect 5358 5013 5479 5015
rect 5358 4893 5370 5013
rect 5426 4893 5479 5013
rect 5358 4891 5479 4893
rect 5370 4883 5426 4891
rect 4673 4626 5569 4638
rect 4673 4570 4685 4626
rect 4741 4570 5503 4626
rect 5559 4570 5569 4626
rect 4673 4558 5569 4570
rect 5856 4400 5912 5343
rect 6396 5155 6452 5469
rect 6580 5413 6636 5611
rect 6568 5411 6648 5413
rect 6568 5355 6580 5411
rect 6636 5355 6648 5411
rect 6568 5353 6648 5355
rect 6580 5155 6636 5353
rect 6764 5297 6820 5611
rect 6897 5413 6965 5743
rect 6897 5411 6977 5413
rect 6897 5355 6909 5411
rect 6965 5355 6977 5411
rect 6897 5353 6977 5355
rect 7164 5411 7234 5423
rect 7164 5355 7166 5411
rect 7222 5355 7490 5411
rect 6752 5295 6832 5297
rect 6752 5239 6764 5295
rect 6820 5239 6832 5295
rect 6752 5237 6832 5239
rect 6764 5155 6820 5237
rect 6384 5145 6464 5155
rect 6384 5089 6396 5145
rect 6452 5089 6464 5145
rect 6384 5079 6464 5089
rect 6568 5145 6648 5155
rect 6568 5089 6580 5145
rect 6636 5089 6648 5145
rect 6568 5079 6648 5089
rect 6752 5145 6832 5155
rect 6752 5089 6764 5145
rect 6820 5089 6832 5145
rect 6752 5079 6832 5089
rect 6897 5023 6965 5353
rect 7164 5345 7234 5355
rect 6856 5015 6965 5023
rect 6844 5013 6965 5015
rect 6844 4893 6856 5013
rect 6912 4893 6965 5013
rect 6844 4891 6965 4893
rect 6856 4883 6912 4891
rect 6159 4626 7055 4638
rect 6159 4570 6171 4626
rect 6227 4570 6989 4626
rect 7045 4570 7055 4626
rect 6159 4558 7055 4570
rect 7166 4401 7222 5345
rect 7330 4509 7410 4519
rect 7330 4453 7342 4509
rect 7398 4453 7410 4509
rect 7330 4451 7410 4453
rect 5854 4398 5924 4400
rect 5854 4342 5856 4398
rect 5912 4342 5924 4398
rect 5854 4330 5924 4342
rect 7154 4399 7234 4401
rect 7154 4343 7166 4399
rect 7222 4343 7234 4399
rect 7154 4331 7234 4343
rect 4818 4291 5564 4303
rect 4818 4235 5186 4291
rect 5242 4235 5564 4291
rect 4818 4223 5564 4235
rect 4818 3970 4874 4223
rect 5186 3970 5242 4223
rect 5508 3970 5564 4223
rect 6304 4292 7050 4304
rect 6304 4236 6672 4292
rect 6728 4236 7050 4292
rect 6304 4224 7050 4236
rect 6304 3971 6360 4224
rect 6672 3971 6728 4224
rect 6994 3971 7050 4224
rect 4806 3968 4886 3970
rect 4806 3848 4818 3968
rect 4874 3848 4886 3968
rect 4806 3846 4886 3848
rect 5174 3968 5254 3970
rect 5174 3848 5186 3968
rect 5242 3848 5254 3968
rect 5174 3846 5254 3848
rect 5496 3968 5576 3970
rect 5496 3847 5508 3968
rect 5564 3847 5576 3968
rect 6292 3969 6372 3971
rect 6292 3849 6304 3969
rect 6360 3849 6372 3969
rect 6292 3847 6372 3849
rect 6660 3969 6740 3971
rect 6660 3849 6672 3969
rect 6728 3849 6740 3969
rect 6660 3847 6740 3849
rect 6982 3969 7062 3971
rect 6982 3848 6994 3969
rect 7050 3848 7062 3969
rect 4818 3838 4874 3846
rect 5186 3838 5242 3846
rect 5496 3845 5576 3847
rect 5508 3837 5564 3845
rect 6304 3839 6360 3847
rect 6672 3839 6728 3847
rect 6982 3846 7062 3848
rect 6994 3838 7050 3846
rect 5002 3670 5058 3678
rect 5370 3670 5426 3678
rect 6488 3671 6544 3679
rect 6856 3671 6912 3679
rect 4990 3668 5479 3670
rect 4990 3548 5002 3668
rect 5058 3548 5370 3668
rect 5426 3548 5479 3668
rect 4990 3546 5479 3548
rect 6476 3669 6965 3671
rect 6476 3549 6488 3669
rect 6544 3549 6856 3669
rect 6912 3549 6965 3669
rect 6476 3547 6965 3549
rect 5002 3538 5058 3546
rect 5370 3538 5479 3546
rect 6488 3539 6544 3547
rect 6856 3539 6965 3547
rect 4898 3472 4978 3482
rect 4898 3416 4910 3472
rect 4966 3416 4978 3472
rect 4898 3406 4978 3416
rect 5082 3472 5162 3482
rect 5082 3416 5094 3472
rect 5150 3416 5162 3472
rect 5082 3406 5162 3416
rect 5266 3472 5346 3482
rect 5266 3416 5278 3472
rect 5334 3416 5346 3472
rect 5266 3406 5346 3416
rect 4910 3324 4966 3406
rect 4898 3322 4978 3324
rect 4898 3266 4910 3322
rect 4966 3266 4978 3322
rect 4898 3264 4978 3266
rect 4226 3090 4296 3102
rect 4226 3034 4238 3090
rect 4294 3034 4296 3090
rect 4226 3022 4296 3034
rect 4910 2950 4966 3264
rect 5094 3208 5150 3406
rect 5082 3206 5162 3208
rect 5082 3150 5094 3206
rect 5150 3150 5162 3206
rect 5082 3148 5162 3150
rect 5094 2950 5150 3148
rect 5278 3092 5334 3406
rect 5411 3208 5479 3538
rect 6384 3473 6464 3483
rect 6384 3417 6396 3473
rect 6452 3417 6464 3473
rect 6384 3407 6464 3417
rect 6568 3473 6648 3483
rect 6568 3417 6580 3473
rect 6636 3417 6648 3473
rect 6568 3407 6648 3417
rect 6752 3473 6832 3483
rect 6752 3417 6764 3473
rect 6820 3417 6832 3473
rect 6752 3407 6832 3417
rect 6396 3325 6452 3407
rect 6384 3323 6464 3325
rect 6384 3267 6396 3323
rect 6452 3267 6464 3323
rect 6384 3265 6464 3267
rect 5411 3206 5491 3208
rect 5411 3150 5423 3206
rect 5479 3150 5491 3206
rect 5411 3148 5491 3150
rect 5678 3206 5748 3218
rect 5678 3150 5680 3206
rect 5736 3150 5748 3206
rect 5266 3090 5346 3092
rect 5266 3034 5278 3090
rect 5334 3034 5346 3090
rect 5266 3032 5346 3034
rect 5278 2950 5334 3032
rect 4898 2940 4978 2950
rect 4898 2884 4910 2940
rect 4966 2884 4978 2940
rect 4898 2874 4978 2884
rect 5082 2940 5162 2950
rect 5082 2884 5094 2940
rect 5150 2884 5162 2940
rect 5082 2874 5162 2884
rect 5266 2940 5346 2950
rect 5266 2884 5278 2940
rect 5334 2884 5346 2940
rect 5266 2874 5346 2884
rect 5411 2818 5479 3148
rect 5678 3140 5748 3150
rect 5370 2810 5479 2818
rect 5358 2808 5479 2810
rect 5358 2688 5370 2808
rect 5426 2688 5479 2808
rect 5358 2686 5479 2688
rect 5370 2678 5426 2686
rect 4673 2421 5569 2433
rect 4673 2365 4685 2421
rect 4741 2365 5503 2421
rect 5559 2365 5569 2421
rect 4673 2353 5569 2365
rect 5680 2196 5736 3140
rect 6396 2951 6452 3265
rect 6580 3209 6636 3407
rect 6568 3207 6648 3209
rect 6568 3151 6580 3207
rect 6636 3151 6648 3207
rect 6568 3149 6648 3151
rect 6580 2951 6636 3149
rect 6764 3093 6820 3407
rect 6897 3209 6965 3539
rect 7342 3217 7398 4451
rect 6897 3207 6977 3209
rect 6897 3151 6909 3207
rect 6965 3151 6977 3207
rect 6897 3149 6977 3151
rect 7340 3207 7410 3217
rect 7570 3207 7626 17250
rect 7706 14992 7762 19504
rect 11760 18739 11816 19501
rect 12038 19089 12108 19101
rect 12038 19033 12050 19089
rect 12106 19033 12108 19089
rect 12038 19031 12108 19033
rect 11758 18737 11828 18739
rect 11758 18681 11760 18737
rect 11816 18681 11828 18737
rect 11758 18679 11828 18681
rect 7996 18561 8066 18573
rect 7996 18505 8008 18561
rect 8064 18505 8066 18561
rect 7996 18503 8066 18505
rect 7704 14990 7774 14992
rect 7704 14934 7706 14990
rect 7762 14934 7774 14990
rect 7704 14922 7774 14934
rect 8008 14087 8064 18503
rect 8860 18277 9606 18289
rect 8860 18221 9228 18277
rect 9284 18221 9606 18277
rect 8860 18209 9606 18221
rect 8860 17956 8916 18209
rect 9228 17956 9284 18209
rect 9550 17956 9606 18209
rect 8848 17954 8928 17956
rect 8848 17834 8860 17954
rect 8916 17834 8928 17954
rect 8848 17832 8928 17834
rect 9216 17954 9296 17956
rect 9216 17834 9228 17954
rect 9284 17834 9296 17954
rect 9216 17832 9296 17834
rect 9538 17954 9618 17956
rect 9538 17833 9550 17954
rect 9606 17833 9618 17954
rect 8860 17824 8916 17832
rect 9228 17824 9284 17832
rect 9538 17831 9618 17833
rect 9550 17823 9606 17831
rect 9044 17656 9100 17664
rect 9412 17656 9468 17664
rect 9032 17654 9521 17656
rect 9032 17534 9044 17654
rect 9100 17534 9412 17654
rect 9468 17534 9521 17654
rect 9032 17532 9521 17534
rect 9044 17524 9100 17532
rect 9412 17524 9521 17532
rect 8940 17458 9020 17468
rect 8940 17402 8952 17458
rect 9008 17402 9020 17458
rect 8940 17392 9020 17402
rect 9124 17458 9204 17468
rect 9124 17402 9136 17458
rect 9192 17402 9204 17458
rect 9124 17392 9204 17402
rect 9308 17458 9388 17468
rect 9308 17402 9320 17458
rect 9376 17402 9388 17458
rect 9308 17392 9388 17402
rect 8952 17310 9008 17392
rect 8940 17308 9020 17310
rect 8940 17252 8952 17308
rect 9008 17252 9020 17308
rect 8940 17250 9020 17252
rect 8268 17192 8338 17204
rect 8268 17136 8280 17192
rect 8336 17136 8338 17192
rect 8268 17124 8338 17136
rect 8132 14987 8202 15001
rect 8132 14931 8144 14987
rect 8200 14931 8202 14987
rect 8132 14919 8202 14931
rect 7996 14085 8066 14087
rect 7996 14029 8008 14085
rect 8064 14029 8066 14085
rect 7996 14017 8066 14029
rect 8144 10591 8200 14919
rect 8280 12678 8336 17124
rect 8952 16936 9008 17250
rect 9136 17194 9192 17392
rect 9124 17192 9204 17194
rect 9124 17136 9136 17192
rect 9192 17136 9204 17192
rect 9124 17134 9204 17136
rect 9136 16936 9192 17134
rect 9320 17078 9376 17392
rect 9453 17194 9521 17524
rect 11600 17308 11670 17320
rect 11600 17252 11612 17308
rect 11668 17252 11670 17308
rect 11600 17250 11670 17252
rect 9453 17192 9533 17194
rect 9453 17136 9465 17192
rect 9521 17136 9533 17192
rect 9453 17134 9533 17136
rect 9720 17192 9790 17204
rect 9720 17136 9722 17192
rect 9778 17136 9790 17192
rect 9308 17076 9388 17078
rect 9308 17020 9320 17076
rect 9376 17020 9388 17076
rect 9308 17018 9388 17020
rect 9320 16936 9376 17018
rect 8940 16926 9020 16936
rect 8940 16870 8952 16926
rect 9008 16870 9020 16926
rect 8940 16860 9020 16870
rect 9124 16926 9204 16936
rect 9124 16870 9136 16926
rect 9192 16870 9204 16926
rect 9124 16860 9204 16870
rect 9308 16926 9388 16936
rect 9308 16870 9320 16926
rect 9376 16870 9388 16926
rect 9308 16860 9388 16870
rect 9453 16804 9521 17134
rect 9720 17126 9790 17136
rect 9412 16796 9521 16804
rect 9400 16794 9521 16796
rect 9400 16674 9412 16794
rect 9468 16674 9521 16794
rect 9400 16672 9521 16674
rect 9412 16664 9468 16672
rect 8715 16407 9613 16419
rect 8715 16351 8727 16407
rect 8783 16351 9545 16407
rect 9601 16351 9613 16407
rect 8715 16339 9613 16351
rect 9722 16182 9778 17126
rect 9886 16289 9966 16299
rect 9886 16233 9898 16289
rect 9954 16233 9966 16289
rect 9886 16231 9966 16233
rect 9720 16179 9790 16182
rect 9720 16125 9722 16179
rect 9778 16125 9790 16179
rect 9720 16113 9790 16125
rect 8860 16072 9606 16084
rect 8860 16016 9228 16072
rect 9284 16016 9606 16072
rect 8860 16004 9606 16016
rect 8860 15751 8916 16004
rect 9228 15751 9284 16004
rect 9550 15751 9606 16004
rect 8848 15749 8928 15751
rect 8848 15629 8860 15749
rect 8916 15629 8928 15749
rect 8848 15627 8928 15629
rect 9216 15749 9296 15751
rect 9216 15629 9228 15749
rect 9284 15629 9296 15749
rect 9216 15627 9296 15629
rect 9538 15749 9618 15751
rect 9538 15628 9550 15749
rect 9606 15628 9618 15749
rect 8860 15619 8916 15627
rect 9228 15619 9284 15627
rect 9538 15626 9618 15628
rect 9550 15618 9606 15626
rect 9044 15451 9100 15459
rect 9412 15451 9468 15459
rect 9032 15449 9521 15451
rect 9032 15329 9044 15449
rect 9100 15329 9412 15449
rect 9468 15329 9521 15449
rect 9032 15327 9521 15329
rect 9044 15319 9100 15327
rect 9412 15319 9521 15327
rect 8940 15253 9020 15263
rect 8940 15197 8952 15253
rect 9008 15197 9020 15253
rect 8940 15187 9020 15197
rect 9124 15253 9204 15263
rect 9124 15197 9136 15253
rect 9192 15197 9204 15253
rect 9124 15187 9204 15197
rect 9308 15253 9388 15263
rect 9308 15197 9320 15253
rect 9376 15197 9388 15253
rect 9308 15187 9388 15197
rect 8952 15105 9008 15187
rect 8940 15103 9020 15105
rect 8940 15047 8952 15103
rect 9008 15047 9020 15103
rect 8940 15045 9020 15047
rect 8952 14731 9008 15045
rect 9136 14989 9192 15187
rect 9124 14987 9204 14989
rect 9124 14931 9136 14987
rect 9192 14931 9204 14987
rect 9124 14929 9204 14931
rect 9136 14731 9192 14929
rect 9320 14873 9376 15187
rect 9453 14989 9521 15319
rect 9898 14997 9954 16231
rect 10346 16072 11092 16084
rect 10346 16016 10714 16072
rect 10770 16016 11092 16072
rect 10346 16004 11092 16016
rect 10346 15751 10402 16004
rect 10714 15751 10770 16004
rect 11036 15751 11092 16004
rect 10334 15749 10414 15751
rect 10334 15629 10346 15749
rect 10402 15629 10414 15749
rect 10334 15627 10414 15629
rect 10702 15749 10782 15751
rect 10702 15629 10714 15749
rect 10770 15629 10782 15749
rect 10702 15627 10782 15629
rect 11024 15749 11104 15751
rect 11024 15628 11036 15749
rect 11092 15628 11104 15749
rect 10346 15619 10402 15627
rect 10714 15619 10770 15627
rect 11024 15626 11104 15628
rect 11036 15618 11092 15626
rect 10530 15451 10586 15459
rect 10898 15451 10954 15459
rect 10518 15449 11007 15451
rect 10518 15329 10530 15449
rect 10586 15329 10898 15449
rect 10954 15329 11007 15449
rect 10518 15327 11007 15329
rect 10530 15319 10586 15327
rect 10898 15319 11007 15327
rect 10426 15253 10506 15263
rect 10426 15197 10438 15253
rect 10494 15197 10506 15253
rect 10426 15187 10506 15197
rect 10610 15253 10690 15263
rect 10610 15197 10622 15253
rect 10678 15197 10690 15253
rect 10610 15187 10690 15197
rect 10794 15253 10874 15263
rect 10794 15197 10806 15253
rect 10862 15197 10874 15253
rect 10794 15187 10874 15197
rect 10438 15105 10494 15187
rect 10426 15103 10506 15105
rect 10426 15047 10438 15103
rect 10494 15047 10506 15103
rect 10426 15045 10506 15047
rect 9453 14987 9533 14989
rect 9453 14931 9465 14987
rect 9521 14931 9533 14987
rect 9453 14929 9533 14931
rect 9896 14987 9956 14997
rect 9896 14931 9898 14987
rect 9954 14931 9956 14987
rect 9308 14871 9388 14873
rect 9308 14815 9320 14871
rect 9376 14815 9388 14871
rect 9308 14813 9388 14815
rect 9320 14731 9376 14813
rect 8940 14721 9020 14731
rect 8940 14665 8952 14721
rect 9008 14665 9020 14721
rect 8940 14655 9020 14665
rect 9124 14721 9204 14731
rect 9124 14665 9136 14721
rect 9192 14665 9204 14721
rect 9124 14655 9204 14665
rect 9308 14721 9388 14731
rect 9308 14665 9320 14721
rect 9376 14665 9388 14721
rect 9308 14655 9388 14665
rect 9453 14599 9521 14929
rect 9896 14919 9956 14931
rect 9412 14591 9521 14599
rect 9400 14589 9521 14591
rect 9400 14469 9412 14589
rect 9468 14469 9521 14589
rect 9400 14467 9521 14469
rect 9412 14459 9468 14467
rect 8715 14202 9611 14214
rect 8715 14146 8727 14202
rect 8783 14146 9545 14202
rect 9601 14146 9611 14202
rect 8715 14134 9611 14146
rect 9898 13976 9954 14919
rect 10438 14731 10494 15045
rect 10622 14989 10678 15187
rect 10610 14987 10690 14989
rect 10610 14931 10622 14987
rect 10678 14931 10690 14987
rect 10610 14929 10690 14931
rect 10622 14731 10678 14929
rect 10806 14873 10862 15187
rect 10939 14989 11007 15319
rect 10939 14987 11019 14989
rect 10939 14931 10951 14987
rect 11007 14931 11019 14987
rect 10939 14929 11019 14931
rect 11206 14987 11276 14999
rect 11206 14931 11208 14987
rect 11264 14931 11532 14987
rect 10794 14871 10874 14873
rect 10794 14815 10806 14871
rect 10862 14815 10874 14871
rect 10794 14813 10874 14815
rect 10806 14731 10862 14813
rect 10426 14721 10506 14731
rect 10426 14665 10438 14721
rect 10494 14665 10506 14721
rect 10426 14655 10506 14665
rect 10610 14721 10690 14731
rect 10610 14665 10622 14721
rect 10678 14665 10690 14721
rect 10610 14655 10690 14665
rect 10794 14721 10874 14731
rect 10794 14665 10806 14721
rect 10862 14665 10874 14721
rect 10794 14655 10874 14665
rect 10939 14599 11007 14929
rect 11206 14921 11276 14931
rect 10898 14591 11007 14599
rect 10886 14589 11007 14591
rect 10886 14469 10898 14589
rect 10954 14469 11007 14589
rect 10886 14467 11007 14469
rect 10898 14459 10954 14467
rect 10201 14202 11097 14214
rect 10201 14146 10213 14202
rect 10269 14146 11031 14202
rect 11087 14146 11097 14202
rect 10201 14134 11097 14146
rect 11208 13977 11264 14921
rect 11372 14085 11452 14095
rect 11372 14029 11384 14085
rect 11440 14029 11452 14085
rect 11372 14027 11452 14029
rect 9896 13974 9966 13976
rect 9896 13918 9898 13974
rect 9954 13918 9966 13974
rect 9896 13906 9966 13918
rect 11196 13975 11276 13977
rect 11196 13919 11208 13975
rect 11264 13919 11276 13975
rect 11196 13907 11276 13919
rect 8860 13867 9606 13879
rect 8860 13811 9228 13867
rect 9284 13811 9606 13867
rect 8860 13799 9606 13811
rect 8860 13546 8916 13799
rect 9228 13546 9284 13799
rect 9550 13546 9606 13799
rect 10346 13868 11092 13880
rect 10346 13812 10714 13868
rect 10770 13812 11092 13868
rect 10346 13800 11092 13812
rect 10346 13547 10402 13800
rect 10714 13547 10770 13800
rect 11036 13547 11092 13800
rect 8848 13544 8928 13546
rect 8848 13424 8860 13544
rect 8916 13424 8928 13544
rect 8848 13422 8928 13424
rect 9216 13544 9296 13546
rect 9216 13424 9228 13544
rect 9284 13424 9296 13544
rect 9216 13422 9296 13424
rect 9538 13544 9618 13546
rect 9538 13423 9550 13544
rect 9606 13423 9618 13544
rect 10334 13545 10414 13547
rect 10334 13425 10346 13545
rect 10402 13425 10414 13545
rect 10334 13423 10414 13425
rect 10702 13545 10782 13547
rect 10702 13425 10714 13545
rect 10770 13425 10782 13545
rect 10702 13423 10782 13425
rect 11024 13545 11104 13547
rect 11024 13424 11036 13545
rect 11092 13424 11104 13545
rect 8860 13414 8916 13422
rect 9228 13414 9284 13422
rect 9538 13421 9618 13423
rect 9550 13413 9606 13421
rect 10346 13415 10402 13423
rect 10714 13415 10770 13423
rect 11024 13422 11104 13424
rect 11036 13414 11092 13422
rect 9044 13246 9100 13254
rect 9412 13246 9468 13254
rect 10530 13247 10586 13255
rect 10898 13247 10954 13255
rect 9032 13244 9521 13246
rect 9032 13124 9044 13244
rect 9100 13124 9412 13244
rect 9468 13124 9521 13244
rect 9032 13122 9521 13124
rect 10518 13245 11007 13247
rect 10518 13125 10530 13245
rect 10586 13125 10898 13245
rect 10954 13125 11007 13245
rect 10518 13123 11007 13125
rect 9044 13114 9100 13122
rect 9412 13114 9521 13122
rect 10530 13115 10586 13123
rect 10898 13115 11007 13123
rect 8940 13048 9020 13058
rect 8940 12992 8952 13048
rect 9008 12992 9020 13048
rect 8940 12982 9020 12992
rect 9124 13048 9204 13058
rect 9124 12992 9136 13048
rect 9192 12992 9204 13048
rect 9124 12982 9204 12992
rect 9308 13048 9388 13058
rect 9308 12992 9320 13048
rect 9376 12992 9388 13048
rect 9308 12982 9388 12992
rect 8952 12900 9008 12982
rect 8940 12898 9020 12900
rect 8940 12842 8952 12898
rect 9008 12842 9020 12898
rect 8940 12840 9020 12842
rect 8268 12666 8338 12678
rect 8268 12610 8280 12666
rect 8336 12610 8338 12666
rect 8268 12598 8338 12610
rect 8952 12526 9008 12840
rect 9136 12784 9192 12982
rect 9124 12782 9204 12784
rect 9124 12726 9136 12782
rect 9192 12726 9204 12782
rect 9124 12724 9204 12726
rect 9136 12526 9192 12724
rect 9320 12668 9376 12982
rect 9453 12784 9521 13114
rect 10426 13049 10506 13059
rect 10426 12993 10438 13049
rect 10494 12993 10506 13049
rect 10426 12983 10506 12993
rect 10610 13049 10690 13059
rect 10610 12993 10622 13049
rect 10678 12993 10690 13049
rect 10610 12983 10690 12993
rect 10794 13049 10874 13059
rect 10794 12993 10806 13049
rect 10862 12993 10874 13049
rect 10794 12983 10874 12993
rect 10438 12901 10494 12983
rect 10426 12899 10506 12901
rect 10426 12843 10438 12899
rect 10494 12843 10506 12899
rect 10426 12841 10506 12843
rect 9453 12782 9533 12784
rect 9453 12726 9465 12782
rect 9521 12726 9533 12782
rect 9453 12724 9533 12726
rect 9720 12782 9790 12794
rect 9720 12726 9722 12782
rect 9778 12726 9790 12782
rect 9308 12666 9388 12668
rect 9308 12610 9320 12666
rect 9376 12610 9388 12666
rect 9308 12608 9388 12610
rect 9320 12526 9376 12608
rect 8940 12516 9020 12526
rect 8940 12460 8952 12516
rect 9008 12460 9020 12516
rect 8940 12450 9020 12460
rect 9124 12516 9204 12526
rect 9124 12460 9136 12516
rect 9192 12460 9204 12516
rect 9124 12450 9204 12460
rect 9308 12516 9388 12526
rect 9308 12460 9320 12516
rect 9376 12460 9388 12516
rect 9308 12450 9388 12460
rect 9453 12394 9521 12724
rect 9720 12716 9790 12726
rect 9412 12386 9521 12394
rect 9400 12384 9521 12386
rect 9400 12264 9412 12384
rect 9468 12264 9521 12384
rect 9400 12262 9521 12264
rect 9412 12254 9468 12262
rect 8715 11997 9611 12009
rect 8715 11941 8727 11997
rect 8783 11941 9545 11997
rect 9601 11941 9611 11997
rect 8715 11929 9611 11941
rect 9722 11772 9778 12716
rect 10438 12527 10494 12841
rect 10622 12785 10678 12983
rect 10610 12783 10690 12785
rect 10610 12727 10622 12783
rect 10678 12727 10690 12783
rect 10610 12725 10690 12727
rect 10622 12527 10678 12725
rect 10806 12669 10862 12983
rect 10939 12785 11007 13115
rect 11384 12793 11440 14027
rect 10939 12783 11019 12785
rect 10939 12727 10951 12783
rect 11007 12727 11019 12783
rect 10939 12725 11019 12727
rect 11382 12783 11452 12793
rect 11382 12727 11384 12783
rect 11440 12727 11532 12783
rect 10794 12667 10874 12669
rect 10794 12611 10806 12667
rect 10862 12611 10874 12667
rect 10794 12609 10874 12611
rect 10806 12527 10862 12609
rect 10426 12517 10506 12527
rect 10426 12461 10438 12517
rect 10494 12461 10506 12517
rect 10426 12451 10506 12461
rect 10610 12517 10690 12527
rect 10610 12461 10622 12517
rect 10678 12461 10690 12517
rect 10610 12451 10690 12461
rect 10794 12517 10874 12527
rect 10794 12461 10806 12517
rect 10862 12461 10874 12517
rect 10794 12451 10874 12461
rect 10939 12395 11007 12725
rect 11382 12715 11452 12727
rect 10898 12387 11007 12395
rect 10886 12385 11007 12387
rect 10886 12265 10898 12385
rect 10954 12265 11007 12385
rect 10886 12263 11007 12265
rect 10898 12255 10954 12263
rect 10201 11998 11097 12010
rect 10201 11942 10213 11998
rect 10269 11942 11031 11998
rect 11087 11942 11097 11998
rect 10201 11930 11097 11942
rect 9886 11879 9966 11889
rect 9886 11823 9898 11879
rect 9954 11823 9966 11879
rect 9886 11821 9966 11823
rect 9720 11769 9790 11772
rect 9720 11715 9722 11769
rect 9778 11715 9790 11769
rect 9720 11703 9790 11715
rect 8860 11662 9606 11674
rect 8860 11606 9228 11662
rect 9284 11606 9606 11662
rect 8860 11594 9606 11606
rect 8860 11341 8916 11594
rect 9228 11341 9284 11594
rect 9550 11341 9606 11594
rect 8848 11339 8928 11341
rect 8848 11219 8860 11339
rect 8916 11219 8928 11339
rect 8848 11217 8928 11219
rect 9216 11339 9296 11341
rect 9216 11219 9228 11339
rect 9284 11219 9296 11339
rect 9216 11217 9296 11219
rect 9538 11339 9618 11341
rect 9538 11218 9550 11339
rect 9606 11218 9618 11339
rect 8860 11209 8916 11217
rect 9228 11209 9284 11217
rect 9538 11216 9618 11218
rect 9550 11208 9606 11216
rect 9044 11041 9100 11049
rect 9412 11041 9468 11049
rect 9032 11039 9521 11041
rect 9032 10919 9044 11039
rect 9100 10919 9412 11039
rect 9468 10919 9521 11039
rect 9032 10917 9521 10919
rect 9044 10909 9100 10917
rect 9412 10909 9521 10917
rect 8940 10843 9020 10853
rect 8940 10787 8952 10843
rect 9008 10787 9020 10843
rect 8940 10777 9020 10787
rect 9124 10843 9204 10853
rect 9124 10787 9136 10843
rect 9192 10787 9204 10843
rect 9124 10777 9204 10787
rect 9308 10843 9388 10853
rect 9308 10787 9320 10843
rect 9376 10787 9388 10843
rect 9308 10777 9388 10787
rect 8952 10695 9008 10777
rect 8940 10693 9020 10695
rect 8940 10637 8952 10693
rect 9008 10637 9020 10693
rect 8940 10635 9020 10637
rect 8132 10577 8202 10591
rect 8132 10521 8144 10577
rect 8200 10521 8202 10577
rect 8132 10509 8202 10521
rect 7830 9674 7900 9686
rect 8144 9678 8200 10509
rect 8952 10321 9008 10635
rect 9136 10579 9192 10777
rect 9124 10577 9204 10579
rect 9124 10521 9136 10577
rect 9192 10521 9204 10577
rect 9124 10519 9204 10521
rect 9136 10321 9192 10519
rect 9320 10463 9376 10777
rect 9453 10579 9521 10909
rect 9898 10589 9954 11821
rect 9453 10577 9533 10579
rect 9453 10521 9465 10577
rect 9521 10521 9533 10577
rect 9453 10519 9533 10521
rect 9896 10577 9956 10589
rect 9896 10521 9898 10577
rect 9954 10521 9956 10577
rect 9308 10461 9388 10463
rect 9308 10405 9320 10461
rect 9376 10405 9388 10461
rect 9308 10403 9388 10405
rect 9320 10321 9376 10403
rect 8940 10311 9020 10321
rect 8940 10255 8952 10311
rect 9008 10255 9020 10311
rect 8940 10245 9020 10255
rect 9124 10311 9204 10321
rect 9124 10255 9136 10311
rect 9192 10255 9204 10311
rect 9124 10245 9204 10255
rect 9308 10311 9388 10321
rect 9308 10255 9320 10311
rect 9376 10255 9388 10311
rect 9308 10245 9388 10255
rect 9453 10189 9521 10519
rect 9896 10509 9956 10521
rect 11328 10461 11398 10473
rect 11328 10405 11340 10461
rect 11396 10405 11398 10461
rect 11328 10393 11398 10405
rect 9412 10181 9521 10189
rect 9400 10179 9521 10181
rect 9400 10059 9412 10179
rect 9468 10059 9521 10179
rect 9400 10057 9521 10059
rect 9412 10049 9468 10057
rect 8715 9792 9613 9804
rect 8715 9736 8727 9792
rect 8783 9736 9545 9792
rect 9601 9736 9613 9792
rect 8715 9724 9613 9736
rect 7830 9618 7842 9674
rect 7898 9618 7900 9674
rect 7830 9616 7900 9618
rect 8142 9674 8202 9678
rect 8142 9618 8144 9674
rect 8200 9618 8202 9674
rect 7842 9004 7898 9616
rect 8142 9606 8202 9618
rect 11340 9514 11396 10393
rect 11340 9404 11396 9414
rect 7694 4509 7764 4521
rect 7694 4453 7706 4509
rect 7762 4453 7764 4509
rect 7694 4441 7764 4453
rect 7340 3151 7342 3207
rect 7398 3151 7626 3207
rect 6752 3091 6832 3093
rect 6752 3035 6764 3091
rect 6820 3035 6832 3091
rect 6752 3033 6832 3035
rect 6764 2951 6820 3033
rect 6384 2941 6464 2951
rect 6384 2885 6396 2941
rect 6452 2885 6464 2941
rect 6384 2875 6464 2885
rect 6568 2941 6648 2951
rect 6568 2885 6580 2941
rect 6636 2885 6648 2941
rect 6568 2875 6648 2885
rect 6752 2941 6832 2951
rect 6752 2885 6764 2941
rect 6820 2885 6832 2941
rect 6752 2875 6832 2885
rect 6897 2819 6965 3149
rect 7340 3139 7410 3151
rect 6856 2811 6965 2819
rect 6844 2809 6965 2811
rect 6844 2689 6856 2809
rect 6912 2689 6965 2809
rect 6844 2687 6965 2689
rect 6856 2679 6912 2687
rect 6159 2422 7055 2434
rect 6159 2366 6171 2422
rect 6227 2366 6989 2422
rect 7045 2366 7055 2422
rect 6159 2354 7055 2366
rect 5844 2303 5924 2313
rect 5844 2247 5856 2303
rect 5912 2247 5924 2303
rect 5844 2245 5924 2247
rect 5678 2193 5748 2196
rect 5678 2139 5680 2193
rect 5736 2139 5748 2193
rect 5678 2127 5748 2139
rect 4818 2086 5564 2098
rect 4818 2030 5186 2086
rect 5242 2030 5564 2086
rect 4818 2018 5564 2030
rect 4818 1765 4874 2018
rect 5186 1765 5242 2018
rect 5508 1765 5564 2018
rect 4806 1763 4886 1765
rect 4806 1643 4818 1763
rect 4874 1643 4886 1763
rect 4806 1641 4886 1643
rect 5174 1763 5254 1765
rect 5174 1643 5186 1763
rect 5242 1643 5254 1763
rect 5174 1641 5254 1643
rect 5496 1763 5576 1765
rect 5496 1642 5508 1763
rect 5564 1642 5576 1763
rect 4818 1633 4874 1641
rect 5186 1633 5242 1641
rect 5496 1640 5576 1642
rect 5508 1632 5564 1640
rect 5002 1465 5058 1473
rect 5370 1465 5426 1473
rect 4990 1463 5479 1465
rect 4990 1343 5002 1463
rect 5058 1343 5370 1463
rect 5426 1343 5479 1463
rect 4990 1341 5479 1343
rect 5002 1333 5058 1341
rect 5370 1333 5479 1341
rect 4898 1267 4978 1277
rect 4898 1211 4910 1267
rect 4966 1211 4978 1267
rect 4898 1201 4978 1211
rect 5082 1267 5162 1277
rect 5082 1211 5094 1267
rect 5150 1211 5162 1267
rect 5082 1201 5162 1211
rect 5266 1267 5346 1277
rect 5266 1211 5278 1267
rect 5334 1211 5346 1267
rect 5266 1201 5346 1211
rect 4910 1119 4966 1201
rect 4898 1117 4978 1119
rect 4898 1061 4910 1117
rect 4966 1061 4978 1117
rect 4898 1059 4978 1061
rect 4090 1001 4160 1015
rect 4090 945 4102 1001
rect 4158 945 4160 1001
rect 4090 933 4160 945
rect 3954 885 4024 897
rect 3954 829 3966 885
rect 4022 829 4024 885
rect 3954 817 4024 829
rect 3818 98 3888 110
rect 4102 102 4158 933
rect 4910 745 4966 1059
rect 5094 1003 5150 1201
rect 5082 1001 5162 1003
rect 5082 945 5094 1001
rect 5150 945 5162 1001
rect 5082 943 5162 945
rect 5094 745 5150 943
rect 5278 887 5334 1201
rect 5411 1003 5479 1333
rect 5856 1013 5912 2245
rect 5411 1001 5491 1003
rect 5411 945 5423 1001
rect 5479 945 5491 1001
rect 5411 943 5491 945
rect 5854 1001 5914 1013
rect 5854 945 5856 1001
rect 5912 945 5914 1001
rect 5266 885 5346 887
rect 5266 829 5278 885
rect 5334 829 5346 885
rect 5266 827 5346 829
rect 5278 745 5334 827
rect 4898 735 4978 745
rect 4898 679 4910 735
rect 4966 679 4978 735
rect 4898 669 4978 679
rect 5082 735 5162 745
rect 5082 679 5094 735
rect 5150 679 5162 735
rect 5082 669 5162 679
rect 5266 735 5346 745
rect 5266 679 5278 735
rect 5334 679 5346 735
rect 5266 669 5346 679
rect 5411 613 5479 943
rect 5854 933 5914 945
rect 5370 605 5479 613
rect 5358 603 5479 605
rect 5358 483 5370 603
rect 5426 483 5479 603
rect 5358 481 5479 483
rect 5370 473 5426 481
rect 4673 216 5571 228
rect 4673 160 4685 216
rect 4741 160 5503 216
rect 5559 160 5571 216
rect 4673 148 5571 160
rect 3818 42 3830 98
rect 3886 42 3888 98
rect 3818 30 3888 42
rect 4100 98 4160 102
rect 4100 42 4102 98
rect 4158 42 4160 98
rect 4100 30 4160 42
rect 3694 -175 3750 -165
rect 7706 -65 7762 4441
rect 7842 110 7898 8904
rect 8860 8701 9606 8713
rect 8860 8645 9228 8701
rect 9284 8645 9606 8701
rect 8860 8633 9606 8645
rect 8860 8380 8916 8633
rect 9228 8380 9284 8633
rect 9550 8380 9606 8633
rect 8848 8378 8928 8380
rect 8848 8258 8860 8378
rect 8916 8258 8928 8378
rect 8848 8256 8928 8258
rect 9216 8378 9296 8380
rect 9216 8258 9228 8378
rect 9284 8258 9296 8378
rect 9216 8256 9296 8258
rect 9538 8378 9618 8380
rect 9538 8257 9550 8378
rect 9606 8257 9618 8378
rect 8860 8248 8916 8256
rect 9228 8248 9284 8256
rect 9538 8255 9618 8257
rect 9550 8247 9606 8255
rect 9044 8080 9100 8088
rect 9412 8080 9468 8088
rect 9032 8078 9521 8080
rect 9032 7958 9044 8078
rect 9100 7958 9412 8078
rect 9468 7958 9521 8078
rect 9032 7956 9521 7958
rect 9044 7948 9100 7956
rect 9412 7948 9521 7956
rect 8940 7882 9020 7892
rect 8940 7826 8952 7882
rect 9008 7826 9020 7882
rect 8940 7816 9020 7826
rect 9124 7882 9204 7892
rect 9124 7826 9136 7882
rect 9192 7826 9204 7882
rect 9124 7816 9204 7826
rect 9308 7882 9388 7892
rect 9308 7826 9320 7882
rect 9376 7826 9388 7882
rect 9308 7816 9388 7826
rect 8052 7732 8138 7744
rect 8952 7734 9008 7816
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 8940 7732 9020 7734
rect 8940 7676 8952 7732
rect 9008 7676 9020 7732
rect 8940 7674 9020 7676
rect 8268 7616 8338 7628
rect 8268 7560 8280 7616
rect 8336 7560 8338 7616
rect 8268 7548 8338 7560
rect 8132 5411 8202 5425
rect 8132 5355 8144 5411
rect 8200 5355 8202 5411
rect 8132 5343 8202 5355
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 7978 897 8034 5165
rect 8144 1015 8200 5343
rect 8280 3102 8336 7548
rect 8952 7360 9008 7674
rect 9136 7618 9192 7816
rect 9124 7616 9204 7618
rect 9124 7560 9136 7616
rect 9192 7560 9204 7616
rect 9124 7558 9204 7560
rect 9136 7360 9192 7558
rect 9320 7502 9376 7816
rect 9453 7618 9521 7948
rect 9453 7616 9533 7618
rect 9453 7560 9465 7616
rect 9521 7560 9533 7616
rect 9453 7558 9533 7560
rect 9720 7616 9790 7628
rect 9720 7560 9722 7616
rect 9778 7560 9790 7616
rect 9308 7500 9388 7502
rect 9308 7444 9320 7500
rect 9376 7444 9388 7500
rect 9308 7442 9388 7444
rect 9320 7360 9376 7442
rect 8940 7350 9020 7360
rect 8940 7294 8952 7350
rect 9008 7294 9020 7350
rect 8940 7284 9020 7294
rect 9124 7350 9204 7360
rect 9124 7294 9136 7350
rect 9192 7294 9204 7350
rect 9124 7284 9204 7294
rect 9308 7350 9388 7360
rect 9308 7294 9320 7350
rect 9376 7294 9388 7350
rect 9308 7284 9388 7294
rect 9453 7228 9521 7558
rect 9720 7550 9790 7560
rect 9412 7220 9521 7228
rect 9400 7218 9521 7220
rect 9400 7098 9412 7218
rect 9468 7098 9521 7218
rect 9400 7096 9521 7098
rect 9412 7088 9468 7096
rect 8715 6831 9613 6843
rect 8715 6775 8727 6831
rect 8783 6775 9545 6831
rect 9601 6775 9613 6831
rect 8715 6763 9613 6775
rect 9722 6606 9778 7550
rect 9886 6713 9966 6723
rect 9886 6657 9898 6713
rect 9954 6657 9966 6713
rect 9886 6655 9966 6657
rect 9720 6603 9790 6606
rect 9720 6549 9722 6603
rect 9778 6549 9790 6603
rect 9720 6537 9790 6549
rect 8860 6496 9606 6508
rect 8860 6440 9228 6496
rect 9284 6440 9606 6496
rect 8860 6428 9606 6440
rect 8860 6175 8916 6428
rect 9228 6175 9284 6428
rect 9550 6175 9606 6428
rect 8848 6173 8928 6175
rect 8848 6053 8860 6173
rect 8916 6053 8928 6173
rect 8848 6051 8928 6053
rect 9216 6173 9296 6175
rect 9216 6053 9228 6173
rect 9284 6053 9296 6173
rect 9216 6051 9296 6053
rect 9538 6173 9618 6175
rect 9538 6052 9550 6173
rect 9606 6052 9618 6173
rect 8860 6043 8916 6051
rect 9228 6043 9284 6051
rect 9538 6050 9618 6052
rect 9550 6042 9606 6050
rect 9044 5875 9100 5883
rect 9412 5875 9468 5883
rect 9032 5873 9521 5875
rect 9032 5753 9044 5873
rect 9100 5753 9412 5873
rect 9468 5753 9521 5873
rect 9032 5751 9521 5753
rect 9044 5743 9100 5751
rect 9412 5743 9521 5751
rect 8940 5677 9020 5687
rect 8940 5621 8952 5677
rect 9008 5621 9020 5677
rect 8940 5611 9020 5621
rect 9124 5677 9204 5687
rect 9124 5621 9136 5677
rect 9192 5621 9204 5677
rect 9124 5611 9204 5621
rect 9308 5677 9388 5687
rect 9308 5621 9320 5677
rect 9376 5621 9388 5677
rect 9308 5611 9388 5621
rect 8952 5529 9008 5611
rect 8940 5527 9020 5529
rect 8940 5471 8952 5527
rect 9008 5471 9020 5527
rect 8940 5469 9020 5471
rect 8952 5155 9008 5469
rect 9136 5413 9192 5611
rect 9124 5411 9204 5413
rect 9124 5355 9136 5411
rect 9192 5355 9204 5411
rect 9124 5353 9204 5355
rect 9136 5155 9192 5353
rect 9320 5297 9376 5611
rect 9453 5413 9521 5743
rect 9898 5421 9954 6655
rect 10346 6496 11092 6508
rect 10346 6440 10714 6496
rect 10770 6440 11092 6496
rect 10346 6428 11092 6440
rect 10346 6175 10402 6428
rect 10714 6175 10770 6428
rect 11036 6175 11092 6428
rect 10334 6173 10414 6175
rect 10334 6053 10346 6173
rect 10402 6053 10414 6173
rect 10334 6051 10414 6053
rect 10702 6173 10782 6175
rect 10702 6053 10714 6173
rect 10770 6053 10782 6173
rect 10702 6051 10782 6053
rect 11024 6173 11104 6175
rect 11024 6052 11036 6173
rect 11092 6052 11104 6173
rect 10346 6043 10402 6051
rect 10714 6043 10770 6051
rect 11024 6050 11104 6052
rect 11036 6042 11092 6050
rect 10530 5875 10586 5883
rect 10898 5875 10954 5883
rect 10518 5873 11007 5875
rect 10518 5753 10530 5873
rect 10586 5753 10898 5873
rect 10954 5753 11007 5873
rect 10518 5751 11007 5753
rect 10530 5743 10586 5751
rect 10898 5743 11007 5751
rect 10426 5677 10506 5687
rect 10426 5621 10438 5677
rect 10494 5621 10506 5677
rect 10426 5611 10506 5621
rect 10610 5677 10690 5687
rect 10610 5621 10622 5677
rect 10678 5621 10690 5677
rect 10610 5611 10690 5621
rect 10794 5677 10874 5687
rect 10794 5621 10806 5677
rect 10862 5621 10874 5677
rect 10794 5611 10874 5621
rect 10438 5529 10494 5611
rect 10426 5527 10506 5529
rect 10426 5471 10438 5527
rect 10494 5471 10506 5527
rect 10426 5469 10506 5471
rect 9453 5411 9533 5413
rect 9453 5355 9465 5411
rect 9521 5355 9533 5411
rect 9453 5353 9533 5355
rect 9896 5411 9956 5421
rect 9896 5355 9898 5411
rect 9954 5355 9956 5411
rect 9308 5295 9388 5297
rect 9308 5239 9320 5295
rect 9376 5239 9388 5295
rect 9308 5237 9388 5239
rect 9320 5155 9376 5237
rect 8940 5145 9020 5155
rect 8940 5089 8952 5145
rect 9008 5089 9020 5145
rect 8940 5079 9020 5089
rect 9124 5145 9204 5155
rect 9124 5089 9136 5145
rect 9192 5089 9204 5145
rect 9124 5079 9204 5089
rect 9308 5145 9388 5155
rect 9308 5089 9320 5145
rect 9376 5089 9388 5145
rect 9308 5079 9388 5089
rect 9453 5023 9521 5353
rect 9896 5343 9956 5355
rect 9412 5015 9521 5023
rect 9400 5013 9521 5015
rect 9400 4893 9412 5013
rect 9468 4893 9521 5013
rect 9400 4891 9521 4893
rect 9412 4883 9468 4891
rect 8715 4626 9611 4638
rect 8715 4570 8727 4626
rect 8783 4570 9545 4626
rect 9601 4570 9611 4626
rect 8715 4558 9611 4570
rect 9898 4400 9954 5343
rect 10438 5155 10494 5469
rect 10622 5413 10678 5611
rect 10610 5411 10690 5413
rect 10610 5355 10622 5411
rect 10678 5355 10690 5411
rect 10610 5353 10690 5355
rect 10622 5155 10678 5353
rect 10806 5297 10862 5611
rect 10939 5413 11007 5743
rect 10939 5411 11019 5413
rect 10939 5355 10951 5411
rect 11007 5355 11019 5411
rect 10939 5353 11019 5355
rect 11206 5411 11276 5423
rect 11206 5355 11208 5411
rect 11264 5355 11532 5411
rect 10794 5295 10874 5297
rect 10794 5239 10806 5295
rect 10862 5239 10874 5295
rect 10794 5237 10874 5239
rect 10806 5155 10862 5237
rect 10426 5145 10506 5155
rect 10426 5089 10438 5145
rect 10494 5089 10506 5145
rect 10426 5079 10506 5089
rect 10610 5145 10690 5155
rect 10610 5089 10622 5145
rect 10678 5089 10690 5145
rect 10610 5079 10690 5089
rect 10794 5145 10874 5155
rect 10794 5089 10806 5145
rect 10862 5089 10874 5145
rect 10794 5079 10874 5089
rect 10939 5023 11007 5353
rect 11206 5345 11276 5355
rect 10898 5015 11007 5023
rect 10886 5013 11007 5015
rect 10886 4893 10898 5013
rect 10954 4893 11007 5013
rect 10886 4891 11007 4893
rect 10898 4883 10954 4891
rect 10201 4626 11097 4638
rect 10201 4570 10213 4626
rect 10269 4570 11031 4626
rect 11087 4570 11097 4626
rect 10201 4558 11097 4570
rect 11208 4401 11264 5345
rect 11372 4509 11452 4519
rect 11372 4453 11384 4509
rect 11440 4453 11452 4509
rect 11372 4451 11452 4453
rect 9896 4398 9966 4400
rect 9896 4342 9898 4398
rect 9954 4342 9966 4398
rect 9896 4330 9966 4342
rect 11196 4399 11276 4401
rect 11196 4343 11208 4399
rect 11264 4343 11276 4399
rect 11196 4331 11276 4343
rect 8860 4291 9606 4303
rect 8860 4235 9228 4291
rect 9284 4235 9606 4291
rect 8860 4223 9606 4235
rect 8860 3970 8916 4223
rect 9228 3970 9284 4223
rect 9550 3970 9606 4223
rect 10346 4292 11092 4304
rect 10346 4236 10714 4292
rect 10770 4236 11092 4292
rect 10346 4224 11092 4236
rect 10346 3971 10402 4224
rect 10714 3971 10770 4224
rect 11036 3971 11092 4224
rect 8848 3968 8928 3970
rect 8848 3848 8860 3968
rect 8916 3848 8928 3968
rect 8848 3846 8928 3848
rect 9216 3968 9296 3970
rect 9216 3848 9228 3968
rect 9284 3848 9296 3968
rect 9216 3846 9296 3848
rect 9538 3968 9618 3970
rect 9538 3847 9550 3968
rect 9606 3847 9618 3968
rect 10334 3969 10414 3971
rect 10334 3849 10346 3969
rect 10402 3849 10414 3969
rect 10334 3847 10414 3849
rect 10702 3969 10782 3971
rect 10702 3849 10714 3969
rect 10770 3849 10782 3969
rect 10702 3847 10782 3849
rect 11024 3969 11104 3971
rect 11024 3848 11036 3969
rect 11092 3848 11104 3969
rect 8860 3838 8916 3846
rect 9228 3838 9284 3846
rect 9538 3845 9618 3847
rect 9550 3837 9606 3845
rect 10346 3839 10402 3847
rect 10714 3839 10770 3847
rect 11024 3846 11104 3848
rect 11036 3838 11092 3846
rect 9044 3670 9100 3678
rect 9412 3670 9468 3678
rect 10530 3671 10586 3679
rect 10898 3671 10954 3679
rect 9032 3668 9521 3670
rect 9032 3548 9044 3668
rect 9100 3548 9412 3668
rect 9468 3548 9521 3668
rect 9032 3546 9521 3548
rect 10518 3669 11007 3671
rect 10518 3549 10530 3669
rect 10586 3549 10898 3669
rect 10954 3549 11007 3669
rect 10518 3547 11007 3549
rect 9044 3538 9100 3546
rect 9412 3538 9521 3546
rect 10530 3539 10586 3547
rect 10898 3539 11007 3547
rect 8940 3472 9020 3482
rect 8940 3416 8952 3472
rect 9008 3416 9020 3472
rect 8940 3406 9020 3416
rect 9124 3472 9204 3482
rect 9124 3416 9136 3472
rect 9192 3416 9204 3472
rect 9124 3406 9204 3416
rect 9308 3472 9388 3482
rect 9308 3416 9320 3472
rect 9376 3416 9388 3472
rect 9308 3406 9388 3416
rect 8952 3324 9008 3406
rect 8940 3322 9020 3324
rect 8940 3266 8952 3322
rect 9008 3266 9020 3322
rect 8940 3264 9020 3266
rect 8268 3090 8338 3102
rect 8268 3034 8280 3090
rect 8336 3034 8338 3090
rect 8268 3022 8338 3034
rect 8952 2950 9008 3264
rect 9136 3208 9192 3406
rect 9124 3206 9204 3208
rect 9124 3150 9136 3206
rect 9192 3150 9204 3206
rect 9124 3148 9204 3150
rect 9136 2950 9192 3148
rect 9320 3092 9376 3406
rect 9453 3208 9521 3538
rect 10426 3473 10506 3483
rect 10426 3417 10438 3473
rect 10494 3417 10506 3473
rect 10426 3407 10506 3417
rect 10610 3473 10690 3483
rect 10610 3417 10622 3473
rect 10678 3417 10690 3473
rect 10610 3407 10690 3417
rect 10794 3473 10874 3483
rect 10794 3417 10806 3473
rect 10862 3417 10874 3473
rect 10794 3407 10874 3417
rect 10438 3325 10494 3407
rect 10426 3323 10506 3325
rect 10426 3267 10438 3323
rect 10494 3267 10506 3323
rect 10426 3265 10506 3267
rect 9453 3206 9533 3208
rect 9453 3150 9465 3206
rect 9521 3150 9533 3206
rect 9453 3148 9533 3150
rect 9720 3206 9790 3218
rect 9720 3150 9722 3206
rect 9778 3150 9790 3206
rect 9308 3090 9388 3092
rect 9308 3034 9320 3090
rect 9376 3034 9388 3090
rect 9308 3032 9388 3034
rect 9320 2950 9376 3032
rect 8940 2940 9020 2950
rect 8940 2884 8952 2940
rect 9008 2884 9020 2940
rect 8940 2874 9020 2884
rect 9124 2940 9204 2950
rect 9124 2884 9136 2940
rect 9192 2884 9204 2940
rect 9124 2874 9204 2884
rect 9308 2940 9388 2950
rect 9308 2884 9320 2940
rect 9376 2884 9388 2940
rect 9308 2874 9388 2884
rect 9453 2818 9521 3148
rect 9720 3140 9790 3150
rect 9412 2810 9521 2818
rect 9400 2808 9521 2810
rect 9400 2688 9412 2808
rect 9468 2688 9521 2808
rect 9400 2686 9521 2688
rect 9412 2678 9468 2686
rect 8715 2421 9611 2433
rect 8715 2365 8727 2421
rect 8783 2365 9545 2421
rect 9601 2365 9611 2421
rect 8715 2353 9611 2365
rect 9722 2196 9778 3140
rect 10438 2951 10494 3265
rect 10622 3209 10678 3407
rect 10610 3207 10690 3209
rect 10610 3151 10622 3207
rect 10678 3151 10690 3207
rect 10610 3149 10690 3151
rect 10622 2951 10678 3149
rect 10806 3093 10862 3407
rect 10939 3209 11007 3539
rect 11384 3217 11440 4451
rect 10939 3207 11019 3209
rect 10939 3151 10951 3207
rect 11007 3151 11019 3207
rect 10939 3149 11019 3151
rect 11382 3207 11452 3217
rect 11612 3207 11668 17250
rect 11760 14999 11816 18679
rect 11758 14987 11828 14999
rect 11758 14931 11760 14987
rect 11816 14931 11828 14987
rect 11758 14919 11828 14931
rect 12050 14087 12106 19031
rect 15856 18563 15912 19501
rect 19898 19091 19954 19501
rect 19896 19089 19966 19091
rect 19896 19033 19898 19089
rect 19954 19033 19966 19089
rect 19896 19031 19966 19033
rect 16080 18913 16150 18925
rect 16080 18857 16092 18913
rect 16148 18857 16150 18913
rect 16080 18855 16150 18857
rect 15854 18561 15924 18563
rect 15854 18505 15856 18561
rect 15912 18505 15924 18561
rect 15854 18503 15924 18505
rect 12902 18277 13648 18289
rect 12902 18221 13270 18277
rect 13326 18221 13648 18277
rect 12902 18209 13648 18221
rect 12902 17956 12958 18209
rect 13270 17956 13326 18209
rect 13592 17956 13648 18209
rect 12890 17954 12970 17956
rect 12890 17834 12902 17954
rect 12958 17834 12970 17954
rect 12890 17832 12970 17834
rect 13258 17954 13338 17956
rect 13258 17834 13270 17954
rect 13326 17834 13338 17954
rect 13258 17832 13338 17834
rect 13580 17954 13660 17956
rect 13580 17833 13592 17954
rect 13648 17833 13660 17954
rect 12902 17824 12958 17832
rect 13270 17824 13326 17832
rect 13580 17831 13660 17833
rect 13592 17823 13648 17831
rect 13086 17656 13142 17664
rect 13454 17656 13510 17664
rect 13074 17654 13563 17656
rect 13074 17534 13086 17654
rect 13142 17534 13454 17654
rect 13510 17534 13563 17654
rect 13074 17532 13563 17534
rect 13086 17524 13142 17532
rect 13454 17524 13563 17532
rect 12982 17458 13062 17468
rect 12982 17402 12994 17458
rect 13050 17402 13062 17458
rect 12982 17392 13062 17402
rect 13166 17458 13246 17468
rect 13166 17402 13178 17458
rect 13234 17402 13246 17458
rect 13166 17392 13246 17402
rect 13350 17458 13430 17468
rect 13350 17402 13362 17458
rect 13418 17402 13430 17458
rect 13350 17392 13430 17402
rect 12994 17310 13050 17392
rect 12982 17308 13062 17310
rect 12982 17252 12994 17308
rect 13050 17252 13062 17308
rect 12982 17250 13062 17252
rect 12310 17192 12380 17204
rect 12310 17136 12322 17192
rect 12378 17136 12380 17192
rect 12310 17124 12380 17136
rect 12174 14987 12244 15001
rect 12174 14931 12186 14987
rect 12242 14931 12244 14987
rect 12174 14919 12244 14931
rect 12038 14085 12108 14087
rect 12038 14029 12050 14085
rect 12106 14029 12108 14085
rect 12038 14017 12108 14029
rect 12186 10591 12242 14919
rect 12322 12678 12378 17124
rect 12994 16936 13050 17250
rect 13178 17194 13234 17392
rect 13166 17192 13246 17194
rect 13166 17136 13178 17192
rect 13234 17136 13246 17192
rect 13166 17134 13246 17136
rect 13178 16936 13234 17134
rect 13362 17078 13418 17392
rect 13495 17194 13563 17524
rect 15642 17308 15712 17320
rect 15642 17252 15654 17308
rect 15710 17252 15712 17308
rect 15642 17250 15712 17252
rect 13495 17192 13575 17194
rect 13495 17136 13507 17192
rect 13563 17136 13575 17192
rect 13495 17134 13575 17136
rect 13762 17192 13832 17204
rect 13762 17136 13764 17192
rect 13820 17136 13832 17192
rect 13350 17076 13430 17078
rect 13350 17020 13362 17076
rect 13418 17020 13430 17076
rect 13350 17018 13430 17020
rect 13362 16936 13418 17018
rect 12982 16926 13062 16936
rect 12982 16870 12994 16926
rect 13050 16870 13062 16926
rect 12982 16860 13062 16870
rect 13166 16926 13246 16936
rect 13166 16870 13178 16926
rect 13234 16870 13246 16926
rect 13166 16860 13246 16870
rect 13350 16926 13430 16936
rect 13350 16870 13362 16926
rect 13418 16870 13430 16926
rect 13350 16860 13430 16870
rect 13495 16804 13563 17134
rect 13762 17126 13832 17136
rect 13454 16796 13563 16804
rect 13442 16794 13563 16796
rect 13442 16674 13454 16794
rect 13510 16674 13563 16794
rect 13442 16672 13563 16674
rect 13454 16664 13510 16672
rect 12757 16407 13655 16419
rect 12757 16351 12769 16407
rect 12825 16351 13587 16407
rect 13643 16351 13655 16407
rect 12757 16339 13655 16351
rect 13764 16182 13820 17126
rect 13928 16289 14008 16299
rect 13928 16233 13940 16289
rect 13996 16233 14008 16289
rect 13928 16231 14008 16233
rect 13762 16179 13832 16182
rect 13762 16125 13764 16179
rect 13820 16125 13832 16179
rect 13762 16113 13832 16125
rect 12902 16072 13648 16084
rect 12902 16016 13270 16072
rect 13326 16016 13648 16072
rect 12902 16004 13648 16016
rect 12902 15751 12958 16004
rect 13270 15751 13326 16004
rect 13592 15751 13648 16004
rect 12890 15749 12970 15751
rect 12890 15629 12902 15749
rect 12958 15629 12970 15749
rect 12890 15627 12970 15629
rect 13258 15749 13338 15751
rect 13258 15629 13270 15749
rect 13326 15629 13338 15749
rect 13258 15627 13338 15629
rect 13580 15749 13660 15751
rect 13580 15628 13592 15749
rect 13648 15628 13660 15749
rect 12902 15619 12958 15627
rect 13270 15619 13326 15627
rect 13580 15626 13660 15628
rect 13592 15618 13648 15626
rect 13086 15451 13142 15459
rect 13454 15451 13510 15459
rect 13074 15449 13563 15451
rect 13074 15329 13086 15449
rect 13142 15329 13454 15449
rect 13510 15329 13563 15449
rect 13074 15327 13563 15329
rect 13086 15319 13142 15327
rect 13454 15319 13563 15327
rect 12982 15253 13062 15263
rect 12982 15197 12994 15253
rect 13050 15197 13062 15253
rect 12982 15187 13062 15197
rect 13166 15253 13246 15263
rect 13166 15197 13178 15253
rect 13234 15197 13246 15253
rect 13166 15187 13246 15197
rect 13350 15253 13430 15263
rect 13350 15197 13362 15253
rect 13418 15197 13430 15253
rect 13350 15187 13430 15197
rect 12994 15105 13050 15187
rect 12982 15103 13062 15105
rect 12982 15047 12994 15103
rect 13050 15047 13062 15103
rect 12982 15045 13062 15047
rect 12994 14731 13050 15045
rect 13178 14989 13234 15187
rect 13166 14987 13246 14989
rect 13166 14931 13178 14987
rect 13234 14931 13246 14987
rect 13166 14929 13246 14931
rect 13178 14731 13234 14929
rect 13362 14873 13418 15187
rect 13495 14989 13563 15319
rect 13940 14997 13996 16231
rect 14388 16072 15134 16084
rect 14388 16016 14756 16072
rect 14812 16016 15134 16072
rect 14388 16004 15134 16016
rect 14388 15751 14444 16004
rect 14756 15751 14812 16004
rect 15078 15751 15134 16004
rect 14376 15749 14456 15751
rect 14376 15629 14388 15749
rect 14444 15629 14456 15749
rect 14376 15627 14456 15629
rect 14744 15749 14824 15751
rect 14744 15629 14756 15749
rect 14812 15629 14824 15749
rect 14744 15627 14824 15629
rect 15066 15749 15146 15751
rect 15066 15628 15078 15749
rect 15134 15628 15146 15749
rect 14388 15619 14444 15627
rect 14756 15619 14812 15627
rect 15066 15626 15146 15628
rect 15078 15618 15134 15626
rect 14572 15451 14628 15459
rect 14940 15451 14996 15459
rect 14560 15449 15049 15451
rect 14560 15329 14572 15449
rect 14628 15329 14940 15449
rect 14996 15329 15049 15449
rect 14560 15327 15049 15329
rect 14572 15319 14628 15327
rect 14940 15319 15049 15327
rect 14468 15253 14548 15263
rect 14468 15197 14480 15253
rect 14536 15197 14548 15253
rect 14468 15187 14548 15197
rect 14652 15253 14732 15263
rect 14652 15197 14664 15253
rect 14720 15197 14732 15253
rect 14652 15187 14732 15197
rect 14836 15253 14916 15263
rect 14836 15197 14848 15253
rect 14904 15197 14916 15253
rect 14836 15187 14916 15197
rect 14480 15105 14536 15187
rect 14468 15103 14548 15105
rect 14468 15047 14480 15103
rect 14536 15047 14548 15103
rect 14468 15045 14548 15047
rect 13495 14987 13575 14989
rect 13495 14931 13507 14987
rect 13563 14931 13575 14987
rect 13495 14929 13575 14931
rect 13938 14987 13998 14997
rect 13938 14931 13940 14987
rect 13996 14931 13998 14987
rect 13350 14871 13430 14873
rect 13350 14815 13362 14871
rect 13418 14815 13430 14871
rect 13350 14813 13430 14815
rect 13362 14731 13418 14813
rect 12982 14721 13062 14731
rect 12982 14665 12994 14721
rect 13050 14665 13062 14721
rect 12982 14655 13062 14665
rect 13166 14721 13246 14731
rect 13166 14665 13178 14721
rect 13234 14665 13246 14721
rect 13166 14655 13246 14665
rect 13350 14721 13430 14731
rect 13350 14665 13362 14721
rect 13418 14665 13430 14721
rect 13350 14655 13430 14665
rect 13495 14599 13563 14929
rect 13938 14919 13998 14931
rect 13454 14591 13563 14599
rect 13442 14589 13563 14591
rect 13442 14469 13454 14589
rect 13510 14469 13563 14589
rect 13442 14467 13563 14469
rect 13454 14459 13510 14467
rect 12757 14202 13653 14214
rect 12757 14146 12769 14202
rect 12825 14146 13587 14202
rect 13643 14146 13653 14202
rect 12757 14134 13653 14146
rect 13940 13976 13996 14919
rect 14480 14731 14536 15045
rect 14664 14989 14720 15187
rect 14652 14987 14732 14989
rect 14652 14931 14664 14987
rect 14720 14931 14732 14987
rect 14652 14929 14732 14931
rect 14664 14731 14720 14929
rect 14848 14873 14904 15187
rect 14981 14989 15049 15319
rect 14981 14987 15061 14989
rect 14981 14931 14993 14987
rect 15049 14931 15061 14987
rect 14981 14929 15061 14931
rect 15248 14987 15318 14999
rect 15248 14931 15250 14987
rect 15306 14931 15574 14987
rect 14836 14871 14916 14873
rect 14836 14815 14848 14871
rect 14904 14815 14916 14871
rect 14836 14813 14916 14815
rect 14848 14731 14904 14813
rect 14468 14721 14548 14731
rect 14468 14665 14480 14721
rect 14536 14665 14548 14721
rect 14468 14655 14548 14665
rect 14652 14721 14732 14731
rect 14652 14665 14664 14721
rect 14720 14665 14732 14721
rect 14652 14655 14732 14665
rect 14836 14721 14916 14731
rect 14836 14665 14848 14721
rect 14904 14665 14916 14721
rect 14836 14655 14916 14665
rect 14981 14599 15049 14929
rect 15248 14921 15318 14931
rect 14940 14591 15049 14599
rect 14928 14589 15049 14591
rect 14928 14469 14940 14589
rect 14996 14469 15049 14589
rect 14928 14467 15049 14469
rect 14940 14459 14996 14467
rect 14243 14202 15139 14214
rect 14243 14146 14255 14202
rect 14311 14146 15073 14202
rect 15129 14146 15139 14202
rect 14243 14134 15139 14146
rect 15250 13977 15306 14921
rect 15414 14085 15494 14095
rect 15414 14029 15426 14085
rect 15482 14029 15494 14085
rect 15414 14027 15494 14029
rect 13938 13974 14008 13976
rect 13938 13918 13940 13974
rect 13996 13918 14008 13974
rect 13938 13906 14008 13918
rect 15238 13975 15318 13977
rect 15238 13919 15250 13975
rect 15306 13919 15318 13975
rect 15238 13907 15318 13919
rect 12902 13867 13648 13879
rect 12902 13811 13270 13867
rect 13326 13811 13648 13867
rect 12902 13799 13648 13811
rect 12902 13546 12958 13799
rect 13270 13546 13326 13799
rect 13592 13546 13648 13799
rect 14388 13868 15134 13880
rect 14388 13812 14756 13868
rect 14812 13812 15134 13868
rect 14388 13800 15134 13812
rect 14388 13547 14444 13800
rect 14756 13547 14812 13800
rect 15078 13547 15134 13800
rect 12890 13544 12970 13546
rect 12890 13424 12902 13544
rect 12958 13424 12970 13544
rect 12890 13422 12970 13424
rect 13258 13544 13338 13546
rect 13258 13424 13270 13544
rect 13326 13424 13338 13544
rect 13258 13422 13338 13424
rect 13580 13544 13660 13546
rect 13580 13423 13592 13544
rect 13648 13423 13660 13544
rect 14376 13545 14456 13547
rect 14376 13425 14388 13545
rect 14444 13425 14456 13545
rect 14376 13423 14456 13425
rect 14744 13545 14824 13547
rect 14744 13425 14756 13545
rect 14812 13425 14824 13545
rect 14744 13423 14824 13425
rect 15066 13545 15146 13547
rect 15066 13424 15078 13545
rect 15134 13424 15146 13545
rect 12902 13414 12958 13422
rect 13270 13414 13326 13422
rect 13580 13421 13660 13423
rect 13592 13413 13648 13421
rect 14388 13415 14444 13423
rect 14756 13415 14812 13423
rect 15066 13422 15146 13424
rect 15078 13414 15134 13422
rect 13086 13246 13142 13254
rect 13454 13246 13510 13254
rect 14572 13247 14628 13255
rect 14940 13247 14996 13255
rect 13074 13244 13563 13246
rect 13074 13124 13086 13244
rect 13142 13124 13454 13244
rect 13510 13124 13563 13244
rect 13074 13122 13563 13124
rect 14560 13245 15049 13247
rect 14560 13125 14572 13245
rect 14628 13125 14940 13245
rect 14996 13125 15049 13245
rect 14560 13123 15049 13125
rect 13086 13114 13142 13122
rect 13454 13114 13563 13122
rect 14572 13115 14628 13123
rect 14940 13115 15049 13123
rect 12982 13048 13062 13058
rect 12982 12992 12994 13048
rect 13050 12992 13062 13048
rect 12982 12982 13062 12992
rect 13166 13048 13246 13058
rect 13166 12992 13178 13048
rect 13234 12992 13246 13048
rect 13166 12982 13246 12992
rect 13350 13048 13430 13058
rect 13350 12992 13362 13048
rect 13418 12992 13430 13048
rect 13350 12982 13430 12992
rect 12994 12900 13050 12982
rect 12982 12898 13062 12900
rect 12982 12842 12994 12898
rect 13050 12842 13062 12898
rect 12982 12840 13062 12842
rect 12310 12666 12380 12678
rect 12310 12610 12322 12666
rect 12378 12610 12380 12666
rect 12310 12598 12380 12610
rect 12994 12526 13050 12840
rect 13178 12784 13234 12982
rect 13166 12782 13246 12784
rect 13166 12726 13178 12782
rect 13234 12726 13246 12782
rect 13166 12724 13246 12726
rect 13178 12526 13234 12724
rect 13362 12668 13418 12982
rect 13495 12784 13563 13114
rect 14468 13049 14548 13059
rect 14468 12993 14480 13049
rect 14536 12993 14548 13049
rect 14468 12983 14548 12993
rect 14652 13049 14732 13059
rect 14652 12993 14664 13049
rect 14720 12993 14732 13049
rect 14652 12983 14732 12993
rect 14836 13049 14916 13059
rect 14836 12993 14848 13049
rect 14904 12993 14916 13049
rect 14836 12983 14916 12993
rect 14480 12901 14536 12983
rect 14468 12899 14548 12901
rect 14468 12843 14480 12899
rect 14536 12843 14548 12899
rect 14468 12841 14548 12843
rect 13495 12782 13575 12784
rect 13495 12726 13507 12782
rect 13563 12726 13575 12782
rect 13495 12724 13575 12726
rect 13762 12782 13832 12794
rect 13762 12726 13764 12782
rect 13820 12726 13832 12782
rect 13350 12666 13430 12668
rect 13350 12610 13362 12666
rect 13418 12610 13430 12666
rect 13350 12608 13430 12610
rect 13362 12526 13418 12608
rect 12982 12516 13062 12526
rect 12982 12460 12994 12516
rect 13050 12460 13062 12516
rect 12982 12450 13062 12460
rect 13166 12516 13246 12526
rect 13166 12460 13178 12516
rect 13234 12460 13246 12516
rect 13166 12450 13246 12460
rect 13350 12516 13430 12526
rect 13350 12460 13362 12516
rect 13418 12460 13430 12516
rect 13350 12450 13430 12460
rect 13495 12394 13563 12724
rect 13762 12716 13832 12726
rect 13454 12386 13563 12394
rect 13442 12384 13563 12386
rect 13442 12264 13454 12384
rect 13510 12264 13563 12384
rect 13442 12262 13563 12264
rect 13454 12254 13510 12262
rect 12757 11997 13653 12009
rect 12757 11941 12769 11997
rect 12825 11941 13587 11997
rect 13643 11941 13653 11997
rect 12757 11929 13653 11941
rect 13764 11772 13820 12716
rect 14480 12527 14536 12841
rect 14664 12785 14720 12983
rect 14652 12783 14732 12785
rect 14652 12727 14664 12783
rect 14720 12727 14732 12783
rect 14652 12725 14732 12727
rect 14664 12527 14720 12725
rect 14848 12669 14904 12983
rect 14981 12785 15049 13115
rect 15426 12793 15482 14027
rect 14981 12783 15061 12785
rect 14981 12727 14993 12783
rect 15049 12727 15061 12783
rect 14981 12725 15061 12727
rect 15424 12783 15494 12793
rect 15424 12727 15426 12783
rect 15482 12727 15574 12783
rect 14836 12667 14916 12669
rect 14836 12611 14848 12667
rect 14904 12611 14916 12667
rect 14836 12609 14916 12611
rect 14848 12527 14904 12609
rect 14468 12517 14548 12527
rect 14468 12461 14480 12517
rect 14536 12461 14548 12517
rect 14468 12451 14548 12461
rect 14652 12517 14732 12527
rect 14652 12461 14664 12517
rect 14720 12461 14732 12517
rect 14652 12451 14732 12461
rect 14836 12517 14916 12527
rect 14836 12461 14848 12517
rect 14904 12461 14916 12517
rect 14836 12451 14916 12461
rect 14981 12395 15049 12725
rect 15424 12715 15494 12727
rect 14940 12387 15049 12395
rect 14928 12385 15049 12387
rect 14928 12265 14940 12385
rect 14996 12265 15049 12385
rect 14928 12263 15049 12265
rect 14940 12255 14996 12263
rect 14243 11998 15139 12010
rect 14243 11942 14255 11998
rect 14311 11942 15073 11998
rect 15129 11942 15139 11998
rect 14243 11930 15139 11942
rect 13928 11879 14008 11889
rect 13928 11823 13940 11879
rect 13996 11823 14008 11879
rect 13928 11821 14008 11823
rect 13762 11769 13832 11772
rect 13762 11715 13764 11769
rect 13820 11715 13832 11769
rect 13762 11703 13832 11715
rect 12902 11662 13648 11674
rect 12902 11606 13270 11662
rect 13326 11606 13648 11662
rect 12902 11594 13648 11606
rect 12902 11341 12958 11594
rect 13270 11341 13326 11594
rect 13592 11341 13648 11594
rect 12890 11339 12970 11341
rect 12890 11219 12902 11339
rect 12958 11219 12970 11339
rect 12890 11217 12970 11219
rect 13258 11339 13338 11341
rect 13258 11219 13270 11339
rect 13326 11219 13338 11339
rect 13258 11217 13338 11219
rect 13580 11339 13660 11341
rect 13580 11218 13592 11339
rect 13648 11218 13660 11339
rect 12902 11209 12958 11217
rect 13270 11209 13326 11217
rect 13580 11216 13660 11218
rect 13592 11208 13648 11216
rect 13086 11041 13142 11049
rect 13454 11041 13510 11049
rect 13074 11039 13563 11041
rect 13074 10919 13086 11039
rect 13142 10919 13454 11039
rect 13510 10919 13563 11039
rect 13074 10917 13563 10919
rect 13086 10909 13142 10917
rect 13454 10909 13563 10917
rect 12982 10843 13062 10853
rect 12982 10787 12994 10843
rect 13050 10787 13062 10843
rect 12982 10777 13062 10787
rect 13166 10843 13246 10853
rect 13166 10787 13178 10843
rect 13234 10787 13246 10843
rect 13166 10777 13246 10787
rect 13350 10843 13430 10853
rect 13350 10787 13362 10843
rect 13418 10787 13430 10843
rect 13350 10777 13430 10787
rect 12994 10695 13050 10777
rect 12982 10693 13062 10695
rect 12982 10637 12994 10693
rect 13050 10637 13062 10693
rect 12982 10635 13062 10637
rect 12174 10577 12244 10591
rect 12174 10521 12186 10577
rect 12242 10521 12244 10577
rect 12174 10509 12244 10521
rect 11872 9674 11942 9686
rect 12186 9678 12242 10509
rect 12994 10321 13050 10635
rect 13178 10579 13234 10777
rect 13166 10577 13246 10579
rect 13166 10521 13178 10577
rect 13234 10521 13246 10577
rect 13166 10519 13246 10521
rect 13178 10321 13234 10519
rect 13362 10463 13418 10777
rect 13495 10579 13563 10909
rect 13940 10589 13996 11821
rect 13495 10577 13575 10579
rect 13495 10521 13507 10577
rect 13563 10521 13575 10577
rect 13495 10519 13575 10521
rect 13938 10577 13998 10589
rect 13938 10521 13940 10577
rect 13996 10521 13998 10577
rect 13350 10461 13430 10463
rect 13350 10405 13362 10461
rect 13418 10405 13430 10461
rect 13350 10403 13430 10405
rect 13362 10321 13418 10403
rect 12982 10311 13062 10321
rect 12982 10255 12994 10311
rect 13050 10255 13062 10311
rect 12982 10245 13062 10255
rect 13166 10311 13246 10321
rect 13166 10255 13178 10311
rect 13234 10255 13246 10311
rect 13166 10245 13246 10255
rect 13350 10311 13430 10321
rect 13350 10255 13362 10311
rect 13418 10255 13430 10311
rect 13350 10245 13430 10255
rect 13495 10189 13563 10519
rect 13938 10509 13998 10521
rect 15370 10461 15440 10473
rect 15370 10405 15382 10461
rect 15438 10405 15440 10461
rect 15370 10393 15440 10405
rect 13454 10181 13563 10189
rect 13442 10179 13563 10181
rect 13442 10059 13454 10179
rect 13510 10059 13563 10179
rect 13442 10057 13563 10059
rect 13454 10049 13510 10057
rect 12757 9792 13655 9804
rect 12757 9736 12769 9792
rect 12825 9736 13587 9792
rect 13643 9736 13655 9792
rect 12757 9724 13655 9736
rect 11872 9618 11884 9674
rect 11940 9618 11942 9674
rect 11872 9616 11942 9618
rect 12184 9674 12244 9678
rect 12184 9618 12186 9674
rect 12242 9618 12244 9674
rect 11884 9004 11940 9616
rect 12184 9606 12244 9618
rect 15382 9514 15438 10393
rect 15382 9404 15438 9414
rect 11736 4509 11806 4521
rect 11736 4453 11748 4509
rect 11804 4453 11806 4509
rect 11736 4441 11806 4453
rect 11382 3151 11384 3207
rect 11440 3151 11668 3207
rect 10794 3091 10874 3093
rect 10794 3035 10806 3091
rect 10862 3035 10874 3091
rect 10794 3033 10874 3035
rect 10806 2951 10862 3033
rect 10426 2941 10506 2951
rect 10426 2885 10438 2941
rect 10494 2885 10506 2941
rect 10426 2875 10506 2885
rect 10610 2941 10690 2951
rect 10610 2885 10622 2941
rect 10678 2885 10690 2941
rect 10610 2875 10690 2885
rect 10794 2941 10874 2951
rect 10794 2885 10806 2941
rect 10862 2885 10874 2941
rect 10794 2875 10874 2885
rect 10939 2819 11007 3149
rect 11382 3139 11452 3151
rect 10898 2811 11007 2819
rect 10886 2809 11007 2811
rect 10886 2689 10898 2809
rect 10954 2689 11007 2809
rect 10886 2687 11007 2689
rect 10898 2679 10954 2687
rect 10201 2422 11097 2434
rect 10201 2366 10213 2422
rect 10269 2366 11031 2422
rect 11087 2366 11097 2422
rect 10201 2354 11097 2366
rect 9886 2303 9966 2313
rect 9886 2247 9898 2303
rect 9954 2247 9966 2303
rect 9886 2245 9966 2247
rect 9720 2193 9790 2196
rect 9720 2139 9722 2193
rect 9778 2139 9790 2193
rect 9720 2127 9790 2139
rect 8860 2086 9606 2098
rect 8860 2030 9228 2086
rect 9284 2030 9606 2086
rect 8860 2018 9606 2030
rect 8860 1765 8916 2018
rect 9228 1765 9284 2018
rect 9550 1765 9606 2018
rect 8848 1763 8928 1765
rect 8848 1643 8860 1763
rect 8916 1643 8928 1763
rect 8848 1641 8928 1643
rect 9216 1763 9296 1765
rect 9216 1643 9228 1763
rect 9284 1643 9296 1763
rect 9216 1641 9296 1643
rect 9538 1763 9618 1765
rect 9538 1642 9550 1763
rect 9606 1642 9618 1763
rect 8860 1633 8916 1641
rect 9228 1633 9284 1641
rect 9538 1640 9618 1642
rect 9550 1632 9606 1640
rect 9044 1465 9100 1473
rect 9412 1465 9468 1473
rect 9032 1463 9521 1465
rect 9032 1343 9044 1463
rect 9100 1343 9412 1463
rect 9468 1343 9521 1463
rect 9032 1341 9521 1343
rect 9044 1333 9100 1341
rect 9412 1333 9521 1341
rect 8940 1267 9020 1277
rect 8940 1211 8952 1267
rect 9008 1211 9020 1267
rect 8940 1201 9020 1211
rect 9124 1267 9204 1277
rect 9124 1211 9136 1267
rect 9192 1211 9204 1267
rect 9124 1201 9204 1211
rect 9308 1267 9388 1277
rect 9308 1211 9320 1267
rect 9376 1211 9388 1267
rect 9308 1201 9388 1211
rect 8952 1119 9008 1201
rect 8940 1117 9020 1119
rect 8940 1061 8952 1117
rect 9008 1061 9020 1117
rect 8940 1059 9020 1061
rect 8132 1001 8202 1015
rect 8132 945 8144 1001
rect 8200 945 8202 1001
rect 8132 933 8202 945
rect 7966 885 8046 897
rect 7966 829 7978 885
rect 8034 829 8046 885
rect 7966 817 8046 829
rect 7830 98 7900 110
rect 8144 102 8200 933
rect 8952 745 9008 1059
rect 9136 1003 9192 1201
rect 9124 1001 9204 1003
rect 9124 945 9136 1001
rect 9192 945 9204 1001
rect 9124 943 9204 945
rect 9136 745 9192 943
rect 9320 887 9376 1201
rect 9453 1003 9521 1333
rect 9898 1013 9954 2245
rect 9453 1001 9533 1003
rect 9453 945 9465 1001
rect 9521 945 9533 1001
rect 9453 943 9533 945
rect 9896 1001 9956 1013
rect 9896 945 9898 1001
rect 9954 945 9956 1001
rect 9308 885 9388 887
rect 9308 829 9320 885
rect 9376 829 9388 885
rect 9308 827 9388 829
rect 9320 745 9376 827
rect 8940 735 9020 745
rect 8940 679 8952 735
rect 9008 679 9020 735
rect 8940 669 9020 679
rect 9124 735 9204 745
rect 9124 679 9136 735
rect 9192 679 9204 735
rect 9124 669 9204 679
rect 9308 735 9388 745
rect 9308 679 9320 735
rect 9376 679 9388 735
rect 9308 669 9388 679
rect 9453 613 9521 943
rect 9896 933 9956 945
rect 9412 605 9521 613
rect 9400 603 9521 605
rect 9400 483 9412 603
rect 9468 483 9521 603
rect 9400 481 9521 483
rect 9412 473 9468 481
rect 8715 216 9613 228
rect 8715 160 8727 216
rect 8783 160 9545 216
rect 9601 160 9613 216
rect 8715 148 9613 160
rect 7830 42 7842 98
rect 7898 42 7900 98
rect 7830 30 7900 42
rect 8142 98 8202 102
rect 8142 42 8144 98
rect 8200 42 8202 98
rect 8142 30 8202 42
rect 7706 -175 7762 -165
rect 11748 -65 11804 4441
rect 11884 110 11940 8904
rect 12902 8701 13648 8713
rect 12902 8645 13270 8701
rect 13326 8645 13648 8701
rect 12902 8633 13648 8645
rect 12902 8380 12958 8633
rect 13270 8380 13326 8633
rect 13592 8380 13648 8633
rect 12890 8378 12970 8380
rect 12890 8258 12902 8378
rect 12958 8258 12970 8378
rect 12890 8256 12970 8258
rect 13258 8378 13338 8380
rect 13258 8258 13270 8378
rect 13326 8258 13338 8378
rect 13258 8256 13338 8258
rect 13580 8378 13660 8380
rect 13580 8257 13592 8378
rect 13648 8257 13660 8378
rect 12902 8248 12958 8256
rect 13270 8248 13326 8256
rect 13580 8255 13660 8257
rect 13592 8247 13648 8255
rect 13086 8080 13142 8088
rect 13454 8080 13510 8088
rect 13074 8078 13563 8080
rect 13074 7958 13086 8078
rect 13142 7958 13454 8078
rect 13510 7958 13563 8078
rect 13074 7956 13563 7958
rect 13086 7948 13142 7956
rect 13454 7948 13563 7956
rect 12982 7882 13062 7892
rect 12982 7826 12994 7882
rect 13050 7826 13062 7882
rect 12982 7816 13062 7826
rect 13166 7882 13246 7892
rect 13166 7826 13178 7882
rect 13234 7826 13246 7882
rect 13166 7816 13246 7826
rect 13350 7882 13430 7892
rect 13350 7826 13362 7882
rect 13418 7826 13430 7882
rect 13350 7816 13430 7826
rect 12094 7732 12180 7744
rect 12994 7734 13050 7816
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 12982 7732 13062 7734
rect 12982 7676 12994 7732
rect 13050 7676 13062 7732
rect 12982 7674 13062 7676
rect 12310 7616 12380 7628
rect 12310 7560 12322 7616
rect 12378 7560 12380 7616
rect 12310 7548 12380 7560
rect 12174 5411 12244 5425
rect 12174 5355 12186 5411
rect 12242 5355 12244 5411
rect 12174 5343 12244 5355
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 12020 897 12076 5165
rect 12186 1015 12242 5343
rect 12322 3102 12378 7548
rect 12994 7360 13050 7674
rect 13178 7618 13234 7816
rect 13166 7616 13246 7618
rect 13166 7560 13178 7616
rect 13234 7560 13246 7616
rect 13166 7558 13246 7560
rect 13178 7360 13234 7558
rect 13362 7502 13418 7816
rect 13495 7618 13563 7948
rect 13495 7616 13575 7618
rect 13495 7560 13507 7616
rect 13563 7560 13575 7616
rect 13495 7558 13575 7560
rect 13762 7616 13832 7628
rect 13762 7560 13764 7616
rect 13820 7560 13832 7616
rect 13350 7500 13430 7502
rect 13350 7444 13362 7500
rect 13418 7444 13430 7500
rect 13350 7442 13430 7444
rect 13362 7360 13418 7442
rect 12982 7350 13062 7360
rect 12982 7294 12994 7350
rect 13050 7294 13062 7350
rect 12982 7284 13062 7294
rect 13166 7350 13246 7360
rect 13166 7294 13178 7350
rect 13234 7294 13246 7350
rect 13166 7284 13246 7294
rect 13350 7350 13430 7360
rect 13350 7294 13362 7350
rect 13418 7294 13430 7350
rect 13350 7284 13430 7294
rect 13495 7228 13563 7558
rect 13762 7550 13832 7560
rect 13454 7220 13563 7228
rect 13442 7218 13563 7220
rect 13442 7098 13454 7218
rect 13510 7098 13563 7218
rect 13442 7096 13563 7098
rect 13454 7088 13510 7096
rect 12757 6831 13655 6843
rect 12757 6775 12769 6831
rect 12825 6775 13587 6831
rect 13643 6775 13655 6831
rect 12757 6763 13655 6775
rect 13764 6606 13820 7550
rect 13928 6713 14008 6723
rect 13928 6657 13940 6713
rect 13996 6657 14008 6713
rect 13928 6655 14008 6657
rect 13762 6603 13832 6606
rect 13762 6549 13764 6603
rect 13820 6549 13832 6603
rect 13762 6537 13832 6549
rect 12902 6496 13648 6508
rect 12902 6440 13270 6496
rect 13326 6440 13648 6496
rect 12902 6428 13648 6440
rect 12902 6175 12958 6428
rect 13270 6175 13326 6428
rect 13592 6175 13648 6428
rect 12890 6173 12970 6175
rect 12890 6053 12902 6173
rect 12958 6053 12970 6173
rect 12890 6051 12970 6053
rect 13258 6173 13338 6175
rect 13258 6053 13270 6173
rect 13326 6053 13338 6173
rect 13258 6051 13338 6053
rect 13580 6173 13660 6175
rect 13580 6052 13592 6173
rect 13648 6052 13660 6173
rect 12902 6043 12958 6051
rect 13270 6043 13326 6051
rect 13580 6050 13660 6052
rect 13592 6042 13648 6050
rect 13086 5875 13142 5883
rect 13454 5875 13510 5883
rect 13074 5873 13563 5875
rect 13074 5753 13086 5873
rect 13142 5753 13454 5873
rect 13510 5753 13563 5873
rect 13074 5751 13563 5753
rect 13086 5743 13142 5751
rect 13454 5743 13563 5751
rect 12982 5677 13062 5687
rect 12982 5621 12994 5677
rect 13050 5621 13062 5677
rect 12982 5611 13062 5621
rect 13166 5677 13246 5687
rect 13166 5621 13178 5677
rect 13234 5621 13246 5677
rect 13166 5611 13246 5621
rect 13350 5677 13430 5687
rect 13350 5621 13362 5677
rect 13418 5621 13430 5677
rect 13350 5611 13430 5621
rect 12994 5529 13050 5611
rect 12982 5527 13062 5529
rect 12982 5471 12994 5527
rect 13050 5471 13062 5527
rect 12982 5469 13062 5471
rect 12994 5155 13050 5469
rect 13178 5413 13234 5611
rect 13166 5411 13246 5413
rect 13166 5355 13178 5411
rect 13234 5355 13246 5411
rect 13166 5353 13246 5355
rect 13178 5155 13234 5353
rect 13362 5297 13418 5611
rect 13495 5413 13563 5743
rect 13940 5421 13996 6655
rect 14388 6496 15134 6508
rect 14388 6440 14756 6496
rect 14812 6440 15134 6496
rect 14388 6428 15134 6440
rect 14388 6175 14444 6428
rect 14756 6175 14812 6428
rect 15078 6175 15134 6428
rect 14376 6173 14456 6175
rect 14376 6053 14388 6173
rect 14444 6053 14456 6173
rect 14376 6051 14456 6053
rect 14744 6173 14824 6175
rect 14744 6053 14756 6173
rect 14812 6053 14824 6173
rect 14744 6051 14824 6053
rect 15066 6173 15146 6175
rect 15066 6052 15078 6173
rect 15134 6052 15146 6173
rect 14388 6043 14444 6051
rect 14756 6043 14812 6051
rect 15066 6050 15146 6052
rect 15078 6042 15134 6050
rect 14572 5875 14628 5883
rect 14940 5875 14996 5883
rect 14560 5873 15049 5875
rect 14560 5753 14572 5873
rect 14628 5753 14940 5873
rect 14996 5753 15049 5873
rect 14560 5751 15049 5753
rect 14572 5743 14628 5751
rect 14940 5743 15049 5751
rect 14468 5677 14548 5687
rect 14468 5621 14480 5677
rect 14536 5621 14548 5677
rect 14468 5611 14548 5621
rect 14652 5677 14732 5687
rect 14652 5621 14664 5677
rect 14720 5621 14732 5677
rect 14652 5611 14732 5621
rect 14836 5677 14916 5687
rect 14836 5621 14848 5677
rect 14904 5621 14916 5677
rect 14836 5611 14916 5621
rect 14480 5529 14536 5611
rect 14468 5527 14548 5529
rect 14468 5471 14480 5527
rect 14536 5471 14548 5527
rect 14468 5469 14548 5471
rect 13495 5411 13575 5413
rect 13495 5355 13507 5411
rect 13563 5355 13575 5411
rect 13495 5353 13575 5355
rect 13938 5411 13998 5421
rect 13938 5355 13940 5411
rect 13996 5355 13998 5411
rect 13350 5295 13430 5297
rect 13350 5239 13362 5295
rect 13418 5239 13430 5295
rect 13350 5237 13430 5239
rect 13362 5155 13418 5237
rect 12982 5145 13062 5155
rect 12982 5089 12994 5145
rect 13050 5089 13062 5145
rect 12982 5079 13062 5089
rect 13166 5145 13246 5155
rect 13166 5089 13178 5145
rect 13234 5089 13246 5145
rect 13166 5079 13246 5089
rect 13350 5145 13430 5155
rect 13350 5089 13362 5145
rect 13418 5089 13430 5145
rect 13350 5079 13430 5089
rect 13495 5023 13563 5353
rect 13938 5343 13998 5355
rect 13454 5015 13563 5023
rect 13442 5013 13563 5015
rect 13442 4893 13454 5013
rect 13510 4893 13563 5013
rect 13442 4891 13563 4893
rect 13454 4883 13510 4891
rect 12757 4626 13653 4638
rect 12757 4570 12769 4626
rect 12825 4570 13587 4626
rect 13643 4570 13653 4626
rect 12757 4558 13653 4570
rect 13940 4400 13996 5343
rect 14480 5155 14536 5469
rect 14664 5413 14720 5611
rect 14652 5411 14732 5413
rect 14652 5355 14664 5411
rect 14720 5355 14732 5411
rect 14652 5353 14732 5355
rect 14664 5155 14720 5353
rect 14848 5297 14904 5611
rect 14981 5413 15049 5743
rect 14981 5411 15061 5413
rect 14981 5355 14993 5411
rect 15049 5355 15061 5411
rect 14981 5353 15061 5355
rect 15248 5411 15318 5423
rect 15248 5355 15250 5411
rect 15306 5355 15574 5411
rect 14836 5295 14916 5297
rect 14836 5239 14848 5295
rect 14904 5239 14916 5295
rect 14836 5237 14916 5239
rect 14848 5155 14904 5237
rect 14468 5145 14548 5155
rect 14468 5089 14480 5145
rect 14536 5089 14548 5145
rect 14468 5079 14548 5089
rect 14652 5145 14732 5155
rect 14652 5089 14664 5145
rect 14720 5089 14732 5145
rect 14652 5079 14732 5089
rect 14836 5145 14916 5155
rect 14836 5089 14848 5145
rect 14904 5089 14916 5145
rect 14836 5079 14916 5089
rect 14981 5023 15049 5353
rect 15248 5345 15318 5355
rect 14940 5015 15049 5023
rect 14928 5013 15049 5015
rect 14928 4893 14940 5013
rect 14996 4893 15049 5013
rect 14928 4891 15049 4893
rect 14940 4883 14996 4891
rect 14243 4626 15139 4638
rect 14243 4570 14255 4626
rect 14311 4570 15073 4626
rect 15129 4570 15139 4626
rect 14243 4558 15139 4570
rect 15250 4401 15306 5345
rect 15414 4509 15494 4519
rect 15414 4453 15426 4509
rect 15482 4453 15494 4509
rect 15414 4451 15494 4453
rect 13938 4398 14008 4400
rect 13938 4342 13940 4398
rect 13996 4342 14008 4398
rect 13938 4330 14008 4342
rect 15238 4399 15318 4401
rect 15238 4343 15250 4399
rect 15306 4343 15318 4399
rect 15238 4331 15318 4343
rect 12902 4291 13648 4303
rect 12902 4235 13270 4291
rect 13326 4235 13648 4291
rect 12902 4223 13648 4235
rect 12902 3970 12958 4223
rect 13270 3970 13326 4223
rect 13592 3970 13648 4223
rect 14388 4292 15134 4304
rect 14388 4236 14756 4292
rect 14812 4236 15134 4292
rect 14388 4224 15134 4236
rect 14388 3971 14444 4224
rect 14756 3971 14812 4224
rect 15078 3971 15134 4224
rect 12890 3968 12970 3970
rect 12890 3848 12902 3968
rect 12958 3848 12970 3968
rect 12890 3846 12970 3848
rect 13258 3968 13338 3970
rect 13258 3848 13270 3968
rect 13326 3848 13338 3968
rect 13258 3846 13338 3848
rect 13580 3968 13660 3970
rect 13580 3847 13592 3968
rect 13648 3847 13660 3968
rect 14376 3969 14456 3971
rect 14376 3849 14388 3969
rect 14444 3849 14456 3969
rect 14376 3847 14456 3849
rect 14744 3969 14824 3971
rect 14744 3849 14756 3969
rect 14812 3849 14824 3969
rect 14744 3847 14824 3849
rect 15066 3969 15146 3971
rect 15066 3848 15078 3969
rect 15134 3848 15146 3969
rect 12902 3838 12958 3846
rect 13270 3838 13326 3846
rect 13580 3845 13660 3847
rect 13592 3837 13648 3845
rect 14388 3839 14444 3847
rect 14756 3839 14812 3847
rect 15066 3846 15146 3848
rect 15078 3838 15134 3846
rect 13086 3670 13142 3678
rect 13454 3670 13510 3678
rect 14572 3671 14628 3679
rect 14940 3671 14996 3679
rect 13074 3668 13563 3670
rect 13074 3548 13086 3668
rect 13142 3548 13454 3668
rect 13510 3548 13563 3668
rect 13074 3546 13563 3548
rect 14560 3669 15049 3671
rect 14560 3549 14572 3669
rect 14628 3549 14940 3669
rect 14996 3549 15049 3669
rect 14560 3547 15049 3549
rect 13086 3538 13142 3546
rect 13454 3538 13563 3546
rect 14572 3539 14628 3547
rect 14940 3539 15049 3547
rect 12982 3472 13062 3482
rect 12982 3416 12994 3472
rect 13050 3416 13062 3472
rect 12982 3406 13062 3416
rect 13166 3472 13246 3482
rect 13166 3416 13178 3472
rect 13234 3416 13246 3472
rect 13166 3406 13246 3416
rect 13350 3472 13430 3482
rect 13350 3416 13362 3472
rect 13418 3416 13430 3472
rect 13350 3406 13430 3416
rect 12994 3324 13050 3406
rect 12982 3322 13062 3324
rect 12982 3266 12994 3322
rect 13050 3266 13062 3322
rect 12982 3264 13062 3266
rect 12310 3090 12380 3102
rect 12310 3034 12322 3090
rect 12378 3034 12380 3090
rect 12310 3022 12380 3034
rect 12994 2950 13050 3264
rect 13178 3208 13234 3406
rect 13166 3206 13246 3208
rect 13166 3150 13178 3206
rect 13234 3150 13246 3206
rect 13166 3148 13246 3150
rect 13178 2950 13234 3148
rect 13362 3092 13418 3406
rect 13495 3208 13563 3538
rect 14468 3473 14548 3483
rect 14468 3417 14480 3473
rect 14536 3417 14548 3473
rect 14468 3407 14548 3417
rect 14652 3473 14732 3483
rect 14652 3417 14664 3473
rect 14720 3417 14732 3473
rect 14652 3407 14732 3417
rect 14836 3473 14916 3483
rect 14836 3417 14848 3473
rect 14904 3417 14916 3473
rect 14836 3407 14916 3417
rect 14480 3325 14536 3407
rect 14468 3323 14548 3325
rect 14468 3267 14480 3323
rect 14536 3267 14548 3323
rect 14468 3265 14548 3267
rect 13495 3206 13575 3208
rect 13495 3150 13507 3206
rect 13563 3150 13575 3206
rect 13495 3148 13575 3150
rect 13762 3206 13832 3218
rect 13762 3150 13764 3206
rect 13820 3150 13832 3206
rect 13350 3090 13430 3092
rect 13350 3034 13362 3090
rect 13418 3034 13430 3090
rect 13350 3032 13430 3034
rect 13362 2950 13418 3032
rect 12982 2940 13062 2950
rect 12982 2884 12994 2940
rect 13050 2884 13062 2940
rect 12982 2874 13062 2884
rect 13166 2940 13246 2950
rect 13166 2884 13178 2940
rect 13234 2884 13246 2940
rect 13166 2874 13246 2884
rect 13350 2940 13430 2950
rect 13350 2884 13362 2940
rect 13418 2884 13430 2940
rect 13350 2874 13430 2884
rect 13495 2818 13563 3148
rect 13762 3140 13832 3150
rect 13454 2810 13563 2818
rect 13442 2808 13563 2810
rect 13442 2688 13454 2808
rect 13510 2688 13563 2808
rect 13442 2686 13563 2688
rect 13454 2678 13510 2686
rect 12757 2421 13653 2433
rect 12757 2365 12769 2421
rect 12825 2365 13587 2421
rect 13643 2365 13653 2421
rect 12757 2353 13653 2365
rect 13764 2196 13820 3140
rect 14480 2951 14536 3265
rect 14664 3209 14720 3407
rect 14652 3207 14732 3209
rect 14652 3151 14664 3207
rect 14720 3151 14732 3207
rect 14652 3149 14732 3151
rect 14664 2951 14720 3149
rect 14848 3093 14904 3407
rect 14981 3209 15049 3539
rect 15426 3217 15482 4451
rect 14981 3207 15061 3209
rect 14981 3151 14993 3207
rect 15049 3151 15061 3207
rect 14981 3149 15061 3151
rect 15424 3207 15494 3217
rect 15654 3207 15710 17250
rect 15856 14999 15912 18503
rect 15854 14987 15924 14999
rect 15854 14931 15856 14987
rect 15912 14931 15924 14987
rect 15854 14919 15924 14931
rect 16092 14087 16148 18855
rect 16944 18277 17690 18289
rect 16944 18221 17312 18277
rect 17368 18221 17690 18277
rect 16944 18209 17690 18221
rect 16944 17956 17000 18209
rect 17312 17956 17368 18209
rect 17634 17956 17690 18209
rect 16932 17954 17012 17956
rect 16932 17834 16944 17954
rect 17000 17834 17012 17954
rect 16932 17832 17012 17834
rect 17300 17954 17380 17956
rect 17300 17834 17312 17954
rect 17368 17834 17380 17954
rect 17300 17832 17380 17834
rect 17622 17954 17702 17956
rect 17622 17833 17634 17954
rect 17690 17833 17702 17954
rect 16944 17824 17000 17832
rect 17312 17824 17368 17832
rect 17622 17831 17702 17833
rect 17634 17823 17690 17831
rect 17128 17656 17184 17664
rect 17496 17656 17552 17664
rect 17116 17654 17605 17656
rect 17116 17534 17128 17654
rect 17184 17534 17496 17654
rect 17552 17534 17605 17654
rect 17116 17532 17605 17534
rect 17128 17524 17184 17532
rect 17496 17524 17605 17532
rect 17024 17458 17104 17468
rect 17024 17402 17036 17458
rect 17092 17402 17104 17458
rect 17024 17392 17104 17402
rect 17208 17458 17288 17468
rect 17208 17402 17220 17458
rect 17276 17402 17288 17458
rect 17208 17392 17288 17402
rect 17392 17458 17472 17468
rect 17392 17402 17404 17458
rect 17460 17402 17472 17458
rect 17392 17392 17472 17402
rect 17036 17310 17092 17392
rect 17024 17308 17104 17310
rect 17024 17252 17036 17308
rect 17092 17252 17104 17308
rect 17024 17250 17104 17252
rect 16352 17192 16422 17204
rect 16352 17136 16364 17192
rect 16420 17136 16422 17192
rect 16352 17124 16422 17136
rect 16216 14987 16286 15001
rect 16216 14931 16228 14987
rect 16284 14931 16286 14987
rect 16216 14919 16286 14931
rect 16080 14085 16150 14087
rect 16080 14029 16092 14085
rect 16148 14029 16150 14085
rect 16080 14017 16150 14029
rect 16228 10591 16284 14919
rect 16364 12678 16420 17124
rect 17036 16936 17092 17250
rect 17220 17194 17276 17392
rect 17208 17192 17288 17194
rect 17208 17136 17220 17192
rect 17276 17136 17288 17192
rect 17208 17134 17288 17136
rect 17220 16936 17276 17134
rect 17404 17078 17460 17392
rect 17537 17194 17605 17524
rect 19684 17308 19754 17320
rect 19684 17252 19696 17308
rect 19752 17252 19754 17308
rect 19684 17250 19754 17252
rect 17537 17192 17617 17194
rect 17537 17136 17549 17192
rect 17605 17136 17617 17192
rect 17537 17134 17617 17136
rect 17804 17192 17874 17204
rect 17804 17136 17806 17192
rect 17862 17136 17874 17192
rect 17392 17076 17472 17078
rect 17392 17020 17404 17076
rect 17460 17020 17472 17076
rect 17392 17018 17472 17020
rect 17404 16936 17460 17018
rect 17024 16926 17104 16936
rect 17024 16870 17036 16926
rect 17092 16870 17104 16926
rect 17024 16860 17104 16870
rect 17208 16926 17288 16936
rect 17208 16870 17220 16926
rect 17276 16870 17288 16926
rect 17208 16860 17288 16870
rect 17392 16926 17472 16936
rect 17392 16870 17404 16926
rect 17460 16870 17472 16926
rect 17392 16860 17472 16870
rect 17537 16804 17605 17134
rect 17804 17126 17874 17136
rect 17496 16796 17605 16804
rect 17484 16794 17605 16796
rect 17484 16674 17496 16794
rect 17552 16674 17605 16794
rect 17484 16672 17605 16674
rect 17496 16664 17552 16672
rect 16799 16407 17697 16419
rect 16799 16351 16811 16407
rect 16867 16351 17629 16407
rect 17685 16351 17697 16407
rect 16799 16339 17697 16351
rect 17806 16182 17862 17126
rect 17970 16289 18050 16299
rect 17970 16233 17982 16289
rect 18038 16233 18050 16289
rect 17970 16231 18050 16233
rect 17804 16179 17874 16182
rect 17804 16125 17806 16179
rect 17862 16125 17874 16179
rect 17804 16113 17874 16125
rect 16944 16072 17690 16084
rect 16944 16016 17312 16072
rect 17368 16016 17690 16072
rect 16944 16004 17690 16016
rect 16944 15751 17000 16004
rect 17312 15751 17368 16004
rect 17634 15751 17690 16004
rect 16932 15749 17012 15751
rect 16932 15629 16944 15749
rect 17000 15629 17012 15749
rect 16932 15627 17012 15629
rect 17300 15749 17380 15751
rect 17300 15629 17312 15749
rect 17368 15629 17380 15749
rect 17300 15627 17380 15629
rect 17622 15749 17702 15751
rect 17622 15628 17634 15749
rect 17690 15628 17702 15749
rect 16944 15619 17000 15627
rect 17312 15619 17368 15627
rect 17622 15626 17702 15628
rect 17634 15618 17690 15626
rect 17128 15451 17184 15459
rect 17496 15451 17552 15459
rect 17116 15449 17605 15451
rect 17116 15329 17128 15449
rect 17184 15329 17496 15449
rect 17552 15329 17605 15449
rect 17116 15327 17605 15329
rect 17128 15319 17184 15327
rect 17496 15319 17605 15327
rect 17024 15253 17104 15263
rect 17024 15197 17036 15253
rect 17092 15197 17104 15253
rect 17024 15187 17104 15197
rect 17208 15253 17288 15263
rect 17208 15197 17220 15253
rect 17276 15197 17288 15253
rect 17208 15187 17288 15197
rect 17392 15253 17472 15263
rect 17392 15197 17404 15253
rect 17460 15197 17472 15253
rect 17392 15187 17472 15197
rect 17036 15105 17092 15187
rect 17024 15103 17104 15105
rect 17024 15047 17036 15103
rect 17092 15047 17104 15103
rect 17024 15045 17104 15047
rect 17036 14731 17092 15045
rect 17220 14989 17276 15187
rect 17208 14987 17288 14989
rect 17208 14931 17220 14987
rect 17276 14931 17288 14987
rect 17208 14929 17288 14931
rect 17220 14731 17276 14929
rect 17404 14873 17460 15187
rect 17537 14989 17605 15319
rect 17982 14997 18038 16231
rect 18430 16072 19176 16084
rect 18430 16016 18798 16072
rect 18854 16016 19176 16072
rect 18430 16004 19176 16016
rect 18430 15751 18486 16004
rect 18798 15751 18854 16004
rect 19120 15751 19176 16004
rect 18418 15749 18498 15751
rect 18418 15629 18430 15749
rect 18486 15629 18498 15749
rect 18418 15627 18498 15629
rect 18786 15749 18866 15751
rect 18786 15629 18798 15749
rect 18854 15629 18866 15749
rect 18786 15627 18866 15629
rect 19108 15749 19188 15751
rect 19108 15628 19120 15749
rect 19176 15628 19188 15749
rect 18430 15619 18486 15627
rect 18798 15619 18854 15627
rect 19108 15626 19188 15628
rect 19120 15618 19176 15626
rect 18614 15451 18670 15459
rect 18982 15451 19038 15459
rect 18602 15449 19091 15451
rect 18602 15329 18614 15449
rect 18670 15329 18982 15449
rect 19038 15329 19091 15449
rect 18602 15327 19091 15329
rect 18614 15319 18670 15327
rect 18982 15319 19091 15327
rect 18510 15253 18590 15263
rect 18510 15197 18522 15253
rect 18578 15197 18590 15253
rect 18510 15187 18590 15197
rect 18694 15253 18774 15263
rect 18694 15197 18706 15253
rect 18762 15197 18774 15253
rect 18694 15187 18774 15197
rect 18878 15253 18958 15263
rect 18878 15197 18890 15253
rect 18946 15197 18958 15253
rect 18878 15187 18958 15197
rect 18522 15105 18578 15187
rect 18510 15103 18590 15105
rect 18510 15047 18522 15103
rect 18578 15047 18590 15103
rect 18510 15045 18590 15047
rect 17537 14987 17617 14989
rect 17537 14931 17549 14987
rect 17605 14931 17617 14987
rect 17537 14929 17617 14931
rect 17980 14987 18040 14997
rect 17980 14931 17982 14987
rect 18038 14931 18040 14987
rect 17392 14871 17472 14873
rect 17392 14815 17404 14871
rect 17460 14815 17472 14871
rect 17392 14813 17472 14815
rect 17404 14731 17460 14813
rect 17024 14721 17104 14731
rect 17024 14665 17036 14721
rect 17092 14665 17104 14721
rect 17024 14655 17104 14665
rect 17208 14721 17288 14731
rect 17208 14665 17220 14721
rect 17276 14665 17288 14721
rect 17208 14655 17288 14665
rect 17392 14721 17472 14731
rect 17392 14665 17404 14721
rect 17460 14665 17472 14721
rect 17392 14655 17472 14665
rect 17537 14599 17605 14929
rect 17980 14919 18040 14931
rect 17496 14591 17605 14599
rect 17484 14589 17605 14591
rect 17484 14469 17496 14589
rect 17552 14469 17605 14589
rect 17484 14467 17605 14469
rect 17496 14459 17552 14467
rect 16799 14202 17695 14214
rect 16799 14146 16811 14202
rect 16867 14146 17629 14202
rect 17685 14146 17695 14202
rect 16799 14134 17695 14146
rect 17982 13976 18038 14919
rect 18522 14731 18578 15045
rect 18706 14989 18762 15187
rect 18694 14987 18774 14989
rect 18694 14931 18706 14987
rect 18762 14931 18774 14987
rect 18694 14929 18774 14931
rect 18706 14731 18762 14929
rect 18890 14873 18946 15187
rect 19023 14989 19091 15319
rect 19023 14987 19103 14989
rect 19023 14931 19035 14987
rect 19091 14931 19103 14987
rect 19023 14929 19103 14931
rect 19290 14987 19360 14999
rect 19290 14931 19292 14987
rect 19348 14931 19616 14987
rect 18878 14871 18958 14873
rect 18878 14815 18890 14871
rect 18946 14815 18958 14871
rect 18878 14813 18958 14815
rect 18890 14731 18946 14813
rect 18510 14721 18590 14731
rect 18510 14665 18522 14721
rect 18578 14665 18590 14721
rect 18510 14655 18590 14665
rect 18694 14721 18774 14731
rect 18694 14665 18706 14721
rect 18762 14665 18774 14721
rect 18694 14655 18774 14665
rect 18878 14721 18958 14731
rect 18878 14665 18890 14721
rect 18946 14665 18958 14721
rect 18878 14655 18958 14665
rect 19023 14599 19091 14929
rect 19290 14921 19360 14931
rect 18982 14591 19091 14599
rect 18970 14589 19091 14591
rect 18970 14469 18982 14589
rect 19038 14469 19091 14589
rect 18970 14467 19091 14469
rect 18982 14459 19038 14467
rect 18285 14202 19181 14214
rect 18285 14146 18297 14202
rect 18353 14146 19115 14202
rect 19171 14146 19181 14202
rect 18285 14134 19181 14146
rect 19292 13977 19348 14921
rect 19456 14085 19536 14095
rect 19456 14029 19468 14085
rect 19524 14029 19536 14085
rect 19456 14027 19536 14029
rect 17980 13974 18050 13976
rect 17980 13918 17982 13974
rect 18038 13918 18050 13974
rect 17980 13906 18050 13918
rect 19280 13975 19360 13977
rect 19280 13919 19292 13975
rect 19348 13919 19360 13975
rect 19280 13907 19360 13919
rect 16944 13867 17690 13879
rect 16944 13811 17312 13867
rect 17368 13811 17690 13867
rect 16944 13799 17690 13811
rect 16944 13546 17000 13799
rect 17312 13546 17368 13799
rect 17634 13546 17690 13799
rect 18430 13868 19176 13880
rect 18430 13812 18798 13868
rect 18854 13812 19176 13868
rect 18430 13800 19176 13812
rect 18430 13547 18486 13800
rect 18798 13547 18854 13800
rect 19120 13547 19176 13800
rect 16932 13544 17012 13546
rect 16932 13424 16944 13544
rect 17000 13424 17012 13544
rect 16932 13422 17012 13424
rect 17300 13544 17380 13546
rect 17300 13424 17312 13544
rect 17368 13424 17380 13544
rect 17300 13422 17380 13424
rect 17622 13544 17702 13546
rect 17622 13423 17634 13544
rect 17690 13423 17702 13544
rect 18418 13545 18498 13547
rect 18418 13425 18430 13545
rect 18486 13425 18498 13545
rect 18418 13423 18498 13425
rect 18786 13545 18866 13547
rect 18786 13425 18798 13545
rect 18854 13425 18866 13545
rect 18786 13423 18866 13425
rect 19108 13545 19188 13547
rect 19108 13424 19120 13545
rect 19176 13424 19188 13545
rect 16944 13414 17000 13422
rect 17312 13414 17368 13422
rect 17622 13421 17702 13423
rect 17634 13413 17690 13421
rect 18430 13415 18486 13423
rect 18798 13415 18854 13423
rect 19108 13422 19188 13424
rect 19120 13414 19176 13422
rect 17128 13246 17184 13254
rect 17496 13246 17552 13254
rect 18614 13247 18670 13255
rect 18982 13247 19038 13255
rect 17116 13244 17605 13246
rect 17116 13124 17128 13244
rect 17184 13124 17496 13244
rect 17552 13124 17605 13244
rect 17116 13122 17605 13124
rect 18602 13245 19091 13247
rect 18602 13125 18614 13245
rect 18670 13125 18982 13245
rect 19038 13125 19091 13245
rect 18602 13123 19091 13125
rect 17128 13114 17184 13122
rect 17496 13114 17605 13122
rect 18614 13115 18670 13123
rect 18982 13115 19091 13123
rect 17024 13048 17104 13058
rect 17024 12992 17036 13048
rect 17092 12992 17104 13048
rect 17024 12982 17104 12992
rect 17208 13048 17288 13058
rect 17208 12992 17220 13048
rect 17276 12992 17288 13048
rect 17208 12982 17288 12992
rect 17392 13048 17472 13058
rect 17392 12992 17404 13048
rect 17460 12992 17472 13048
rect 17392 12982 17472 12992
rect 17036 12900 17092 12982
rect 17024 12898 17104 12900
rect 17024 12842 17036 12898
rect 17092 12842 17104 12898
rect 17024 12840 17104 12842
rect 16352 12666 16422 12678
rect 16352 12610 16364 12666
rect 16420 12610 16422 12666
rect 16352 12598 16422 12610
rect 17036 12526 17092 12840
rect 17220 12784 17276 12982
rect 17208 12782 17288 12784
rect 17208 12726 17220 12782
rect 17276 12726 17288 12782
rect 17208 12724 17288 12726
rect 17220 12526 17276 12724
rect 17404 12668 17460 12982
rect 17537 12784 17605 13114
rect 18510 13049 18590 13059
rect 18510 12993 18522 13049
rect 18578 12993 18590 13049
rect 18510 12983 18590 12993
rect 18694 13049 18774 13059
rect 18694 12993 18706 13049
rect 18762 12993 18774 13049
rect 18694 12983 18774 12993
rect 18878 13049 18958 13059
rect 18878 12993 18890 13049
rect 18946 12993 18958 13049
rect 18878 12983 18958 12993
rect 18522 12901 18578 12983
rect 18510 12899 18590 12901
rect 18510 12843 18522 12899
rect 18578 12843 18590 12899
rect 18510 12841 18590 12843
rect 17537 12782 17617 12784
rect 17537 12726 17549 12782
rect 17605 12726 17617 12782
rect 17537 12724 17617 12726
rect 17804 12782 17874 12794
rect 17804 12726 17806 12782
rect 17862 12726 17874 12782
rect 17392 12666 17472 12668
rect 17392 12610 17404 12666
rect 17460 12610 17472 12666
rect 17392 12608 17472 12610
rect 17404 12526 17460 12608
rect 17024 12516 17104 12526
rect 17024 12460 17036 12516
rect 17092 12460 17104 12516
rect 17024 12450 17104 12460
rect 17208 12516 17288 12526
rect 17208 12460 17220 12516
rect 17276 12460 17288 12516
rect 17208 12450 17288 12460
rect 17392 12516 17472 12526
rect 17392 12460 17404 12516
rect 17460 12460 17472 12516
rect 17392 12450 17472 12460
rect 17537 12394 17605 12724
rect 17804 12716 17874 12726
rect 17496 12386 17605 12394
rect 17484 12384 17605 12386
rect 17484 12264 17496 12384
rect 17552 12264 17605 12384
rect 17484 12262 17605 12264
rect 17496 12254 17552 12262
rect 16799 11997 17695 12009
rect 16799 11941 16811 11997
rect 16867 11941 17629 11997
rect 17685 11941 17695 11997
rect 16799 11929 17695 11941
rect 17806 11772 17862 12716
rect 18522 12527 18578 12841
rect 18706 12785 18762 12983
rect 18694 12783 18774 12785
rect 18694 12727 18706 12783
rect 18762 12727 18774 12783
rect 18694 12725 18774 12727
rect 18706 12527 18762 12725
rect 18890 12669 18946 12983
rect 19023 12785 19091 13115
rect 19468 12793 19524 14027
rect 19023 12783 19103 12785
rect 19023 12727 19035 12783
rect 19091 12727 19103 12783
rect 19023 12725 19103 12727
rect 19466 12783 19536 12793
rect 19466 12727 19468 12783
rect 19524 12727 19616 12783
rect 18878 12667 18958 12669
rect 18878 12611 18890 12667
rect 18946 12611 18958 12667
rect 18878 12609 18958 12611
rect 18890 12527 18946 12609
rect 18510 12517 18590 12527
rect 18510 12461 18522 12517
rect 18578 12461 18590 12517
rect 18510 12451 18590 12461
rect 18694 12517 18774 12527
rect 18694 12461 18706 12517
rect 18762 12461 18774 12517
rect 18694 12451 18774 12461
rect 18878 12517 18958 12527
rect 18878 12461 18890 12517
rect 18946 12461 18958 12517
rect 18878 12451 18958 12461
rect 19023 12395 19091 12725
rect 19466 12715 19536 12727
rect 18982 12387 19091 12395
rect 18970 12385 19091 12387
rect 18970 12265 18982 12385
rect 19038 12265 19091 12385
rect 18970 12263 19091 12265
rect 18982 12255 19038 12263
rect 18285 11998 19181 12010
rect 18285 11942 18297 11998
rect 18353 11942 19115 11998
rect 19171 11942 19181 11998
rect 18285 11930 19181 11942
rect 17970 11879 18050 11889
rect 17970 11823 17982 11879
rect 18038 11823 18050 11879
rect 17970 11821 18050 11823
rect 17804 11769 17874 11772
rect 17804 11715 17806 11769
rect 17862 11715 17874 11769
rect 17804 11703 17874 11715
rect 16944 11662 17690 11674
rect 16944 11606 17312 11662
rect 17368 11606 17690 11662
rect 16944 11594 17690 11606
rect 16944 11341 17000 11594
rect 17312 11341 17368 11594
rect 17634 11341 17690 11594
rect 16932 11339 17012 11341
rect 16932 11219 16944 11339
rect 17000 11219 17012 11339
rect 16932 11217 17012 11219
rect 17300 11339 17380 11341
rect 17300 11219 17312 11339
rect 17368 11219 17380 11339
rect 17300 11217 17380 11219
rect 17622 11339 17702 11341
rect 17622 11218 17634 11339
rect 17690 11218 17702 11339
rect 16944 11209 17000 11217
rect 17312 11209 17368 11217
rect 17622 11216 17702 11218
rect 17634 11208 17690 11216
rect 17128 11041 17184 11049
rect 17496 11041 17552 11049
rect 17116 11039 17605 11041
rect 17116 10919 17128 11039
rect 17184 10919 17496 11039
rect 17552 10919 17605 11039
rect 17116 10917 17605 10919
rect 17128 10909 17184 10917
rect 17496 10909 17605 10917
rect 17024 10843 17104 10853
rect 17024 10787 17036 10843
rect 17092 10787 17104 10843
rect 17024 10777 17104 10787
rect 17208 10843 17288 10853
rect 17208 10787 17220 10843
rect 17276 10787 17288 10843
rect 17208 10777 17288 10787
rect 17392 10843 17472 10853
rect 17392 10787 17404 10843
rect 17460 10787 17472 10843
rect 17392 10777 17472 10787
rect 17036 10695 17092 10777
rect 17024 10693 17104 10695
rect 17024 10637 17036 10693
rect 17092 10637 17104 10693
rect 17024 10635 17104 10637
rect 16216 10577 16286 10591
rect 16216 10521 16228 10577
rect 16284 10521 16286 10577
rect 16216 10509 16286 10521
rect 15914 9674 15984 9686
rect 16228 9678 16284 10509
rect 17036 10321 17092 10635
rect 17220 10579 17276 10777
rect 17208 10577 17288 10579
rect 17208 10521 17220 10577
rect 17276 10521 17288 10577
rect 17208 10519 17288 10521
rect 17220 10321 17276 10519
rect 17404 10463 17460 10777
rect 17537 10579 17605 10909
rect 17982 10589 18038 11821
rect 17537 10577 17617 10579
rect 17537 10521 17549 10577
rect 17605 10521 17617 10577
rect 17537 10519 17617 10521
rect 17980 10577 18040 10589
rect 17980 10521 17982 10577
rect 18038 10521 18040 10577
rect 17392 10461 17472 10463
rect 17392 10405 17404 10461
rect 17460 10405 17472 10461
rect 17392 10403 17472 10405
rect 17404 10321 17460 10403
rect 17024 10311 17104 10321
rect 17024 10255 17036 10311
rect 17092 10255 17104 10311
rect 17024 10245 17104 10255
rect 17208 10311 17288 10321
rect 17208 10255 17220 10311
rect 17276 10255 17288 10311
rect 17208 10245 17288 10255
rect 17392 10311 17472 10321
rect 17392 10255 17404 10311
rect 17460 10255 17472 10311
rect 17392 10245 17472 10255
rect 17537 10189 17605 10519
rect 17980 10509 18040 10521
rect 19412 10461 19482 10473
rect 19412 10405 19424 10461
rect 19480 10405 19482 10461
rect 19412 10393 19482 10405
rect 17496 10181 17605 10189
rect 17484 10179 17605 10181
rect 17484 10059 17496 10179
rect 17552 10059 17605 10179
rect 17484 10057 17605 10059
rect 17496 10049 17552 10057
rect 16799 9792 17697 9804
rect 16799 9736 16811 9792
rect 16867 9736 17629 9792
rect 17685 9736 17697 9792
rect 16799 9724 17697 9736
rect 15914 9618 15926 9674
rect 15982 9618 15984 9674
rect 15914 9616 15984 9618
rect 16226 9674 16286 9678
rect 16226 9618 16228 9674
rect 16284 9618 16286 9674
rect 15926 9004 15982 9616
rect 16226 9606 16286 9618
rect 19424 9514 19480 10393
rect 19424 9404 19480 9414
rect 15778 4509 15848 4521
rect 15778 4453 15790 4509
rect 15846 4453 15848 4509
rect 15778 4441 15848 4453
rect 15424 3151 15426 3207
rect 15482 3151 15710 3207
rect 14836 3091 14916 3093
rect 14836 3035 14848 3091
rect 14904 3035 14916 3091
rect 14836 3033 14916 3035
rect 14848 2951 14904 3033
rect 14468 2941 14548 2951
rect 14468 2885 14480 2941
rect 14536 2885 14548 2941
rect 14468 2875 14548 2885
rect 14652 2941 14732 2951
rect 14652 2885 14664 2941
rect 14720 2885 14732 2941
rect 14652 2875 14732 2885
rect 14836 2941 14916 2951
rect 14836 2885 14848 2941
rect 14904 2885 14916 2941
rect 14836 2875 14916 2885
rect 14981 2819 15049 3149
rect 15424 3139 15494 3151
rect 14940 2811 15049 2819
rect 14928 2809 15049 2811
rect 14928 2689 14940 2809
rect 14996 2689 15049 2809
rect 14928 2687 15049 2689
rect 14940 2679 14996 2687
rect 14243 2422 15139 2434
rect 14243 2366 14255 2422
rect 14311 2366 15073 2422
rect 15129 2366 15139 2422
rect 14243 2354 15139 2366
rect 13928 2303 14008 2313
rect 13928 2247 13940 2303
rect 13996 2247 14008 2303
rect 13928 2245 14008 2247
rect 13762 2193 13832 2196
rect 13762 2139 13764 2193
rect 13820 2139 13832 2193
rect 13762 2127 13832 2139
rect 12902 2086 13648 2098
rect 12902 2030 13270 2086
rect 13326 2030 13648 2086
rect 12902 2018 13648 2030
rect 12902 1765 12958 2018
rect 13270 1765 13326 2018
rect 13592 1765 13648 2018
rect 12890 1763 12970 1765
rect 12890 1643 12902 1763
rect 12958 1643 12970 1763
rect 12890 1641 12970 1643
rect 13258 1763 13338 1765
rect 13258 1643 13270 1763
rect 13326 1643 13338 1763
rect 13258 1641 13338 1643
rect 13580 1763 13660 1765
rect 13580 1642 13592 1763
rect 13648 1642 13660 1763
rect 12902 1633 12958 1641
rect 13270 1633 13326 1641
rect 13580 1640 13660 1642
rect 13592 1632 13648 1640
rect 13086 1465 13142 1473
rect 13454 1465 13510 1473
rect 13074 1463 13563 1465
rect 13074 1343 13086 1463
rect 13142 1343 13454 1463
rect 13510 1343 13563 1463
rect 13074 1341 13563 1343
rect 13086 1333 13142 1341
rect 13454 1333 13563 1341
rect 12982 1267 13062 1277
rect 12982 1211 12994 1267
rect 13050 1211 13062 1267
rect 12982 1201 13062 1211
rect 13166 1267 13246 1277
rect 13166 1211 13178 1267
rect 13234 1211 13246 1267
rect 13166 1201 13246 1211
rect 13350 1267 13430 1277
rect 13350 1211 13362 1267
rect 13418 1211 13430 1267
rect 13350 1201 13430 1211
rect 12994 1119 13050 1201
rect 12982 1117 13062 1119
rect 12982 1061 12994 1117
rect 13050 1061 13062 1117
rect 12982 1059 13062 1061
rect 12174 1001 12244 1015
rect 12174 945 12186 1001
rect 12242 945 12244 1001
rect 12174 933 12244 945
rect 12008 885 12088 897
rect 12008 829 12020 885
rect 12076 829 12088 885
rect 12008 817 12088 829
rect 11872 98 11942 110
rect 12186 102 12242 933
rect 12994 745 13050 1059
rect 13178 1003 13234 1201
rect 13166 1001 13246 1003
rect 13166 945 13178 1001
rect 13234 945 13246 1001
rect 13166 943 13246 945
rect 13178 745 13234 943
rect 13362 887 13418 1201
rect 13495 1003 13563 1333
rect 13940 1013 13996 2245
rect 13495 1001 13575 1003
rect 13495 945 13507 1001
rect 13563 945 13575 1001
rect 13495 943 13575 945
rect 13938 1001 13998 1013
rect 13938 945 13940 1001
rect 13996 945 13998 1001
rect 13350 885 13430 887
rect 13350 829 13362 885
rect 13418 829 13430 885
rect 13350 827 13430 829
rect 13362 745 13418 827
rect 12982 735 13062 745
rect 12982 679 12994 735
rect 13050 679 13062 735
rect 12982 669 13062 679
rect 13166 735 13246 745
rect 13166 679 13178 735
rect 13234 679 13246 735
rect 13166 669 13246 679
rect 13350 735 13430 745
rect 13350 679 13362 735
rect 13418 679 13430 735
rect 13350 669 13430 679
rect 13495 613 13563 943
rect 13938 933 13998 945
rect 13454 605 13563 613
rect 13442 603 13563 605
rect 13442 483 13454 603
rect 13510 483 13563 603
rect 13442 481 13563 483
rect 13454 473 13510 481
rect 12757 216 13655 228
rect 12757 160 12769 216
rect 12825 160 13587 216
rect 13643 160 13655 216
rect 12757 148 13655 160
rect 11872 42 11884 98
rect 11940 42 11942 98
rect 11872 30 11942 42
rect 12184 98 12244 102
rect 12184 42 12186 98
rect 12242 42 12244 98
rect 12184 30 12244 42
rect 11748 -175 11804 -165
rect 15790 -65 15846 4441
rect 15926 110 15982 8904
rect 16944 8701 17690 8713
rect 16944 8645 17312 8701
rect 17368 8645 17690 8701
rect 16944 8633 17690 8645
rect 16944 8380 17000 8633
rect 17312 8380 17368 8633
rect 17634 8380 17690 8633
rect 16932 8378 17012 8380
rect 16932 8258 16944 8378
rect 17000 8258 17012 8378
rect 16932 8256 17012 8258
rect 17300 8378 17380 8380
rect 17300 8258 17312 8378
rect 17368 8258 17380 8378
rect 17300 8256 17380 8258
rect 17622 8378 17702 8380
rect 17622 8257 17634 8378
rect 17690 8257 17702 8378
rect 16944 8248 17000 8256
rect 17312 8248 17368 8256
rect 17622 8255 17702 8257
rect 17634 8247 17690 8255
rect 17128 8080 17184 8088
rect 17496 8080 17552 8088
rect 17116 8078 17605 8080
rect 17116 7958 17128 8078
rect 17184 7958 17496 8078
rect 17552 7958 17605 8078
rect 17116 7956 17605 7958
rect 17128 7948 17184 7956
rect 17496 7948 17605 7956
rect 17024 7882 17104 7892
rect 17024 7826 17036 7882
rect 17092 7826 17104 7882
rect 17024 7816 17104 7826
rect 17208 7882 17288 7892
rect 17208 7826 17220 7882
rect 17276 7826 17288 7882
rect 17208 7816 17288 7826
rect 17392 7882 17472 7892
rect 17392 7826 17404 7882
rect 17460 7826 17472 7882
rect 17392 7816 17472 7826
rect 16136 7732 16222 7744
rect 17036 7734 17092 7816
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 17024 7732 17104 7734
rect 17024 7676 17036 7732
rect 17092 7676 17104 7732
rect 17024 7674 17104 7676
rect 16352 7616 16422 7628
rect 16352 7560 16364 7616
rect 16420 7560 16422 7616
rect 16352 7548 16422 7560
rect 16216 5411 16286 5425
rect 16216 5355 16228 5411
rect 16284 5355 16286 5411
rect 16216 5343 16286 5355
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 16062 897 16118 5165
rect 16228 1015 16284 5343
rect 16364 3102 16420 7548
rect 17036 7360 17092 7674
rect 17220 7618 17276 7816
rect 17208 7616 17288 7618
rect 17208 7560 17220 7616
rect 17276 7560 17288 7616
rect 17208 7558 17288 7560
rect 17220 7360 17276 7558
rect 17404 7502 17460 7816
rect 17537 7618 17605 7948
rect 17537 7616 17617 7618
rect 17537 7560 17549 7616
rect 17605 7560 17617 7616
rect 17537 7558 17617 7560
rect 17804 7616 17874 7628
rect 17804 7560 17806 7616
rect 17862 7560 17874 7616
rect 17392 7500 17472 7502
rect 17392 7444 17404 7500
rect 17460 7444 17472 7500
rect 17392 7442 17472 7444
rect 17404 7360 17460 7442
rect 17024 7350 17104 7360
rect 17024 7294 17036 7350
rect 17092 7294 17104 7350
rect 17024 7284 17104 7294
rect 17208 7350 17288 7360
rect 17208 7294 17220 7350
rect 17276 7294 17288 7350
rect 17208 7284 17288 7294
rect 17392 7350 17472 7360
rect 17392 7294 17404 7350
rect 17460 7294 17472 7350
rect 17392 7284 17472 7294
rect 17537 7228 17605 7558
rect 17804 7550 17874 7560
rect 17496 7220 17605 7228
rect 17484 7218 17605 7220
rect 17484 7098 17496 7218
rect 17552 7098 17605 7218
rect 17484 7096 17605 7098
rect 17496 7088 17552 7096
rect 16799 6831 17697 6843
rect 16799 6775 16811 6831
rect 16867 6775 17629 6831
rect 17685 6775 17697 6831
rect 16799 6763 17697 6775
rect 17806 6606 17862 7550
rect 17970 6713 18050 6723
rect 17970 6657 17982 6713
rect 18038 6657 18050 6713
rect 17970 6655 18050 6657
rect 17804 6603 17874 6606
rect 17804 6549 17806 6603
rect 17862 6549 17874 6603
rect 17804 6537 17874 6549
rect 16944 6496 17690 6508
rect 16944 6440 17312 6496
rect 17368 6440 17690 6496
rect 16944 6428 17690 6440
rect 16944 6175 17000 6428
rect 17312 6175 17368 6428
rect 17634 6175 17690 6428
rect 16932 6173 17012 6175
rect 16932 6053 16944 6173
rect 17000 6053 17012 6173
rect 16932 6051 17012 6053
rect 17300 6173 17380 6175
rect 17300 6053 17312 6173
rect 17368 6053 17380 6173
rect 17300 6051 17380 6053
rect 17622 6173 17702 6175
rect 17622 6052 17634 6173
rect 17690 6052 17702 6173
rect 16944 6043 17000 6051
rect 17312 6043 17368 6051
rect 17622 6050 17702 6052
rect 17634 6042 17690 6050
rect 17128 5875 17184 5883
rect 17496 5875 17552 5883
rect 17116 5873 17605 5875
rect 17116 5753 17128 5873
rect 17184 5753 17496 5873
rect 17552 5753 17605 5873
rect 17116 5751 17605 5753
rect 17128 5743 17184 5751
rect 17496 5743 17605 5751
rect 17024 5677 17104 5687
rect 17024 5621 17036 5677
rect 17092 5621 17104 5677
rect 17024 5611 17104 5621
rect 17208 5677 17288 5687
rect 17208 5621 17220 5677
rect 17276 5621 17288 5677
rect 17208 5611 17288 5621
rect 17392 5677 17472 5687
rect 17392 5621 17404 5677
rect 17460 5621 17472 5677
rect 17392 5611 17472 5621
rect 17036 5529 17092 5611
rect 17024 5527 17104 5529
rect 17024 5471 17036 5527
rect 17092 5471 17104 5527
rect 17024 5469 17104 5471
rect 17036 5155 17092 5469
rect 17220 5413 17276 5611
rect 17208 5411 17288 5413
rect 17208 5355 17220 5411
rect 17276 5355 17288 5411
rect 17208 5353 17288 5355
rect 17220 5155 17276 5353
rect 17404 5297 17460 5611
rect 17537 5413 17605 5743
rect 17982 5421 18038 6655
rect 18430 6496 19176 6508
rect 18430 6440 18798 6496
rect 18854 6440 19176 6496
rect 18430 6428 19176 6440
rect 18430 6175 18486 6428
rect 18798 6175 18854 6428
rect 19120 6175 19176 6428
rect 18418 6173 18498 6175
rect 18418 6053 18430 6173
rect 18486 6053 18498 6173
rect 18418 6051 18498 6053
rect 18786 6173 18866 6175
rect 18786 6053 18798 6173
rect 18854 6053 18866 6173
rect 18786 6051 18866 6053
rect 19108 6173 19188 6175
rect 19108 6052 19120 6173
rect 19176 6052 19188 6173
rect 18430 6043 18486 6051
rect 18798 6043 18854 6051
rect 19108 6050 19188 6052
rect 19120 6042 19176 6050
rect 18614 5875 18670 5883
rect 18982 5875 19038 5883
rect 18602 5873 19091 5875
rect 18602 5753 18614 5873
rect 18670 5753 18982 5873
rect 19038 5753 19091 5873
rect 18602 5751 19091 5753
rect 18614 5743 18670 5751
rect 18982 5743 19091 5751
rect 18510 5677 18590 5687
rect 18510 5621 18522 5677
rect 18578 5621 18590 5677
rect 18510 5611 18590 5621
rect 18694 5677 18774 5687
rect 18694 5621 18706 5677
rect 18762 5621 18774 5677
rect 18694 5611 18774 5621
rect 18878 5677 18958 5687
rect 18878 5621 18890 5677
rect 18946 5621 18958 5677
rect 18878 5611 18958 5621
rect 18522 5529 18578 5611
rect 18510 5527 18590 5529
rect 18510 5471 18522 5527
rect 18578 5471 18590 5527
rect 18510 5469 18590 5471
rect 17537 5411 17617 5413
rect 17537 5355 17549 5411
rect 17605 5355 17617 5411
rect 17537 5353 17617 5355
rect 17980 5411 18040 5421
rect 17980 5355 17982 5411
rect 18038 5355 18040 5411
rect 17392 5295 17472 5297
rect 17392 5239 17404 5295
rect 17460 5239 17472 5295
rect 17392 5237 17472 5239
rect 17404 5155 17460 5237
rect 17024 5145 17104 5155
rect 17024 5089 17036 5145
rect 17092 5089 17104 5145
rect 17024 5079 17104 5089
rect 17208 5145 17288 5155
rect 17208 5089 17220 5145
rect 17276 5089 17288 5145
rect 17208 5079 17288 5089
rect 17392 5145 17472 5155
rect 17392 5089 17404 5145
rect 17460 5089 17472 5145
rect 17392 5079 17472 5089
rect 17537 5023 17605 5353
rect 17980 5343 18040 5355
rect 17496 5015 17605 5023
rect 17484 5013 17605 5015
rect 17484 4893 17496 5013
rect 17552 4893 17605 5013
rect 17484 4891 17605 4893
rect 17496 4883 17552 4891
rect 16799 4626 17695 4638
rect 16799 4570 16811 4626
rect 16867 4570 17629 4626
rect 17685 4570 17695 4626
rect 16799 4558 17695 4570
rect 17982 4400 18038 5343
rect 18522 5155 18578 5469
rect 18706 5413 18762 5611
rect 18694 5411 18774 5413
rect 18694 5355 18706 5411
rect 18762 5355 18774 5411
rect 18694 5353 18774 5355
rect 18706 5155 18762 5353
rect 18890 5297 18946 5611
rect 19023 5413 19091 5743
rect 19023 5411 19103 5413
rect 19023 5355 19035 5411
rect 19091 5355 19103 5411
rect 19023 5353 19103 5355
rect 19290 5411 19360 5423
rect 19290 5355 19292 5411
rect 19348 5355 19616 5411
rect 18878 5295 18958 5297
rect 18878 5239 18890 5295
rect 18946 5239 18958 5295
rect 18878 5237 18958 5239
rect 18890 5155 18946 5237
rect 18510 5145 18590 5155
rect 18510 5089 18522 5145
rect 18578 5089 18590 5145
rect 18510 5079 18590 5089
rect 18694 5145 18774 5155
rect 18694 5089 18706 5145
rect 18762 5089 18774 5145
rect 18694 5079 18774 5089
rect 18878 5145 18958 5155
rect 18878 5089 18890 5145
rect 18946 5089 18958 5145
rect 18878 5079 18958 5089
rect 19023 5023 19091 5353
rect 19290 5345 19360 5355
rect 18982 5015 19091 5023
rect 18970 5013 19091 5015
rect 18970 4893 18982 5013
rect 19038 4893 19091 5013
rect 18970 4891 19091 4893
rect 18982 4883 19038 4891
rect 18285 4626 19181 4638
rect 18285 4570 18297 4626
rect 18353 4570 19115 4626
rect 19171 4570 19181 4626
rect 18285 4558 19181 4570
rect 19292 4401 19348 5345
rect 19456 4509 19536 4519
rect 19456 4453 19468 4509
rect 19524 4453 19536 4509
rect 19456 4451 19536 4453
rect 17980 4398 18050 4400
rect 17980 4342 17982 4398
rect 18038 4342 18050 4398
rect 17980 4330 18050 4342
rect 19280 4399 19360 4401
rect 19280 4343 19292 4399
rect 19348 4343 19360 4399
rect 19280 4331 19360 4343
rect 16944 4291 17690 4303
rect 16944 4235 17312 4291
rect 17368 4235 17690 4291
rect 16944 4223 17690 4235
rect 16944 3970 17000 4223
rect 17312 3970 17368 4223
rect 17634 3970 17690 4223
rect 18430 4292 19176 4304
rect 18430 4236 18798 4292
rect 18854 4236 19176 4292
rect 18430 4224 19176 4236
rect 18430 3971 18486 4224
rect 18798 3971 18854 4224
rect 19120 3971 19176 4224
rect 16932 3968 17012 3970
rect 16932 3848 16944 3968
rect 17000 3848 17012 3968
rect 16932 3846 17012 3848
rect 17300 3968 17380 3970
rect 17300 3848 17312 3968
rect 17368 3848 17380 3968
rect 17300 3846 17380 3848
rect 17622 3968 17702 3970
rect 17622 3847 17634 3968
rect 17690 3847 17702 3968
rect 18418 3969 18498 3971
rect 18418 3849 18430 3969
rect 18486 3849 18498 3969
rect 18418 3847 18498 3849
rect 18786 3969 18866 3971
rect 18786 3849 18798 3969
rect 18854 3849 18866 3969
rect 18786 3847 18866 3849
rect 19108 3969 19188 3971
rect 19108 3848 19120 3969
rect 19176 3848 19188 3969
rect 16944 3838 17000 3846
rect 17312 3838 17368 3846
rect 17622 3845 17702 3847
rect 17634 3837 17690 3845
rect 18430 3839 18486 3847
rect 18798 3839 18854 3847
rect 19108 3846 19188 3848
rect 19120 3838 19176 3846
rect 17128 3670 17184 3678
rect 17496 3670 17552 3678
rect 18614 3671 18670 3679
rect 18982 3671 19038 3679
rect 17116 3668 17605 3670
rect 17116 3548 17128 3668
rect 17184 3548 17496 3668
rect 17552 3548 17605 3668
rect 17116 3546 17605 3548
rect 18602 3669 19091 3671
rect 18602 3549 18614 3669
rect 18670 3549 18982 3669
rect 19038 3549 19091 3669
rect 18602 3547 19091 3549
rect 17128 3538 17184 3546
rect 17496 3538 17605 3546
rect 18614 3539 18670 3547
rect 18982 3539 19091 3547
rect 17024 3472 17104 3482
rect 17024 3416 17036 3472
rect 17092 3416 17104 3472
rect 17024 3406 17104 3416
rect 17208 3472 17288 3482
rect 17208 3416 17220 3472
rect 17276 3416 17288 3472
rect 17208 3406 17288 3416
rect 17392 3472 17472 3482
rect 17392 3416 17404 3472
rect 17460 3416 17472 3472
rect 17392 3406 17472 3416
rect 17036 3324 17092 3406
rect 17024 3322 17104 3324
rect 17024 3266 17036 3322
rect 17092 3266 17104 3322
rect 17024 3264 17104 3266
rect 16352 3090 16422 3102
rect 16352 3034 16364 3090
rect 16420 3034 16422 3090
rect 16352 3022 16422 3034
rect 17036 2950 17092 3264
rect 17220 3208 17276 3406
rect 17208 3206 17288 3208
rect 17208 3150 17220 3206
rect 17276 3150 17288 3206
rect 17208 3148 17288 3150
rect 17220 2950 17276 3148
rect 17404 3092 17460 3406
rect 17537 3208 17605 3538
rect 18510 3473 18590 3483
rect 18510 3417 18522 3473
rect 18578 3417 18590 3473
rect 18510 3407 18590 3417
rect 18694 3473 18774 3483
rect 18694 3417 18706 3473
rect 18762 3417 18774 3473
rect 18694 3407 18774 3417
rect 18878 3473 18958 3483
rect 18878 3417 18890 3473
rect 18946 3417 18958 3473
rect 18878 3407 18958 3417
rect 18522 3325 18578 3407
rect 18510 3323 18590 3325
rect 18510 3267 18522 3323
rect 18578 3267 18590 3323
rect 18510 3265 18590 3267
rect 17537 3206 17617 3208
rect 17537 3150 17549 3206
rect 17605 3150 17617 3206
rect 17537 3148 17617 3150
rect 17804 3206 17874 3218
rect 17804 3150 17806 3206
rect 17862 3150 17874 3206
rect 17392 3090 17472 3092
rect 17392 3034 17404 3090
rect 17460 3034 17472 3090
rect 17392 3032 17472 3034
rect 17404 2950 17460 3032
rect 17024 2940 17104 2950
rect 17024 2884 17036 2940
rect 17092 2884 17104 2940
rect 17024 2874 17104 2884
rect 17208 2940 17288 2950
rect 17208 2884 17220 2940
rect 17276 2884 17288 2940
rect 17208 2874 17288 2884
rect 17392 2940 17472 2950
rect 17392 2884 17404 2940
rect 17460 2884 17472 2940
rect 17392 2874 17472 2884
rect 17537 2818 17605 3148
rect 17804 3140 17874 3150
rect 17496 2810 17605 2818
rect 17484 2808 17605 2810
rect 17484 2688 17496 2808
rect 17552 2688 17605 2808
rect 17484 2686 17605 2688
rect 17496 2678 17552 2686
rect 16799 2421 17695 2433
rect 16799 2365 16811 2421
rect 16867 2365 17629 2421
rect 17685 2365 17695 2421
rect 16799 2353 17695 2365
rect 17806 2196 17862 3140
rect 18522 2951 18578 3265
rect 18706 3209 18762 3407
rect 18694 3207 18774 3209
rect 18694 3151 18706 3207
rect 18762 3151 18774 3207
rect 18694 3149 18774 3151
rect 18706 2951 18762 3149
rect 18890 3093 18946 3407
rect 19023 3209 19091 3539
rect 19468 3217 19524 4451
rect 19023 3207 19103 3209
rect 19023 3151 19035 3207
rect 19091 3151 19103 3207
rect 19023 3149 19103 3151
rect 19466 3207 19536 3217
rect 19696 3207 19752 17250
rect 19898 14999 19954 19031
rect 23940 18915 23996 19504
rect 23938 18913 24008 18915
rect 23938 18857 23940 18913
rect 23996 18857 24008 18913
rect 23938 18855 24008 18857
rect 20122 18737 20192 18749
rect 20122 18681 20134 18737
rect 20190 18681 20192 18737
rect 20122 18679 20192 18681
rect 19896 14987 19966 14999
rect 19896 14931 19898 14987
rect 19954 14931 19966 14987
rect 19896 14919 19966 14931
rect 20134 14087 20190 18679
rect 20986 18277 21732 18289
rect 20986 18221 21354 18277
rect 21410 18221 21732 18277
rect 20986 18209 21732 18221
rect 20986 17956 21042 18209
rect 21354 17956 21410 18209
rect 21676 17956 21732 18209
rect 20974 17954 21054 17956
rect 20974 17834 20986 17954
rect 21042 17834 21054 17954
rect 20974 17832 21054 17834
rect 21342 17954 21422 17956
rect 21342 17834 21354 17954
rect 21410 17834 21422 17954
rect 21342 17832 21422 17834
rect 21664 17954 21744 17956
rect 21664 17833 21676 17954
rect 21732 17833 21744 17954
rect 20986 17824 21042 17832
rect 21354 17824 21410 17832
rect 21664 17831 21744 17833
rect 21676 17823 21732 17831
rect 21170 17656 21226 17664
rect 21538 17656 21594 17664
rect 21158 17654 21647 17656
rect 21158 17534 21170 17654
rect 21226 17534 21538 17654
rect 21594 17534 21647 17654
rect 21158 17532 21647 17534
rect 21170 17524 21226 17532
rect 21538 17524 21647 17532
rect 21066 17458 21146 17468
rect 21066 17402 21078 17458
rect 21134 17402 21146 17458
rect 21066 17392 21146 17402
rect 21250 17458 21330 17468
rect 21250 17402 21262 17458
rect 21318 17402 21330 17458
rect 21250 17392 21330 17402
rect 21434 17458 21514 17468
rect 21434 17402 21446 17458
rect 21502 17402 21514 17458
rect 21434 17392 21514 17402
rect 21078 17310 21134 17392
rect 21066 17308 21146 17310
rect 21066 17252 21078 17308
rect 21134 17252 21146 17308
rect 21066 17250 21146 17252
rect 20394 17192 20464 17204
rect 20394 17136 20406 17192
rect 20462 17136 20464 17192
rect 20394 17124 20464 17136
rect 20258 14987 20328 15001
rect 20258 14931 20270 14987
rect 20326 14931 20328 14987
rect 20258 14919 20328 14931
rect 20122 14085 20192 14087
rect 20122 14029 20134 14085
rect 20190 14029 20192 14085
rect 20122 14017 20192 14029
rect 20270 10591 20326 14919
rect 20406 12678 20462 17124
rect 21078 16936 21134 17250
rect 21262 17194 21318 17392
rect 21250 17192 21330 17194
rect 21250 17136 21262 17192
rect 21318 17136 21330 17192
rect 21250 17134 21330 17136
rect 21262 16936 21318 17134
rect 21446 17078 21502 17392
rect 21579 17194 21647 17524
rect 23726 17308 23796 17320
rect 23726 17252 23738 17308
rect 23794 17252 23796 17308
rect 23726 17250 23796 17252
rect 21579 17192 21659 17194
rect 21579 17136 21591 17192
rect 21647 17136 21659 17192
rect 21579 17134 21659 17136
rect 21846 17192 21916 17204
rect 21846 17136 21848 17192
rect 21904 17136 21916 17192
rect 21434 17076 21514 17078
rect 21434 17020 21446 17076
rect 21502 17020 21514 17076
rect 21434 17018 21514 17020
rect 21446 16936 21502 17018
rect 21066 16926 21146 16936
rect 21066 16870 21078 16926
rect 21134 16870 21146 16926
rect 21066 16860 21146 16870
rect 21250 16926 21330 16936
rect 21250 16870 21262 16926
rect 21318 16870 21330 16926
rect 21250 16860 21330 16870
rect 21434 16926 21514 16936
rect 21434 16870 21446 16926
rect 21502 16870 21514 16926
rect 21434 16860 21514 16870
rect 21579 16804 21647 17134
rect 21846 17126 21916 17136
rect 21538 16796 21647 16804
rect 21526 16794 21647 16796
rect 21526 16674 21538 16794
rect 21594 16674 21647 16794
rect 21526 16672 21647 16674
rect 21538 16664 21594 16672
rect 20841 16407 21739 16419
rect 20841 16351 20853 16407
rect 20909 16351 21671 16407
rect 21727 16351 21739 16407
rect 20841 16339 21739 16351
rect 21848 16182 21904 17126
rect 22012 16289 22092 16299
rect 22012 16233 22024 16289
rect 22080 16233 22092 16289
rect 22012 16231 22092 16233
rect 21846 16179 21916 16182
rect 21846 16125 21848 16179
rect 21904 16125 21916 16179
rect 21846 16113 21916 16125
rect 20986 16072 21732 16084
rect 20986 16016 21354 16072
rect 21410 16016 21732 16072
rect 20986 16004 21732 16016
rect 20986 15751 21042 16004
rect 21354 15751 21410 16004
rect 21676 15751 21732 16004
rect 20974 15749 21054 15751
rect 20974 15629 20986 15749
rect 21042 15629 21054 15749
rect 20974 15627 21054 15629
rect 21342 15749 21422 15751
rect 21342 15629 21354 15749
rect 21410 15629 21422 15749
rect 21342 15627 21422 15629
rect 21664 15749 21744 15751
rect 21664 15628 21676 15749
rect 21732 15628 21744 15749
rect 20986 15619 21042 15627
rect 21354 15619 21410 15627
rect 21664 15626 21744 15628
rect 21676 15618 21732 15626
rect 21170 15451 21226 15459
rect 21538 15451 21594 15459
rect 21158 15449 21647 15451
rect 21158 15329 21170 15449
rect 21226 15329 21538 15449
rect 21594 15329 21647 15449
rect 21158 15327 21647 15329
rect 21170 15319 21226 15327
rect 21538 15319 21647 15327
rect 21066 15253 21146 15263
rect 21066 15197 21078 15253
rect 21134 15197 21146 15253
rect 21066 15187 21146 15197
rect 21250 15253 21330 15263
rect 21250 15197 21262 15253
rect 21318 15197 21330 15253
rect 21250 15187 21330 15197
rect 21434 15253 21514 15263
rect 21434 15197 21446 15253
rect 21502 15197 21514 15253
rect 21434 15187 21514 15197
rect 21078 15105 21134 15187
rect 21066 15103 21146 15105
rect 21066 15047 21078 15103
rect 21134 15047 21146 15103
rect 21066 15045 21146 15047
rect 21078 14731 21134 15045
rect 21262 14989 21318 15187
rect 21250 14987 21330 14989
rect 21250 14931 21262 14987
rect 21318 14931 21330 14987
rect 21250 14929 21330 14931
rect 21262 14731 21318 14929
rect 21446 14873 21502 15187
rect 21579 14989 21647 15319
rect 22024 14997 22080 16231
rect 22472 16072 23218 16084
rect 22472 16016 22840 16072
rect 22896 16016 23218 16072
rect 22472 16004 23218 16016
rect 22472 15751 22528 16004
rect 22840 15751 22896 16004
rect 23162 15751 23218 16004
rect 22460 15749 22540 15751
rect 22460 15629 22472 15749
rect 22528 15629 22540 15749
rect 22460 15627 22540 15629
rect 22828 15749 22908 15751
rect 22828 15629 22840 15749
rect 22896 15629 22908 15749
rect 22828 15627 22908 15629
rect 23150 15749 23230 15751
rect 23150 15628 23162 15749
rect 23218 15628 23230 15749
rect 22472 15619 22528 15627
rect 22840 15619 22896 15627
rect 23150 15626 23230 15628
rect 23162 15618 23218 15626
rect 22656 15451 22712 15459
rect 23024 15451 23080 15459
rect 22644 15449 23133 15451
rect 22644 15329 22656 15449
rect 22712 15329 23024 15449
rect 23080 15329 23133 15449
rect 22644 15327 23133 15329
rect 22656 15319 22712 15327
rect 23024 15319 23133 15327
rect 22552 15253 22632 15263
rect 22552 15197 22564 15253
rect 22620 15197 22632 15253
rect 22552 15187 22632 15197
rect 22736 15253 22816 15263
rect 22736 15197 22748 15253
rect 22804 15197 22816 15253
rect 22736 15187 22816 15197
rect 22920 15253 23000 15263
rect 22920 15197 22932 15253
rect 22988 15197 23000 15253
rect 22920 15187 23000 15197
rect 22564 15105 22620 15187
rect 22552 15103 22632 15105
rect 22552 15047 22564 15103
rect 22620 15047 22632 15103
rect 22552 15045 22632 15047
rect 21579 14987 21659 14989
rect 21579 14931 21591 14987
rect 21647 14931 21659 14987
rect 21579 14929 21659 14931
rect 22022 14987 22082 14997
rect 22022 14931 22024 14987
rect 22080 14931 22082 14987
rect 21434 14871 21514 14873
rect 21434 14815 21446 14871
rect 21502 14815 21514 14871
rect 21434 14813 21514 14815
rect 21446 14731 21502 14813
rect 21066 14721 21146 14731
rect 21066 14665 21078 14721
rect 21134 14665 21146 14721
rect 21066 14655 21146 14665
rect 21250 14721 21330 14731
rect 21250 14665 21262 14721
rect 21318 14665 21330 14721
rect 21250 14655 21330 14665
rect 21434 14721 21514 14731
rect 21434 14665 21446 14721
rect 21502 14665 21514 14721
rect 21434 14655 21514 14665
rect 21579 14599 21647 14929
rect 22022 14919 22082 14931
rect 21538 14591 21647 14599
rect 21526 14589 21647 14591
rect 21526 14469 21538 14589
rect 21594 14469 21647 14589
rect 21526 14467 21647 14469
rect 21538 14459 21594 14467
rect 20841 14202 21737 14214
rect 20841 14146 20853 14202
rect 20909 14146 21671 14202
rect 21727 14146 21737 14202
rect 20841 14134 21737 14146
rect 22024 13976 22080 14919
rect 22564 14731 22620 15045
rect 22748 14989 22804 15187
rect 22736 14987 22816 14989
rect 22736 14931 22748 14987
rect 22804 14931 22816 14987
rect 22736 14929 22816 14931
rect 22748 14731 22804 14929
rect 22932 14873 22988 15187
rect 23065 14989 23133 15319
rect 23065 14987 23145 14989
rect 23065 14931 23077 14987
rect 23133 14931 23145 14987
rect 23065 14929 23145 14931
rect 23332 14987 23402 14999
rect 23332 14931 23334 14987
rect 23390 14931 23658 14987
rect 22920 14871 23000 14873
rect 22920 14815 22932 14871
rect 22988 14815 23000 14871
rect 22920 14813 23000 14815
rect 22932 14731 22988 14813
rect 22552 14721 22632 14731
rect 22552 14665 22564 14721
rect 22620 14665 22632 14721
rect 22552 14655 22632 14665
rect 22736 14721 22816 14731
rect 22736 14665 22748 14721
rect 22804 14665 22816 14721
rect 22736 14655 22816 14665
rect 22920 14721 23000 14731
rect 22920 14665 22932 14721
rect 22988 14665 23000 14721
rect 22920 14655 23000 14665
rect 23065 14599 23133 14929
rect 23332 14921 23402 14931
rect 23024 14591 23133 14599
rect 23012 14589 23133 14591
rect 23012 14469 23024 14589
rect 23080 14469 23133 14589
rect 23012 14467 23133 14469
rect 23024 14459 23080 14467
rect 22327 14202 23223 14214
rect 22327 14146 22339 14202
rect 22395 14146 23157 14202
rect 23213 14146 23223 14202
rect 22327 14134 23223 14146
rect 23334 13977 23390 14921
rect 23498 14085 23578 14095
rect 23498 14029 23510 14085
rect 23566 14029 23578 14085
rect 23498 14027 23578 14029
rect 22022 13974 22092 13976
rect 22022 13918 22024 13974
rect 22080 13918 22092 13974
rect 22022 13906 22092 13918
rect 23322 13975 23402 13977
rect 23322 13919 23334 13975
rect 23390 13919 23402 13975
rect 23322 13907 23402 13919
rect 20986 13867 21732 13879
rect 20986 13811 21354 13867
rect 21410 13811 21732 13867
rect 20986 13799 21732 13811
rect 20986 13546 21042 13799
rect 21354 13546 21410 13799
rect 21676 13546 21732 13799
rect 22472 13868 23218 13880
rect 22472 13812 22840 13868
rect 22896 13812 23218 13868
rect 22472 13800 23218 13812
rect 22472 13547 22528 13800
rect 22840 13547 22896 13800
rect 23162 13547 23218 13800
rect 20974 13544 21054 13546
rect 20974 13424 20986 13544
rect 21042 13424 21054 13544
rect 20974 13422 21054 13424
rect 21342 13544 21422 13546
rect 21342 13424 21354 13544
rect 21410 13424 21422 13544
rect 21342 13422 21422 13424
rect 21664 13544 21744 13546
rect 21664 13423 21676 13544
rect 21732 13423 21744 13544
rect 22460 13545 22540 13547
rect 22460 13425 22472 13545
rect 22528 13425 22540 13545
rect 22460 13423 22540 13425
rect 22828 13545 22908 13547
rect 22828 13425 22840 13545
rect 22896 13425 22908 13545
rect 22828 13423 22908 13425
rect 23150 13545 23230 13547
rect 23150 13424 23162 13545
rect 23218 13424 23230 13545
rect 20986 13414 21042 13422
rect 21354 13414 21410 13422
rect 21664 13421 21744 13423
rect 21676 13413 21732 13421
rect 22472 13415 22528 13423
rect 22840 13415 22896 13423
rect 23150 13422 23230 13424
rect 23162 13414 23218 13422
rect 21170 13246 21226 13254
rect 21538 13246 21594 13254
rect 22656 13247 22712 13255
rect 23024 13247 23080 13255
rect 21158 13244 21647 13246
rect 21158 13124 21170 13244
rect 21226 13124 21538 13244
rect 21594 13124 21647 13244
rect 21158 13122 21647 13124
rect 22644 13245 23133 13247
rect 22644 13125 22656 13245
rect 22712 13125 23024 13245
rect 23080 13125 23133 13245
rect 22644 13123 23133 13125
rect 21170 13114 21226 13122
rect 21538 13114 21647 13122
rect 22656 13115 22712 13123
rect 23024 13115 23133 13123
rect 21066 13048 21146 13058
rect 21066 12992 21078 13048
rect 21134 12992 21146 13048
rect 21066 12982 21146 12992
rect 21250 13048 21330 13058
rect 21250 12992 21262 13048
rect 21318 12992 21330 13048
rect 21250 12982 21330 12992
rect 21434 13048 21514 13058
rect 21434 12992 21446 13048
rect 21502 12992 21514 13048
rect 21434 12982 21514 12992
rect 21078 12900 21134 12982
rect 21066 12898 21146 12900
rect 21066 12842 21078 12898
rect 21134 12842 21146 12898
rect 21066 12840 21146 12842
rect 20394 12666 20464 12678
rect 20394 12610 20406 12666
rect 20462 12610 20464 12666
rect 20394 12598 20464 12610
rect 21078 12526 21134 12840
rect 21262 12784 21318 12982
rect 21250 12782 21330 12784
rect 21250 12726 21262 12782
rect 21318 12726 21330 12782
rect 21250 12724 21330 12726
rect 21262 12526 21318 12724
rect 21446 12668 21502 12982
rect 21579 12784 21647 13114
rect 22552 13049 22632 13059
rect 22552 12993 22564 13049
rect 22620 12993 22632 13049
rect 22552 12983 22632 12993
rect 22736 13049 22816 13059
rect 22736 12993 22748 13049
rect 22804 12993 22816 13049
rect 22736 12983 22816 12993
rect 22920 13049 23000 13059
rect 22920 12993 22932 13049
rect 22988 12993 23000 13049
rect 22920 12983 23000 12993
rect 22564 12901 22620 12983
rect 22552 12899 22632 12901
rect 22552 12843 22564 12899
rect 22620 12843 22632 12899
rect 22552 12841 22632 12843
rect 21579 12782 21659 12784
rect 21579 12726 21591 12782
rect 21647 12726 21659 12782
rect 21579 12724 21659 12726
rect 21846 12782 21916 12794
rect 21846 12726 21848 12782
rect 21904 12726 21916 12782
rect 21434 12666 21514 12668
rect 21434 12610 21446 12666
rect 21502 12610 21514 12666
rect 21434 12608 21514 12610
rect 21446 12526 21502 12608
rect 21066 12516 21146 12526
rect 21066 12460 21078 12516
rect 21134 12460 21146 12516
rect 21066 12450 21146 12460
rect 21250 12516 21330 12526
rect 21250 12460 21262 12516
rect 21318 12460 21330 12516
rect 21250 12450 21330 12460
rect 21434 12516 21514 12526
rect 21434 12460 21446 12516
rect 21502 12460 21514 12516
rect 21434 12450 21514 12460
rect 21579 12394 21647 12724
rect 21846 12716 21916 12726
rect 21538 12386 21647 12394
rect 21526 12384 21647 12386
rect 21526 12264 21538 12384
rect 21594 12264 21647 12384
rect 21526 12262 21647 12264
rect 21538 12254 21594 12262
rect 20841 11997 21737 12009
rect 20841 11941 20853 11997
rect 20909 11941 21671 11997
rect 21727 11941 21737 11997
rect 20841 11929 21737 11941
rect 21848 11772 21904 12716
rect 22564 12527 22620 12841
rect 22748 12785 22804 12983
rect 22736 12783 22816 12785
rect 22736 12727 22748 12783
rect 22804 12727 22816 12783
rect 22736 12725 22816 12727
rect 22748 12527 22804 12725
rect 22932 12669 22988 12983
rect 23065 12785 23133 13115
rect 23510 12793 23566 14027
rect 23065 12783 23145 12785
rect 23065 12727 23077 12783
rect 23133 12727 23145 12783
rect 23065 12725 23145 12727
rect 23508 12783 23578 12793
rect 23508 12727 23510 12783
rect 23566 12727 23658 12783
rect 22920 12667 23000 12669
rect 22920 12611 22932 12667
rect 22988 12611 23000 12667
rect 22920 12609 23000 12611
rect 22932 12527 22988 12609
rect 22552 12517 22632 12527
rect 22552 12461 22564 12517
rect 22620 12461 22632 12517
rect 22552 12451 22632 12461
rect 22736 12517 22816 12527
rect 22736 12461 22748 12517
rect 22804 12461 22816 12517
rect 22736 12451 22816 12461
rect 22920 12517 23000 12527
rect 22920 12461 22932 12517
rect 22988 12461 23000 12517
rect 22920 12451 23000 12461
rect 23065 12395 23133 12725
rect 23508 12715 23578 12727
rect 23024 12387 23133 12395
rect 23012 12385 23133 12387
rect 23012 12265 23024 12385
rect 23080 12265 23133 12385
rect 23012 12263 23133 12265
rect 23024 12255 23080 12263
rect 22327 11998 23223 12010
rect 22327 11942 22339 11998
rect 22395 11942 23157 11998
rect 23213 11942 23223 11998
rect 22327 11930 23223 11942
rect 22012 11879 22092 11889
rect 22012 11823 22024 11879
rect 22080 11823 22092 11879
rect 22012 11821 22092 11823
rect 21846 11769 21916 11772
rect 21846 11715 21848 11769
rect 21904 11715 21916 11769
rect 21846 11703 21916 11715
rect 20986 11662 21732 11674
rect 20986 11606 21354 11662
rect 21410 11606 21732 11662
rect 20986 11594 21732 11606
rect 20986 11341 21042 11594
rect 21354 11341 21410 11594
rect 21676 11341 21732 11594
rect 20974 11339 21054 11341
rect 20974 11219 20986 11339
rect 21042 11219 21054 11339
rect 20974 11217 21054 11219
rect 21342 11339 21422 11341
rect 21342 11219 21354 11339
rect 21410 11219 21422 11339
rect 21342 11217 21422 11219
rect 21664 11339 21744 11341
rect 21664 11218 21676 11339
rect 21732 11218 21744 11339
rect 20986 11209 21042 11217
rect 21354 11209 21410 11217
rect 21664 11216 21744 11218
rect 21676 11208 21732 11216
rect 21170 11041 21226 11049
rect 21538 11041 21594 11049
rect 21158 11039 21647 11041
rect 21158 10919 21170 11039
rect 21226 10919 21538 11039
rect 21594 10919 21647 11039
rect 21158 10917 21647 10919
rect 21170 10909 21226 10917
rect 21538 10909 21647 10917
rect 21066 10843 21146 10853
rect 21066 10787 21078 10843
rect 21134 10787 21146 10843
rect 21066 10777 21146 10787
rect 21250 10843 21330 10853
rect 21250 10787 21262 10843
rect 21318 10787 21330 10843
rect 21250 10777 21330 10787
rect 21434 10843 21514 10853
rect 21434 10787 21446 10843
rect 21502 10787 21514 10843
rect 21434 10777 21514 10787
rect 21078 10695 21134 10777
rect 21066 10693 21146 10695
rect 21066 10637 21078 10693
rect 21134 10637 21146 10693
rect 21066 10635 21146 10637
rect 20258 10577 20328 10591
rect 20258 10521 20270 10577
rect 20326 10521 20328 10577
rect 20258 10509 20328 10521
rect 19956 9674 20026 9686
rect 20270 9678 20326 10509
rect 21078 10321 21134 10635
rect 21262 10579 21318 10777
rect 21250 10577 21330 10579
rect 21250 10521 21262 10577
rect 21318 10521 21330 10577
rect 21250 10519 21330 10521
rect 21262 10321 21318 10519
rect 21446 10463 21502 10777
rect 21579 10579 21647 10909
rect 22024 10589 22080 11821
rect 21579 10577 21659 10579
rect 21579 10521 21591 10577
rect 21647 10521 21659 10577
rect 21579 10519 21659 10521
rect 22022 10577 22082 10589
rect 22022 10521 22024 10577
rect 22080 10521 22082 10577
rect 21434 10461 21514 10463
rect 21434 10405 21446 10461
rect 21502 10405 21514 10461
rect 21434 10403 21514 10405
rect 21446 10321 21502 10403
rect 21066 10311 21146 10321
rect 21066 10255 21078 10311
rect 21134 10255 21146 10311
rect 21066 10245 21146 10255
rect 21250 10311 21330 10321
rect 21250 10255 21262 10311
rect 21318 10255 21330 10311
rect 21250 10245 21330 10255
rect 21434 10311 21514 10321
rect 21434 10255 21446 10311
rect 21502 10255 21514 10311
rect 21434 10245 21514 10255
rect 21579 10189 21647 10519
rect 22022 10509 22082 10521
rect 23454 10461 23524 10473
rect 23454 10405 23466 10461
rect 23522 10405 23524 10461
rect 23454 10393 23524 10405
rect 21538 10181 21647 10189
rect 21526 10179 21647 10181
rect 21526 10059 21538 10179
rect 21594 10059 21647 10179
rect 21526 10057 21647 10059
rect 21538 10049 21594 10057
rect 20841 9792 21739 9804
rect 20841 9736 20853 9792
rect 20909 9736 21671 9792
rect 21727 9736 21739 9792
rect 20841 9724 21739 9736
rect 19956 9618 19968 9674
rect 20024 9618 20026 9674
rect 19956 9616 20026 9618
rect 20268 9674 20328 9678
rect 20268 9618 20270 9674
rect 20326 9618 20328 9674
rect 19968 9004 20024 9616
rect 20268 9606 20328 9618
rect 23466 9514 23522 10393
rect 23466 9404 23522 9414
rect 19820 4509 19890 4521
rect 19820 4453 19832 4509
rect 19888 4453 19890 4509
rect 19820 4441 19890 4453
rect 19466 3151 19468 3207
rect 19524 3151 19752 3207
rect 18878 3091 18958 3093
rect 18878 3035 18890 3091
rect 18946 3035 18958 3091
rect 18878 3033 18958 3035
rect 18890 2951 18946 3033
rect 18510 2941 18590 2951
rect 18510 2885 18522 2941
rect 18578 2885 18590 2941
rect 18510 2875 18590 2885
rect 18694 2941 18774 2951
rect 18694 2885 18706 2941
rect 18762 2885 18774 2941
rect 18694 2875 18774 2885
rect 18878 2941 18958 2951
rect 18878 2885 18890 2941
rect 18946 2885 18958 2941
rect 18878 2875 18958 2885
rect 19023 2819 19091 3149
rect 19466 3139 19536 3151
rect 18982 2811 19091 2819
rect 18970 2809 19091 2811
rect 18970 2689 18982 2809
rect 19038 2689 19091 2809
rect 18970 2687 19091 2689
rect 18982 2679 19038 2687
rect 18285 2422 19181 2434
rect 18285 2366 18297 2422
rect 18353 2366 19115 2422
rect 19171 2366 19181 2422
rect 18285 2354 19181 2366
rect 17970 2303 18050 2313
rect 17970 2247 17982 2303
rect 18038 2247 18050 2303
rect 17970 2245 18050 2247
rect 17804 2193 17874 2196
rect 17804 2139 17806 2193
rect 17862 2139 17874 2193
rect 17804 2127 17874 2139
rect 16944 2086 17690 2098
rect 16944 2030 17312 2086
rect 17368 2030 17690 2086
rect 16944 2018 17690 2030
rect 16944 1765 17000 2018
rect 17312 1765 17368 2018
rect 17634 1765 17690 2018
rect 16932 1763 17012 1765
rect 16932 1643 16944 1763
rect 17000 1643 17012 1763
rect 16932 1641 17012 1643
rect 17300 1763 17380 1765
rect 17300 1643 17312 1763
rect 17368 1643 17380 1763
rect 17300 1641 17380 1643
rect 17622 1763 17702 1765
rect 17622 1642 17634 1763
rect 17690 1642 17702 1763
rect 16944 1633 17000 1641
rect 17312 1633 17368 1641
rect 17622 1640 17702 1642
rect 17634 1632 17690 1640
rect 17128 1465 17184 1473
rect 17496 1465 17552 1473
rect 17116 1463 17605 1465
rect 17116 1343 17128 1463
rect 17184 1343 17496 1463
rect 17552 1343 17605 1463
rect 17116 1341 17605 1343
rect 17128 1333 17184 1341
rect 17496 1333 17605 1341
rect 17024 1267 17104 1277
rect 17024 1211 17036 1267
rect 17092 1211 17104 1267
rect 17024 1201 17104 1211
rect 17208 1267 17288 1277
rect 17208 1211 17220 1267
rect 17276 1211 17288 1267
rect 17208 1201 17288 1211
rect 17392 1267 17472 1277
rect 17392 1211 17404 1267
rect 17460 1211 17472 1267
rect 17392 1201 17472 1211
rect 17036 1119 17092 1201
rect 17024 1117 17104 1119
rect 17024 1061 17036 1117
rect 17092 1061 17104 1117
rect 17024 1059 17104 1061
rect 16216 1001 16286 1015
rect 16216 945 16228 1001
rect 16284 945 16286 1001
rect 16216 933 16286 945
rect 16050 885 16130 897
rect 16050 829 16062 885
rect 16118 829 16130 885
rect 16050 817 16130 829
rect 15914 98 15984 110
rect 16228 102 16284 933
rect 17036 745 17092 1059
rect 17220 1003 17276 1201
rect 17208 1001 17288 1003
rect 17208 945 17220 1001
rect 17276 945 17288 1001
rect 17208 943 17288 945
rect 17220 745 17276 943
rect 17404 887 17460 1201
rect 17537 1003 17605 1333
rect 17982 1013 18038 2245
rect 17537 1001 17617 1003
rect 17537 945 17549 1001
rect 17605 945 17617 1001
rect 17537 943 17617 945
rect 17980 1001 18040 1013
rect 17980 945 17982 1001
rect 18038 945 18040 1001
rect 17392 885 17472 887
rect 17392 829 17404 885
rect 17460 829 17472 885
rect 17392 827 17472 829
rect 17404 745 17460 827
rect 17024 735 17104 745
rect 17024 679 17036 735
rect 17092 679 17104 735
rect 17024 669 17104 679
rect 17208 735 17288 745
rect 17208 679 17220 735
rect 17276 679 17288 735
rect 17208 669 17288 679
rect 17392 735 17472 745
rect 17392 679 17404 735
rect 17460 679 17472 735
rect 17392 669 17472 679
rect 17537 613 17605 943
rect 17980 933 18040 945
rect 17496 605 17605 613
rect 17484 603 17605 605
rect 17484 483 17496 603
rect 17552 483 17605 603
rect 17484 481 17605 483
rect 17496 473 17552 481
rect 16799 216 17697 228
rect 16799 160 16811 216
rect 16867 160 17629 216
rect 17685 160 17697 216
rect 16799 148 17697 160
rect 15914 42 15926 98
rect 15982 42 15984 98
rect 15914 30 15984 42
rect 16226 98 16286 102
rect 16226 42 16228 98
rect 16284 42 16286 98
rect 16226 30 16286 42
rect 15790 -175 15846 -165
rect 19832 -65 19888 4441
rect 19968 110 20024 8904
rect 20986 8701 21732 8713
rect 20986 8645 21354 8701
rect 21410 8645 21732 8701
rect 20986 8633 21732 8645
rect 20986 8380 21042 8633
rect 21354 8380 21410 8633
rect 21676 8380 21732 8633
rect 20974 8378 21054 8380
rect 20974 8258 20986 8378
rect 21042 8258 21054 8378
rect 20974 8256 21054 8258
rect 21342 8378 21422 8380
rect 21342 8258 21354 8378
rect 21410 8258 21422 8378
rect 21342 8256 21422 8258
rect 21664 8378 21744 8380
rect 21664 8257 21676 8378
rect 21732 8257 21744 8378
rect 20986 8248 21042 8256
rect 21354 8248 21410 8256
rect 21664 8255 21744 8257
rect 21676 8247 21732 8255
rect 21170 8080 21226 8088
rect 21538 8080 21594 8088
rect 21158 8078 21647 8080
rect 21158 7958 21170 8078
rect 21226 7958 21538 8078
rect 21594 7958 21647 8078
rect 21158 7956 21647 7958
rect 21170 7948 21226 7956
rect 21538 7948 21647 7956
rect 21066 7882 21146 7892
rect 21066 7826 21078 7882
rect 21134 7826 21146 7882
rect 21066 7816 21146 7826
rect 21250 7882 21330 7892
rect 21250 7826 21262 7882
rect 21318 7826 21330 7882
rect 21250 7816 21330 7826
rect 21434 7882 21514 7892
rect 21434 7826 21446 7882
rect 21502 7826 21514 7882
rect 21434 7816 21514 7826
rect 20178 7732 20264 7744
rect 21078 7734 21134 7816
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 21066 7732 21146 7734
rect 21066 7676 21078 7732
rect 21134 7676 21146 7732
rect 21066 7674 21146 7676
rect 20394 7616 20464 7628
rect 20394 7560 20406 7616
rect 20462 7560 20464 7616
rect 20394 7548 20464 7560
rect 20258 5411 20328 5425
rect 20258 5355 20270 5411
rect 20326 5355 20328 5411
rect 20258 5343 20328 5355
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 20104 897 20160 5165
rect 20270 1015 20326 5343
rect 20406 3102 20462 7548
rect 21078 7360 21134 7674
rect 21262 7618 21318 7816
rect 21250 7616 21330 7618
rect 21250 7560 21262 7616
rect 21318 7560 21330 7616
rect 21250 7558 21330 7560
rect 21262 7360 21318 7558
rect 21446 7502 21502 7816
rect 21579 7618 21647 7948
rect 21579 7616 21659 7618
rect 21579 7560 21591 7616
rect 21647 7560 21659 7616
rect 21579 7558 21659 7560
rect 21846 7616 21916 7628
rect 21846 7560 21848 7616
rect 21904 7560 21916 7616
rect 21434 7500 21514 7502
rect 21434 7444 21446 7500
rect 21502 7444 21514 7500
rect 21434 7442 21514 7444
rect 21446 7360 21502 7442
rect 21066 7350 21146 7360
rect 21066 7294 21078 7350
rect 21134 7294 21146 7350
rect 21066 7284 21146 7294
rect 21250 7350 21330 7360
rect 21250 7294 21262 7350
rect 21318 7294 21330 7350
rect 21250 7284 21330 7294
rect 21434 7350 21514 7360
rect 21434 7294 21446 7350
rect 21502 7294 21514 7350
rect 21434 7284 21514 7294
rect 21579 7228 21647 7558
rect 21846 7550 21916 7560
rect 21538 7220 21647 7228
rect 21526 7218 21647 7220
rect 21526 7098 21538 7218
rect 21594 7098 21647 7218
rect 21526 7096 21647 7098
rect 21538 7088 21594 7096
rect 20841 6831 21739 6843
rect 20841 6775 20853 6831
rect 20909 6775 21671 6831
rect 21727 6775 21739 6831
rect 20841 6763 21739 6775
rect 21848 6606 21904 7550
rect 22012 6713 22092 6723
rect 22012 6657 22024 6713
rect 22080 6657 22092 6713
rect 22012 6655 22092 6657
rect 21846 6603 21916 6606
rect 21846 6549 21848 6603
rect 21904 6549 21916 6603
rect 21846 6537 21916 6549
rect 20986 6496 21732 6508
rect 20986 6440 21354 6496
rect 21410 6440 21732 6496
rect 20986 6428 21732 6440
rect 20986 6175 21042 6428
rect 21354 6175 21410 6428
rect 21676 6175 21732 6428
rect 20974 6173 21054 6175
rect 20974 6053 20986 6173
rect 21042 6053 21054 6173
rect 20974 6051 21054 6053
rect 21342 6173 21422 6175
rect 21342 6053 21354 6173
rect 21410 6053 21422 6173
rect 21342 6051 21422 6053
rect 21664 6173 21744 6175
rect 21664 6052 21676 6173
rect 21732 6052 21744 6173
rect 20986 6043 21042 6051
rect 21354 6043 21410 6051
rect 21664 6050 21744 6052
rect 21676 6042 21732 6050
rect 21170 5875 21226 5883
rect 21538 5875 21594 5883
rect 21158 5873 21647 5875
rect 21158 5753 21170 5873
rect 21226 5753 21538 5873
rect 21594 5753 21647 5873
rect 21158 5751 21647 5753
rect 21170 5743 21226 5751
rect 21538 5743 21647 5751
rect 21066 5677 21146 5687
rect 21066 5621 21078 5677
rect 21134 5621 21146 5677
rect 21066 5611 21146 5621
rect 21250 5677 21330 5687
rect 21250 5621 21262 5677
rect 21318 5621 21330 5677
rect 21250 5611 21330 5621
rect 21434 5677 21514 5687
rect 21434 5621 21446 5677
rect 21502 5621 21514 5677
rect 21434 5611 21514 5621
rect 21078 5529 21134 5611
rect 21066 5527 21146 5529
rect 21066 5471 21078 5527
rect 21134 5471 21146 5527
rect 21066 5469 21146 5471
rect 21078 5155 21134 5469
rect 21262 5413 21318 5611
rect 21250 5411 21330 5413
rect 21250 5355 21262 5411
rect 21318 5355 21330 5411
rect 21250 5353 21330 5355
rect 21262 5155 21318 5353
rect 21446 5297 21502 5611
rect 21579 5413 21647 5743
rect 22024 5421 22080 6655
rect 22472 6496 23218 6508
rect 22472 6440 22840 6496
rect 22896 6440 23218 6496
rect 22472 6428 23218 6440
rect 22472 6175 22528 6428
rect 22840 6175 22896 6428
rect 23162 6175 23218 6428
rect 22460 6173 22540 6175
rect 22460 6053 22472 6173
rect 22528 6053 22540 6173
rect 22460 6051 22540 6053
rect 22828 6173 22908 6175
rect 22828 6053 22840 6173
rect 22896 6053 22908 6173
rect 22828 6051 22908 6053
rect 23150 6173 23230 6175
rect 23150 6052 23162 6173
rect 23218 6052 23230 6173
rect 22472 6043 22528 6051
rect 22840 6043 22896 6051
rect 23150 6050 23230 6052
rect 23162 6042 23218 6050
rect 22656 5875 22712 5883
rect 23024 5875 23080 5883
rect 22644 5873 23133 5875
rect 22644 5753 22656 5873
rect 22712 5753 23024 5873
rect 23080 5753 23133 5873
rect 22644 5751 23133 5753
rect 22656 5743 22712 5751
rect 23024 5743 23133 5751
rect 22552 5677 22632 5687
rect 22552 5621 22564 5677
rect 22620 5621 22632 5677
rect 22552 5611 22632 5621
rect 22736 5677 22816 5687
rect 22736 5621 22748 5677
rect 22804 5621 22816 5677
rect 22736 5611 22816 5621
rect 22920 5677 23000 5687
rect 22920 5621 22932 5677
rect 22988 5621 23000 5677
rect 22920 5611 23000 5621
rect 22564 5529 22620 5611
rect 22552 5527 22632 5529
rect 22552 5471 22564 5527
rect 22620 5471 22632 5527
rect 22552 5469 22632 5471
rect 21579 5411 21659 5413
rect 21579 5355 21591 5411
rect 21647 5355 21659 5411
rect 21579 5353 21659 5355
rect 22022 5411 22082 5421
rect 22022 5355 22024 5411
rect 22080 5355 22082 5411
rect 21434 5295 21514 5297
rect 21434 5239 21446 5295
rect 21502 5239 21514 5295
rect 21434 5237 21514 5239
rect 21446 5155 21502 5237
rect 21066 5145 21146 5155
rect 21066 5089 21078 5145
rect 21134 5089 21146 5145
rect 21066 5079 21146 5089
rect 21250 5145 21330 5155
rect 21250 5089 21262 5145
rect 21318 5089 21330 5145
rect 21250 5079 21330 5089
rect 21434 5145 21514 5155
rect 21434 5089 21446 5145
rect 21502 5089 21514 5145
rect 21434 5079 21514 5089
rect 21579 5023 21647 5353
rect 22022 5343 22082 5355
rect 21538 5015 21647 5023
rect 21526 5013 21647 5015
rect 21526 4893 21538 5013
rect 21594 4893 21647 5013
rect 21526 4891 21647 4893
rect 21538 4883 21594 4891
rect 20841 4626 21737 4638
rect 20841 4570 20853 4626
rect 20909 4570 21671 4626
rect 21727 4570 21737 4626
rect 20841 4558 21737 4570
rect 22024 4400 22080 5343
rect 22564 5155 22620 5469
rect 22748 5413 22804 5611
rect 22736 5411 22816 5413
rect 22736 5355 22748 5411
rect 22804 5355 22816 5411
rect 22736 5353 22816 5355
rect 22748 5155 22804 5353
rect 22932 5297 22988 5611
rect 23065 5413 23133 5743
rect 23065 5411 23145 5413
rect 23065 5355 23077 5411
rect 23133 5355 23145 5411
rect 23065 5353 23145 5355
rect 23332 5411 23402 5423
rect 23332 5355 23334 5411
rect 23390 5355 23658 5411
rect 22920 5295 23000 5297
rect 22920 5239 22932 5295
rect 22988 5239 23000 5295
rect 22920 5237 23000 5239
rect 22932 5155 22988 5237
rect 22552 5145 22632 5155
rect 22552 5089 22564 5145
rect 22620 5089 22632 5145
rect 22552 5079 22632 5089
rect 22736 5145 22816 5155
rect 22736 5089 22748 5145
rect 22804 5089 22816 5145
rect 22736 5079 22816 5089
rect 22920 5145 23000 5155
rect 22920 5089 22932 5145
rect 22988 5089 23000 5145
rect 22920 5079 23000 5089
rect 23065 5023 23133 5353
rect 23332 5345 23402 5355
rect 23024 5015 23133 5023
rect 23012 5013 23133 5015
rect 23012 4893 23024 5013
rect 23080 4893 23133 5013
rect 23012 4891 23133 4893
rect 23024 4883 23080 4891
rect 22327 4626 23223 4638
rect 22327 4570 22339 4626
rect 22395 4570 23157 4626
rect 23213 4570 23223 4626
rect 22327 4558 23223 4570
rect 23334 4401 23390 5345
rect 23498 4509 23578 4519
rect 23498 4453 23510 4509
rect 23566 4453 23578 4509
rect 23498 4451 23578 4453
rect 22022 4398 22092 4400
rect 22022 4342 22024 4398
rect 22080 4342 22092 4398
rect 22022 4330 22092 4342
rect 23322 4399 23402 4401
rect 23322 4343 23334 4399
rect 23390 4343 23402 4399
rect 23322 4331 23402 4343
rect 20986 4291 21732 4303
rect 20986 4235 21354 4291
rect 21410 4235 21732 4291
rect 20986 4223 21732 4235
rect 20986 3970 21042 4223
rect 21354 3970 21410 4223
rect 21676 3970 21732 4223
rect 22472 4292 23218 4304
rect 22472 4236 22840 4292
rect 22896 4236 23218 4292
rect 22472 4224 23218 4236
rect 22472 3971 22528 4224
rect 22840 3971 22896 4224
rect 23162 3971 23218 4224
rect 20974 3968 21054 3970
rect 20974 3848 20986 3968
rect 21042 3848 21054 3968
rect 20974 3846 21054 3848
rect 21342 3968 21422 3970
rect 21342 3848 21354 3968
rect 21410 3848 21422 3968
rect 21342 3846 21422 3848
rect 21664 3968 21744 3970
rect 21664 3847 21676 3968
rect 21732 3847 21744 3968
rect 22460 3969 22540 3971
rect 22460 3849 22472 3969
rect 22528 3849 22540 3969
rect 22460 3847 22540 3849
rect 22828 3969 22908 3971
rect 22828 3849 22840 3969
rect 22896 3849 22908 3969
rect 22828 3847 22908 3849
rect 23150 3969 23230 3971
rect 23150 3848 23162 3969
rect 23218 3848 23230 3969
rect 20986 3838 21042 3846
rect 21354 3838 21410 3846
rect 21664 3845 21744 3847
rect 21676 3837 21732 3845
rect 22472 3839 22528 3847
rect 22840 3839 22896 3847
rect 23150 3846 23230 3848
rect 23162 3838 23218 3846
rect 21170 3670 21226 3678
rect 21538 3670 21594 3678
rect 22656 3671 22712 3679
rect 23024 3671 23080 3679
rect 21158 3668 21647 3670
rect 21158 3548 21170 3668
rect 21226 3548 21538 3668
rect 21594 3548 21647 3668
rect 21158 3546 21647 3548
rect 22644 3669 23133 3671
rect 22644 3549 22656 3669
rect 22712 3549 23024 3669
rect 23080 3549 23133 3669
rect 22644 3547 23133 3549
rect 21170 3538 21226 3546
rect 21538 3538 21647 3546
rect 22656 3539 22712 3547
rect 23024 3539 23133 3547
rect 21066 3472 21146 3482
rect 21066 3416 21078 3472
rect 21134 3416 21146 3472
rect 21066 3406 21146 3416
rect 21250 3472 21330 3482
rect 21250 3416 21262 3472
rect 21318 3416 21330 3472
rect 21250 3406 21330 3416
rect 21434 3472 21514 3482
rect 21434 3416 21446 3472
rect 21502 3416 21514 3472
rect 21434 3406 21514 3416
rect 21078 3324 21134 3406
rect 21066 3322 21146 3324
rect 21066 3266 21078 3322
rect 21134 3266 21146 3322
rect 21066 3264 21146 3266
rect 20394 3090 20464 3102
rect 20394 3034 20406 3090
rect 20462 3034 20464 3090
rect 20394 3022 20464 3034
rect 21078 2950 21134 3264
rect 21262 3208 21318 3406
rect 21250 3206 21330 3208
rect 21250 3150 21262 3206
rect 21318 3150 21330 3206
rect 21250 3148 21330 3150
rect 21262 2950 21318 3148
rect 21446 3092 21502 3406
rect 21579 3208 21647 3538
rect 22552 3473 22632 3483
rect 22552 3417 22564 3473
rect 22620 3417 22632 3473
rect 22552 3407 22632 3417
rect 22736 3473 22816 3483
rect 22736 3417 22748 3473
rect 22804 3417 22816 3473
rect 22736 3407 22816 3417
rect 22920 3473 23000 3483
rect 22920 3417 22932 3473
rect 22988 3417 23000 3473
rect 22920 3407 23000 3417
rect 22564 3325 22620 3407
rect 22552 3323 22632 3325
rect 22552 3267 22564 3323
rect 22620 3267 22632 3323
rect 22552 3265 22632 3267
rect 21579 3206 21659 3208
rect 21579 3150 21591 3206
rect 21647 3150 21659 3206
rect 21579 3148 21659 3150
rect 21846 3206 21916 3218
rect 21846 3150 21848 3206
rect 21904 3150 21916 3206
rect 21434 3090 21514 3092
rect 21434 3034 21446 3090
rect 21502 3034 21514 3090
rect 21434 3032 21514 3034
rect 21446 2950 21502 3032
rect 21066 2940 21146 2950
rect 21066 2884 21078 2940
rect 21134 2884 21146 2940
rect 21066 2874 21146 2884
rect 21250 2940 21330 2950
rect 21250 2884 21262 2940
rect 21318 2884 21330 2940
rect 21250 2874 21330 2884
rect 21434 2940 21514 2950
rect 21434 2884 21446 2940
rect 21502 2884 21514 2940
rect 21434 2874 21514 2884
rect 21579 2818 21647 3148
rect 21846 3140 21916 3150
rect 21538 2810 21647 2818
rect 21526 2808 21647 2810
rect 21526 2688 21538 2808
rect 21594 2688 21647 2808
rect 21526 2686 21647 2688
rect 21538 2678 21594 2686
rect 20841 2421 21737 2433
rect 20841 2365 20853 2421
rect 20909 2365 21671 2421
rect 21727 2365 21737 2421
rect 20841 2353 21737 2365
rect 21848 2196 21904 3140
rect 22564 2951 22620 3265
rect 22748 3209 22804 3407
rect 22736 3207 22816 3209
rect 22736 3151 22748 3207
rect 22804 3151 22816 3207
rect 22736 3149 22816 3151
rect 22748 2951 22804 3149
rect 22932 3093 22988 3407
rect 23065 3209 23133 3539
rect 23510 3217 23566 4451
rect 23065 3207 23145 3209
rect 23065 3151 23077 3207
rect 23133 3151 23145 3207
rect 23065 3149 23145 3151
rect 23508 3207 23578 3217
rect 23738 3207 23794 17250
rect 23940 14999 23996 18855
rect 27982 18739 28038 19501
rect 27980 18737 28050 18739
rect 27980 18681 27982 18737
rect 28038 18681 28050 18737
rect 27980 18679 28050 18681
rect 24164 18561 24234 18573
rect 24164 18505 24176 18561
rect 24232 18505 24234 18561
rect 24164 18503 24234 18505
rect 23938 14987 24008 14999
rect 23938 14931 23940 14987
rect 23996 14931 24008 14987
rect 23938 14919 24008 14931
rect 24176 14087 24232 18503
rect 25028 18277 25774 18289
rect 25028 18221 25396 18277
rect 25452 18221 25774 18277
rect 25028 18209 25774 18221
rect 25028 17956 25084 18209
rect 25396 17956 25452 18209
rect 25718 17956 25774 18209
rect 25016 17954 25096 17956
rect 25016 17834 25028 17954
rect 25084 17834 25096 17954
rect 25016 17832 25096 17834
rect 25384 17954 25464 17956
rect 25384 17834 25396 17954
rect 25452 17834 25464 17954
rect 25384 17832 25464 17834
rect 25706 17954 25786 17956
rect 25706 17833 25718 17954
rect 25774 17833 25786 17954
rect 25028 17824 25084 17832
rect 25396 17824 25452 17832
rect 25706 17831 25786 17833
rect 25718 17823 25774 17831
rect 25212 17656 25268 17664
rect 25580 17656 25636 17664
rect 25200 17654 25689 17656
rect 25200 17534 25212 17654
rect 25268 17534 25580 17654
rect 25636 17534 25689 17654
rect 25200 17532 25689 17534
rect 25212 17524 25268 17532
rect 25580 17524 25689 17532
rect 25108 17458 25188 17468
rect 25108 17402 25120 17458
rect 25176 17402 25188 17458
rect 25108 17392 25188 17402
rect 25292 17458 25372 17468
rect 25292 17402 25304 17458
rect 25360 17402 25372 17458
rect 25292 17392 25372 17402
rect 25476 17458 25556 17468
rect 25476 17402 25488 17458
rect 25544 17402 25556 17458
rect 25476 17392 25556 17402
rect 25120 17310 25176 17392
rect 25108 17308 25188 17310
rect 25108 17252 25120 17308
rect 25176 17252 25188 17308
rect 25108 17250 25188 17252
rect 24436 17192 24506 17204
rect 24436 17136 24448 17192
rect 24504 17136 24506 17192
rect 24436 17124 24506 17136
rect 24300 14987 24370 15001
rect 24300 14931 24312 14987
rect 24368 14931 24370 14987
rect 24300 14919 24370 14931
rect 24164 14085 24234 14087
rect 24164 14029 24176 14085
rect 24232 14029 24234 14085
rect 24164 14017 24234 14029
rect 24312 10591 24368 14919
rect 24448 12678 24504 17124
rect 25120 16936 25176 17250
rect 25304 17194 25360 17392
rect 25292 17192 25372 17194
rect 25292 17136 25304 17192
rect 25360 17136 25372 17192
rect 25292 17134 25372 17136
rect 25304 16936 25360 17134
rect 25488 17078 25544 17392
rect 25621 17194 25689 17524
rect 27768 17308 27848 17320
rect 27768 17252 27780 17308
rect 27836 17252 27848 17308
rect 27768 17250 27848 17252
rect 25621 17192 25701 17194
rect 25621 17136 25633 17192
rect 25689 17136 25701 17192
rect 25621 17134 25701 17136
rect 25888 17192 25958 17204
rect 25888 17136 25890 17192
rect 25946 17136 25958 17192
rect 25476 17076 25556 17078
rect 25476 17020 25488 17076
rect 25544 17020 25556 17076
rect 25476 17018 25556 17020
rect 25488 16936 25544 17018
rect 25108 16926 25188 16936
rect 25108 16870 25120 16926
rect 25176 16870 25188 16926
rect 25108 16860 25188 16870
rect 25292 16926 25372 16936
rect 25292 16870 25304 16926
rect 25360 16870 25372 16926
rect 25292 16860 25372 16870
rect 25476 16926 25556 16936
rect 25476 16870 25488 16926
rect 25544 16870 25556 16926
rect 25476 16860 25556 16870
rect 25621 16804 25689 17134
rect 25888 17126 25958 17136
rect 25580 16796 25689 16804
rect 25568 16794 25689 16796
rect 25568 16674 25580 16794
rect 25636 16674 25689 16794
rect 25568 16672 25689 16674
rect 25580 16664 25636 16672
rect 24883 16407 25781 16419
rect 24883 16351 24895 16407
rect 24951 16351 25713 16407
rect 25769 16351 25781 16407
rect 24883 16339 25781 16351
rect 25890 16182 25946 17126
rect 26054 16289 26134 16299
rect 26054 16233 26066 16289
rect 26122 16233 26134 16289
rect 26054 16231 26134 16233
rect 25888 16179 25958 16182
rect 25888 16125 25890 16179
rect 25946 16125 25958 16179
rect 25888 16113 25958 16125
rect 25028 16072 25774 16084
rect 25028 16016 25396 16072
rect 25452 16016 25774 16072
rect 25028 16004 25774 16016
rect 25028 15751 25084 16004
rect 25396 15751 25452 16004
rect 25718 15751 25774 16004
rect 25016 15749 25096 15751
rect 25016 15629 25028 15749
rect 25084 15629 25096 15749
rect 25016 15627 25096 15629
rect 25384 15749 25464 15751
rect 25384 15629 25396 15749
rect 25452 15629 25464 15749
rect 25384 15627 25464 15629
rect 25706 15749 25786 15751
rect 25706 15628 25718 15749
rect 25774 15628 25786 15749
rect 25028 15619 25084 15627
rect 25396 15619 25452 15627
rect 25706 15626 25786 15628
rect 25718 15618 25774 15626
rect 25212 15451 25268 15459
rect 25580 15451 25636 15459
rect 25200 15449 25689 15451
rect 25200 15329 25212 15449
rect 25268 15329 25580 15449
rect 25636 15329 25689 15449
rect 25200 15327 25689 15329
rect 25212 15319 25268 15327
rect 25580 15319 25689 15327
rect 25108 15253 25188 15263
rect 25108 15197 25120 15253
rect 25176 15197 25188 15253
rect 25108 15187 25188 15197
rect 25292 15253 25372 15263
rect 25292 15197 25304 15253
rect 25360 15197 25372 15253
rect 25292 15187 25372 15197
rect 25476 15253 25556 15263
rect 25476 15197 25488 15253
rect 25544 15197 25556 15253
rect 25476 15187 25556 15197
rect 25120 15105 25176 15187
rect 25108 15103 25188 15105
rect 25108 15047 25120 15103
rect 25176 15047 25188 15103
rect 25108 15045 25188 15047
rect 25120 14731 25176 15045
rect 25304 14989 25360 15187
rect 25292 14987 25372 14989
rect 25292 14931 25304 14987
rect 25360 14931 25372 14987
rect 25292 14929 25372 14931
rect 25304 14731 25360 14929
rect 25488 14873 25544 15187
rect 25621 14989 25689 15319
rect 26066 14997 26122 16231
rect 26514 16072 27260 16084
rect 26514 16016 26882 16072
rect 26938 16016 27260 16072
rect 26514 16004 27260 16016
rect 26514 15751 26570 16004
rect 26882 15751 26938 16004
rect 27204 15751 27260 16004
rect 26502 15749 26582 15751
rect 26502 15629 26514 15749
rect 26570 15629 26582 15749
rect 26502 15627 26582 15629
rect 26870 15749 26950 15751
rect 26870 15629 26882 15749
rect 26938 15629 26950 15749
rect 26870 15627 26950 15629
rect 27192 15749 27272 15751
rect 27192 15628 27204 15749
rect 27260 15628 27272 15749
rect 26514 15619 26570 15627
rect 26882 15619 26938 15627
rect 27192 15626 27272 15628
rect 27204 15618 27260 15626
rect 26698 15451 26754 15459
rect 27066 15451 27122 15459
rect 26686 15449 27175 15451
rect 26686 15329 26698 15449
rect 26754 15329 27066 15449
rect 27122 15329 27175 15449
rect 26686 15327 27175 15329
rect 26698 15319 26754 15327
rect 27066 15319 27175 15327
rect 26594 15253 26674 15263
rect 26594 15197 26606 15253
rect 26662 15197 26674 15253
rect 26594 15187 26674 15197
rect 26778 15253 26858 15263
rect 26778 15197 26790 15253
rect 26846 15197 26858 15253
rect 26778 15187 26858 15197
rect 26962 15253 27042 15263
rect 26962 15197 26974 15253
rect 27030 15197 27042 15253
rect 26962 15187 27042 15197
rect 26606 15105 26662 15187
rect 26594 15103 26674 15105
rect 26594 15047 26606 15103
rect 26662 15047 26674 15103
rect 26594 15045 26674 15047
rect 25621 14987 25701 14989
rect 25621 14931 25633 14987
rect 25689 14931 25701 14987
rect 25621 14929 25701 14931
rect 26064 14987 26124 14997
rect 26064 14931 26066 14987
rect 26122 14931 26124 14987
rect 25476 14871 25556 14873
rect 25476 14815 25488 14871
rect 25544 14815 25556 14871
rect 25476 14813 25556 14815
rect 25488 14731 25544 14813
rect 25108 14721 25188 14731
rect 25108 14665 25120 14721
rect 25176 14665 25188 14721
rect 25108 14655 25188 14665
rect 25292 14721 25372 14731
rect 25292 14665 25304 14721
rect 25360 14665 25372 14721
rect 25292 14655 25372 14665
rect 25476 14721 25556 14731
rect 25476 14665 25488 14721
rect 25544 14665 25556 14721
rect 25476 14655 25556 14665
rect 25621 14599 25689 14929
rect 26064 14919 26124 14931
rect 25580 14591 25689 14599
rect 25568 14589 25689 14591
rect 25568 14469 25580 14589
rect 25636 14469 25689 14589
rect 25568 14467 25689 14469
rect 25580 14459 25636 14467
rect 24883 14202 25779 14214
rect 24883 14146 24895 14202
rect 24951 14146 25713 14202
rect 25769 14146 25779 14202
rect 24883 14134 25779 14146
rect 26066 13976 26122 14919
rect 26606 14731 26662 15045
rect 26790 14989 26846 15187
rect 26778 14987 26858 14989
rect 26778 14931 26790 14987
rect 26846 14931 26858 14987
rect 26778 14929 26858 14931
rect 26790 14731 26846 14929
rect 26974 14873 27030 15187
rect 27107 14989 27175 15319
rect 27107 14987 27187 14989
rect 27107 14931 27119 14987
rect 27175 14931 27187 14987
rect 27107 14929 27187 14931
rect 27374 14987 27444 14999
rect 27374 14931 27376 14987
rect 27432 14931 27700 14987
rect 26962 14871 27042 14873
rect 26962 14815 26974 14871
rect 27030 14815 27042 14871
rect 26962 14813 27042 14815
rect 26974 14731 27030 14813
rect 26594 14721 26674 14731
rect 26594 14665 26606 14721
rect 26662 14665 26674 14721
rect 26594 14655 26674 14665
rect 26778 14721 26858 14731
rect 26778 14665 26790 14721
rect 26846 14665 26858 14721
rect 26778 14655 26858 14665
rect 26962 14721 27042 14731
rect 26962 14665 26974 14721
rect 27030 14665 27042 14721
rect 26962 14655 27042 14665
rect 27107 14599 27175 14929
rect 27374 14921 27444 14931
rect 27066 14591 27175 14599
rect 27054 14589 27175 14591
rect 27054 14469 27066 14589
rect 27122 14469 27175 14589
rect 27054 14467 27175 14469
rect 27066 14459 27122 14467
rect 26369 14202 27265 14214
rect 26369 14146 26381 14202
rect 26437 14146 27199 14202
rect 27255 14146 27265 14202
rect 26369 14134 27265 14146
rect 27376 13977 27432 14921
rect 27540 14085 27620 14095
rect 27540 14029 27552 14085
rect 27608 14029 27620 14085
rect 27540 14027 27620 14029
rect 26064 13974 26134 13976
rect 26064 13918 26066 13974
rect 26122 13918 26134 13974
rect 26064 13906 26134 13918
rect 27364 13975 27444 13977
rect 27364 13919 27376 13975
rect 27432 13919 27444 13975
rect 27364 13907 27444 13919
rect 25028 13867 25774 13879
rect 25028 13811 25396 13867
rect 25452 13811 25774 13867
rect 25028 13799 25774 13811
rect 25028 13546 25084 13799
rect 25396 13546 25452 13799
rect 25718 13546 25774 13799
rect 26514 13868 27260 13880
rect 26514 13812 26882 13868
rect 26938 13812 27260 13868
rect 26514 13800 27260 13812
rect 26514 13547 26570 13800
rect 26882 13547 26938 13800
rect 27204 13547 27260 13800
rect 25016 13544 25096 13546
rect 25016 13424 25028 13544
rect 25084 13424 25096 13544
rect 25016 13422 25096 13424
rect 25384 13544 25464 13546
rect 25384 13424 25396 13544
rect 25452 13424 25464 13544
rect 25384 13422 25464 13424
rect 25706 13544 25786 13546
rect 25706 13423 25718 13544
rect 25774 13423 25786 13544
rect 26502 13545 26582 13547
rect 26502 13425 26514 13545
rect 26570 13425 26582 13545
rect 26502 13423 26582 13425
rect 26870 13545 26950 13547
rect 26870 13425 26882 13545
rect 26938 13425 26950 13545
rect 26870 13423 26950 13425
rect 27192 13545 27272 13547
rect 27192 13424 27204 13545
rect 27260 13424 27272 13545
rect 25028 13414 25084 13422
rect 25396 13414 25452 13422
rect 25706 13421 25786 13423
rect 25718 13413 25774 13421
rect 26514 13415 26570 13423
rect 26882 13415 26938 13423
rect 27192 13422 27272 13424
rect 27204 13414 27260 13422
rect 25212 13246 25268 13254
rect 25580 13246 25636 13254
rect 26698 13247 26754 13255
rect 27066 13247 27122 13255
rect 25200 13244 25689 13246
rect 25200 13124 25212 13244
rect 25268 13124 25580 13244
rect 25636 13124 25689 13244
rect 25200 13122 25689 13124
rect 26686 13245 27175 13247
rect 26686 13125 26698 13245
rect 26754 13125 27066 13245
rect 27122 13125 27175 13245
rect 26686 13123 27175 13125
rect 25212 13114 25268 13122
rect 25580 13114 25689 13122
rect 26698 13115 26754 13123
rect 27066 13115 27175 13123
rect 25108 13048 25188 13058
rect 25108 12992 25120 13048
rect 25176 12992 25188 13048
rect 25108 12982 25188 12992
rect 25292 13048 25372 13058
rect 25292 12992 25304 13048
rect 25360 12992 25372 13048
rect 25292 12982 25372 12992
rect 25476 13048 25556 13058
rect 25476 12992 25488 13048
rect 25544 12992 25556 13048
rect 25476 12982 25556 12992
rect 25120 12900 25176 12982
rect 25108 12898 25188 12900
rect 25108 12842 25120 12898
rect 25176 12842 25188 12898
rect 25108 12840 25188 12842
rect 24436 12666 24506 12678
rect 24436 12610 24448 12666
rect 24504 12610 24506 12666
rect 24436 12598 24506 12610
rect 25120 12526 25176 12840
rect 25304 12784 25360 12982
rect 25292 12782 25372 12784
rect 25292 12726 25304 12782
rect 25360 12726 25372 12782
rect 25292 12724 25372 12726
rect 25304 12526 25360 12724
rect 25488 12668 25544 12982
rect 25621 12784 25689 13114
rect 26594 13049 26674 13059
rect 26594 12993 26606 13049
rect 26662 12993 26674 13049
rect 26594 12983 26674 12993
rect 26778 13049 26858 13059
rect 26778 12993 26790 13049
rect 26846 12993 26858 13049
rect 26778 12983 26858 12993
rect 26962 13049 27042 13059
rect 26962 12993 26974 13049
rect 27030 12993 27042 13049
rect 26962 12983 27042 12993
rect 26606 12901 26662 12983
rect 26594 12899 26674 12901
rect 26594 12843 26606 12899
rect 26662 12843 26674 12899
rect 26594 12841 26674 12843
rect 25621 12782 25701 12784
rect 25621 12726 25633 12782
rect 25689 12726 25701 12782
rect 25621 12724 25701 12726
rect 25888 12782 25958 12794
rect 25888 12726 25890 12782
rect 25946 12726 25958 12782
rect 25476 12666 25556 12668
rect 25476 12610 25488 12666
rect 25544 12610 25556 12666
rect 25476 12608 25556 12610
rect 25488 12526 25544 12608
rect 25108 12516 25188 12526
rect 25108 12460 25120 12516
rect 25176 12460 25188 12516
rect 25108 12450 25188 12460
rect 25292 12516 25372 12526
rect 25292 12460 25304 12516
rect 25360 12460 25372 12516
rect 25292 12450 25372 12460
rect 25476 12516 25556 12526
rect 25476 12460 25488 12516
rect 25544 12460 25556 12516
rect 25476 12450 25556 12460
rect 25621 12394 25689 12724
rect 25888 12716 25958 12726
rect 25580 12386 25689 12394
rect 25568 12384 25689 12386
rect 25568 12264 25580 12384
rect 25636 12264 25689 12384
rect 25568 12262 25689 12264
rect 25580 12254 25636 12262
rect 24883 11997 25779 12009
rect 24883 11941 24895 11997
rect 24951 11941 25713 11997
rect 25769 11941 25779 11997
rect 24883 11929 25779 11941
rect 25890 11772 25946 12716
rect 26606 12527 26662 12841
rect 26790 12785 26846 12983
rect 26778 12783 26858 12785
rect 26778 12727 26790 12783
rect 26846 12727 26858 12783
rect 26778 12725 26858 12727
rect 26790 12527 26846 12725
rect 26974 12669 27030 12983
rect 27107 12785 27175 13115
rect 27552 12793 27608 14027
rect 27107 12783 27187 12785
rect 27107 12727 27119 12783
rect 27175 12727 27187 12783
rect 27107 12725 27187 12727
rect 27550 12783 27620 12793
rect 27550 12727 27552 12783
rect 27608 12727 27700 12783
rect 26962 12667 27042 12669
rect 26962 12611 26974 12667
rect 27030 12611 27042 12667
rect 26962 12609 27042 12611
rect 26974 12527 27030 12609
rect 26594 12517 26674 12527
rect 26594 12461 26606 12517
rect 26662 12461 26674 12517
rect 26594 12451 26674 12461
rect 26778 12517 26858 12527
rect 26778 12461 26790 12517
rect 26846 12461 26858 12517
rect 26778 12451 26858 12461
rect 26962 12517 27042 12527
rect 26962 12461 26974 12517
rect 27030 12461 27042 12517
rect 26962 12451 27042 12461
rect 27107 12395 27175 12725
rect 27550 12715 27620 12727
rect 27066 12387 27175 12395
rect 27054 12385 27175 12387
rect 27054 12265 27066 12385
rect 27122 12265 27175 12385
rect 27054 12263 27175 12265
rect 27066 12255 27122 12263
rect 26369 11998 27265 12010
rect 26369 11942 26381 11998
rect 26437 11942 27199 11998
rect 27255 11942 27265 11998
rect 26369 11930 27265 11942
rect 26054 11879 26134 11889
rect 26054 11823 26066 11879
rect 26122 11823 26134 11879
rect 26054 11821 26134 11823
rect 25888 11769 25958 11772
rect 25888 11715 25890 11769
rect 25946 11715 25958 11769
rect 25888 11703 25958 11715
rect 25028 11662 25774 11674
rect 25028 11606 25396 11662
rect 25452 11606 25774 11662
rect 25028 11594 25774 11606
rect 25028 11341 25084 11594
rect 25396 11341 25452 11594
rect 25718 11341 25774 11594
rect 25016 11339 25096 11341
rect 25016 11219 25028 11339
rect 25084 11219 25096 11339
rect 25016 11217 25096 11219
rect 25384 11339 25464 11341
rect 25384 11219 25396 11339
rect 25452 11219 25464 11339
rect 25384 11217 25464 11219
rect 25706 11339 25786 11341
rect 25706 11218 25718 11339
rect 25774 11218 25786 11339
rect 25028 11209 25084 11217
rect 25396 11209 25452 11217
rect 25706 11216 25786 11218
rect 25718 11208 25774 11216
rect 25212 11041 25268 11049
rect 25580 11041 25636 11049
rect 25200 11039 25689 11041
rect 25200 10919 25212 11039
rect 25268 10919 25580 11039
rect 25636 10919 25689 11039
rect 25200 10917 25689 10919
rect 25212 10909 25268 10917
rect 25580 10909 25689 10917
rect 25108 10843 25188 10853
rect 25108 10787 25120 10843
rect 25176 10787 25188 10843
rect 25108 10777 25188 10787
rect 25292 10843 25372 10853
rect 25292 10787 25304 10843
rect 25360 10787 25372 10843
rect 25292 10777 25372 10787
rect 25476 10843 25556 10853
rect 25476 10787 25488 10843
rect 25544 10787 25556 10843
rect 25476 10777 25556 10787
rect 25120 10695 25176 10777
rect 25108 10693 25188 10695
rect 25108 10637 25120 10693
rect 25176 10637 25188 10693
rect 25108 10635 25188 10637
rect 24300 10577 24370 10591
rect 24300 10521 24312 10577
rect 24368 10521 24370 10577
rect 24300 10509 24370 10521
rect 23998 9674 24068 9686
rect 24312 9678 24368 10509
rect 25120 10321 25176 10635
rect 25304 10579 25360 10777
rect 25292 10577 25372 10579
rect 25292 10521 25304 10577
rect 25360 10521 25372 10577
rect 25292 10519 25372 10521
rect 25304 10321 25360 10519
rect 25488 10463 25544 10777
rect 25621 10579 25689 10909
rect 26066 10589 26122 11821
rect 25621 10577 25701 10579
rect 25621 10521 25633 10577
rect 25689 10521 25701 10577
rect 25621 10519 25701 10521
rect 26064 10577 26124 10589
rect 26064 10521 26066 10577
rect 26122 10521 26124 10577
rect 25476 10461 25556 10463
rect 25476 10405 25488 10461
rect 25544 10405 25556 10461
rect 25476 10403 25556 10405
rect 25488 10321 25544 10403
rect 25108 10311 25188 10321
rect 25108 10255 25120 10311
rect 25176 10255 25188 10311
rect 25108 10245 25188 10255
rect 25292 10311 25372 10321
rect 25292 10255 25304 10311
rect 25360 10255 25372 10311
rect 25292 10245 25372 10255
rect 25476 10311 25556 10321
rect 25476 10255 25488 10311
rect 25544 10255 25556 10311
rect 25476 10245 25556 10255
rect 25621 10189 25689 10519
rect 26064 10509 26124 10521
rect 25580 10181 25689 10189
rect 25568 10179 25689 10181
rect 25568 10059 25580 10179
rect 25636 10059 25689 10179
rect 25568 10057 25689 10059
rect 25580 10049 25636 10057
rect 24883 9792 25781 9804
rect 24883 9736 24895 9792
rect 24951 9736 25713 9792
rect 25769 9736 25781 9792
rect 24883 9724 25781 9736
rect 23998 9618 24010 9674
rect 24066 9618 24068 9674
rect 23998 9616 24068 9618
rect 24310 9674 24370 9678
rect 24310 9618 24312 9674
rect 24368 9618 24370 9674
rect 24010 9004 24066 9616
rect 24310 9606 24370 9618
rect 23862 4509 23932 4521
rect 23862 4453 23874 4509
rect 23930 4453 23932 4509
rect 23862 4441 23932 4453
rect 23508 3151 23510 3207
rect 23566 3151 23794 3207
rect 22920 3091 23000 3093
rect 22920 3035 22932 3091
rect 22988 3035 23000 3091
rect 22920 3033 23000 3035
rect 22932 2951 22988 3033
rect 22552 2941 22632 2951
rect 22552 2885 22564 2941
rect 22620 2885 22632 2941
rect 22552 2875 22632 2885
rect 22736 2941 22816 2951
rect 22736 2885 22748 2941
rect 22804 2885 22816 2941
rect 22736 2875 22816 2885
rect 22920 2941 23000 2951
rect 22920 2885 22932 2941
rect 22988 2885 23000 2941
rect 22920 2875 23000 2885
rect 23065 2819 23133 3149
rect 23508 3139 23578 3151
rect 23024 2811 23133 2819
rect 23012 2809 23133 2811
rect 23012 2689 23024 2809
rect 23080 2689 23133 2809
rect 23012 2687 23133 2689
rect 23024 2679 23080 2687
rect 22327 2422 23223 2434
rect 22327 2366 22339 2422
rect 22395 2366 23157 2422
rect 23213 2366 23223 2422
rect 22327 2354 23223 2366
rect 22012 2303 22092 2313
rect 22012 2247 22024 2303
rect 22080 2247 22092 2303
rect 22012 2245 22092 2247
rect 21846 2193 21916 2196
rect 21846 2139 21848 2193
rect 21904 2139 21916 2193
rect 21846 2127 21916 2139
rect 20986 2086 21732 2098
rect 20986 2030 21354 2086
rect 21410 2030 21732 2086
rect 20986 2018 21732 2030
rect 20986 1765 21042 2018
rect 21354 1765 21410 2018
rect 21676 1765 21732 2018
rect 20974 1763 21054 1765
rect 20974 1643 20986 1763
rect 21042 1643 21054 1763
rect 20974 1641 21054 1643
rect 21342 1763 21422 1765
rect 21342 1643 21354 1763
rect 21410 1643 21422 1763
rect 21342 1641 21422 1643
rect 21664 1763 21744 1765
rect 21664 1642 21676 1763
rect 21732 1642 21744 1763
rect 20986 1633 21042 1641
rect 21354 1633 21410 1641
rect 21664 1640 21744 1642
rect 21676 1632 21732 1640
rect 21170 1465 21226 1473
rect 21538 1465 21594 1473
rect 21158 1463 21647 1465
rect 21158 1343 21170 1463
rect 21226 1343 21538 1463
rect 21594 1343 21647 1463
rect 21158 1341 21647 1343
rect 21170 1333 21226 1341
rect 21538 1333 21647 1341
rect 21066 1267 21146 1277
rect 21066 1211 21078 1267
rect 21134 1211 21146 1267
rect 21066 1201 21146 1211
rect 21250 1267 21330 1277
rect 21250 1211 21262 1267
rect 21318 1211 21330 1267
rect 21250 1201 21330 1211
rect 21434 1267 21514 1277
rect 21434 1211 21446 1267
rect 21502 1211 21514 1267
rect 21434 1201 21514 1211
rect 21078 1119 21134 1201
rect 21066 1117 21146 1119
rect 21066 1061 21078 1117
rect 21134 1061 21146 1117
rect 21066 1059 21146 1061
rect 20258 1001 20328 1015
rect 20258 945 20270 1001
rect 20326 945 20328 1001
rect 20258 933 20328 945
rect 20092 885 20172 897
rect 20092 829 20104 885
rect 20160 829 20172 885
rect 20092 817 20172 829
rect 19956 98 20026 110
rect 20270 102 20326 933
rect 21078 745 21134 1059
rect 21262 1003 21318 1201
rect 21250 1001 21330 1003
rect 21250 945 21262 1001
rect 21318 945 21330 1001
rect 21250 943 21330 945
rect 21262 745 21318 943
rect 21446 887 21502 1201
rect 21579 1003 21647 1333
rect 22024 1013 22080 2245
rect 21579 1001 21659 1003
rect 21579 945 21591 1001
rect 21647 945 21659 1001
rect 21579 943 21659 945
rect 22022 1001 22082 1013
rect 22022 945 22024 1001
rect 22080 945 22082 1001
rect 21434 885 21514 887
rect 21434 829 21446 885
rect 21502 829 21514 885
rect 21434 827 21514 829
rect 21446 745 21502 827
rect 21066 735 21146 745
rect 21066 679 21078 735
rect 21134 679 21146 735
rect 21066 669 21146 679
rect 21250 735 21330 745
rect 21250 679 21262 735
rect 21318 679 21330 735
rect 21250 669 21330 679
rect 21434 735 21514 745
rect 21434 679 21446 735
rect 21502 679 21514 735
rect 21434 669 21514 679
rect 21579 613 21647 943
rect 22022 933 22082 945
rect 21538 605 21647 613
rect 21526 603 21647 605
rect 21526 483 21538 603
rect 21594 483 21647 603
rect 21526 481 21647 483
rect 21538 473 21594 481
rect 20841 216 21739 228
rect 20841 160 20853 216
rect 20909 160 21671 216
rect 21727 160 21739 216
rect 20841 148 21739 160
rect 19956 42 19968 98
rect 20024 42 20026 98
rect 19956 30 20026 42
rect 20268 98 20328 102
rect 20268 42 20270 98
rect 20326 42 20328 98
rect 20268 30 20328 42
rect 19832 -175 19888 -165
rect 23874 -65 23930 4441
rect 24010 110 24066 8904
rect 25028 8701 25774 8713
rect 25028 8645 25396 8701
rect 25452 8645 25774 8701
rect 25028 8633 25774 8645
rect 25028 8380 25084 8633
rect 25396 8380 25452 8633
rect 25718 8380 25774 8633
rect 25016 8378 25096 8380
rect 25016 8258 25028 8378
rect 25084 8258 25096 8378
rect 25016 8256 25096 8258
rect 25384 8378 25464 8380
rect 25384 8258 25396 8378
rect 25452 8258 25464 8378
rect 25384 8256 25464 8258
rect 25706 8378 25786 8380
rect 25706 8257 25718 8378
rect 25774 8257 25786 8378
rect 25028 8248 25084 8256
rect 25396 8248 25452 8256
rect 25706 8255 25786 8257
rect 25718 8247 25774 8255
rect 25212 8080 25268 8088
rect 25580 8080 25636 8088
rect 25200 8078 25689 8080
rect 25200 7958 25212 8078
rect 25268 7958 25580 8078
rect 25636 7958 25689 8078
rect 25200 7956 25689 7958
rect 25212 7948 25268 7956
rect 25580 7948 25689 7956
rect 25108 7882 25188 7892
rect 25108 7826 25120 7882
rect 25176 7826 25188 7882
rect 25108 7816 25188 7826
rect 25292 7882 25372 7892
rect 25292 7826 25304 7882
rect 25360 7826 25372 7882
rect 25292 7816 25372 7826
rect 25476 7882 25556 7892
rect 25476 7826 25488 7882
rect 25544 7826 25556 7882
rect 25476 7816 25556 7826
rect 24220 7732 24306 7744
rect 25120 7734 25176 7816
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 25108 7732 25188 7734
rect 25108 7676 25120 7732
rect 25176 7676 25188 7732
rect 25108 7674 25188 7676
rect 24436 7616 24506 7628
rect 24436 7560 24448 7616
rect 24504 7560 24506 7616
rect 24436 7548 24506 7560
rect 24300 5411 24370 5425
rect 24300 5355 24312 5411
rect 24368 5355 24370 5411
rect 24300 5343 24370 5355
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect 24146 897 24202 5165
rect 24312 1015 24368 5343
rect 24448 3102 24504 7548
rect 25120 7360 25176 7674
rect 25304 7618 25360 7816
rect 25292 7616 25372 7618
rect 25292 7560 25304 7616
rect 25360 7560 25372 7616
rect 25292 7558 25372 7560
rect 25304 7360 25360 7558
rect 25488 7502 25544 7816
rect 25621 7618 25689 7948
rect 25621 7616 25701 7618
rect 25621 7560 25633 7616
rect 25689 7560 25701 7616
rect 25621 7558 25701 7560
rect 25888 7616 25958 7628
rect 25888 7560 25890 7616
rect 25946 7560 25958 7616
rect 25476 7500 25556 7502
rect 25476 7444 25488 7500
rect 25544 7444 25556 7500
rect 25476 7442 25556 7444
rect 25488 7360 25544 7442
rect 25108 7350 25188 7360
rect 25108 7294 25120 7350
rect 25176 7294 25188 7350
rect 25108 7284 25188 7294
rect 25292 7350 25372 7360
rect 25292 7294 25304 7350
rect 25360 7294 25372 7350
rect 25292 7284 25372 7294
rect 25476 7350 25556 7360
rect 25476 7294 25488 7350
rect 25544 7294 25556 7350
rect 25476 7284 25556 7294
rect 25621 7228 25689 7558
rect 25888 7550 25958 7560
rect 25580 7220 25689 7228
rect 25568 7218 25689 7220
rect 25568 7098 25580 7218
rect 25636 7098 25689 7218
rect 25568 7096 25689 7098
rect 25580 7088 25636 7096
rect 24883 6831 25781 6843
rect 24883 6775 24895 6831
rect 24951 6775 25713 6831
rect 25769 6775 25781 6831
rect 24883 6763 25781 6775
rect 25890 6606 25946 7550
rect 26054 6713 26134 6723
rect 26054 6657 26066 6713
rect 26122 6657 26134 6713
rect 26054 6655 26134 6657
rect 25888 6603 25958 6606
rect 25888 6549 25890 6603
rect 25946 6549 25958 6603
rect 25888 6537 25958 6549
rect 25028 6496 25774 6508
rect 25028 6440 25396 6496
rect 25452 6440 25774 6496
rect 25028 6428 25774 6440
rect 25028 6175 25084 6428
rect 25396 6175 25452 6428
rect 25718 6175 25774 6428
rect 25016 6173 25096 6175
rect 25016 6053 25028 6173
rect 25084 6053 25096 6173
rect 25016 6051 25096 6053
rect 25384 6173 25464 6175
rect 25384 6053 25396 6173
rect 25452 6053 25464 6173
rect 25384 6051 25464 6053
rect 25706 6173 25786 6175
rect 25706 6052 25718 6173
rect 25774 6052 25786 6173
rect 25028 6043 25084 6051
rect 25396 6043 25452 6051
rect 25706 6050 25786 6052
rect 25718 6042 25774 6050
rect 25212 5875 25268 5883
rect 25580 5875 25636 5883
rect 25200 5873 25689 5875
rect 25200 5753 25212 5873
rect 25268 5753 25580 5873
rect 25636 5753 25689 5873
rect 25200 5751 25689 5753
rect 25212 5743 25268 5751
rect 25580 5743 25689 5751
rect 25108 5677 25188 5687
rect 25108 5621 25120 5677
rect 25176 5621 25188 5677
rect 25108 5611 25188 5621
rect 25292 5677 25372 5687
rect 25292 5621 25304 5677
rect 25360 5621 25372 5677
rect 25292 5611 25372 5621
rect 25476 5677 25556 5687
rect 25476 5621 25488 5677
rect 25544 5621 25556 5677
rect 25476 5611 25556 5621
rect 25120 5529 25176 5611
rect 25108 5527 25188 5529
rect 25108 5471 25120 5527
rect 25176 5471 25188 5527
rect 25108 5469 25188 5471
rect 25120 5155 25176 5469
rect 25304 5413 25360 5611
rect 25292 5411 25372 5413
rect 25292 5355 25304 5411
rect 25360 5355 25372 5411
rect 25292 5353 25372 5355
rect 25304 5155 25360 5353
rect 25488 5297 25544 5611
rect 25621 5413 25689 5743
rect 26066 5421 26122 6655
rect 26514 6496 27260 6508
rect 26514 6440 26882 6496
rect 26938 6440 27260 6496
rect 26514 6428 27260 6440
rect 26514 6175 26570 6428
rect 26882 6175 26938 6428
rect 27204 6175 27260 6428
rect 26502 6173 26582 6175
rect 26502 6053 26514 6173
rect 26570 6053 26582 6173
rect 26502 6051 26582 6053
rect 26870 6173 26950 6175
rect 26870 6053 26882 6173
rect 26938 6053 26950 6173
rect 26870 6051 26950 6053
rect 27192 6173 27272 6175
rect 27192 6052 27204 6173
rect 27260 6052 27272 6173
rect 26514 6043 26570 6051
rect 26882 6043 26938 6051
rect 27192 6050 27272 6052
rect 27204 6042 27260 6050
rect 26698 5875 26754 5883
rect 27066 5875 27122 5883
rect 26686 5873 27175 5875
rect 26686 5753 26698 5873
rect 26754 5753 27066 5873
rect 27122 5753 27175 5873
rect 26686 5751 27175 5753
rect 26698 5743 26754 5751
rect 27066 5743 27175 5751
rect 26594 5677 26674 5687
rect 26594 5621 26606 5677
rect 26662 5621 26674 5677
rect 26594 5611 26674 5621
rect 26778 5677 26858 5687
rect 26778 5621 26790 5677
rect 26846 5621 26858 5677
rect 26778 5611 26858 5621
rect 26962 5677 27042 5687
rect 26962 5621 26974 5677
rect 27030 5621 27042 5677
rect 26962 5611 27042 5621
rect 26606 5529 26662 5611
rect 26594 5527 26674 5529
rect 26594 5471 26606 5527
rect 26662 5471 26674 5527
rect 26594 5469 26674 5471
rect 25621 5411 25701 5413
rect 25621 5355 25633 5411
rect 25689 5355 25701 5411
rect 25621 5353 25701 5355
rect 26064 5411 26124 5421
rect 26064 5355 26066 5411
rect 26122 5355 26124 5411
rect 25476 5295 25556 5297
rect 25476 5239 25488 5295
rect 25544 5239 25556 5295
rect 25476 5237 25556 5239
rect 25488 5155 25544 5237
rect 25108 5145 25188 5155
rect 25108 5089 25120 5145
rect 25176 5089 25188 5145
rect 25108 5079 25188 5089
rect 25292 5145 25372 5155
rect 25292 5089 25304 5145
rect 25360 5089 25372 5145
rect 25292 5079 25372 5089
rect 25476 5145 25556 5155
rect 25476 5089 25488 5145
rect 25544 5089 25556 5145
rect 25476 5079 25556 5089
rect 25621 5023 25689 5353
rect 26064 5343 26124 5355
rect 25580 5015 25689 5023
rect 25568 5013 25689 5015
rect 25568 4893 25580 5013
rect 25636 4893 25689 5013
rect 25568 4891 25689 4893
rect 25580 4883 25636 4891
rect 24883 4626 25779 4638
rect 24883 4570 24895 4626
rect 24951 4570 25713 4626
rect 25769 4570 25779 4626
rect 24883 4558 25779 4570
rect 26066 4400 26122 5343
rect 26606 5155 26662 5469
rect 26790 5413 26846 5611
rect 26778 5411 26858 5413
rect 26778 5355 26790 5411
rect 26846 5355 26858 5411
rect 26778 5353 26858 5355
rect 26790 5155 26846 5353
rect 26974 5297 27030 5611
rect 27107 5413 27175 5743
rect 27107 5411 27187 5413
rect 27107 5355 27119 5411
rect 27175 5355 27187 5411
rect 27107 5353 27187 5355
rect 27374 5411 27444 5423
rect 27374 5355 27376 5411
rect 27432 5355 27700 5411
rect 26962 5295 27042 5297
rect 26962 5239 26974 5295
rect 27030 5239 27042 5295
rect 26962 5237 27042 5239
rect 26974 5155 27030 5237
rect 26594 5145 26674 5155
rect 26594 5089 26606 5145
rect 26662 5089 26674 5145
rect 26594 5079 26674 5089
rect 26778 5145 26858 5155
rect 26778 5089 26790 5145
rect 26846 5089 26858 5145
rect 26778 5079 26858 5089
rect 26962 5145 27042 5155
rect 26962 5089 26974 5145
rect 27030 5089 27042 5145
rect 26962 5079 27042 5089
rect 27107 5023 27175 5353
rect 27374 5345 27444 5355
rect 27066 5015 27175 5023
rect 27054 5013 27175 5015
rect 27054 4893 27066 5013
rect 27122 4893 27175 5013
rect 27054 4891 27175 4893
rect 27066 4883 27122 4891
rect 26369 4626 27265 4638
rect 26369 4570 26381 4626
rect 26437 4570 27199 4626
rect 27255 4570 27265 4626
rect 26369 4558 27265 4570
rect 27376 4401 27432 5345
rect 27540 4509 27620 4519
rect 27540 4453 27552 4509
rect 27608 4453 27620 4509
rect 27540 4451 27620 4453
rect 26064 4398 26134 4400
rect 26064 4342 26066 4398
rect 26122 4342 26134 4398
rect 26064 4330 26134 4342
rect 27364 4399 27444 4401
rect 27364 4343 27376 4399
rect 27432 4343 27444 4399
rect 27364 4331 27444 4343
rect 25028 4291 25774 4303
rect 25028 4235 25396 4291
rect 25452 4235 25774 4291
rect 25028 4223 25774 4235
rect 25028 3970 25084 4223
rect 25396 3970 25452 4223
rect 25718 3970 25774 4223
rect 26514 4292 27260 4304
rect 26514 4236 26882 4292
rect 26938 4236 27260 4292
rect 26514 4224 27260 4236
rect 26514 3971 26570 4224
rect 26882 3971 26938 4224
rect 27204 3971 27260 4224
rect 25016 3968 25096 3970
rect 25016 3848 25028 3968
rect 25084 3848 25096 3968
rect 25016 3846 25096 3848
rect 25384 3968 25464 3970
rect 25384 3848 25396 3968
rect 25452 3848 25464 3968
rect 25384 3846 25464 3848
rect 25706 3968 25786 3970
rect 25706 3847 25718 3968
rect 25774 3847 25786 3968
rect 26502 3969 26582 3971
rect 26502 3849 26514 3969
rect 26570 3849 26582 3969
rect 26502 3847 26582 3849
rect 26870 3969 26950 3971
rect 26870 3849 26882 3969
rect 26938 3849 26950 3969
rect 26870 3847 26950 3849
rect 27192 3969 27272 3971
rect 27192 3848 27204 3969
rect 27260 3848 27272 3969
rect 25028 3838 25084 3846
rect 25396 3838 25452 3846
rect 25706 3845 25786 3847
rect 25718 3837 25774 3845
rect 26514 3839 26570 3847
rect 26882 3839 26938 3847
rect 27192 3846 27272 3848
rect 27204 3838 27260 3846
rect 25212 3670 25268 3678
rect 25580 3670 25636 3678
rect 26698 3671 26754 3679
rect 27066 3671 27122 3679
rect 25200 3668 25689 3670
rect 25200 3548 25212 3668
rect 25268 3548 25580 3668
rect 25636 3548 25689 3668
rect 25200 3546 25689 3548
rect 26686 3669 27175 3671
rect 26686 3549 26698 3669
rect 26754 3549 27066 3669
rect 27122 3549 27175 3669
rect 26686 3547 27175 3549
rect 25212 3538 25268 3546
rect 25580 3538 25689 3546
rect 26698 3539 26754 3547
rect 27066 3539 27175 3547
rect 25108 3472 25188 3482
rect 25108 3416 25120 3472
rect 25176 3416 25188 3472
rect 25108 3406 25188 3416
rect 25292 3472 25372 3482
rect 25292 3416 25304 3472
rect 25360 3416 25372 3472
rect 25292 3406 25372 3416
rect 25476 3472 25556 3482
rect 25476 3416 25488 3472
rect 25544 3416 25556 3472
rect 25476 3406 25556 3416
rect 25120 3324 25176 3406
rect 25108 3322 25188 3324
rect 25108 3266 25120 3322
rect 25176 3266 25188 3322
rect 25108 3264 25188 3266
rect 24436 3090 24506 3102
rect 24436 3034 24448 3090
rect 24504 3034 24506 3090
rect 24436 3022 24506 3034
rect 25120 2950 25176 3264
rect 25304 3208 25360 3406
rect 25292 3206 25372 3208
rect 25292 3150 25304 3206
rect 25360 3150 25372 3206
rect 25292 3148 25372 3150
rect 25304 2950 25360 3148
rect 25488 3092 25544 3406
rect 25621 3208 25689 3538
rect 26594 3473 26674 3483
rect 26594 3417 26606 3473
rect 26662 3417 26674 3473
rect 26594 3407 26674 3417
rect 26778 3473 26858 3483
rect 26778 3417 26790 3473
rect 26846 3417 26858 3473
rect 26778 3407 26858 3417
rect 26962 3473 27042 3483
rect 26962 3417 26974 3473
rect 27030 3417 27042 3473
rect 26962 3407 27042 3417
rect 26606 3325 26662 3407
rect 26594 3323 26674 3325
rect 26594 3267 26606 3323
rect 26662 3267 26674 3323
rect 26594 3265 26674 3267
rect 25621 3206 25701 3208
rect 25621 3150 25633 3206
rect 25689 3150 25701 3206
rect 25621 3148 25701 3150
rect 25888 3206 25958 3218
rect 25888 3150 25890 3206
rect 25946 3150 25958 3206
rect 25476 3090 25556 3092
rect 25476 3034 25488 3090
rect 25544 3034 25556 3090
rect 25476 3032 25556 3034
rect 25488 2950 25544 3032
rect 25108 2940 25188 2950
rect 25108 2884 25120 2940
rect 25176 2884 25188 2940
rect 25108 2874 25188 2884
rect 25292 2940 25372 2950
rect 25292 2884 25304 2940
rect 25360 2884 25372 2940
rect 25292 2874 25372 2884
rect 25476 2940 25556 2950
rect 25476 2884 25488 2940
rect 25544 2884 25556 2940
rect 25476 2874 25556 2884
rect 25621 2818 25689 3148
rect 25888 3140 25958 3150
rect 25580 2810 25689 2818
rect 25568 2808 25689 2810
rect 25568 2688 25580 2808
rect 25636 2688 25689 2808
rect 25568 2686 25689 2688
rect 25580 2678 25636 2686
rect 24883 2421 25779 2433
rect 24883 2365 24895 2421
rect 24951 2365 25713 2421
rect 25769 2365 25779 2421
rect 24883 2353 25779 2365
rect 25890 2196 25946 3140
rect 26606 2951 26662 3265
rect 26790 3209 26846 3407
rect 26778 3207 26858 3209
rect 26778 3151 26790 3207
rect 26846 3151 26858 3207
rect 26778 3149 26858 3151
rect 26790 2951 26846 3149
rect 26974 3093 27030 3407
rect 27107 3209 27175 3539
rect 27552 3217 27608 4451
rect 27107 3207 27187 3209
rect 27107 3151 27119 3207
rect 27175 3151 27187 3207
rect 27107 3149 27187 3151
rect 27550 3207 27620 3217
rect 27780 3207 27836 17250
rect 27982 14999 28038 18679
rect 32022 18561 32092 18573
rect 32022 18505 32024 18561
rect 32080 18505 32092 18561
rect 32022 18503 32092 18505
rect 29070 18277 29816 18289
rect 29070 18221 29438 18277
rect 29494 18221 29816 18277
rect 29070 18209 29816 18221
rect 29070 17956 29126 18209
rect 29438 17956 29494 18209
rect 29760 17956 29816 18209
rect 29058 17954 29138 17956
rect 29058 17834 29070 17954
rect 29126 17834 29138 17954
rect 29058 17832 29138 17834
rect 29426 17954 29506 17956
rect 29426 17834 29438 17954
rect 29494 17834 29506 17954
rect 29426 17832 29506 17834
rect 29748 17954 29828 17956
rect 29748 17833 29760 17954
rect 29816 17833 29828 17954
rect 29070 17824 29126 17832
rect 29438 17824 29494 17832
rect 29748 17831 29828 17833
rect 29760 17823 29816 17831
rect 29254 17656 29310 17664
rect 29622 17656 29678 17664
rect 29242 17654 29731 17656
rect 29242 17534 29254 17654
rect 29310 17534 29622 17654
rect 29678 17534 29731 17654
rect 29242 17532 29731 17534
rect 29254 17524 29310 17532
rect 29622 17524 29731 17532
rect 29150 17458 29230 17468
rect 29150 17402 29162 17458
rect 29218 17402 29230 17458
rect 29150 17392 29230 17402
rect 29334 17458 29414 17468
rect 29334 17402 29346 17458
rect 29402 17402 29414 17458
rect 29334 17392 29414 17402
rect 29518 17458 29598 17468
rect 29518 17402 29530 17458
rect 29586 17402 29598 17458
rect 29518 17392 29598 17402
rect 29162 17310 29218 17392
rect 29150 17308 29230 17310
rect 29150 17252 29162 17308
rect 29218 17252 29230 17308
rect 29150 17250 29230 17252
rect 28478 17192 28548 17204
rect 28478 17136 28490 17192
rect 28546 17136 28548 17192
rect 28478 17124 28548 17136
rect 27980 14987 28050 14999
rect 27980 14931 27982 14987
rect 28038 14931 28050 14987
rect 27980 14919 28050 14931
rect 28342 14987 28412 15001
rect 28342 14931 28354 14987
rect 28410 14931 28412 14987
rect 28342 14919 28412 14931
rect 28162 14085 28240 14097
rect 28162 14029 28173 14085
rect 28229 14029 28240 14085
rect 28162 14017 28240 14029
rect 28354 10591 28410 14919
rect 28490 12678 28546 17124
rect 29162 16936 29218 17250
rect 29346 17194 29402 17392
rect 29334 17192 29414 17194
rect 29334 17136 29346 17192
rect 29402 17136 29414 17192
rect 29334 17134 29414 17136
rect 29346 16936 29402 17134
rect 29530 17078 29586 17392
rect 29663 17194 29731 17524
rect 29663 17192 29743 17194
rect 29663 17136 29675 17192
rect 29731 17136 29743 17192
rect 29663 17134 29743 17136
rect 29930 17192 30000 17204
rect 29930 17136 29932 17192
rect 29988 17136 30000 17192
rect 29518 17076 29598 17078
rect 29518 17020 29530 17076
rect 29586 17020 29598 17076
rect 29518 17018 29598 17020
rect 29530 16936 29586 17018
rect 29150 16926 29230 16936
rect 29150 16870 29162 16926
rect 29218 16870 29230 16926
rect 29150 16860 29230 16870
rect 29334 16926 29414 16936
rect 29334 16870 29346 16926
rect 29402 16870 29414 16926
rect 29334 16860 29414 16870
rect 29518 16926 29598 16936
rect 29518 16870 29530 16926
rect 29586 16870 29598 16926
rect 29518 16860 29598 16870
rect 29663 16804 29731 17134
rect 29930 17126 30000 17136
rect 29622 16796 29731 16804
rect 29610 16794 29731 16796
rect 29610 16674 29622 16794
rect 29678 16674 29731 16794
rect 29610 16672 29731 16674
rect 29622 16664 29678 16672
rect 28925 16407 29823 16419
rect 28925 16351 28937 16407
rect 28993 16351 29755 16407
rect 29811 16351 29823 16407
rect 28925 16339 29823 16351
rect 29932 16182 29988 17126
rect 30096 16289 30176 16299
rect 30096 16233 30108 16289
rect 30164 16233 30176 16289
rect 30096 16231 30176 16233
rect 29930 16179 30000 16182
rect 29930 16125 29932 16179
rect 29988 16125 30000 16179
rect 29930 16113 30000 16125
rect 29070 16072 29816 16084
rect 29070 16016 29438 16072
rect 29494 16016 29816 16072
rect 29070 16004 29816 16016
rect 29070 15751 29126 16004
rect 29438 15751 29494 16004
rect 29760 15751 29816 16004
rect 29058 15749 29138 15751
rect 29058 15629 29070 15749
rect 29126 15629 29138 15749
rect 29058 15627 29138 15629
rect 29426 15749 29506 15751
rect 29426 15629 29438 15749
rect 29494 15629 29506 15749
rect 29426 15627 29506 15629
rect 29748 15749 29828 15751
rect 29748 15628 29760 15749
rect 29816 15628 29828 15749
rect 29070 15619 29126 15627
rect 29438 15619 29494 15627
rect 29748 15626 29828 15628
rect 29760 15618 29816 15626
rect 29254 15451 29310 15459
rect 29622 15451 29678 15459
rect 29242 15449 29731 15451
rect 29242 15329 29254 15449
rect 29310 15329 29622 15449
rect 29678 15329 29731 15449
rect 29242 15327 29731 15329
rect 29254 15319 29310 15327
rect 29622 15319 29731 15327
rect 29150 15253 29230 15263
rect 29150 15197 29162 15253
rect 29218 15197 29230 15253
rect 29150 15187 29230 15197
rect 29334 15253 29414 15263
rect 29334 15197 29346 15253
rect 29402 15197 29414 15253
rect 29334 15187 29414 15197
rect 29518 15253 29598 15263
rect 29518 15197 29530 15253
rect 29586 15197 29598 15253
rect 29518 15187 29598 15197
rect 29162 15105 29218 15187
rect 29150 15103 29230 15105
rect 29150 15047 29162 15103
rect 29218 15047 29230 15103
rect 29150 15045 29230 15047
rect 29162 14731 29218 15045
rect 29346 14989 29402 15187
rect 29334 14987 29414 14989
rect 29334 14931 29346 14987
rect 29402 14931 29414 14987
rect 29334 14929 29414 14931
rect 29346 14731 29402 14929
rect 29530 14873 29586 15187
rect 29663 14989 29731 15319
rect 30108 14997 30164 16231
rect 30556 16072 31302 16084
rect 30556 16016 30924 16072
rect 30980 16016 31302 16072
rect 30556 16004 31302 16016
rect 30556 15751 30612 16004
rect 30924 15751 30980 16004
rect 31246 15751 31302 16004
rect 30544 15749 30624 15751
rect 30544 15629 30556 15749
rect 30612 15629 30624 15749
rect 30544 15627 30624 15629
rect 30912 15749 30992 15751
rect 30912 15629 30924 15749
rect 30980 15629 30992 15749
rect 30912 15627 30992 15629
rect 31234 15749 31314 15751
rect 31234 15628 31246 15749
rect 31302 15628 31314 15749
rect 30556 15619 30612 15627
rect 30924 15619 30980 15627
rect 31234 15626 31314 15628
rect 31246 15618 31302 15626
rect 30740 15451 30796 15459
rect 31108 15451 31164 15459
rect 30728 15449 31217 15451
rect 30728 15329 30740 15449
rect 30796 15329 31108 15449
rect 31164 15329 31217 15449
rect 30728 15327 31217 15329
rect 30740 15319 30796 15327
rect 31108 15319 31217 15327
rect 30636 15253 30716 15263
rect 30636 15197 30648 15253
rect 30704 15197 30716 15253
rect 30636 15187 30716 15197
rect 30820 15253 30900 15263
rect 30820 15197 30832 15253
rect 30888 15197 30900 15253
rect 30820 15187 30900 15197
rect 31004 15253 31084 15263
rect 31004 15197 31016 15253
rect 31072 15197 31084 15253
rect 31004 15187 31084 15197
rect 30648 15105 30704 15187
rect 30636 15103 30716 15105
rect 30636 15047 30648 15103
rect 30704 15047 30716 15103
rect 30636 15045 30716 15047
rect 29663 14987 29743 14989
rect 29663 14931 29675 14987
rect 29731 14931 29743 14987
rect 29663 14929 29743 14931
rect 30106 14987 30166 14997
rect 30106 14931 30108 14987
rect 30164 14931 30166 14987
rect 29518 14871 29598 14873
rect 29518 14815 29530 14871
rect 29586 14815 29598 14871
rect 29518 14813 29598 14815
rect 29530 14731 29586 14813
rect 29150 14721 29230 14731
rect 29150 14665 29162 14721
rect 29218 14665 29230 14721
rect 29150 14655 29230 14665
rect 29334 14721 29414 14731
rect 29334 14665 29346 14721
rect 29402 14665 29414 14721
rect 29334 14655 29414 14665
rect 29518 14721 29598 14731
rect 29518 14665 29530 14721
rect 29586 14665 29598 14721
rect 29518 14655 29598 14665
rect 29663 14599 29731 14929
rect 30106 14919 30166 14931
rect 29622 14591 29731 14599
rect 29610 14589 29731 14591
rect 29610 14469 29622 14589
rect 29678 14469 29731 14589
rect 29610 14467 29731 14469
rect 29622 14459 29678 14467
rect 28925 14202 29821 14214
rect 28925 14146 28937 14202
rect 28993 14146 29755 14202
rect 29811 14146 29821 14202
rect 28925 14134 29821 14146
rect 30108 13976 30164 14919
rect 30648 14731 30704 15045
rect 30832 14989 30888 15187
rect 30820 14987 30900 14989
rect 30820 14931 30832 14987
rect 30888 14931 30900 14987
rect 30820 14929 30900 14931
rect 30832 14731 30888 14929
rect 31016 14873 31072 15187
rect 31149 14989 31217 15319
rect 32024 14999 32080 18503
rect 31149 14987 31229 14989
rect 31149 14931 31161 14987
rect 31217 14931 31229 14987
rect 31149 14929 31229 14931
rect 31416 14987 31486 14999
rect 32022 14987 32092 14999
rect 31416 14931 31418 14987
rect 31474 14931 31742 14987
rect 32022 14931 32024 14987
rect 32080 14931 32092 14987
rect 31004 14871 31084 14873
rect 31004 14815 31016 14871
rect 31072 14815 31084 14871
rect 31004 14813 31084 14815
rect 31016 14731 31072 14813
rect 30636 14721 30716 14731
rect 30636 14665 30648 14721
rect 30704 14665 30716 14721
rect 30636 14655 30716 14665
rect 30820 14721 30900 14731
rect 30820 14665 30832 14721
rect 30888 14665 30900 14721
rect 30820 14655 30900 14665
rect 31004 14721 31084 14731
rect 31004 14665 31016 14721
rect 31072 14665 31084 14721
rect 31004 14655 31084 14665
rect 31149 14599 31217 14929
rect 31416 14921 31486 14931
rect 31108 14591 31217 14599
rect 31096 14589 31217 14591
rect 31096 14469 31108 14589
rect 31164 14469 31217 14589
rect 31096 14467 31217 14469
rect 31108 14459 31164 14467
rect 30411 14202 31307 14214
rect 30411 14146 30423 14202
rect 30479 14146 31241 14202
rect 31297 14146 31307 14202
rect 30411 14134 31307 14146
rect 31418 13977 31474 14921
rect 32022 14919 32092 14931
rect 31582 14085 31662 14095
rect 31582 14029 31594 14085
rect 31650 14029 31662 14085
rect 31582 14027 31662 14029
rect 30106 13974 30176 13976
rect 30106 13918 30108 13974
rect 30164 13918 30176 13974
rect 30106 13906 30176 13918
rect 31406 13975 31486 13977
rect 31406 13919 31418 13975
rect 31474 13919 31486 13975
rect 31406 13907 31486 13919
rect 29070 13867 29816 13879
rect 29070 13811 29438 13867
rect 29494 13811 29816 13867
rect 29070 13799 29816 13811
rect 29070 13546 29126 13799
rect 29438 13546 29494 13799
rect 29760 13546 29816 13799
rect 30556 13868 31302 13880
rect 30556 13812 30924 13868
rect 30980 13812 31302 13868
rect 30556 13800 31302 13812
rect 30556 13547 30612 13800
rect 30924 13547 30980 13800
rect 31246 13547 31302 13800
rect 29058 13544 29138 13546
rect 29058 13424 29070 13544
rect 29126 13424 29138 13544
rect 29058 13422 29138 13424
rect 29426 13544 29506 13546
rect 29426 13424 29438 13544
rect 29494 13424 29506 13544
rect 29426 13422 29506 13424
rect 29748 13544 29828 13546
rect 29748 13423 29760 13544
rect 29816 13423 29828 13544
rect 30544 13545 30624 13547
rect 30544 13425 30556 13545
rect 30612 13425 30624 13545
rect 30544 13423 30624 13425
rect 30912 13545 30992 13547
rect 30912 13425 30924 13545
rect 30980 13425 30992 13545
rect 30912 13423 30992 13425
rect 31234 13545 31314 13547
rect 31234 13424 31246 13545
rect 31302 13424 31314 13545
rect 29070 13414 29126 13422
rect 29438 13414 29494 13422
rect 29748 13421 29828 13423
rect 29760 13413 29816 13421
rect 30556 13415 30612 13423
rect 30924 13415 30980 13423
rect 31234 13422 31314 13424
rect 31246 13414 31302 13422
rect 29254 13246 29310 13254
rect 29622 13246 29678 13254
rect 30740 13247 30796 13255
rect 31108 13247 31164 13255
rect 29242 13244 29731 13246
rect 29242 13124 29254 13244
rect 29310 13124 29622 13244
rect 29678 13124 29731 13244
rect 29242 13122 29731 13124
rect 30728 13245 31217 13247
rect 30728 13125 30740 13245
rect 30796 13125 31108 13245
rect 31164 13125 31217 13245
rect 30728 13123 31217 13125
rect 29254 13114 29310 13122
rect 29622 13114 29731 13122
rect 30740 13115 30796 13123
rect 31108 13115 31217 13123
rect 29150 13048 29230 13058
rect 29150 12992 29162 13048
rect 29218 12992 29230 13048
rect 29150 12982 29230 12992
rect 29334 13048 29414 13058
rect 29334 12992 29346 13048
rect 29402 12992 29414 13048
rect 29334 12982 29414 12992
rect 29518 13048 29598 13058
rect 29518 12992 29530 13048
rect 29586 12992 29598 13048
rect 29518 12982 29598 12992
rect 29162 12900 29218 12982
rect 29150 12898 29230 12900
rect 29150 12842 29162 12898
rect 29218 12842 29230 12898
rect 29150 12840 29230 12842
rect 28478 12666 28548 12678
rect 28478 12610 28490 12666
rect 28546 12610 28548 12666
rect 28478 12598 28548 12610
rect 29162 12526 29218 12840
rect 29346 12784 29402 12982
rect 29334 12782 29414 12784
rect 29334 12726 29346 12782
rect 29402 12726 29414 12782
rect 29334 12724 29414 12726
rect 29346 12526 29402 12724
rect 29530 12668 29586 12982
rect 29663 12784 29731 13114
rect 30636 13049 30716 13059
rect 30636 12993 30648 13049
rect 30704 12993 30716 13049
rect 30636 12983 30716 12993
rect 30820 13049 30900 13059
rect 30820 12993 30832 13049
rect 30888 12993 30900 13049
rect 30820 12983 30900 12993
rect 31004 13049 31084 13059
rect 31004 12993 31016 13049
rect 31072 12993 31084 13049
rect 31004 12983 31084 12993
rect 30648 12901 30704 12983
rect 30636 12899 30716 12901
rect 30636 12843 30648 12899
rect 30704 12843 30716 12899
rect 30636 12841 30716 12843
rect 29663 12782 29743 12784
rect 29663 12726 29675 12782
rect 29731 12726 29743 12782
rect 29663 12724 29743 12726
rect 29930 12782 30000 12794
rect 29930 12726 29932 12782
rect 29988 12726 30000 12782
rect 29518 12666 29598 12668
rect 29518 12610 29530 12666
rect 29586 12610 29598 12666
rect 29518 12608 29598 12610
rect 29530 12526 29586 12608
rect 29150 12516 29230 12526
rect 29150 12460 29162 12516
rect 29218 12460 29230 12516
rect 29150 12450 29230 12460
rect 29334 12516 29414 12526
rect 29334 12460 29346 12516
rect 29402 12460 29414 12516
rect 29334 12450 29414 12460
rect 29518 12516 29598 12526
rect 29518 12460 29530 12516
rect 29586 12460 29598 12516
rect 29518 12450 29598 12460
rect 29663 12394 29731 12724
rect 29930 12716 30000 12726
rect 29622 12386 29731 12394
rect 29610 12384 29731 12386
rect 29610 12264 29622 12384
rect 29678 12264 29731 12384
rect 29610 12262 29731 12264
rect 29622 12254 29678 12262
rect 28925 11997 29821 12009
rect 28925 11941 28937 11997
rect 28993 11941 29755 11997
rect 29811 11941 29821 11997
rect 28925 11929 29821 11941
rect 29932 11772 29988 12716
rect 30648 12527 30704 12841
rect 30832 12785 30888 12983
rect 30820 12783 30900 12785
rect 30820 12727 30832 12783
rect 30888 12727 30900 12783
rect 30820 12725 30900 12727
rect 30832 12527 30888 12725
rect 31016 12669 31072 12983
rect 31149 12785 31217 13115
rect 31594 12793 31650 14027
rect 31149 12783 31229 12785
rect 31149 12727 31161 12783
rect 31217 12727 31229 12783
rect 31149 12725 31229 12727
rect 31592 12783 31662 12793
rect 31592 12727 31594 12783
rect 31650 12727 31742 12783
rect 31004 12667 31084 12669
rect 31004 12611 31016 12667
rect 31072 12611 31084 12667
rect 31004 12609 31084 12611
rect 31016 12527 31072 12609
rect 30636 12517 30716 12527
rect 30636 12461 30648 12517
rect 30704 12461 30716 12517
rect 30636 12451 30716 12461
rect 30820 12517 30900 12527
rect 30820 12461 30832 12517
rect 30888 12461 30900 12517
rect 30820 12451 30900 12461
rect 31004 12517 31084 12527
rect 31004 12461 31016 12517
rect 31072 12461 31084 12517
rect 31004 12451 31084 12461
rect 31149 12395 31217 12725
rect 31592 12715 31662 12727
rect 31108 12387 31217 12395
rect 31096 12385 31217 12387
rect 31096 12265 31108 12385
rect 31164 12265 31217 12385
rect 31096 12263 31217 12265
rect 31108 12255 31164 12263
rect 30411 11998 31307 12010
rect 30411 11942 30423 11998
rect 30479 11942 31241 11998
rect 31297 11942 31307 11998
rect 30411 11930 31307 11942
rect 30096 11879 30176 11889
rect 30096 11823 30108 11879
rect 30164 11823 30176 11879
rect 30096 11821 30176 11823
rect 29930 11769 30000 11772
rect 29930 11715 29932 11769
rect 29988 11715 30000 11769
rect 29930 11703 30000 11715
rect 29070 11662 29816 11674
rect 29070 11606 29438 11662
rect 29494 11606 29816 11662
rect 29070 11594 29816 11606
rect 29070 11341 29126 11594
rect 29438 11341 29494 11594
rect 29760 11341 29816 11594
rect 29058 11339 29138 11341
rect 29058 11219 29070 11339
rect 29126 11219 29138 11339
rect 29058 11217 29138 11219
rect 29426 11339 29506 11341
rect 29426 11219 29438 11339
rect 29494 11219 29506 11339
rect 29426 11217 29506 11219
rect 29748 11339 29828 11341
rect 29748 11218 29760 11339
rect 29816 11218 29828 11339
rect 29070 11209 29126 11217
rect 29438 11209 29494 11217
rect 29748 11216 29828 11218
rect 29760 11208 29816 11216
rect 29254 11041 29310 11049
rect 29622 11041 29678 11049
rect 29242 11039 29731 11041
rect 29242 10919 29254 11039
rect 29310 10919 29622 11039
rect 29678 10919 29731 11039
rect 29242 10917 29731 10919
rect 29254 10909 29310 10917
rect 29622 10909 29731 10917
rect 29150 10843 29230 10853
rect 29150 10787 29162 10843
rect 29218 10787 29230 10843
rect 29150 10777 29230 10787
rect 29334 10843 29414 10853
rect 29334 10787 29346 10843
rect 29402 10787 29414 10843
rect 29334 10777 29414 10787
rect 29518 10843 29598 10853
rect 29518 10787 29530 10843
rect 29586 10787 29598 10843
rect 29518 10777 29598 10787
rect 29162 10695 29218 10777
rect 29150 10693 29230 10695
rect 29150 10637 29162 10693
rect 29218 10637 29230 10693
rect 29150 10635 29230 10637
rect 28342 10577 28412 10591
rect 28342 10521 28354 10577
rect 28410 10521 28412 10577
rect 28342 10509 28412 10521
rect 28162 10461 28240 10473
rect 28162 10405 28173 10461
rect 28229 10405 28240 10461
rect 28162 10393 28240 10405
rect 28040 9674 28110 9686
rect 28354 9678 28410 10509
rect 29162 10321 29218 10635
rect 29346 10579 29402 10777
rect 29334 10577 29414 10579
rect 29334 10521 29346 10577
rect 29402 10521 29414 10577
rect 29334 10519 29414 10521
rect 29346 10321 29402 10519
rect 29530 10463 29586 10777
rect 29663 10579 29731 10909
rect 30108 10589 30164 11821
rect 29663 10577 29743 10579
rect 29663 10521 29675 10577
rect 29731 10521 29743 10577
rect 29663 10519 29743 10521
rect 30106 10577 30166 10589
rect 30106 10521 30108 10577
rect 30164 10521 30166 10577
rect 29518 10461 29598 10463
rect 29518 10405 29530 10461
rect 29586 10405 29598 10461
rect 29518 10403 29598 10405
rect 29530 10321 29586 10403
rect 29150 10311 29230 10321
rect 29150 10255 29162 10311
rect 29218 10255 29230 10311
rect 29150 10245 29230 10255
rect 29334 10311 29414 10321
rect 29334 10255 29346 10311
rect 29402 10255 29414 10311
rect 29334 10245 29414 10255
rect 29518 10311 29598 10321
rect 29518 10255 29530 10311
rect 29586 10255 29598 10311
rect 29518 10245 29598 10255
rect 29663 10189 29731 10519
rect 30106 10509 30166 10521
rect 29622 10181 29731 10189
rect 29610 10179 29731 10181
rect 29610 10059 29622 10179
rect 29678 10059 29731 10179
rect 29610 10057 29731 10059
rect 29622 10049 29678 10057
rect 28925 9792 29823 9804
rect 28925 9736 28937 9792
rect 28993 9736 29755 9792
rect 29811 9736 29823 9792
rect 28925 9724 29823 9736
rect 28040 9618 28052 9674
rect 28108 9618 28110 9674
rect 28040 9606 28110 9618
rect 28352 9674 28412 9678
rect 28352 9618 28354 9674
rect 28410 9618 28412 9674
rect 28352 9606 28412 9618
rect 28052 9004 28108 9606
rect 28052 8894 28108 8904
rect 27550 3151 27552 3207
rect 27608 3151 27836 3207
rect 26962 3091 27042 3093
rect 26962 3035 26974 3091
rect 27030 3035 27042 3091
rect 26962 3033 27042 3035
rect 26974 2951 27030 3033
rect 26594 2941 26674 2951
rect 26594 2885 26606 2941
rect 26662 2885 26674 2941
rect 26594 2875 26674 2885
rect 26778 2941 26858 2951
rect 26778 2885 26790 2941
rect 26846 2885 26858 2941
rect 26778 2875 26858 2885
rect 26962 2941 27042 2951
rect 26962 2885 26974 2941
rect 27030 2885 27042 2941
rect 26962 2875 27042 2885
rect 27107 2819 27175 3149
rect 27550 3139 27620 3151
rect 27066 2811 27175 2819
rect 27054 2809 27175 2811
rect 27054 2689 27066 2809
rect 27122 2689 27175 2809
rect 27054 2687 27175 2689
rect 27066 2679 27122 2687
rect 26369 2422 27265 2434
rect 26369 2366 26381 2422
rect 26437 2366 27199 2422
rect 27255 2366 27265 2422
rect 26369 2354 27265 2366
rect 26054 2303 26134 2313
rect 26054 2247 26066 2303
rect 26122 2247 26134 2303
rect 26054 2245 26134 2247
rect 25888 2193 25958 2196
rect 25888 2139 25890 2193
rect 25946 2139 25958 2193
rect 25888 2127 25958 2139
rect 25028 2086 25774 2098
rect 25028 2030 25396 2086
rect 25452 2030 25774 2086
rect 25028 2018 25774 2030
rect 25028 1765 25084 2018
rect 25396 1765 25452 2018
rect 25718 1765 25774 2018
rect 25016 1763 25096 1765
rect 25016 1643 25028 1763
rect 25084 1643 25096 1763
rect 25016 1641 25096 1643
rect 25384 1763 25464 1765
rect 25384 1643 25396 1763
rect 25452 1643 25464 1763
rect 25384 1641 25464 1643
rect 25706 1763 25786 1765
rect 25706 1642 25718 1763
rect 25774 1642 25786 1763
rect 25028 1633 25084 1641
rect 25396 1633 25452 1641
rect 25706 1640 25786 1642
rect 25718 1632 25774 1640
rect 25212 1465 25268 1473
rect 25580 1465 25636 1473
rect 25200 1463 25689 1465
rect 25200 1343 25212 1463
rect 25268 1343 25580 1463
rect 25636 1343 25689 1463
rect 25200 1341 25689 1343
rect 25212 1333 25268 1341
rect 25580 1333 25689 1341
rect 25108 1267 25188 1277
rect 25108 1211 25120 1267
rect 25176 1211 25188 1267
rect 25108 1201 25188 1211
rect 25292 1267 25372 1277
rect 25292 1211 25304 1267
rect 25360 1211 25372 1267
rect 25292 1201 25372 1211
rect 25476 1267 25556 1277
rect 25476 1211 25488 1267
rect 25544 1211 25556 1267
rect 25476 1201 25556 1211
rect 25120 1119 25176 1201
rect 25108 1117 25188 1119
rect 25108 1061 25120 1117
rect 25176 1061 25188 1117
rect 25108 1059 25188 1061
rect 24300 1001 24370 1015
rect 24300 945 24312 1001
rect 24368 945 24370 1001
rect 24300 933 24370 945
rect 24134 885 24214 897
rect 24134 829 24146 885
rect 24202 829 24214 885
rect 24134 817 24214 829
rect 23998 98 24068 110
rect 24312 102 24368 933
rect 25120 745 25176 1059
rect 25304 1003 25360 1201
rect 25292 1001 25372 1003
rect 25292 945 25304 1001
rect 25360 945 25372 1001
rect 25292 943 25372 945
rect 25304 745 25360 943
rect 25488 887 25544 1201
rect 25621 1003 25689 1333
rect 26066 1013 26122 2245
rect 25621 1001 25701 1003
rect 25621 945 25633 1001
rect 25689 945 25701 1001
rect 25621 943 25701 945
rect 26064 1001 26124 1013
rect 26064 945 26066 1001
rect 26122 945 26124 1001
rect 25476 885 25556 887
rect 25476 829 25488 885
rect 25544 829 25556 885
rect 25476 827 25556 829
rect 25488 745 25544 827
rect 25108 735 25188 745
rect 25108 679 25120 735
rect 25176 679 25188 735
rect 25108 669 25188 679
rect 25292 735 25372 745
rect 25292 679 25304 735
rect 25360 679 25372 735
rect 25292 669 25372 679
rect 25476 735 25556 745
rect 25476 679 25488 735
rect 25544 679 25556 735
rect 25476 669 25556 679
rect 25621 613 25689 943
rect 26064 933 26124 945
rect 25580 605 25689 613
rect 25568 603 25689 605
rect 25568 483 25580 603
rect 25636 483 25689 603
rect 25568 481 25689 483
rect 25580 473 25636 481
rect 24883 216 25781 228
rect 24883 160 24895 216
rect 24951 160 25713 216
rect 25769 160 25781 216
rect 24883 148 25781 160
rect 23998 42 24010 98
rect 24066 42 24068 98
rect 23998 30 24068 42
rect 24310 98 24370 102
rect 24310 42 24312 98
rect 24368 42 24370 98
rect 24310 30 24370 42
rect 23874 -175 23930 -165
<< via2 >>
rect -46 9414 10 9514
rect 3286 9414 3342 9514
rect -46 8904 10 9004
rect 1174 8645 1230 8701
rect 673 6775 729 6831
rect 1491 6775 1547 6831
rect 1174 6440 1230 6496
rect 2660 6440 2716 6496
rect 673 4570 729 4626
rect 1491 4570 1547 4626
rect 2159 4570 2215 4626
rect 2977 4570 3033 4626
rect 1174 4235 1230 4291
rect 2660 4236 2716 4292
rect 673 2365 729 2421
rect 1491 2365 1547 2421
rect 5186 18224 5242 18280
rect 4685 16354 4741 16410
rect 5503 16354 5559 16410
rect 5186 16019 5242 16075
rect 6672 16019 6728 16075
rect 4685 14149 4741 14205
rect 5503 14149 5559 14205
rect 6171 14149 6227 14205
rect 6989 14149 7045 14205
rect 5186 13814 5242 13870
rect 6672 13815 6728 13871
rect 4685 11944 4741 12000
rect 5503 11944 5559 12000
rect 6171 11945 6227 12001
rect 6989 11945 7045 12001
rect 5186 11609 5242 11665
rect 4685 9739 4741 9795
rect 5503 9739 5559 9795
rect 7298 9414 7354 9514
rect 3830 8907 3886 9007
rect 2159 2366 2215 2422
rect 2977 2366 3033 2422
rect 1174 2030 1230 2086
rect -109 829 -53 885
rect 673 160 729 216
rect 1491 160 1547 216
rect -109 42 -53 98
rect -318 -165 -262 -65
rect 5186 8645 5242 8701
rect 4022 7676 4078 7732
rect 4685 6775 4741 6831
rect 5503 6775 5559 6831
rect 5186 6440 5242 6496
rect 6672 6440 6728 6496
rect 4685 4570 4741 4626
rect 5503 4570 5559 4626
rect 6171 4570 6227 4626
rect 6989 4570 7045 4626
rect 5186 4235 5242 4291
rect 6672 4236 6728 4292
rect 4685 2365 4741 2421
rect 5503 2365 5559 2421
rect 9228 18221 9284 18277
rect 8727 16351 8783 16407
rect 9545 16351 9601 16407
rect 9228 16016 9284 16072
rect 10714 16016 10770 16072
rect 8727 14146 8783 14202
rect 9545 14146 9601 14202
rect 10213 14146 10269 14202
rect 11031 14146 11087 14202
rect 9228 13811 9284 13867
rect 10714 13812 10770 13868
rect 8727 11941 8783 11997
rect 9545 11941 9601 11997
rect 10213 11942 10269 11998
rect 11031 11942 11087 11998
rect 9228 11606 9284 11662
rect 8727 9736 8783 9792
rect 9545 9736 9601 9792
rect 11340 9414 11396 9514
rect 7842 8904 7898 9004
rect 6171 2366 6227 2422
rect 6989 2366 7045 2422
rect 5186 2030 5242 2086
rect 4685 160 4741 216
rect 5503 160 5559 216
rect 3694 -165 3750 -65
rect 9228 8645 9284 8701
rect 8064 7676 8120 7732
rect 8727 6775 8783 6831
rect 9545 6775 9601 6831
rect 9228 6440 9284 6496
rect 10714 6440 10770 6496
rect 8727 4570 8783 4626
rect 9545 4570 9601 4626
rect 10213 4570 10269 4626
rect 11031 4570 11087 4626
rect 9228 4235 9284 4291
rect 10714 4236 10770 4292
rect 8727 2365 8783 2421
rect 9545 2365 9601 2421
rect 13270 18221 13326 18277
rect 12769 16351 12825 16407
rect 13587 16351 13643 16407
rect 13270 16016 13326 16072
rect 14756 16016 14812 16072
rect 12769 14146 12825 14202
rect 13587 14146 13643 14202
rect 14255 14146 14311 14202
rect 15073 14146 15129 14202
rect 13270 13811 13326 13867
rect 14756 13812 14812 13868
rect 12769 11941 12825 11997
rect 13587 11941 13643 11997
rect 14255 11942 14311 11998
rect 15073 11942 15129 11998
rect 13270 11606 13326 11662
rect 12769 9736 12825 9792
rect 13587 9736 13643 9792
rect 15382 9414 15438 9514
rect 11884 8904 11940 9004
rect 10213 2366 10269 2422
rect 11031 2366 11087 2422
rect 9228 2030 9284 2086
rect 8727 160 8783 216
rect 9545 160 9601 216
rect 7706 -165 7762 -65
rect 13270 8645 13326 8701
rect 12106 7676 12162 7732
rect 12769 6775 12825 6831
rect 13587 6775 13643 6831
rect 13270 6440 13326 6496
rect 14756 6440 14812 6496
rect 12769 4570 12825 4626
rect 13587 4570 13643 4626
rect 14255 4570 14311 4626
rect 15073 4570 15129 4626
rect 13270 4235 13326 4291
rect 14756 4236 14812 4292
rect 12769 2365 12825 2421
rect 13587 2365 13643 2421
rect 17312 18221 17368 18277
rect 16811 16351 16867 16407
rect 17629 16351 17685 16407
rect 17312 16016 17368 16072
rect 18798 16016 18854 16072
rect 16811 14146 16867 14202
rect 17629 14146 17685 14202
rect 18297 14146 18353 14202
rect 19115 14146 19171 14202
rect 17312 13811 17368 13867
rect 18798 13812 18854 13868
rect 16811 11941 16867 11997
rect 17629 11941 17685 11997
rect 18297 11942 18353 11998
rect 19115 11942 19171 11998
rect 17312 11606 17368 11662
rect 16811 9736 16867 9792
rect 17629 9736 17685 9792
rect 19424 9414 19480 9514
rect 15926 8904 15982 9004
rect 14255 2366 14311 2422
rect 15073 2366 15129 2422
rect 13270 2030 13326 2086
rect 12769 160 12825 216
rect 13587 160 13643 216
rect 11748 -165 11804 -65
rect 17312 8645 17368 8701
rect 16148 7676 16204 7732
rect 16811 6775 16867 6831
rect 17629 6775 17685 6831
rect 17312 6440 17368 6496
rect 18798 6440 18854 6496
rect 16811 4570 16867 4626
rect 17629 4570 17685 4626
rect 18297 4570 18353 4626
rect 19115 4570 19171 4626
rect 17312 4235 17368 4291
rect 18798 4236 18854 4292
rect 16811 2365 16867 2421
rect 17629 2365 17685 2421
rect 21354 18221 21410 18277
rect 20853 16351 20909 16407
rect 21671 16351 21727 16407
rect 21354 16016 21410 16072
rect 22840 16016 22896 16072
rect 20853 14146 20909 14202
rect 21671 14146 21727 14202
rect 22339 14146 22395 14202
rect 23157 14146 23213 14202
rect 21354 13811 21410 13867
rect 22840 13812 22896 13868
rect 20853 11941 20909 11997
rect 21671 11941 21727 11997
rect 22339 11942 22395 11998
rect 23157 11942 23213 11998
rect 21354 11606 21410 11662
rect 20853 9736 20909 9792
rect 21671 9736 21727 9792
rect 23466 9414 23522 9514
rect 19968 8904 20024 9004
rect 18297 2366 18353 2422
rect 19115 2366 19171 2422
rect 17312 2030 17368 2086
rect 16811 160 16867 216
rect 17629 160 17685 216
rect 15790 -165 15846 -65
rect 21354 8645 21410 8701
rect 20190 7676 20246 7732
rect 20853 6775 20909 6831
rect 21671 6775 21727 6831
rect 21354 6440 21410 6496
rect 22840 6440 22896 6496
rect 20853 4570 20909 4626
rect 21671 4570 21727 4626
rect 22339 4570 22395 4626
rect 23157 4570 23213 4626
rect 21354 4235 21410 4291
rect 22840 4236 22896 4292
rect 20853 2365 20909 2421
rect 21671 2365 21727 2421
rect 25396 18221 25452 18277
rect 24895 16351 24951 16407
rect 25713 16351 25769 16407
rect 25396 16016 25452 16072
rect 26882 16016 26938 16072
rect 24895 14146 24951 14202
rect 25713 14146 25769 14202
rect 26381 14146 26437 14202
rect 27199 14146 27255 14202
rect 25396 13811 25452 13867
rect 26882 13812 26938 13868
rect 24895 11941 24951 11997
rect 25713 11941 25769 11997
rect 26381 11942 26437 11998
rect 27199 11942 27255 11998
rect 25396 11606 25452 11662
rect 24895 9736 24951 9792
rect 25713 9736 25769 9792
rect 24010 8904 24066 9004
rect 22339 2366 22395 2422
rect 23157 2366 23213 2422
rect 21354 2030 21410 2086
rect 20853 160 20909 216
rect 21671 160 21727 216
rect 19832 -165 19888 -65
rect 25396 8645 25452 8701
rect 24232 7676 24288 7732
rect 24895 6775 24951 6831
rect 25713 6775 25769 6831
rect 25396 6440 25452 6496
rect 26882 6440 26938 6496
rect 24895 4570 24951 4626
rect 25713 4570 25769 4626
rect 26381 4570 26437 4626
rect 27199 4570 27255 4626
rect 25396 4235 25452 4291
rect 26882 4236 26938 4292
rect 24895 2365 24951 2421
rect 25713 2365 25769 2421
rect 29438 18221 29494 18277
rect 28173 14029 28229 14085
rect 28937 16351 28993 16407
rect 29755 16351 29811 16407
rect 29438 16016 29494 16072
rect 30924 16016 30980 16072
rect 28937 14146 28993 14202
rect 29755 14146 29811 14202
rect 30423 14146 30479 14202
rect 31241 14146 31297 14202
rect 29438 13811 29494 13867
rect 30924 13812 30980 13868
rect 28937 11941 28993 11997
rect 29755 11941 29811 11997
rect 30423 11942 30479 11998
rect 31241 11942 31297 11998
rect 29438 11606 29494 11662
rect 28173 10405 28229 10461
rect 28937 9736 28993 9792
rect 29755 9736 29811 9792
rect 28052 8904 28108 9004
rect 26381 2366 26437 2422
rect 27199 2366 27255 2422
rect 25396 2030 25452 2086
rect 24895 160 24951 216
rect 25713 160 25769 216
rect 23874 -165 23930 -65
<< metal3 >>
rect 5174 18280 5260 18284
rect 5174 18224 5186 18280
rect 5242 18224 5260 18280
rect 5174 18212 5260 18224
rect 9216 18277 9302 18281
rect 9216 18221 9228 18277
rect 9284 18221 9302 18277
rect 9216 18209 9302 18221
rect 13258 18277 13344 18281
rect 13258 18221 13270 18277
rect 13326 18221 13344 18277
rect 13258 18209 13344 18221
rect 17300 18277 17386 18281
rect 17300 18221 17312 18277
rect 17368 18221 17386 18277
rect 17300 18209 17386 18221
rect 21342 18277 21428 18281
rect 21342 18221 21354 18277
rect 21410 18221 21428 18277
rect 21342 18209 21428 18221
rect 25384 18277 25470 18281
rect 25384 18221 25396 18277
rect 25452 18221 25470 18277
rect 25384 18209 25470 18221
rect 29426 18277 29512 18281
rect 29426 18221 29438 18277
rect 29494 18221 29512 18277
rect 29426 18209 29512 18221
rect 4673 16410 4753 16422
rect 4673 16354 4685 16410
rect 4741 16354 4753 16410
rect 4673 16342 4753 16354
rect 5491 16410 5571 16422
rect 5491 16354 5503 16410
rect 5559 16354 5571 16410
rect 5491 16342 5571 16354
rect 8715 16407 8795 16419
rect 8715 16351 8727 16407
rect 8783 16351 8795 16407
rect 8715 16339 8795 16351
rect 9533 16407 9613 16419
rect 9533 16351 9545 16407
rect 9601 16351 9613 16407
rect 9533 16339 9613 16351
rect 12757 16407 12837 16419
rect 12757 16351 12769 16407
rect 12825 16351 12837 16407
rect 12757 16339 12837 16351
rect 13575 16407 13655 16419
rect 13575 16351 13587 16407
rect 13643 16351 13655 16407
rect 13575 16339 13655 16351
rect 16799 16407 16879 16419
rect 16799 16351 16811 16407
rect 16867 16351 16879 16407
rect 16799 16339 16879 16351
rect 17617 16407 17697 16419
rect 17617 16351 17629 16407
rect 17685 16351 17697 16407
rect 17617 16339 17697 16351
rect 20841 16407 20921 16419
rect 20841 16351 20853 16407
rect 20909 16351 20921 16407
rect 20841 16339 20921 16351
rect 21659 16407 21739 16419
rect 21659 16351 21671 16407
rect 21727 16351 21739 16407
rect 21659 16339 21739 16351
rect 24883 16407 24963 16419
rect 24883 16351 24895 16407
rect 24951 16351 24963 16407
rect 24883 16339 24963 16351
rect 25701 16407 25781 16419
rect 25701 16351 25713 16407
rect 25769 16351 25781 16407
rect 25701 16339 25781 16351
rect 28925 16407 29005 16419
rect 28925 16351 28937 16407
rect 28993 16351 29005 16407
rect 28925 16339 29005 16351
rect 29743 16407 29823 16419
rect 29743 16351 29755 16407
rect 29811 16351 29823 16407
rect 29743 16339 29823 16351
rect 5174 16075 5260 16079
rect 5174 16019 5186 16075
rect 5242 16019 5260 16075
rect 5174 16007 5260 16019
rect 6660 16075 6746 16079
rect 6660 16019 6672 16075
rect 6728 16019 6746 16075
rect 6660 16007 6746 16019
rect 9216 16072 9302 16076
rect 9216 16016 9228 16072
rect 9284 16016 9302 16072
rect 9216 16004 9302 16016
rect 10702 16072 10788 16076
rect 10702 16016 10714 16072
rect 10770 16016 10788 16072
rect 10702 16004 10788 16016
rect 13258 16072 13344 16076
rect 13258 16016 13270 16072
rect 13326 16016 13344 16072
rect 13258 16004 13344 16016
rect 14744 16072 14830 16076
rect 14744 16016 14756 16072
rect 14812 16016 14830 16072
rect 14744 16004 14830 16016
rect 17300 16072 17386 16076
rect 17300 16016 17312 16072
rect 17368 16016 17386 16072
rect 17300 16004 17386 16016
rect 18786 16072 18872 16076
rect 18786 16016 18798 16072
rect 18854 16016 18872 16072
rect 18786 16004 18872 16016
rect 21342 16072 21428 16076
rect 21342 16016 21354 16072
rect 21410 16016 21428 16072
rect 21342 16004 21428 16016
rect 22828 16072 22914 16076
rect 22828 16016 22840 16072
rect 22896 16016 22914 16072
rect 22828 16004 22914 16016
rect 25384 16072 25470 16076
rect 25384 16016 25396 16072
rect 25452 16016 25470 16072
rect 25384 16004 25470 16016
rect 26870 16072 26956 16076
rect 26870 16016 26882 16072
rect 26938 16016 26956 16072
rect 26870 16004 26956 16016
rect 29426 16072 29512 16076
rect 29426 16016 29438 16072
rect 29494 16016 29512 16072
rect 29426 16004 29512 16016
rect 30912 16072 30998 16076
rect 30912 16016 30924 16072
rect 30980 16016 30998 16072
rect 30912 16004 30998 16016
rect 4673 14205 4753 14217
rect 4673 14149 4685 14205
rect 4741 14149 4753 14205
rect 4673 14137 4753 14149
rect 5491 14205 5571 14217
rect 5491 14149 5503 14205
rect 5559 14149 5571 14205
rect 5491 14137 5571 14149
rect 6159 14205 6239 14217
rect 6159 14149 6171 14205
rect 6227 14149 6239 14205
rect 6159 14137 6239 14149
rect 6977 14205 7057 14217
rect 6977 14149 6989 14205
rect 7045 14149 7057 14205
rect 6977 14137 7057 14149
rect 8715 14202 8795 14214
rect 8715 14146 8727 14202
rect 8783 14146 8795 14202
rect 8715 14134 8795 14146
rect 9533 14202 9613 14214
rect 9533 14146 9545 14202
rect 9601 14146 9613 14202
rect 9533 14134 9613 14146
rect 10201 14202 10281 14214
rect 10201 14146 10213 14202
rect 10269 14146 10281 14202
rect 10201 14134 10281 14146
rect 11019 14202 11099 14214
rect 11019 14146 11031 14202
rect 11087 14146 11099 14202
rect 11019 14134 11099 14146
rect 12757 14202 12837 14214
rect 12757 14146 12769 14202
rect 12825 14146 12837 14202
rect 12757 14134 12837 14146
rect 13575 14202 13655 14214
rect 13575 14146 13587 14202
rect 13643 14146 13655 14202
rect 13575 14134 13655 14146
rect 14243 14202 14323 14214
rect 14243 14146 14255 14202
rect 14311 14146 14323 14202
rect 14243 14134 14323 14146
rect 15061 14202 15141 14214
rect 15061 14146 15073 14202
rect 15129 14146 15141 14202
rect 15061 14134 15141 14146
rect 16799 14202 16879 14214
rect 16799 14146 16811 14202
rect 16867 14146 16879 14202
rect 16799 14134 16879 14146
rect 17617 14202 17697 14214
rect 17617 14146 17629 14202
rect 17685 14146 17697 14202
rect 17617 14134 17697 14146
rect 18285 14202 18365 14214
rect 18285 14146 18297 14202
rect 18353 14146 18365 14202
rect 18285 14134 18365 14146
rect 19103 14202 19183 14214
rect 19103 14146 19115 14202
rect 19171 14146 19183 14202
rect 19103 14134 19183 14146
rect 20841 14202 20921 14214
rect 20841 14146 20853 14202
rect 20909 14146 20921 14202
rect 20841 14134 20921 14146
rect 21659 14202 21739 14214
rect 21659 14146 21671 14202
rect 21727 14146 21739 14202
rect 21659 14134 21739 14146
rect 22327 14202 22407 14214
rect 22327 14146 22339 14202
rect 22395 14146 22407 14202
rect 22327 14134 22407 14146
rect 23145 14202 23225 14214
rect 23145 14146 23157 14202
rect 23213 14146 23225 14202
rect 23145 14134 23225 14146
rect 24883 14202 24963 14214
rect 24883 14146 24895 14202
rect 24951 14146 24963 14202
rect 24883 14134 24963 14146
rect 25701 14202 25781 14214
rect 25701 14146 25713 14202
rect 25769 14146 25781 14202
rect 25701 14134 25781 14146
rect 26369 14202 26449 14214
rect 26369 14146 26381 14202
rect 26437 14146 26449 14202
rect 26369 14134 26449 14146
rect 27187 14202 27267 14214
rect 27187 14146 27199 14202
rect 27255 14146 27267 14202
rect 27187 14134 27267 14146
rect 28925 14202 29005 14214
rect 28925 14146 28937 14202
rect 28993 14146 29005 14202
rect 28925 14134 29005 14146
rect 29743 14202 29823 14214
rect 29743 14146 29755 14202
rect 29811 14146 29823 14202
rect 29743 14134 29823 14146
rect 30411 14202 30491 14214
rect 30411 14146 30423 14202
rect 30479 14146 30491 14202
rect 30411 14134 30491 14146
rect 31229 14202 31309 14214
rect 31229 14146 31241 14202
rect 31297 14146 31309 14202
rect 31229 14134 31309 14146
rect 28162 14085 28240 14097
rect 28162 14029 28173 14085
rect 28229 14029 28240 14085
rect 28162 14017 28240 14029
rect 5174 13870 5260 13874
rect 5174 13814 5186 13870
rect 5242 13814 5260 13870
rect 5174 13802 5260 13814
rect 6660 13871 6746 13875
rect 6660 13815 6672 13871
rect 6728 13815 6746 13871
rect 6660 13803 6746 13815
rect 9216 13867 9302 13871
rect 9216 13811 9228 13867
rect 9284 13811 9302 13867
rect 9216 13799 9302 13811
rect 10702 13868 10788 13872
rect 10702 13812 10714 13868
rect 10770 13812 10788 13868
rect 10702 13800 10788 13812
rect 13258 13867 13344 13871
rect 13258 13811 13270 13867
rect 13326 13811 13344 13867
rect 13258 13799 13344 13811
rect 14744 13868 14830 13872
rect 14744 13812 14756 13868
rect 14812 13812 14830 13868
rect 14744 13800 14830 13812
rect 17300 13867 17386 13871
rect 17300 13811 17312 13867
rect 17368 13811 17386 13867
rect 17300 13799 17386 13811
rect 18786 13868 18872 13872
rect 18786 13812 18798 13868
rect 18854 13812 18872 13868
rect 18786 13800 18872 13812
rect 21342 13867 21428 13871
rect 21342 13811 21354 13867
rect 21410 13811 21428 13867
rect 21342 13799 21428 13811
rect 22828 13868 22914 13872
rect 22828 13812 22840 13868
rect 22896 13812 22914 13868
rect 22828 13800 22914 13812
rect 25384 13867 25470 13871
rect 25384 13811 25396 13867
rect 25452 13811 25470 13867
rect 25384 13799 25470 13811
rect 26870 13868 26956 13872
rect 26870 13812 26882 13868
rect 26938 13812 26956 13868
rect 26870 13800 26956 13812
rect 29426 13867 29512 13871
rect 29426 13811 29438 13867
rect 29494 13811 29512 13867
rect 29426 13799 29512 13811
rect 30912 13868 30998 13872
rect 30912 13812 30924 13868
rect 30980 13812 30998 13868
rect 30912 13800 30998 13812
rect 4673 12000 4753 12012
rect 4673 11944 4685 12000
rect 4741 11944 4753 12000
rect 4673 11932 4753 11944
rect 5491 12000 5571 12012
rect 5491 11944 5503 12000
rect 5559 11944 5571 12000
rect 5491 11932 5571 11944
rect 6159 12001 6239 12013
rect 6159 11945 6171 12001
rect 6227 11945 6239 12001
rect 6159 11933 6239 11945
rect 6977 12001 7057 12013
rect 6977 11945 6989 12001
rect 7045 11945 7057 12001
rect 6977 11933 7057 11945
rect 8715 11997 8795 12009
rect 8715 11941 8727 11997
rect 8783 11941 8795 11997
rect 8715 11929 8795 11941
rect 9533 11997 9613 12009
rect 9533 11941 9545 11997
rect 9601 11941 9613 11997
rect 9533 11929 9613 11941
rect 10201 11998 10281 12010
rect 10201 11942 10213 11998
rect 10269 11942 10281 11998
rect 10201 11930 10281 11942
rect 11019 11998 11099 12010
rect 11019 11942 11031 11998
rect 11087 11942 11099 11998
rect 11019 11930 11099 11942
rect 12757 11997 12837 12009
rect 12757 11941 12769 11997
rect 12825 11941 12837 11997
rect 12757 11929 12837 11941
rect 13575 11997 13655 12009
rect 13575 11941 13587 11997
rect 13643 11941 13655 11997
rect 13575 11929 13655 11941
rect 14243 11998 14323 12010
rect 14243 11942 14255 11998
rect 14311 11942 14323 11998
rect 14243 11930 14323 11942
rect 15061 11998 15141 12010
rect 15061 11942 15073 11998
rect 15129 11942 15141 11998
rect 15061 11930 15141 11942
rect 16799 11997 16879 12009
rect 16799 11941 16811 11997
rect 16867 11941 16879 11997
rect 16799 11929 16879 11941
rect 17617 11997 17697 12009
rect 17617 11941 17629 11997
rect 17685 11941 17697 11997
rect 17617 11929 17697 11941
rect 18285 11998 18365 12010
rect 18285 11942 18297 11998
rect 18353 11942 18365 11998
rect 18285 11930 18365 11942
rect 19103 11998 19183 12010
rect 19103 11942 19115 11998
rect 19171 11942 19183 11998
rect 19103 11930 19183 11942
rect 20841 11997 20921 12009
rect 20841 11941 20853 11997
rect 20909 11941 20921 11997
rect 20841 11929 20921 11941
rect 21659 11997 21739 12009
rect 21659 11941 21671 11997
rect 21727 11941 21739 11997
rect 21659 11929 21739 11941
rect 22327 11998 22407 12010
rect 22327 11942 22339 11998
rect 22395 11942 22407 11998
rect 22327 11930 22407 11942
rect 23145 11998 23225 12010
rect 23145 11942 23157 11998
rect 23213 11942 23225 11998
rect 23145 11930 23225 11942
rect 24883 11997 24963 12009
rect 24883 11941 24895 11997
rect 24951 11941 24963 11997
rect 24883 11929 24963 11941
rect 25701 11997 25781 12009
rect 25701 11941 25713 11997
rect 25769 11941 25781 11997
rect 25701 11929 25781 11941
rect 26369 11998 26449 12010
rect 26369 11942 26381 11998
rect 26437 11942 26449 11998
rect 26369 11930 26449 11942
rect 27187 11998 27267 12010
rect 27187 11942 27199 11998
rect 27255 11942 27267 11998
rect 27187 11930 27267 11942
rect 28925 11997 29005 12009
rect 28925 11941 28937 11997
rect 28993 11941 29005 11997
rect 28925 11929 29005 11941
rect 29743 11997 29823 12009
rect 29743 11941 29755 11997
rect 29811 11941 29823 11997
rect 29743 11929 29823 11941
rect 30411 11998 30491 12010
rect 30411 11942 30423 11998
rect 30479 11942 30491 11998
rect 30411 11930 30491 11942
rect 31229 11998 31309 12010
rect 31229 11942 31241 11998
rect 31297 11942 31309 11998
rect 31229 11930 31309 11942
rect 5174 11665 5260 11669
rect 5174 11609 5186 11665
rect 5242 11609 5260 11665
rect 5174 11597 5260 11609
rect 9216 11662 9302 11666
rect 9216 11606 9228 11662
rect 9284 11606 9302 11662
rect 9216 11594 9302 11606
rect 13258 11662 13344 11666
rect 13258 11606 13270 11662
rect 13326 11606 13344 11662
rect 13258 11594 13344 11606
rect 17300 11662 17386 11666
rect 17300 11606 17312 11662
rect 17368 11606 17386 11662
rect 17300 11594 17386 11606
rect 21342 11662 21428 11666
rect 21342 11606 21354 11662
rect 21410 11606 21428 11662
rect 21342 11594 21428 11606
rect 25384 11662 25470 11666
rect 25384 11606 25396 11662
rect 25452 11606 25470 11662
rect 25384 11594 25470 11606
rect 29426 11662 29512 11666
rect 29426 11606 29438 11662
rect 29494 11606 29512 11662
rect 29426 11594 29512 11606
rect 28162 10461 28240 10473
rect 28162 10405 28173 10461
rect 28229 10405 28240 10461
rect 28162 10393 28240 10405
rect 4673 9795 4753 9807
rect 4673 9739 4685 9795
rect 4741 9739 4753 9795
rect 4673 9727 4753 9739
rect 5491 9795 5571 9807
rect 5491 9739 5503 9795
rect 5559 9739 5571 9795
rect 5491 9727 5571 9739
rect 8715 9792 8795 9804
rect 8715 9736 8727 9792
rect 8783 9736 8795 9792
rect 8715 9724 8795 9736
rect 9533 9792 9613 9804
rect 9533 9736 9545 9792
rect 9601 9736 9613 9792
rect 9533 9724 9613 9736
rect 12757 9792 12837 9804
rect 12757 9736 12769 9792
rect 12825 9736 12837 9792
rect 12757 9724 12837 9736
rect 13575 9792 13655 9804
rect 13575 9736 13587 9792
rect 13643 9736 13655 9792
rect 13575 9724 13655 9736
rect 16799 9792 16879 9804
rect 16799 9736 16811 9792
rect 16867 9736 16879 9792
rect 16799 9724 16879 9736
rect 17617 9792 17697 9804
rect 17617 9736 17629 9792
rect 17685 9736 17697 9792
rect 17617 9724 17697 9736
rect 20841 9792 20921 9804
rect 20841 9736 20853 9792
rect 20909 9736 20921 9792
rect 20841 9724 20921 9736
rect 21659 9792 21739 9804
rect 21659 9736 21671 9792
rect 21727 9736 21739 9792
rect 21659 9724 21739 9736
rect 24883 9792 24963 9804
rect 24883 9736 24895 9792
rect 24951 9736 24963 9792
rect 24883 9724 24963 9736
rect 25701 9792 25781 9804
rect 25701 9736 25713 9792
rect 25769 9736 25781 9792
rect 25701 9724 25781 9736
rect 28925 9792 29005 9804
rect 28925 9736 28937 9792
rect 28993 9736 29005 9792
rect 28925 9724 29005 9736
rect 29743 9792 29823 9804
rect 29743 9736 29755 9792
rect 29811 9736 29823 9792
rect 29743 9724 29823 9736
rect -56 9414 -46 9514
rect 10 9414 3286 9514
rect 3342 9414 7298 9514
rect 7354 9414 11340 9514
rect 11396 9414 15382 9514
rect 15438 9414 19424 9514
rect 19480 9414 23466 9514
rect 23522 9414 23532 9514
rect 3820 9004 3830 9007
rect -56 8904 -46 9004
rect 10 8907 3830 9004
rect 3886 9004 3896 9007
rect 3886 8907 7842 9004
rect 10 8904 7842 8907
rect 7898 8904 11884 9004
rect 11940 8904 15926 9004
rect 15982 8904 19968 9004
rect 20024 8904 24010 9004
rect 24066 8904 28052 9004
rect 28108 8904 28118 9004
rect 1162 8701 1248 8705
rect 1162 8645 1174 8701
rect 1230 8645 1248 8701
rect 1162 8633 1248 8645
rect 5174 8701 5260 8705
rect 5174 8645 5186 8701
rect 5242 8645 5260 8701
rect 5174 8633 5260 8645
rect 9216 8701 9302 8705
rect 9216 8645 9228 8701
rect 9284 8645 9302 8701
rect 9216 8633 9302 8645
rect 13258 8701 13344 8705
rect 13258 8645 13270 8701
rect 13326 8645 13344 8701
rect 13258 8633 13344 8645
rect 17300 8701 17386 8705
rect 17300 8645 17312 8701
rect 17368 8645 17386 8701
rect 17300 8633 17386 8645
rect 21342 8701 21428 8705
rect 21342 8645 21354 8701
rect 21410 8645 21428 8701
rect 21342 8633 21428 8645
rect 25384 8701 25470 8705
rect 25384 8645 25396 8701
rect 25452 8645 25470 8701
rect 25384 8633 25470 8645
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 661 6831 741 6843
rect 661 6775 673 6831
rect 729 6775 741 6831
rect 661 6763 741 6775
rect 1479 6831 1559 6843
rect 1479 6775 1491 6831
rect 1547 6775 1559 6831
rect 1479 6763 1559 6775
rect 4673 6831 4753 6843
rect 4673 6775 4685 6831
rect 4741 6775 4753 6831
rect 4673 6763 4753 6775
rect 5491 6831 5571 6843
rect 5491 6775 5503 6831
rect 5559 6775 5571 6831
rect 5491 6763 5571 6775
rect 8715 6831 8795 6843
rect 8715 6775 8727 6831
rect 8783 6775 8795 6831
rect 8715 6763 8795 6775
rect 9533 6831 9613 6843
rect 9533 6775 9545 6831
rect 9601 6775 9613 6831
rect 9533 6763 9613 6775
rect 12757 6831 12837 6843
rect 12757 6775 12769 6831
rect 12825 6775 12837 6831
rect 12757 6763 12837 6775
rect 13575 6831 13655 6843
rect 13575 6775 13587 6831
rect 13643 6775 13655 6831
rect 13575 6763 13655 6775
rect 16799 6831 16879 6843
rect 16799 6775 16811 6831
rect 16867 6775 16879 6831
rect 16799 6763 16879 6775
rect 17617 6831 17697 6843
rect 17617 6775 17629 6831
rect 17685 6775 17697 6831
rect 17617 6763 17697 6775
rect 20841 6831 20921 6843
rect 20841 6775 20853 6831
rect 20909 6775 20921 6831
rect 20841 6763 20921 6775
rect 21659 6831 21739 6843
rect 21659 6775 21671 6831
rect 21727 6775 21739 6831
rect 21659 6763 21739 6775
rect 24883 6831 24963 6843
rect 24883 6775 24895 6831
rect 24951 6775 24963 6831
rect 24883 6763 24963 6775
rect 25701 6831 25781 6843
rect 25701 6775 25713 6831
rect 25769 6775 25781 6831
rect 25701 6763 25781 6775
rect 1162 6496 1248 6500
rect 1162 6440 1174 6496
rect 1230 6440 1248 6496
rect 1162 6428 1248 6440
rect 2648 6496 2734 6500
rect 2648 6440 2660 6496
rect 2716 6440 2734 6496
rect 2648 6428 2734 6440
rect 5174 6496 5260 6500
rect 5174 6440 5186 6496
rect 5242 6440 5260 6496
rect 5174 6428 5260 6440
rect 6660 6496 6746 6500
rect 6660 6440 6672 6496
rect 6728 6440 6746 6496
rect 6660 6428 6746 6440
rect 9216 6496 9302 6500
rect 9216 6440 9228 6496
rect 9284 6440 9302 6496
rect 9216 6428 9302 6440
rect 10702 6496 10788 6500
rect 10702 6440 10714 6496
rect 10770 6440 10788 6496
rect 10702 6428 10788 6440
rect 13258 6496 13344 6500
rect 13258 6440 13270 6496
rect 13326 6440 13344 6496
rect 13258 6428 13344 6440
rect 14744 6496 14830 6500
rect 14744 6440 14756 6496
rect 14812 6440 14830 6496
rect 14744 6428 14830 6440
rect 17300 6496 17386 6500
rect 17300 6440 17312 6496
rect 17368 6440 17386 6496
rect 17300 6428 17386 6440
rect 18786 6496 18872 6500
rect 18786 6440 18798 6496
rect 18854 6440 18872 6496
rect 18786 6428 18872 6440
rect 21342 6496 21428 6500
rect 21342 6440 21354 6496
rect 21410 6440 21428 6496
rect 21342 6428 21428 6440
rect 22828 6496 22914 6500
rect 22828 6440 22840 6496
rect 22896 6440 22914 6496
rect 22828 6428 22914 6440
rect 25384 6496 25470 6500
rect 25384 6440 25396 6496
rect 25452 6440 25470 6496
rect 25384 6428 25470 6440
rect 26870 6496 26956 6500
rect 26870 6440 26882 6496
rect 26938 6440 26956 6496
rect 26870 6428 26956 6440
rect 661 4626 741 4638
rect 661 4570 673 4626
rect 729 4570 741 4626
rect 661 4558 741 4570
rect 1479 4626 1559 4638
rect 1479 4570 1491 4626
rect 1547 4570 1559 4626
rect 1479 4558 1559 4570
rect 2147 4626 2227 4638
rect 2147 4570 2159 4626
rect 2215 4570 2227 4626
rect 2147 4558 2227 4570
rect 2965 4626 3045 4638
rect 2965 4570 2977 4626
rect 3033 4570 3045 4626
rect 2965 4558 3045 4570
rect 4673 4626 4753 4638
rect 4673 4570 4685 4626
rect 4741 4570 4753 4626
rect 4673 4558 4753 4570
rect 5491 4626 5571 4638
rect 5491 4570 5503 4626
rect 5559 4570 5571 4626
rect 5491 4558 5571 4570
rect 6159 4626 6239 4638
rect 6159 4570 6171 4626
rect 6227 4570 6239 4626
rect 6159 4558 6239 4570
rect 6977 4626 7057 4638
rect 6977 4570 6989 4626
rect 7045 4570 7057 4626
rect 6977 4558 7057 4570
rect 8715 4626 8795 4638
rect 8715 4570 8727 4626
rect 8783 4570 8795 4626
rect 8715 4558 8795 4570
rect 9533 4626 9613 4638
rect 9533 4570 9545 4626
rect 9601 4570 9613 4626
rect 9533 4558 9613 4570
rect 10201 4626 10281 4638
rect 10201 4570 10213 4626
rect 10269 4570 10281 4626
rect 10201 4558 10281 4570
rect 11019 4626 11099 4638
rect 11019 4570 11031 4626
rect 11087 4570 11099 4626
rect 11019 4558 11099 4570
rect 12757 4626 12837 4638
rect 12757 4570 12769 4626
rect 12825 4570 12837 4626
rect 12757 4558 12837 4570
rect 13575 4626 13655 4638
rect 13575 4570 13587 4626
rect 13643 4570 13655 4626
rect 13575 4558 13655 4570
rect 14243 4626 14323 4638
rect 14243 4570 14255 4626
rect 14311 4570 14323 4626
rect 14243 4558 14323 4570
rect 15061 4626 15141 4638
rect 15061 4570 15073 4626
rect 15129 4570 15141 4626
rect 15061 4558 15141 4570
rect 16799 4626 16879 4638
rect 16799 4570 16811 4626
rect 16867 4570 16879 4626
rect 16799 4558 16879 4570
rect 17617 4626 17697 4638
rect 17617 4570 17629 4626
rect 17685 4570 17697 4626
rect 17617 4558 17697 4570
rect 18285 4626 18365 4638
rect 18285 4570 18297 4626
rect 18353 4570 18365 4626
rect 18285 4558 18365 4570
rect 19103 4626 19183 4638
rect 19103 4570 19115 4626
rect 19171 4570 19183 4626
rect 19103 4558 19183 4570
rect 20841 4626 20921 4638
rect 20841 4570 20853 4626
rect 20909 4570 20921 4626
rect 20841 4558 20921 4570
rect 21659 4626 21739 4638
rect 21659 4570 21671 4626
rect 21727 4570 21739 4626
rect 21659 4558 21739 4570
rect 22327 4626 22407 4638
rect 22327 4570 22339 4626
rect 22395 4570 22407 4626
rect 22327 4558 22407 4570
rect 23145 4626 23225 4638
rect 23145 4570 23157 4626
rect 23213 4570 23225 4626
rect 23145 4558 23225 4570
rect 24883 4626 24963 4638
rect 24883 4570 24895 4626
rect 24951 4570 24963 4626
rect 24883 4558 24963 4570
rect 25701 4626 25781 4638
rect 25701 4570 25713 4626
rect 25769 4570 25781 4626
rect 25701 4558 25781 4570
rect 26369 4626 26449 4638
rect 26369 4570 26381 4626
rect 26437 4570 26449 4626
rect 26369 4558 26449 4570
rect 27187 4626 27267 4638
rect 27187 4570 27199 4626
rect 27255 4570 27267 4626
rect 27187 4558 27267 4570
rect 1162 4291 1248 4295
rect 1162 4235 1174 4291
rect 1230 4235 1248 4291
rect 1162 4223 1248 4235
rect 2648 4292 2734 4296
rect 2648 4236 2660 4292
rect 2716 4236 2734 4292
rect 2648 4224 2734 4236
rect 5174 4291 5260 4295
rect 5174 4235 5186 4291
rect 5242 4235 5260 4291
rect 5174 4223 5260 4235
rect 6660 4292 6746 4296
rect 6660 4236 6672 4292
rect 6728 4236 6746 4292
rect 6660 4224 6746 4236
rect 9216 4291 9302 4295
rect 9216 4235 9228 4291
rect 9284 4235 9302 4291
rect 9216 4223 9302 4235
rect 10702 4292 10788 4296
rect 10702 4236 10714 4292
rect 10770 4236 10788 4292
rect 10702 4224 10788 4236
rect 13258 4291 13344 4295
rect 13258 4235 13270 4291
rect 13326 4235 13344 4291
rect 13258 4223 13344 4235
rect 14744 4292 14830 4296
rect 14744 4236 14756 4292
rect 14812 4236 14830 4292
rect 14744 4224 14830 4236
rect 17300 4291 17386 4295
rect 17300 4235 17312 4291
rect 17368 4235 17386 4291
rect 17300 4223 17386 4235
rect 18786 4292 18872 4296
rect 18786 4236 18798 4292
rect 18854 4236 18872 4292
rect 18786 4224 18872 4236
rect 21342 4291 21428 4295
rect 21342 4235 21354 4291
rect 21410 4235 21428 4291
rect 21342 4223 21428 4235
rect 22828 4292 22914 4296
rect 22828 4236 22840 4292
rect 22896 4236 22914 4292
rect 22828 4224 22914 4236
rect 25384 4291 25470 4295
rect 25384 4235 25396 4291
rect 25452 4235 25470 4291
rect 25384 4223 25470 4235
rect 26870 4292 26956 4296
rect 26870 4236 26882 4292
rect 26938 4236 26956 4292
rect 26870 4224 26956 4236
rect 661 2421 741 2433
rect 661 2365 673 2421
rect 729 2365 741 2421
rect 661 2353 741 2365
rect 1479 2421 1559 2433
rect 1479 2365 1491 2421
rect 1547 2365 1559 2421
rect 1479 2353 1559 2365
rect 2147 2422 2227 2434
rect 2147 2366 2159 2422
rect 2215 2366 2227 2422
rect 2147 2354 2227 2366
rect 2965 2422 3045 2434
rect 2965 2366 2977 2422
rect 3033 2366 3045 2422
rect 2965 2354 3045 2366
rect 4673 2421 4753 2433
rect 4673 2365 4685 2421
rect 4741 2365 4753 2421
rect 4673 2353 4753 2365
rect 5491 2421 5571 2433
rect 5491 2365 5503 2421
rect 5559 2365 5571 2421
rect 5491 2353 5571 2365
rect 6159 2422 6239 2434
rect 6159 2366 6171 2422
rect 6227 2366 6239 2422
rect 6159 2354 6239 2366
rect 6977 2422 7057 2434
rect 6977 2366 6989 2422
rect 7045 2366 7057 2422
rect 6977 2354 7057 2366
rect 8715 2421 8795 2433
rect 8715 2365 8727 2421
rect 8783 2365 8795 2421
rect 8715 2353 8795 2365
rect 9533 2421 9613 2433
rect 9533 2365 9545 2421
rect 9601 2365 9613 2421
rect 9533 2353 9613 2365
rect 10201 2422 10281 2434
rect 10201 2366 10213 2422
rect 10269 2366 10281 2422
rect 10201 2354 10281 2366
rect 11019 2422 11099 2434
rect 11019 2366 11031 2422
rect 11087 2366 11099 2422
rect 11019 2354 11099 2366
rect 12757 2421 12837 2433
rect 12757 2365 12769 2421
rect 12825 2365 12837 2421
rect 12757 2353 12837 2365
rect 13575 2421 13655 2433
rect 13575 2365 13587 2421
rect 13643 2365 13655 2421
rect 13575 2353 13655 2365
rect 14243 2422 14323 2434
rect 14243 2366 14255 2422
rect 14311 2366 14323 2422
rect 14243 2354 14323 2366
rect 15061 2422 15141 2434
rect 15061 2366 15073 2422
rect 15129 2366 15141 2422
rect 15061 2354 15141 2366
rect 16799 2421 16879 2433
rect 16799 2365 16811 2421
rect 16867 2365 16879 2421
rect 16799 2353 16879 2365
rect 17617 2421 17697 2433
rect 17617 2365 17629 2421
rect 17685 2365 17697 2421
rect 17617 2353 17697 2365
rect 18285 2422 18365 2434
rect 18285 2366 18297 2422
rect 18353 2366 18365 2422
rect 18285 2354 18365 2366
rect 19103 2422 19183 2434
rect 19103 2366 19115 2422
rect 19171 2366 19183 2422
rect 19103 2354 19183 2366
rect 20841 2421 20921 2433
rect 20841 2365 20853 2421
rect 20909 2365 20921 2421
rect 20841 2353 20921 2365
rect 21659 2421 21739 2433
rect 21659 2365 21671 2421
rect 21727 2365 21739 2421
rect 21659 2353 21739 2365
rect 22327 2422 22407 2434
rect 22327 2366 22339 2422
rect 22395 2366 22407 2422
rect 22327 2354 22407 2366
rect 23145 2422 23225 2434
rect 23145 2366 23157 2422
rect 23213 2366 23225 2422
rect 23145 2354 23225 2366
rect 24883 2421 24963 2433
rect 24883 2365 24895 2421
rect 24951 2365 24963 2421
rect 24883 2353 24963 2365
rect 25701 2421 25781 2433
rect 25701 2365 25713 2421
rect 25769 2365 25781 2421
rect 25701 2353 25781 2365
rect 26369 2422 26449 2434
rect 26369 2366 26381 2422
rect 26437 2366 26449 2422
rect 26369 2354 26449 2366
rect 27187 2422 27267 2434
rect 27187 2366 27199 2422
rect 27255 2366 27267 2422
rect 27187 2354 27267 2366
rect 1162 2086 1248 2090
rect 1162 2030 1174 2086
rect 1230 2030 1248 2086
rect 1162 2018 1248 2030
rect 5174 2086 5260 2090
rect 5174 2030 5186 2086
rect 5242 2030 5260 2086
rect 5174 2018 5260 2030
rect 9216 2086 9302 2090
rect 9216 2030 9228 2086
rect 9284 2030 9302 2086
rect 9216 2018 9302 2030
rect 13258 2086 13344 2090
rect 13258 2030 13270 2086
rect 13326 2030 13344 2086
rect 13258 2018 13344 2030
rect 17300 2086 17386 2090
rect 17300 2030 17312 2086
rect 17368 2030 17386 2086
rect 17300 2018 17386 2030
rect 21342 2086 21428 2090
rect 21342 2030 21354 2086
rect 21410 2030 21428 2086
rect 21342 2018 21428 2030
rect 25384 2086 25470 2090
rect 25384 2030 25396 2086
rect 25452 2030 25470 2086
rect 25384 2018 25470 2030
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect 661 216 741 228
rect 661 160 673 216
rect 729 160 741 216
rect 661 148 741 160
rect 1479 216 1559 228
rect 1479 160 1491 216
rect 1547 160 1559 216
rect 1479 148 1559 160
rect 4673 216 4753 228
rect 4673 160 4685 216
rect 4741 160 4753 216
rect 4673 148 4753 160
rect 5491 216 5571 228
rect 5491 160 5503 216
rect 5559 160 5571 216
rect 5491 148 5571 160
rect 8715 216 8795 228
rect 8715 160 8727 216
rect 8783 160 8795 216
rect 8715 148 8795 160
rect 9533 216 9613 228
rect 9533 160 9545 216
rect 9601 160 9613 216
rect 9533 148 9613 160
rect 12757 216 12837 228
rect 12757 160 12769 216
rect 12825 160 12837 216
rect 12757 148 12837 160
rect 13575 216 13655 228
rect 13575 160 13587 216
rect 13643 160 13655 216
rect 13575 148 13655 160
rect 16799 216 16879 228
rect 16799 160 16811 216
rect 16867 160 16879 216
rect 16799 148 16879 160
rect 17617 216 17697 228
rect 17617 160 17629 216
rect 17685 160 17697 216
rect 17617 148 17697 160
rect 20841 216 20921 228
rect 20841 160 20853 216
rect 20909 160 20921 216
rect 20841 148 20921 160
rect 21659 216 21739 228
rect 21659 160 21671 216
rect 21727 160 21739 216
rect 21659 148 21739 160
rect 24883 216 24963 228
rect 24883 160 24895 216
rect 24951 160 24963 216
rect 24883 148 24963 160
rect 25701 216 25781 228
rect 25701 160 25713 216
rect 25769 160 25781 216
rect 25701 148 25781 160
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect -328 -165 -318 -65
rect -262 -165 3694 -65
rect 3750 -165 7706 -65
rect 7762 -165 11748 -65
rect 11804 -165 15790 -65
rect 15846 -165 19832 -65
rect 19888 -165 23874 -65
rect 23930 -165 23940 -65
<< via3 >>
rect 5186 18224 5242 18280
rect 9228 18221 9284 18277
rect 13270 18221 13326 18277
rect 17312 18221 17368 18277
rect 21354 18221 21410 18277
rect 25396 18221 25452 18277
rect 29438 18221 29494 18277
rect 4685 16354 4741 16410
rect 5503 16354 5559 16410
rect 8727 16351 8783 16407
rect 9545 16351 9601 16407
rect 12769 16351 12825 16407
rect 13587 16351 13643 16407
rect 16811 16351 16867 16407
rect 17629 16351 17685 16407
rect 20853 16351 20909 16407
rect 21671 16351 21727 16407
rect 24895 16351 24951 16407
rect 25713 16351 25769 16407
rect 28937 16351 28993 16407
rect 29755 16351 29811 16407
rect 5186 16019 5242 16075
rect 6672 16019 6728 16075
rect 9228 16016 9284 16072
rect 10714 16016 10770 16072
rect 13270 16016 13326 16072
rect 14756 16016 14812 16072
rect 17312 16016 17368 16072
rect 18798 16016 18854 16072
rect 21354 16016 21410 16072
rect 22840 16016 22896 16072
rect 25396 16016 25452 16072
rect 26882 16016 26938 16072
rect 29438 16016 29494 16072
rect 30924 16016 30980 16072
rect 4685 14149 4741 14205
rect 5503 14149 5559 14205
rect 6171 14149 6227 14205
rect 6989 14149 7045 14205
rect 8727 14146 8783 14202
rect 9545 14146 9601 14202
rect 10213 14146 10269 14202
rect 11031 14146 11087 14202
rect 12769 14146 12825 14202
rect 13587 14146 13643 14202
rect 14255 14146 14311 14202
rect 15073 14146 15129 14202
rect 16811 14146 16867 14202
rect 17629 14146 17685 14202
rect 18297 14146 18353 14202
rect 19115 14146 19171 14202
rect 20853 14146 20909 14202
rect 21671 14146 21727 14202
rect 22339 14146 22395 14202
rect 23157 14146 23213 14202
rect 24895 14146 24951 14202
rect 25713 14146 25769 14202
rect 26381 14146 26437 14202
rect 27199 14146 27255 14202
rect 28937 14146 28993 14202
rect 29755 14146 29811 14202
rect 30423 14146 30479 14202
rect 31241 14146 31297 14202
rect 28173 14029 28229 14085
rect 5186 13814 5242 13870
rect 6672 13815 6728 13871
rect 9228 13811 9284 13867
rect 10714 13812 10770 13868
rect 13270 13811 13326 13867
rect 14756 13812 14812 13868
rect 17312 13811 17368 13867
rect 18798 13812 18854 13868
rect 21354 13811 21410 13867
rect 22840 13812 22896 13868
rect 25396 13811 25452 13867
rect 26882 13812 26938 13868
rect 29438 13811 29494 13867
rect 30924 13812 30980 13868
rect 4685 11944 4741 12000
rect 5503 11944 5559 12000
rect 6171 11945 6227 12001
rect 6989 11945 7045 12001
rect 8727 11941 8783 11997
rect 9545 11941 9601 11997
rect 10213 11942 10269 11998
rect 11031 11942 11087 11998
rect 12769 11941 12825 11997
rect 13587 11941 13643 11997
rect 14255 11942 14311 11998
rect 15073 11942 15129 11998
rect 16811 11941 16867 11997
rect 17629 11941 17685 11997
rect 18297 11942 18353 11998
rect 19115 11942 19171 11998
rect 20853 11941 20909 11997
rect 21671 11941 21727 11997
rect 22339 11942 22395 11998
rect 23157 11942 23213 11998
rect 24895 11941 24951 11997
rect 25713 11941 25769 11997
rect 26381 11942 26437 11998
rect 27199 11942 27255 11998
rect 28937 11941 28993 11997
rect 29755 11941 29811 11997
rect 30423 11942 30479 11998
rect 31241 11942 31297 11998
rect 5186 11609 5242 11665
rect 9228 11606 9284 11662
rect 13270 11606 13326 11662
rect 17312 11606 17368 11662
rect 21354 11606 21410 11662
rect 25396 11606 25452 11662
rect 29438 11606 29494 11662
rect 28173 10405 28229 10461
rect 4685 9739 4741 9795
rect 5503 9739 5559 9795
rect 8727 9736 8783 9792
rect 9545 9736 9601 9792
rect 12769 9736 12825 9792
rect 13587 9736 13643 9792
rect 16811 9736 16867 9792
rect 17629 9736 17685 9792
rect 20853 9736 20909 9792
rect 21671 9736 21727 9792
rect 24895 9736 24951 9792
rect 25713 9736 25769 9792
rect 28937 9736 28993 9792
rect 29755 9736 29811 9792
rect 1174 8645 1230 8701
rect 5186 8645 5242 8701
rect 9228 8645 9284 8701
rect 13270 8645 13326 8701
rect 17312 8645 17368 8701
rect 21354 8645 21410 8701
rect 25396 8645 25452 8701
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect 673 6775 729 6831
rect 1491 6775 1547 6831
rect 4685 6775 4741 6831
rect 5503 6775 5559 6831
rect 8727 6775 8783 6831
rect 9545 6775 9601 6831
rect 12769 6775 12825 6831
rect 13587 6775 13643 6831
rect 16811 6775 16867 6831
rect 17629 6775 17685 6831
rect 20853 6775 20909 6831
rect 21671 6775 21727 6831
rect 24895 6775 24951 6831
rect 25713 6775 25769 6831
rect 1174 6440 1230 6496
rect 2660 6440 2716 6496
rect 5186 6440 5242 6496
rect 6672 6440 6728 6496
rect 9228 6440 9284 6496
rect 10714 6440 10770 6496
rect 13270 6440 13326 6496
rect 14756 6440 14812 6496
rect 17312 6440 17368 6496
rect 18798 6440 18854 6496
rect 21354 6440 21410 6496
rect 22840 6440 22896 6496
rect 25396 6440 25452 6496
rect 26882 6440 26938 6496
rect 673 4570 729 4626
rect 1491 4570 1547 4626
rect 2159 4570 2215 4626
rect 2977 4570 3033 4626
rect 4685 4570 4741 4626
rect 5503 4570 5559 4626
rect 6171 4570 6227 4626
rect 6989 4570 7045 4626
rect 8727 4570 8783 4626
rect 9545 4570 9601 4626
rect 10213 4570 10269 4626
rect 11031 4570 11087 4626
rect 12769 4570 12825 4626
rect 13587 4570 13643 4626
rect 14255 4570 14311 4626
rect 15073 4570 15129 4626
rect 16811 4570 16867 4626
rect 17629 4570 17685 4626
rect 18297 4570 18353 4626
rect 19115 4570 19171 4626
rect 20853 4570 20909 4626
rect 21671 4570 21727 4626
rect 22339 4570 22395 4626
rect 23157 4570 23213 4626
rect 24895 4570 24951 4626
rect 25713 4570 25769 4626
rect 26381 4570 26437 4626
rect 27199 4570 27255 4626
rect 1174 4235 1230 4291
rect 2660 4236 2716 4292
rect 5186 4235 5242 4291
rect 6672 4236 6728 4292
rect 9228 4235 9284 4291
rect 10714 4236 10770 4292
rect 13270 4235 13326 4291
rect 14756 4236 14812 4292
rect 17312 4235 17368 4291
rect 18798 4236 18854 4292
rect 21354 4235 21410 4291
rect 22840 4236 22896 4292
rect 25396 4235 25452 4291
rect 26882 4236 26938 4292
rect 673 2365 729 2421
rect 1491 2365 1547 2421
rect 2159 2366 2215 2422
rect 2977 2366 3033 2422
rect 4685 2365 4741 2421
rect 5503 2365 5559 2421
rect 6171 2366 6227 2422
rect 6989 2366 7045 2422
rect 8727 2365 8783 2421
rect 9545 2365 9601 2421
rect 10213 2366 10269 2422
rect 11031 2366 11087 2422
rect 12769 2365 12825 2421
rect 13587 2365 13643 2421
rect 14255 2366 14311 2422
rect 15073 2366 15129 2422
rect 16811 2365 16867 2421
rect 17629 2365 17685 2421
rect 18297 2366 18353 2422
rect 19115 2366 19171 2422
rect 20853 2365 20909 2421
rect 21671 2365 21727 2421
rect 22339 2366 22395 2422
rect 23157 2366 23213 2422
rect 24895 2365 24951 2421
rect 25713 2365 25769 2421
rect 26381 2366 26437 2422
rect 27199 2366 27255 2422
rect 1174 2030 1230 2086
rect 5186 2030 5242 2086
rect 9228 2030 9284 2086
rect 13270 2030 13326 2086
rect 17312 2030 17368 2086
rect 21354 2030 21410 2086
rect 25396 2030 25452 2086
rect -109 829 -53 885
rect 673 160 729 216
rect 1491 160 1547 216
rect 4685 160 4741 216
rect 5503 160 5559 216
rect 8727 160 8783 216
rect 9545 160 9601 216
rect 12769 160 12825 216
rect 13587 160 13643 216
rect 16811 160 16867 216
rect 17629 160 17685 216
rect 20853 160 20909 216
rect 21671 160 21727 216
rect 24895 160 24951 216
rect 25713 160 25769 216
rect -109 42 -53 98
<< metal4 >>
rect 5174 18280 5260 18284
rect 5174 18224 5186 18280
rect 5242 18224 5260 18280
rect 5174 18212 5260 18224
rect 7460 18076 8202 18385
rect 9216 18277 9302 18281
rect 9216 18221 9228 18277
rect 9284 18221 9302 18277
rect 9216 18209 9302 18221
rect 4160 18073 8202 18076
rect 11502 18073 12244 18385
rect 13258 18277 13344 18281
rect 13258 18221 13270 18277
rect 13326 18221 13344 18277
rect 13258 18209 13344 18221
rect 15544 18073 16286 18385
rect 17300 18277 17386 18281
rect 17300 18221 17312 18277
rect 17368 18221 17386 18277
rect 17300 18209 17386 18221
rect 19586 18073 20328 18385
rect 21342 18277 21428 18281
rect 21342 18221 21354 18277
rect 21410 18221 21428 18277
rect 21342 18209 21428 18221
rect 23628 18073 24370 18385
rect 25384 18277 25470 18281
rect 25384 18221 25396 18277
rect 25452 18221 25470 18277
rect 25384 18209 25470 18221
rect 27670 18073 28412 18385
rect 29426 18277 29512 18281
rect 29426 18221 29438 18277
rect 29494 18221 29512 18277
rect 29426 18209 29512 18221
rect 4160 16410 31712 18073
rect 4160 16354 4685 16410
rect 4741 16354 5503 16410
rect 5559 16407 31712 16410
rect 5559 16354 8727 16407
rect 4160 16351 8727 16354
rect 8783 16351 9545 16407
rect 9601 16351 12769 16407
rect 12825 16351 13587 16407
rect 13643 16351 16811 16407
rect 16867 16351 17629 16407
rect 17685 16351 20853 16407
rect 20909 16351 21671 16407
rect 21727 16351 24895 16407
rect 24951 16351 25713 16407
rect 25769 16351 28937 16407
rect 28993 16351 29755 16407
rect 29811 16351 31712 16407
rect 4160 16236 31712 16351
rect 4160 15871 4992 16236
rect 5174 16075 5260 16079
rect 5174 16019 5186 16075
rect 5242 16019 5260 16075
rect 5174 16007 5260 16019
rect 5442 15871 6478 16236
rect 6928 16233 31712 16236
rect 6660 16075 6746 16079
rect 6660 16019 6672 16075
rect 6728 16019 6746 16075
rect 6660 16007 6746 16019
rect 6928 15871 9034 16233
rect 9216 16072 9302 16076
rect 9216 16016 9228 16072
rect 9284 16016 9302 16072
rect 9216 16004 9302 16016
rect 4160 15868 9034 15871
rect 9484 15868 10520 16233
rect 10702 16072 10788 16076
rect 10702 16016 10714 16072
rect 10770 16016 10788 16072
rect 10702 16004 10788 16016
rect 10970 15868 13076 16233
rect 13258 16072 13344 16076
rect 13258 16016 13270 16072
rect 13326 16016 13344 16072
rect 13258 16004 13344 16016
rect 13526 15868 14562 16233
rect 14744 16072 14830 16076
rect 14744 16016 14756 16072
rect 14812 16016 14830 16072
rect 14744 16004 14830 16016
rect 15012 15868 17118 16233
rect 17300 16072 17386 16076
rect 17300 16016 17312 16072
rect 17368 16016 17386 16072
rect 17300 16004 17386 16016
rect 17568 15868 18604 16233
rect 18786 16072 18872 16076
rect 18786 16016 18798 16072
rect 18854 16016 18872 16072
rect 18786 16004 18872 16016
rect 19054 15868 21160 16233
rect 21342 16072 21428 16076
rect 21342 16016 21354 16072
rect 21410 16016 21428 16072
rect 21342 16004 21428 16016
rect 21610 15868 22646 16233
rect 22828 16072 22914 16076
rect 22828 16016 22840 16072
rect 22896 16016 22914 16072
rect 22828 16004 22914 16016
rect 23096 15868 25202 16233
rect 25384 16072 25470 16076
rect 25384 16016 25396 16072
rect 25452 16016 25470 16072
rect 25384 16004 25470 16016
rect 25652 15868 26688 16233
rect 26870 16072 26956 16076
rect 26870 16016 26882 16072
rect 26938 16016 26956 16072
rect 26870 16004 26956 16016
rect 27138 15868 29244 16233
rect 29426 16072 29512 16076
rect 29426 16016 29438 16072
rect 29494 16016 29512 16072
rect 29426 16004 29512 16016
rect 29694 15868 30730 16233
rect 30912 16072 30998 16076
rect 30912 16016 30924 16072
rect 30980 16016 30998 16072
rect 30912 16004 30998 16016
rect 31180 15868 31712 16233
rect 4160 14205 31712 15868
rect 4160 14149 4685 14205
rect 4741 14149 5503 14205
rect 5559 14149 6171 14205
rect 6227 14149 6989 14205
rect 7045 14202 31712 14205
rect 7045 14149 8727 14202
rect 4160 14146 8727 14149
rect 8783 14146 9545 14202
rect 9601 14146 10213 14202
rect 10269 14146 11031 14202
rect 11087 14146 12769 14202
rect 12825 14146 13587 14202
rect 13643 14146 14255 14202
rect 14311 14146 15073 14202
rect 15129 14146 16811 14202
rect 16867 14146 17629 14202
rect 17685 14146 18297 14202
rect 18353 14146 19115 14202
rect 19171 14146 20853 14202
rect 20909 14146 21671 14202
rect 21727 14146 22339 14202
rect 22395 14146 23157 14202
rect 23213 14146 24895 14202
rect 24951 14146 25713 14202
rect 25769 14146 26381 14202
rect 26437 14146 27199 14202
rect 27255 14146 28937 14202
rect 28993 14146 29755 14202
rect 29811 14146 30423 14202
rect 30479 14146 31241 14202
rect 31297 14146 31712 14202
rect 4160 14085 31712 14146
rect 4160 14031 28173 14085
rect 4160 13666 4992 14031
rect 5174 13870 5260 13874
rect 5174 13814 5186 13870
rect 5242 13814 5260 13870
rect 5174 13802 5260 13814
rect 5442 13666 6478 14031
rect 6928 14029 28173 14031
rect 28229 14029 31712 14085
rect 6928 14028 31712 14029
rect 6660 13871 6746 13875
rect 6660 13815 6672 13871
rect 6728 13815 6746 13871
rect 6660 13803 6746 13815
rect 6928 13666 9034 14028
rect 9216 13867 9302 13871
rect 9216 13811 9228 13867
rect 9284 13811 9302 13867
rect 9216 13799 9302 13811
rect 4160 13663 9034 13666
rect 9484 13663 10520 14028
rect 10702 13868 10788 13872
rect 10702 13812 10714 13868
rect 10770 13812 10788 13868
rect 10702 13800 10788 13812
rect 10970 13663 13076 14028
rect 13258 13867 13344 13871
rect 13258 13811 13270 13867
rect 13326 13811 13344 13867
rect 13258 13799 13344 13811
rect 13526 13663 14562 14028
rect 14744 13868 14830 13872
rect 14744 13812 14756 13868
rect 14812 13812 14830 13868
rect 14744 13800 14830 13812
rect 15012 13663 17118 14028
rect 17300 13867 17386 13871
rect 17300 13811 17312 13867
rect 17368 13811 17386 13867
rect 17300 13799 17386 13811
rect 17568 13663 18604 14028
rect 18786 13868 18872 13872
rect 18786 13812 18798 13868
rect 18854 13812 18872 13868
rect 18786 13800 18872 13812
rect 19054 13663 21160 14028
rect 21342 13867 21428 13871
rect 21342 13811 21354 13867
rect 21410 13811 21428 13867
rect 21342 13799 21428 13811
rect 21610 13663 22646 14028
rect 22828 13868 22914 13872
rect 22828 13812 22840 13868
rect 22896 13812 22914 13868
rect 22828 13800 22914 13812
rect 23096 13663 25202 14028
rect 25384 13867 25470 13871
rect 25384 13811 25396 13867
rect 25452 13811 25470 13867
rect 25384 13799 25470 13811
rect 25652 13663 26688 14028
rect 26870 13868 26956 13872
rect 26870 13812 26882 13868
rect 26938 13812 26956 13868
rect 26870 13800 26956 13812
rect 27138 13663 29244 14028
rect 29426 13867 29512 13871
rect 29426 13811 29438 13867
rect 29494 13811 29512 13867
rect 29426 13799 29512 13811
rect 29694 13663 30730 14028
rect 30912 13868 30998 13872
rect 30912 13812 30924 13868
rect 30980 13812 30998 13868
rect 30912 13800 30998 13812
rect 31180 13663 31712 14028
rect 4160 12001 31712 13663
rect 4160 12000 6171 12001
rect 4160 11944 4685 12000
rect 4741 11944 5503 12000
rect 5559 11945 6171 12000
rect 6227 11945 6989 12001
rect 7045 11998 31712 12001
rect 7045 11997 10213 11998
rect 7045 11945 8727 11997
rect 5559 11944 8727 11945
rect 4160 11941 8727 11944
rect 8783 11941 9545 11997
rect 9601 11942 10213 11997
rect 10269 11942 11031 11998
rect 11087 11997 14255 11998
rect 11087 11942 12769 11997
rect 9601 11941 12769 11942
rect 12825 11941 13587 11997
rect 13643 11942 14255 11997
rect 14311 11942 15073 11998
rect 15129 11997 18297 11998
rect 15129 11942 16811 11997
rect 13643 11941 16811 11942
rect 16867 11941 17629 11997
rect 17685 11942 18297 11997
rect 18353 11942 19115 11998
rect 19171 11997 22339 11998
rect 19171 11942 20853 11997
rect 17685 11941 20853 11942
rect 20909 11941 21671 11997
rect 21727 11942 22339 11997
rect 22395 11942 23157 11998
rect 23213 11997 26381 11998
rect 23213 11942 24895 11997
rect 21727 11941 24895 11942
rect 24951 11941 25713 11997
rect 25769 11942 26381 11997
rect 26437 11942 27199 11998
rect 27255 11997 30423 11998
rect 27255 11942 28937 11997
rect 25769 11941 28937 11942
rect 28993 11941 29755 11997
rect 29811 11942 30423 11997
rect 30479 11942 31241 11998
rect 31297 11942 31712 11998
rect 29811 11941 31712 11942
rect 4160 11826 31712 11941
rect 4160 11461 4992 11826
rect 5442 11823 31712 11826
rect 5174 11665 5260 11669
rect 5174 11609 5186 11665
rect 5242 11609 5260 11665
rect 5174 11597 5260 11609
rect 5442 11461 9034 11823
rect 9216 11662 9302 11666
rect 9216 11606 9228 11662
rect 9284 11606 9302 11662
rect 9216 11594 9302 11606
rect 4160 11458 9034 11461
rect 9484 11458 13076 11823
rect 13258 11662 13344 11666
rect 13258 11606 13270 11662
rect 13326 11606 13344 11662
rect 13258 11594 13344 11606
rect 13526 11458 17118 11823
rect 17300 11662 17386 11666
rect 17300 11606 17312 11662
rect 17368 11606 17386 11662
rect 17300 11594 17386 11606
rect 17568 11458 21160 11823
rect 21342 11662 21428 11666
rect 21342 11606 21354 11662
rect 21410 11606 21428 11662
rect 21342 11594 21428 11606
rect 21610 11458 25202 11823
rect 25384 11662 25470 11666
rect 25384 11606 25396 11662
rect 25452 11606 25470 11662
rect 25384 11594 25470 11606
rect 25652 11458 29244 11823
rect 29426 11662 29512 11666
rect 29426 11606 29438 11662
rect 29494 11606 29512 11662
rect 29426 11594 29512 11606
rect 29694 11458 31712 11823
rect 4160 10461 31712 11458
rect 4160 10405 28173 10461
rect 28229 10405 31712 10461
rect 4160 9795 31712 10405
rect 4160 9739 4685 9795
rect 4741 9739 5503 9795
rect 5559 9792 31712 9795
rect 5559 9739 8727 9792
rect 4160 9736 8727 9739
rect 8783 9736 9545 9792
rect 9601 9736 12769 9792
rect 12825 9736 13587 9792
rect 13643 9736 16811 9792
rect 16867 9736 17629 9792
rect 17685 9736 20853 9792
rect 20909 9736 21671 9792
rect 21727 9736 24895 9792
rect 24951 9736 25713 9792
rect 25769 9736 28937 9792
rect 28993 9736 29755 9792
rect 29811 9736 31712 9792
rect 4160 9609 31712 9736
rect 4100 9606 31712 9609
rect 4100 8809 27730 9606
rect 1162 8701 1248 8705
rect 1162 8645 1174 8701
rect 1230 8645 1248 8701
rect 1162 8633 1248 8645
rect 3448 8497 4160 8809
rect 5174 8701 5260 8705
rect 5174 8645 5186 8701
rect 5242 8645 5260 8701
rect 5174 8633 5260 8645
rect 7460 8497 8202 8809
rect 9216 8701 9302 8705
rect 9216 8645 9228 8701
rect 9284 8645 9302 8701
rect 9216 8633 9302 8645
rect 11502 8497 12244 8809
rect 13258 8701 13344 8705
rect 13258 8645 13270 8701
rect 13326 8645 13344 8701
rect 13258 8633 13344 8645
rect 15544 8497 16286 8809
rect 17300 8701 17386 8705
rect 17300 8645 17312 8701
rect 17368 8645 17386 8701
rect 17300 8633 17386 8645
rect 19586 8497 20328 8809
rect 21342 8701 21428 8705
rect 21342 8645 21354 8701
rect 21410 8645 21428 8701
rect 21342 8633 21428 8645
rect 23628 8497 24370 8809
rect 25384 8701 25470 8705
rect 25384 8645 25396 8701
rect 25452 8645 25470 8701
rect 25384 8633 25470 8645
rect 148 7824 27670 8497
rect 148 7584 3930 7824
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 4160 7584 7972 7824
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 8202 7584 12014 7824
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 12244 7584 16056 7824
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 16286 7584 20098 7824
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 20328 7584 24140 7824
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 24370 7584 27670 7824
rect 148 6831 27670 7584
rect 148 6775 673 6831
rect 729 6775 1491 6831
rect 1547 6775 4685 6831
rect 4741 6775 5503 6831
rect 5559 6775 8727 6831
rect 8783 6775 9545 6831
rect 9601 6775 12769 6831
rect 12825 6775 13587 6831
rect 13643 6775 16811 6831
rect 16867 6775 17629 6831
rect 17685 6775 20853 6831
rect 20909 6775 21671 6831
rect 21727 6775 24895 6831
rect 24951 6775 25713 6831
rect 25769 6775 27670 6831
rect 148 6657 27670 6775
rect 148 6292 980 6657
rect 1162 6496 1248 6500
rect 1162 6440 1174 6496
rect 1230 6440 1248 6496
rect 1162 6428 1248 6440
rect 1430 6292 2466 6657
rect 2648 6496 2734 6500
rect 2648 6440 2660 6496
rect 2716 6440 2734 6496
rect 2648 6428 2734 6440
rect 2916 6292 4992 6657
rect 5174 6496 5260 6500
rect 5174 6440 5186 6496
rect 5242 6440 5260 6496
rect 5174 6428 5260 6440
rect 5442 6292 6478 6657
rect 6660 6496 6746 6500
rect 6660 6440 6672 6496
rect 6728 6440 6746 6496
rect 6660 6428 6746 6440
rect 6928 6292 9034 6657
rect 9216 6496 9302 6500
rect 9216 6440 9228 6496
rect 9284 6440 9302 6496
rect 9216 6428 9302 6440
rect 9484 6292 10520 6657
rect 10702 6496 10788 6500
rect 10702 6440 10714 6496
rect 10770 6440 10788 6496
rect 10702 6428 10788 6440
rect 10970 6292 13076 6657
rect 13258 6496 13344 6500
rect 13258 6440 13270 6496
rect 13326 6440 13344 6496
rect 13258 6428 13344 6440
rect 13526 6292 14562 6657
rect 14744 6496 14830 6500
rect 14744 6440 14756 6496
rect 14812 6440 14830 6496
rect 14744 6428 14830 6440
rect 15012 6292 17118 6657
rect 17300 6496 17386 6500
rect 17300 6440 17312 6496
rect 17368 6440 17386 6496
rect 17300 6428 17386 6440
rect 17568 6292 18604 6657
rect 18786 6496 18872 6500
rect 18786 6440 18798 6496
rect 18854 6440 18872 6496
rect 18786 6428 18872 6440
rect 19054 6292 21160 6657
rect 21342 6496 21428 6500
rect 21342 6440 21354 6496
rect 21410 6440 21428 6496
rect 21342 6428 21428 6440
rect 21610 6292 22646 6657
rect 22828 6496 22914 6500
rect 22828 6440 22840 6496
rect 22896 6440 22914 6496
rect 22828 6428 22914 6440
rect 23096 6292 25202 6657
rect 25384 6496 25470 6500
rect 25384 6440 25396 6496
rect 25452 6440 25470 6496
rect 25384 6428 25470 6440
rect 25652 6292 26688 6657
rect 26870 6496 26956 6500
rect 26870 6440 26882 6496
rect 26938 6440 26956 6496
rect 26870 6428 26956 6440
rect 27138 6292 27670 6657
rect 148 4626 27670 6292
rect 148 4570 673 4626
rect 729 4570 1491 4626
rect 1547 4570 2159 4626
rect 2215 4570 2977 4626
rect 3033 4570 4685 4626
rect 4741 4570 5503 4626
rect 5559 4570 6171 4626
rect 6227 4570 6989 4626
rect 7045 4570 8727 4626
rect 8783 4570 9545 4626
rect 9601 4570 10213 4626
rect 10269 4570 11031 4626
rect 11087 4570 12769 4626
rect 12825 4570 13587 4626
rect 13643 4570 14255 4626
rect 14311 4570 15073 4626
rect 15129 4570 16811 4626
rect 16867 4570 17629 4626
rect 17685 4570 18297 4626
rect 18353 4570 19115 4626
rect 19171 4570 20853 4626
rect 20909 4570 21671 4626
rect 21727 4570 22339 4626
rect 22395 4570 23157 4626
rect 23213 4570 24895 4626
rect 24951 4570 25713 4626
rect 25769 4570 26381 4626
rect 26437 4570 27199 4626
rect 27255 4570 27670 4626
rect 148 4452 27670 4570
rect 148 4087 980 4452
rect 1162 4291 1248 4295
rect 1162 4235 1174 4291
rect 1230 4235 1248 4291
rect 1162 4223 1248 4235
rect 1430 4087 2466 4452
rect 2648 4292 2734 4296
rect 2648 4236 2660 4292
rect 2716 4236 2734 4292
rect 2648 4224 2734 4236
rect 2916 4087 4992 4452
rect 5174 4291 5260 4295
rect 5174 4235 5186 4291
rect 5242 4235 5260 4291
rect 5174 4223 5260 4235
rect 5442 4087 6478 4452
rect 6660 4292 6746 4296
rect 6660 4236 6672 4292
rect 6728 4236 6746 4292
rect 6660 4224 6746 4236
rect 6928 4087 9034 4452
rect 9216 4291 9302 4295
rect 9216 4235 9228 4291
rect 9284 4235 9302 4291
rect 9216 4223 9302 4235
rect 9484 4087 10520 4452
rect 10702 4292 10788 4296
rect 10702 4236 10714 4292
rect 10770 4236 10788 4292
rect 10702 4224 10788 4236
rect 10970 4087 13076 4452
rect 13258 4291 13344 4295
rect 13258 4235 13270 4291
rect 13326 4235 13344 4291
rect 13258 4223 13344 4235
rect 13526 4087 14562 4452
rect 14744 4292 14830 4296
rect 14744 4236 14756 4292
rect 14812 4236 14830 4292
rect 14744 4224 14830 4236
rect 15012 4087 17118 4452
rect 17300 4291 17386 4295
rect 17300 4235 17312 4291
rect 17368 4235 17386 4291
rect 17300 4223 17386 4235
rect 17568 4087 18604 4452
rect 18786 4292 18872 4296
rect 18786 4236 18798 4292
rect 18854 4236 18872 4292
rect 18786 4224 18872 4236
rect 19054 4087 21160 4452
rect 21342 4291 21428 4295
rect 21342 4235 21354 4291
rect 21410 4235 21428 4291
rect 21342 4223 21428 4235
rect 21610 4087 22646 4452
rect 22828 4292 22914 4296
rect 22828 4236 22840 4292
rect 22896 4236 22914 4292
rect 22828 4224 22914 4236
rect 23096 4087 25202 4452
rect 25384 4291 25470 4295
rect 25384 4235 25396 4291
rect 25452 4235 25470 4291
rect 25384 4223 25470 4235
rect 25652 4087 26688 4452
rect 26870 4292 26956 4296
rect 26870 4236 26882 4292
rect 26938 4236 26956 4292
rect 26870 4224 26956 4236
rect 27138 4087 27670 4452
rect 148 2422 27670 4087
rect 148 2421 2159 2422
rect 148 2365 673 2421
rect 729 2365 1491 2421
rect 1547 2366 2159 2421
rect 2215 2366 2977 2422
rect 3033 2421 6171 2422
rect 3033 2366 4685 2421
rect 1547 2365 4685 2366
rect 4741 2365 5503 2421
rect 5559 2366 6171 2421
rect 6227 2366 6989 2422
rect 7045 2421 10213 2422
rect 7045 2366 8727 2421
rect 5559 2365 8727 2366
rect 8783 2365 9545 2421
rect 9601 2366 10213 2421
rect 10269 2366 11031 2422
rect 11087 2421 14255 2422
rect 11087 2366 12769 2421
rect 9601 2365 12769 2366
rect 12825 2365 13587 2421
rect 13643 2366 14255 2421
rect 14311 2366 15073 2422
rect 15129 2421 18297 2422
rect 15129 2366 16811 2421
rect 13643 2365 16811 2366
rect 16867 2365 17629 2421
rect 17685 2366 18297 2421
rect 18353 2366 19115 2422
rect 19171 2421 22339 2422
rect 19171 2366 20853 2421
rect 17685 2365 20853 2366
rect 20909 2365 21671 2421
rect 21727 2366 22339 2421
rect 22395 2366 23157 2422
rect 23213 2421 26381 2422
rect 23213 2366 24895 2421
rect 21727 2365 24895 2366
rect 24951 2365 25713 2421
rect 25769 2366 26381 2421
rect 26437 2366 27199 2422
rect 27255 2366 27670 2422
rect 25769 2365 27670 2366
rect 148 2247 27670 2365
rect 148 1882 980 2247
rect 1162 2086 1248 2090
rect 1162 2030 1174 2086
rect 1230 2030 1248 2086
rect 1162 2018 1248 2030
rect 1430 1882 4992 2247
rect 5174 2086 5260 2090
rect 5174 2030 5186 2086
rect 5242 2030 5260 2086
rect 5174 2018 5260 2030
rect 5442 1882 9034 2247
rect 9216 2086 9302 2090
rect 9216 2030 9228 2086
rect 9284 2030 9302 2086
rect 9216 2018 9302 2030
rect 9484 1882 13076 2247
rect 13258 2086 13344 2090
rect 13258 2030 13270 2086
rect 13326 2030 13344 2086
rect 13258 2018 13344 2030
rect 13526 1882 17118 2247
rect 17300 2086 17386 2090
rect 17300 2030 17312 2086
rect 17368 2030 17386 2086
rect 17300 2018 17386 2030
rect 17568 1882 21160 2247
rect 21342 2086 21428 2090
rect 21342 2030 21354 2086
rect 21410 2030 21428 2086
rect 21342 2018 21428 2030
rect 21610 1882 25202 2247
rect 25384 2086 25470 2090
rect 25384 2030 25396 2086
rect 25452 2030 25470 2086
rect 25384 2018 25470 2030
rect 25652 1882 27670 2247
rect 148 897 27670 1882
rect -121 885 27670 897
rect -121 829 -109 885
rect -53 829 27670 885
rect -121 737 27670 829
rect 148 216 27670 737
rect 148 160 673 216
rect 729 160 1491 216
rect 1547 160 4685 216
rect 4741 160 5503 216
rect 5559 160 8727 216
rect 8783 160 9545 216
rect 9601 160 12769 216
rect 12825 160 13587 216
rect 13643 160 16811 216
rect 16867 160 17629 216
rect 17685 160 20853 216
rect 20909 160 21671 216
rect 21727 160 24895 216
rect 24951 160 25713 216
rect 25769 160 27670 216
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect 148 30 27670 160
<< via4 >>
rect 5186 18224 5242 18280
rect 9228 18221 9284 18277
rect 13270 18221 13326 18277
rect 17312 18221 17368 18277
rect 21354 18221 21410 18277
rect 25396 18221 25452 18277
rect 29438 18221 29494 18277
rect 5186 16019 5242 16075
rect 6672 16019 6728 16075
rect 9228 16016 9284 16072
rect 10714 16016 10770 16072
rect 13270 16016 13326 16072
rect 14756 16016 14812 16072
rect 17312 16016 17368 16072
rect 18798 16016 18854 16072
rect 21354 16016 21410 16072
rect 22840 16016 22896 16072
rect 25396 16016 25452 16072
rect 26882 16016 26938 16072
rect 29438 16016 29494 16072
rect 30924 16016 30980 16072
rect 5186 13814 5242 13870
rect 6672 13815 6728 13871
rect 9228 13811 9284 13867
rect 10714 13812 10770 13868
rect 13270 13811 13326 13867
rect 14756 13812 14812 13868
rect 17312 13811 17368 13867
rect 18798 13812 18854 13868
rect 21354 13811 21410 13867
rect 22840 13812 22896 13868
rect 25396 13811 25452 13867
rect 26882 13812 26938 13868
rect 29438 13811 29494 13867
rect 30924 13812 30980 13868
rect 5186 11609 5242 11665
rect 9228 11606 9284 11662
rect 13270 11606 13326 11662
rect 17312 11606 17368 11662
rect 21354 11606 21410 11662
rect 25396 11606 25452 11662
rect 29438 11606 29494 11662
rect 1174 8645 1230 8701
rect 5186 8645 5242 8701
rect 9228 8645 9284 8701
rect 13270 8645 13326 8701
rect 17312 8645 17368 8701
rect 21354 8645 21410 8701
rect 25396 8645 25452 8701
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect 1174 6440 1230 6496
rect 2660 6440 2716 6496
rect 5186 6440 5242 6496
rect 6672 6440 6728 6496
rect 9228 6440 9284 6496
rect 10714 6440 10770 6496
rect 13270 6440 13326 6496
rect 14756 6440 14812 6496
rect 17312 6440 17368 6496
rect 18798 6440 18854 6496
rect 21354 6440 21410 6496
rect 22840 6440 22896 6496
rect 25396 6440 25452 6496
rect 26882 6440 26938 6496
rect 1174 4235 1230 4291
rect 2660 4236 2716 4292
rect 5186 4235 5242 4291
rect 6672 4236 6728 4292
rect 9228 4235 9284 4291
rect 10714 4236 10770 4292
rect 13270 4235 13326 4291
rect 14756 4236 14812 4292
rect 17312 4235 17368 4291
rect 18798 4236 18854 4292
rect 21354 4235 21410 4291
rect 22840 4236 22896 4292
rect 25396 4235 25452 4291
rect 26882 4236 26938 4292
rect 1174 2030 1230 2086
rect 5186 2030 5242 2086
rect 9228 2030 9284 2086
rect 13270 2030 13326 2086
rect 17312 2030 17368 2086
rect 21354 2030 21410 2086
rect 25396 2030 25452 2086
rect -109 42 -53 98
<< metal5 >>
rect 4160 18385 7460 18388
rect 4160 18280 31712 18385
rect 4160 18224 5186 18280
rect 5242 18277 31712 18280
rect 5242 18224 9228 18277
rect 4160 18221 9228 18224
rect 9284 18221 13270 18277
rect 13326 18221 17312 18277
rect 17368 18221 21354 18277
rect 21410 18221 25396 18277
rect 25452 18221 29438 18277
rect 29494 18221 31712 18277
rect 4160 16075 31712 18221
rect 4160 16019 5186 16075
rect 5242 16019 6672 16075
rect 6728 16072 31712 16075
rect 6728 16019 9228 16072
rect 4160 16016 9228 16019
rect 9284 16016 10714 16072
rect 10770 16016 13270 16072
rect 13326 16016 14756 16072
rect 14812 16016 17312 16072
rect 17368 16016 18798 16072
rect 18854 16016 21354 16072
rect 21410 16016 22840 16072
rect 22896 16016 25396 16072
rect 25452 16016 26882 16072
rect 26938 16016 29438 16072
rect 29494 16016 30924 16072
rect 30980 16016 31712 16072
rect 4160 14177 31712 16016
rect 4160 13937 28082 14177
rect 28320 13937 31712 14177
rect 4160 13871 31712 13937
rect 4160 13870 6672 13871
rect 4160 13814 5186 13870
rect 5242 13815 6672 13870
rect 6728 13868 31712 13871
rect 6728 13867 10714 13868
rect 6728 13815 9228 13867
rect 5242 13814 9228 13815
rect 4160 13811 9228 13814
rect 9284 13812 10714 13867
rect 10770 13867 14756 13868
rect 10770 13812 13270 13867
rect 9284 13811 13270 13812
rect 13326 13812 14756 13867
rect 14812 13867 18798 13868
rect 14812 13812 17312 13867
rect 13326 13811 17312 13812
rect 17368 13812 18798 13867
rect 18854 13867 22840 13868
rect 18854 13812 21354 13867
rect 17368 13811 21354 13812
rect 21410 13812 22840 13867
rect 22896 13867 26882 13868
rect 22896 13812 25396 13867
rect 21410 13811 25396 13812
rect 25452 13812 26882 13867
rect 26938 13867 30924 13868
rect 26938 13812 29438 13867
rect 25452 13811 29438 13812
rect 29494 13812 30924 13867
rect 30980 13812 31712 13868
rect 29494 13811 31712 13812
rect 4160 11665 31712 13811
rect 4160 11609 5186 11665
rect 5242 11662 31712 11665
rect 5242 11609 9228 11662
rect 4160 11606 9228 11609
rect 9284 11606 13270 11662
rect 13326 11606 17312 11662
rect 17368 11606 21354 11662
rect 21410 11606 25396 11662
rect 25452 11606 29438 11662
rect 29494 11606 31712 11662
rect 4160 10553 31712 11606
rect 4160 10313 28080 10553
rect 28322 10313 31712 10553
rect 4160 9609 31712 10313
rect 4100 9606 31712 9609
rect 4100 8809 27730 9606
rect 148 8701 27670 8809
rect 148 8645 1174 8701
rect 1230 8645 5186 8701
rect 5242 8645 9228 8701
rect 9284 8645 13270 8701
rect 13326 8645 17312 8701
rect 17368 8645 21354 8701
rect 21410 8645 25396 8701
rect 25452 8645 27670 8701
rect 148 7732 27670 8645
rect 148 7676 4022 7732
rect 4078 7676 8064 7732
rect 8120 7676 12106 7732
rect 12162 7676 16148 7732
rect 16204 7676 20190 7732
rect 20246 7676 24232 7732
rect 24288 7676 27670 7732
rect 148 6496 27670 7676
rect 148 6440 1174 6496
rect 1230 6440 2660 6496
rect 2716 6440 5186 6496
rect 5242 6440 6672 6496
rect 6728 6440 9228 6496
rect 9284 6440 10714 6496
rect 10770 6440 13270 6496
rect 13326 6440 14756 6496
rect 14812 6440 17312 6496
rect 17368 6440 18798 6496
rect 18854 6440 21354 6496
rect 21410 6440 22840 6496
rect 22896 6440 25396 6496
rect 25452 6440 26882 6496
rect 26938 6440 27670 6496
rect 148 4292 27670 6440
rect 148 4291 2660 4292
rect 148 4235 1174 4291
rect 1230 4236 2660 4291
rect 2716 4291 6672 4292
rect 2716 4236 5186 4291
rect 1230 4235 5186 4236
rect 5242 4236 6672 4291
rect 6728 4291 10714 4292
rect 6728 4236 9228 4291
rect 5242 4235 9228 4236
rect 9284 4236 10714 4291
rect 10770 4291 14756 4292
rect 10770 4236 13270 4291
rect 9284 4235 13270 4236
rect 13326 4236 14756 4291
rect 14812 4291 18798 4292
rect 14812 4236 17312 4291
rect 13326 4235 17312 4236
rect 17368 4236 18798 4291
rect 18854 4291 22840 4292
rect 18854 4236 21354 4291
rect 17368 4235 21354 4236
rect 21410 4236 22840 4291
rect 22896 4291 26882 4292
rect 22896 4236 25396 4291
rect 21410 4235 25396 4236
rect 25452 4236 26882 4291
rect 26938 4236 27670 4292
rect 25452 4235 27670 4236
rect 148 2086 27670 4235
rect 148 2030 1174 2086
rect 1230 2030 5186 2086
rect 5242 2030 9228 2086
rect 9284 2030 13270 2086
rect 13326 2030 17312 2086
rect 17368 2030 21354 2086
rect 21410 2030 25396 2086
rect 25452 2030 27670 2086
rect 148 190 27670 2030
rect -121 98 27670 190
rect -121 42 -109 98
rect -53 42 27670 98
rect -121 30 27670 42
<< labels >>
rlabel metal2 -473 -113 -473 -113 7 clk
port 2 w
rlabel metal2 -201 8954 -201 8954 7 reset
port 3 w
rlabel metal2 -201 9462 -201 9462 7 comp_in
port 4 w
rlabel metal2 7734 19504 7734 19504 1 d5
port 5 n
rlabel metal2 11789 19501 11789 19501 1 d4
port 6 n
rlabel metal2 15885 19501 15885 19501 1 d3
port 7 n
rlabel metal2 19926 19501 19926 19501 1 d2
port 8 n
rlabel metal2 23968 19504 23968 19504 1 d1
port 9 n
rlabel metal2 28012 19501 28012 19501 1 d0
port 10 n
rlabel metal5 19630 18385 19630 18385 1 vdd
port 0 n
rlabel metal4 15578 30 15578 30 5 vss
port 1 s
rlabel metal1 4022 7704 4022 7704 7 dffrs_0.setb
rlabel metal1 4022 4481 4022 4481 7 dffrs_0.clk
rlabel metal1 4022 856 4022 856 7 dffrs_0.d
rlabel metal1 4039 69 4039 69 7 dffrs_0.resetb
rlabel metal2 7490 5383 7490 5383 3 dffrs_0.Q
rlabel metal2 7490 3178 7490 3178 3 dffrs_0.Qb
rlabel metal5 6130 8809 6130 8809 1 dffrs_0.vdd
rlabel metal4 6238 30 6238 30 5 dffrs_0.vss
rlabel metal2 5186 2098 5186 2098 1 dffrs_0.nand3_8.VDD
rlabel metal1 5596 972 5596 972 3 dffrs_0.nand3_8.Z
rlabel metal1 4510 854 4510 854 7 dffrs_0.nand3_8.A
rlabel metal1 4510 973 4510 973 7 dffrs_0.nand3_8.B
rlabel metal1 4510 1089 4510 1089 7 dffrs_0.nand3_8.C
rlabel metal2 5114 148 5114 148 5 dffrs_0.nand3_8.VSS
rlabel metal2 6672 4304 6672 4304 1 dffrs_0.nand3_7.VDD
rlabel metal1 7082 3178 7082 3178 3 dffrs_0.nand3_7.Z
rlabel metal1 5996 3060 5996 3060 7 dffrs_0.nand3_7.A
rlabel metal1 5996 3179 5996 3179 7 dffrs_0.nand3_7.B
rlabel metal1 5996 3295 5996 3295 7 dffrs_0.nand3_7.C
rlabel metal2 6600 2354 6600 2354 5 dffrs_0.nand3_7.VSS
rlabel metal2 5186 4303 5186 4303 1 dffrs_0.nand3_6.VDD
rlabel metal1 5596 3177 5596 3177 3 dffrs_0.nand3_6.Z
rlabel metal1 4510 3059 4510 3059 7 dffrs_0.nand3_6.A
rlabel metal1 4510 3178 4510 3178 7 dffrs_0.nand3_6.B
rlabel metal1 4510 3294 4510 3294 7 dffrs_0.nand3_6.C
rlabel metal2 5114 2353 5114 2353 5 dffrs_0.nand3_6.VSS
rlabel metal2 6672 6508 6672 6508 1 dffrs_0.nand3_2.VDD
rlabel metal1 7082 5382 7082 5382 3 dffrs_0.nand3_2.Z
rlabel metal1 5996 5264 5996 5264 7 dffrs_0.nand3_2.A
rlabel metal1 5996 5383 5996 5383 7 dffrs_0.nand3_2.B
rlabel metal1 5996 5499 5996 5499 7 dffrs_0.nand3_2.C
rlabel metal2 6600 4558 6600 4558 5 dffrs_0.nand3_2.VSS
rlabel metal2 5186 6508 5186 6508 1 dffrs_0.nand3_1.VDD
rlabel metal1 5596 5382 5596 5382 3 dffrs_0.nand3_1.Z
rlabel metal1 4510 5264 4510 5264 7 dffrs_0.nand3_1.A
rlabel metal1 4510 5383 4510 5383 7 dffrs_0.nand3_1.B
rlabel metal1 4510 5499 4510 5499 7 dffrs_0.nand3_1.C
rlabel metal2 5114 4558 5114 4558 5 dffrs_0.nand3_1.VSS
rlabel metal2 5186 8713 5186 8713 1 dffrs_0.nand3_0.VDD
rlabel metal1 5596 7587 5596 7587 3 dffrs_0.nand3_0.Z
rlabel metal1 4510 7469 4510 7469 7 dffrs_0.nand3_0.A
rlabel metal1 4510 7588 4510 7588 7 dffrs_0.nand3_0.B
rlabel metal1 4510 7704 4510 7704 7 dffrs_0.nand3_0.C
rlabel metal2 5114 6763 5114 6763 5 dffrs_0.nand3_0.VSS
rlabel metal1 10 7704 10 7704 7 dffrs_13.setb
rlabel metal1 10 4481 10 4481 7 dffrs_13.clk
rlabel metal1 10 856 10 856 7 dffrs_13.d
rlabel metal1 27 69 27 69 7 dffrs_13.resetb
rlabel metal2 3478 5383 3478 5383 3 dffrs_13.Q
rlabel metal2 3478 3178 3478 3178 3 dffrs_13.Qb
rlabel metal5 2118 8809 2118 8809 1 dffrs_13.vdd
rlabel metal4 2226 30 2226 30 5 dffrs_13.vss
rlabel metal2 1174 2098 1174 2098 1 dffrs_13.nand3_8.VDD
rlabel metal1 1584 972 1584 972 3 dffrs_13.nand3_8.Z
rlabel metal1 498 854 498 854 7 dffrs_13.nand3_8.A
rlabel metal1 498 973 498 973 7 dffrs_13.nand3_8.B
rlabel metal1 498 1089 498 1089 7 dffrs_13.nand3_8.C
rlabel metal2 1102 148 1102 148 5 dffrs_13.nand3_8.VSS
rlabel metal2 2660 4304 2660 4304 1 dffrs_13.nand3_7.VDD
rlabel metal1 3070 3178 3070 3178 3 dffrs_13.nand3_7.Z
rlabel metal1 1984 3060 1984 3060 7 dffrs_13.nand3_7.A
rlabel metal1 1984 3179 1984 3179 7 dffrs_13.nand3_7.B
rlabel metal1 1984 3295 1984 3295 7 dffrs_13.nand3_7.C
rlabel metal2 2588 2354 2588 2354 5 dffrs_13.nand3_7.VSS
rlabel metal2 1174 4303 1174 4303 1 dffrs_13.nand3_6.VDD
rlabel metal1 1584 3177 1584 3177 3 dffrs_13.nand3_6.Z
rlabel metal1 498 3059 498 3059 7 dffrs_13.nand3_6.A
rlabel metal1 498 3178 498 3178 7 dffrs_13.nand3_6.B
rlabel metal1 498 3294 498 3294 7 dffrs_13.nand3_6.C
rlabel metal2 1102 2353 1102 2353 5 dffrs_13.nand3_6.VSS
rlabel metal2 2660 6508 2660 6508 1 dffrs_13.nand3_2.VDD
rlabel metal1 3070 5382 3070 5382 3 dffrs_13.nand3_2.Z
rlabel metal1 1984 5264 1984 5264 7 dffrs_13.nand3_2.A
rlabel metal1 1984 5383 1984 5383 7 dffrs_13.nand3_2.B
rlabel metal1 1984 5499 1984 5499 7 dffrs_13.nand3_2.C
rlabel metal2 2588 4558 2588 4558 5 dffrs_13.nand3_2.VSS
rlabel metal2 1174 6508 1174 6508 1 dffrs_13.nand3_1.VDD
rlabel metal1 1584 5382 1584 5382 3 dffrs_13.nand3_1.Z
rlabel metal1 498 5264 498 5264 7 dffrs_13.nand3_1.A
rlabel metal1 498 5383 498 5383 7 dffrs_13.nand3_1.B
rlabel metal1 498 5499 498 5499 7 dffrs_13.nand3_1.C
rlabel metal2 1102 4558 1102 4558 5 dffrs_13.nand3_1.VSS
rlabel metal2 1174 8713 1174 8713 1 dffrs_13.nand3_0.VDD
rlabel metal1 1584 7587 1584 7587 3 dffrs_13.nand3_0.Z
rlabel metal1 498 7469 498 7469 7 dffrs_13.nand3_0.A
rlabel metal1 498 7588 498 7588 7 dffrs_13.nand3_0.B
rlabel metal1 498 7704 498 7704 7 dffrs_13.nand3_0.C
rlabel metal2 1102 6763 1102 6763 5 dffrs_13.nand3_0.VSS
rlabel metal1 12106 7704 12106 7704 7 dffrs_2.setb
rlabel metal1 12106 4481 12106 4481 7 dffrs_2.clk
rlabel metal1 12106 856 12106 856 7 dffrs_2.d
rlabel metal1 12123 69 12123 69 7 dffrs_2.resetb
rlabel metal2 15574 5383 15574 5383 3 dffrs_2.Q
rlabel metal2 15574 3178 15574 3178 3 dffrs_2.Qb
rlabel metal5 14214 8809 14214 8809 1 dffrs_2.vdd
rlabel metal4 14322 30 14322 30 5 dffrs_2.vss
rlabel metal2 13270 2098 13270 2098 1 dffrs_2.nand3_8.VDD
rlabel metal1 13680 972 13680 972 3 dffrs_2.nand3_8.Z
rlabel metal1 12594 854 12594 854 7 dffrs_2.nand3_8.A
rlabel metal1 12594 973 12594 973 7 dffrs_2.nand3_8.B
rlabel metal1 12594 1089 12594 1089 7 dffrs_2.nand3_8.C
rlabel metal2 13198 148 13198 148 5 dffrs_2.nand3_8.VSS
rlabel metal2 14756 4304 14756 4304 1 dffrs_2.nand3_7.VDD
rlabel metal1 15166 3178 15166 3178 3 dffrs_2.nand3_7.Z
rlabel metal1 14080 3060 14080 3060 7 dffrs_2.nand3_7.A
rlabel metal1 14080 3179 14080 3179 7 dffrs_2.nand3_7.B
rlabel metal1 14080 3295 14080 3295 7 dffrs_2.nand3_7.C
rlabel metal2 14684 2354 14684 2354 5 dffrs_2.nand3_7.VSS
rlabel metal2 13270 4303 13270 4303 1 dffrs_2.nand3_6.VDD
rlabel metal1 13680 3177 13680 3177 3 dffrs_2.nand3_6.Z
rlabel metal1 12594 3059 12594 3059 7 dffrs_2.nand3_6.A
rlabel metal1 12594 3178 12594 3178 7 dffrs_2.nand3_6.B
rlabel metal1 12594 3294 12594 3294 7 dffrs_2.nand3_6.C
rlabel metal2 13198 2353 13198 2353 5 dffrs_2.nand3_6.VSS
rlabel metal2 14756 6508 14756 6508 1 dffrs_2.nand3_2.VDD
rlabel metal1 15166 5382 15166 5382 3 dffrs_2.nand3_2.Z
rlabel metal1 14080 5264 14080 5264 7 dffrs_2.nand3_2.A
rlabel metal1 14080 5383 14080 5383 7 dffrs_2.nand3_2.B
rlabel metal1 14080 5499 14080 5499 7 dffrs_2.nand3_2.C
rlabel metal2 14684 4558 14684 4558 5 dffrs_2.nand3_2.VSS
rlabel metal2 13270 6508 13270 6508 1 dffrs_2.nand3_1.VDD
rlabel metal1 13680 5382 13680 5382 3 dffrs_2.nand3_1.Z
rlabel metal1 12594 5264 12594 5264 7 dffrs_2.nand3_1.A
rlabel metal1 12594 5383 12594 5383 7 dffrs_2.nand3_1.B
rlabel metal1 12594 5499 12594 5499 7 dffrs_2.nand3_1.C
rlabel metal2 13198 4558 13198 4558 5 dffrs_2.nand3_1.VSS
rlabel metal2 13270 8713 13270 8713 1 dffrs_2.nand3_0.VDD
rlabel metal1 13680 7587 13680 7587 3 dffrs_2.nand3_0.Z
rlabel metal1 12594 7469 12594 7469 7 dffrs_2.nand3_0.A
rlabel metal1 12594 7588 12594 7588 7 dffrs_2.nand3_0.B
rlabel metal1 12594 7704 12594 7704 7 dffrs_2.nand3_0.C
rlabel metal2 13198 6763 13198 6763 5 dffrs_2.nand3_0.VSS
rlabel metal1 8064 7704 8064 7704 7 dffrs_1.setb
rlabel metal1 8064 4481 8064 4481 7 dffrs_1.clk
rlabel metal1 8064 856 8064 856 7 dffrs_1.d
rlabel metal1 8081 69 8081 69 7 dffrs_1.resetb
rlabel metal2 11532 5383 11532 5383 3 dffrs_1.Q
rlabel metal2 11532 3178 11532 3178 3 dffrs_1.Qb
rlabel metal5 10172 8809 10172 8809 1 dffrs_1.vdd
rlabel metal4 10280 30 10280 30 5 dffrs_1.vss
rlabel metal2 9228 2098 9228 2098 1 dffrs_1.nand3_8.VDD
rlabel metal1 9638 972 9638 972 3 dffrs_1.nand3_8.Z
rlabel metal1 8552 854 8552 854 7 dffrs_1.nand3_8.A
rlabel metal1 8552 973 8552 973 7 dffrs_1.nand3_8.B
rlabel metal1 8552 1089 8552 1089 7 dffrs_1.nand3_8.C
rlabel metal2 9156 148 9156 148 5 dffrs_1.nand3_8.VSS
rlabel metal2 10714 4304 10714 4304 1 dffrs_1.nand3_7.VDD
rlabel metal1 11124 3178 11124 3178 3 dffrs_1.nand3_7.Z
rlabel metal1 10038 3060 10038 3060 7 dffrs_1.nand3_7.A
rlabel metal1 10038 3179 10038 3179 7 dffrs_1.nand3_7.B
rlabel metal1 10038 3295 10038 3295 7 dffrs_1.nand3_7.C
rlabel metal2 10642 2354 10642 2354 5 dffrs_1.nand3_7.VSS
rlabel metal2 9228 4303 9228 4303 1 dffrs_1.nand3_6.VDD
rlabel metal1 9638 3177 9638 3177 3 dffrs_1.nand3_6.Z
rlabel metal1 8552 3059 8552 3059 7 dffrs_1.nand3_6.A
rlabel metal1 8552 3178 8552 3178 7 dffrs_1.nand3_6.B
rlabel metal1 8552 3294 8552 3294 7 dffrs_1.nand3_6.C
rlabel metal2 9156 2353 9156 2353 5 dffrs_1.nand3_6.VSS
rlabel metal2 10714 6508 10714 6508 1 dffrs_1.nand3_2.VDD
rlabel metal1 11124 5382 11124 5382 3 dffrs_1.nand3_2.Z
rlabel metal1 10038 5264 10038 5264 7 dffrs_1.nand3_2.A
rlabel metal1 10038 5383 10038 5383 7 dffrs_1.nand3_2.B
rlabel metal1 10038 5499 10038 5499 7 dffrs_1.nand3_2.C
rlabel metal2 10642 4558 10642 4558 5 dffrs_1.nand3_2.VSS
rlabel metal2 9228 6508 9228 6508 1 dffrs_1.nand3_1.VDD
rlabel metal1 9638 5382 9638 5382 3 dffrs_1.nand3_1.Z
rlabel metal1 8552 5264 8552 5264 7 dffrs_1.nand3_1.A
rlabel metal1 8552 5383 8552 5383 7 dffrs_1.nand3_1.B
rlabel metal1 8552 5499 8552 5499 7 dffrs_1.nand3_1.C
rlabel metal2 9156 4558 9156 4558 5 dffrs_1.nand3_1.VSS
rlabel metal2 9228 8713 9228 8713 1 dffrs_1.nand3_0.VDD
rlabel metal1 9638 7587 9638 7587 3 dffrs_1.nand3_0.Z
rlabel metal1 8552 7469 8552 7469 7 dffrs_1.nand3_0.A
rlabel metal1 8552 7588 8552 7588 7 dffrs_1.nand3_0.B
rlabel metal1 8552 7704 8552 7704 7 dffrs_1.nand3_0.C
rlabel metal2 9156 6763 9156 6763 5 dffrs_1.nand3_0.VSS
rlabel metal1 20190 7704 20190 7704 7 dffrs_4.setb
rlabel metal1 20190 4481 20190 4481 7 dffrs_4.clk
rlabel metal1 20190 856 20190 856 7 dffrs_4.d
rlabel metal1 20207 69 20207 69 7 dffrs_4.resetb
rlabel metal2 23658 5383 23658 5383 3 dffrs_4.Q
rlabel metal2 23658 3178 23658 3178 3 dffrs_4.Qb
rlabel metal5 22298 8809 22298 8809 1 dffrs_4.vdd
rlabel metal4 22406 30 22406 30 5 dffrs_4.vss
rlabel metal2 21354 2098 21354 2098 1 dffrs_4.nand3_8.VDD
rlabel metal1 21764 972 21764 972 3 dffrs_4.nand3_8.Z
rlabel metal1 20678 854 20678 854 7 dffrs_4.nand3_8.A
rlabel metal1 20678 973 20678 973 7 dffrs_4.nand3_8.B
rlabel metal1 20678 1089 20678 1089 7 dffrs_4.nand3_8.C
rlabel metal2 21282 148 21282 148 5 dffrs_4.nand3_8.VSS
rlabel metal2 22840 4304 22840 4304 1 dffrs_4.nand3_7.VDD
rlabel metal1 23250 3178 23250 3178 3 dffrs_4.nand3_7.Z
rlabel metal1 22164 3060 22164 3060 7 dffrs_4.nand3_7.A
rlabel metal1 22164 3179 22164 3179 7 dffrs_4.nand3_7.B
rlabel metal1 22164 3295 22164 3295 7 dffrs_4.nand3_7.C
rlabel metal2 22768 2354 22768 2354 5 dffrs_4.nand3_7.VSS
rlabel metal2 21354 4303 21354 4303 1 dffrs_4.nand3_6.VDD
rlabel metal1 21764 3177 21764 3177 3 dffrs_4.nand3_6.Z
rlabel metal1 20678 3059 20678 3059 7 dffrs_4.nand3_6.A
rlabel metal1 20678 3178 20678 3178 7 dffrs_4.nand3_6.B
rlabel metal1 20678 3294 20678 3294 7 dffrs_4.nand3_6.C
rlabel metal2 21282 2353 21282 2353 5 dffrs_4.nand3_6.VSS
rlabel metal2 22840 6508 22840 6508 1 dffrs_4.nand3_2.VDD
rlabel metal1 23250 5382 23250 5382 3 dffrs_4.nand3_2.Z
rlabel metal1 22164 5264 22164 5264 7 dffrs_4.nand3_2.A
rlabel metal1 22164 5383 22164 5383 7 dffrs_4.nand3_2.B
rlabel metal1 22164 5499 22164 5499 7 dffrs_4.nand3_2.C
rlabel metal2 22768 4558 22768 4558 5 dffrs_4.nand3_2.VSS
rlabel metal2 21354 6508 21354 6508 1 dffrs_4.nand3_1.VDD
rlabel metal1 21764 5382 21764 5382 3 dffrs_4.nand3_1.Z
rlabel metal1 20678 5264 20678 5264 7 dffrs_4.nand3_1.A
rlabel metal1 20678 5383 20678 5383 7 dffrs_4.nand3_1.B
rlabel metal1 20678 5499 20678 5499 7 dffrs_4.nand3_1.C
rlabel metal2 21282 4558 21282 4558 5 dffrs_4.nand3_1.VSS
rlabel metal2 21354 8713 21354 8713 1 dffrs_4.nand3_0.VDD
rlabel metal1 21764 7587 21764 7587 3 dffrs_4.nand3_0.Z
rlabel metal1 20678 7469 20678 7469 7 dffrs_4.nand3_0.A
rlabel metal1 20678 7588 20678 7588 7 dffrs_4.nand3_0.B
rlabel metal1 20678 7704 20678 7704 7 dffrs_4.nand3_0.C
rlabel metal2 21282 6763 21282 6763 5 dffrs_4.nand3_0.VSS
rlabel metal1 16148 7704 16148 7704 7 dffrs_3.setb
rlabel metal1 16148 4481 16148 4481 7 dffrs_3.clk
rlabel metal1 16148 856 16148 856 7 dffrs_3.d
rlabel metal1 16165 69 16165 69 7 dffrs_3.resetb
rlabel metal2 19616 5383 19616 5383 3 dffrs_3.Q
rlabel metal2 19616 3178 19616 3178 3 dffrs_3.Qb
rlabel metal5 18256 8809 18256 8809 1 dffrs_3.vdd
rlabel metal4 18364 30 18364 30 5 dffrs_3.vss
rlabel metal2 17312 2098 17312 2098 1 dffrs_3.nand3_8.VDD
rlabel metal1 17722 972 17722 972 3 dffrs_3.nand3_8.Z
rlabel metal1 16636 854 16636 854 7 dffrs_3.nand3_8.A
rlabel metal1 16636 973 16636 973 7 dffrs_3.nand3_8.B
rlabel metal1 16636 1089 16636 1089 7 dffrs_3.nand3_8.C
rlabel metal2 17240 148 17240 148 5 dffrs_3.nand3_8.VSS
rlabel metal2 18798 4304 18798 4304 1 dffrs_3.nand3_7.VDD
rlabel metal1 19208 3178 19208 3178 3 dffrs_3.nand3_7.Z
rlabel metal1 18122 3060 18122 3060 7 dffrs_3.nand3_7.A
rlabel metal1 18122 3179 18122 3179 7 dffrs_3.nand3_7.B
rlabel metal1 18122 3295 18122 3295 7 dffrs_3.nand3_7.C
rlabel metal2 18726 2354 18726 2354 5 dffrs_3.nand3_7.VSS
rlabel metal2 17312 4303 17312 4303 1 dffrs_3.nand3_6.VDD
rlabel metal1 17722 3177 17722 3177 3 dffrs_3.nand3_6.Z
rlabel metal1 16636 3059 16636 3059 7 dffrs_3.nand3_6.A
rlabel metal1 16636 3178 16636 3178 7 dffrs_3.nand3_6.B
rlabel metal1 16636 3294 16636 3294 7 dffrs_3.nand3_6.C
rlabel metal2 17240 2353 17240 2353 5 dffrs_3.nand3_6.VSS
rlabel metal2 18798 6508 18798 6508 1 dffrs_3.nand3_2.VDD
rlabel metal1 19208 5382 19208 5382 3 dffrs_3.nand3_2.Z
rlabel metal1 18122 5264 18122 5264 7 dffrs_3.nand3_2.A
rlabel metal1 18122 5383 18122 5383 7 dffrs_3.nand3_2.B
rlabel metal1 18122 5499 18122 5499 7 dffrs_3.nand3_2.C
rlabel metal2 18726 4558 18726 4558 5 dffrs_3.nand3_2.VSS
rlabel metal2 17312 6508 17312 6508 1 dffrs_3.nand3_1.VDD
rlabel metal1 17722 5382 17722 5382 3 dffrs_3.nand3_1.Z
rlabel metal1 16636 5264 16636 5264 7 dffrs_3.nand3_1.A
rlabel metal1 16636 5383 16636 5383 7 dffrs_3.nand3_1.B
rlabel metal1 16636 5499 16636 5499 7 dffrs_3.nand3_1.C
rlabel metal2 17240 4558 17240 4558 5 dffrs_3.nand3_1.VSS
rlabel metal2 17312 8713 17312 8713 1 dffrs_3.nand3_0.VDD
rlabel metal1 17722 7587 17722 7587 3 dffrs_3.nand3_0.Z
rlabel metal1 16636 7469 16636 7469 7 dffrs_3.nand3_0.A
rlabel metal1 16636 7588 16636 7588 7 dffrs_3.nand3_0.B
rlabel metal1 16636 7704 16636 7704 7 dffrs_3.nand3_0.C
rlabel metal2 17240 6763 17240 6763 5 dffrs_3.nand3_0.VSS
rlabel metal1 24232 7704 24232 7704 7 dffrs_5.setb
rlabel metal1 24232 4481 24232 4481 7 dffrs_5.clk
rlabel metal1 24232 856 24232 856 7 dffrs_5.d
rlabel metal1 24249 69 24249 69 7 dffrs_5.resetb
rlabel metal2 27700 5383 27700 5383 3 dffrs_5.Q
rlabel metal2 27700 3178 27700 3178 3 dffrs_5.Qb
rlabel metal5 26340 8809 26340 8809 1 dffrs_5.vdd
rlabel metal4 26448 30 26448 30 5 dffrs_5.vss
rlabel metal2 25396 2098 25396 2098 1 dffrs_5.nand3_8.VDD
rlabel metal1 25806 972 25806 972 3 dffrs_5.nand3_8.Z
rlabel metal1 24720 854 24720 854 7 dffrs_5.nand3_8.A
rlabel metal1 24720 973 24720 973 7 dffrs_5.nand3_8.B
rlabel metal1 24720 1089 24720 1089 7 dffrs_5.nand3_8.C
rlabel metal2 25324 148 25324 148 5 dffrs_5.nand3_8.VSS
rlabel metal2 26882 4304 26882 4304 1 dffrs_5.nand3_7.VDD
rlabel metal1 27292 3178 27292 3178 3 dffrs_5.nand3_7.Z
rlabel metal1 26206 3060 26206 3060 7 dffrs_5.nand3_7.A
rlabel metal1 26206 3179 26206 3179 7 dffrs_5.nand3_7.B
rlabel metal1 26206 3295 26206 3295 7 dffrs_5.nand3_7.C
rlabel metal2 26810 2354 26810 2354 5 dffrs_5.nand3_7.VSS
rlabel metal2 25396 4303 25396 4303 1 dffrs_5.nand3_6.VDD
rlabel metal1 25806 3177 25806 3177 3 dffrs_5.nand3_6.Z
rlabel metal1 24720 3059 24720 3059 7 dffrs_5.nand3_6.A
rlabel metal1 24720 3178 24720 3178 7 dffrs_5.nand3_6.B
rlabel metal1 24720 3294 24720 3294 7 dffrs_5.nand3_6.C
rlabel metal2 25324 2353 25324 2353 5 dffrs_5.nand3_6.VSS
rlabel metal2 26882 6508 26882 6508 1 dffrs_5.nand3_2.VDD
rlabel metal1 27292 5382 27292 5382 3 dffrs_5.nand3_2.Z
rlabel metal1 26206 5264 26206 5264 7 dffrs_5.nand3_2.A
rlabel metal1 26206 5383 26206 5383 7 dffrs_5.nand3_2.B
rlabel metal1 26206 5499 26206 5499 7 dffrs_5.nand3_2.C
rlabel metal2 26810 4558 26810 4558 5 dffrs_5.nand3_2.VSS
rlabel metal2 25396 6508 25396 6508 1 dffrs_5.nand3_1.VDD
rlabel metal1 25806 5382 25806 5382 3 dffrs_5.nand3_1.Z
rlabel metal1 24720 5264 24720 5264 7 dffrs_5.nand3_1.A
rlabel metal1 24720 5383 24720 5383 7 dffrs_5.nand3_1.B
rlabel metal1 24720 5499 24720 5499 7 dffrs_5.nand3_1.C
rlabel metal2 25324 4558 25324 4558 5 dffrs_5.nand3_1.VSS
rlabel metal2 25396 8713 25396 8713 1 dffrs_5.nand3_0.VDD
rlabel metal1 25806 7587 25806 7587 3 dffrs_5.nand3_0.Z
rlabel metal1 24720 7469 24720 7469 7 dffrs_5.nand3_0.A
rlabel metal1 24720 7588 24720 7588 7 dffrs_5.nand3_0.B
rlabel metal1 24720 7704 24720 7704 7 dffrs_5.nand3_0.C
rlabel metal2 25324 6763 25324 6763 5 dffrs_5.nand3_0.VSS
rlabel metal1 4022 17283 4022 17283 7 dffrs_14.setb
rlabel metal1 4022 14060 4022 14060 7 dffrs_14.clk
rlabel metal1 4022 10435 4022 10435 7 dffrs_14.d
rlabel metal1 4039 9648 4039 9648 7 dffrs_14.resetb
rlabel metal2 7490 14962 7490 14962 3 dffrs_14.Q
rlabel metal2 7490 12757 7490 12757 3 dffrs_14.Qb
rlabel metal5 6130 18388 6130 18388 1 dffrs_14.vdd
rlabel metal4 6238 9609 6238 9609 5 dffrs_14.vss
rlabel metal2 5186 11677 5186 11677 1 dffrs_14.nand3_8.VDD
rlabel metal1 5596 10551 5596 10551 3 dffrs_14.nand3_8.Z
rlabel metal1 4510 10433 4510 10433 7 dffrs_14.nand3_8.A
rlabel metal1 4510 10552 4510 10552 7 dffrs_14.nand3_8.B
rlabel metal1 4510 10668 4510 10668 7 dffrs_14.nand3_8.C
rlabel metal2 5114 9727 5114 9727 5 dffrs_14.nand3_8.VSS
rlabel metal2 6672 13883 6672 13883 1 dffrs_14.nand3_7.VDD
rlabel metal1 7082 12757 7082 12757 3 dffrs_14.nand3_7.Z
rlabel metal1 5996 12639 5996 12639 7 dffrs_14.nand3_7.A
rlabel metal1 5996 12758 5996 12758 7 dffrs_14.nand3_7.B
rlabel metal1 5996 12874 5996 12874 7 dffrs_14.nand3_7.C
rlabel metal2 6600 11933 6600 11933 5 dffrs_14.nand3_7.VSS
rlabel metal2 5186 13882 5186 13882 1 dffrs_14.nand3_6.VDD
rlabel metal1 5596 12756 5596 12756 3 dffrs_14.nand3_6.Z
rlabel metal1 4510 12638 4510 12638 7 dffrs_14.nand3_6.A
rlabel metal1 4510 12757 4510 12757 7 dffrs_14.nand3_6.B
rlabel metal1 4510 12873 4510 12873 7 dffrs_14.nand3_6.C
rlabel metal2 5114 11932 5114 11932 5 dffrs_14.nand3_6.VSS
rlabel metal2 6672 16087 6672 16087 1 dffrs_14.nand3_2.VDD
rlabel metal1 7082 14961 7082 14961 3 dffrs_14.nand3_2.Z
rlabel metal1 5996 14843 5996 14843 7 dffrs_14.nand3_2.A
rlabel metal1 5996 14962 5996 14962 7 dffrs_14.nand3_2.B
rlabel metal1 5996 15078 5996 15078 7 dffrs_14.nand3_2.C
rlabel metal2 6600 14137 6600 14137 5 dffrs_14.nand3_2.VSS
rlabel metal2 5186 16087 5186 16087 1 dffrs_14.nand3_1.VDD
rlabel metal1 5596 14961 5596 14961 3 dffrs_14.nand3_1.Z
rlabel metal1 4510 14843 4510 14843 7 dffrs_14.nand3_1.A
rlabel metal1 4510 14962 4510 14962 7 dffrs_14.nand3_1.B
rlabel metal1 4510 15078 4510 15078 7 dffrs_14.nand3_1.C
rlabel metal2 5114 14137 5114 14137 5 dffrs_14.nand3_1.VSS
rlabel metal2 5186 18292 5186 18292 1 dffrs_14.nand3_0.VDD
rlabel metal1 5596 17166 5596 17166 3 dffrs_14.nand3_0.Z
rlabel metal1 4510 17048 4510 17048 7 dffrs_14.nand3_0.A
rlabel metal1 4510 17167 4510 17167 7 dffrs_14.nand3_0.B
rlabel metal1 4510 17283 4510 17283 7 dffrs_14.nand3_0.C
rlabel metal2 5114 16342 5114 16342 5 dffrs_14.nand3_0.VSS
rlabel metal1 12106 17280 12106 17280 7 dffrs_8.setb
rlabel metal1 12106 14057 12106 14057 7 dffrs_8.clk
rlabel metal1 12106 10432 12106 10432 7 dffrs_8.d
rlabel metal1 12123 9645 12123 9645 7 dffrs_8.resetb
rlabel metal2 15574 14959 15574 14959 3 dffrs_8.Q
rlabel metal2 15574 12754 15574 12754 3 dffrs_8.Qb
rlabel metal5 14214 18385 14214 18385 1 dffrs_8.vdd
rlabel metal4 14322 9606 14322 9606 5 dffrs_8.vss
rlabel metal2 13270 11674 13270 11674 1 dffrs_8.nand3_8.VDD
rlabel metal1 13680 10548 13680 10548 3 dffrs_8.nand3_8.Z
rlabel metal1 12594 10430 12594 10430 7 dffrs_8.nand3_8.A
rlabel metal1 12594 10549 12594 10549 7 dffrs_8.nand3_8.B
rlabel metal1 12594 10665 12594 10665 7 dffrs_8.nand3_8.C
rlabel metal2 13198 9724 13198 9724 5 dffrs_8.nand3_8.VSS
rlabel metal2 14756 13880 14756 13880 1 dffrs_8.nand3_7.VDD
rlabel metal1 15166 12754 15166 12754 3 dffrs_8.nand3_7.Z
rlabel metal1 14080 12636 14080 12636 7 dffrs_8.nand3_7.A
rlabel metal1 14080 12755 14080 12755 7 dffrs_8.nand3_7.B
rlabel metal1 14080 12871 14080 12871 7 dffrs_8.nand3_7.C
rlabel metal2 14684 11930 14684 11930 5 dffrs_8.nand3_7.VSS
rlabel metal2 13270 13879 13270 13879 1 dffrs_8.nand3_6.VDD
rlabel metal1 13680 12753 13680 12753 3 dffrs_8.nand3_6.Z
rlabel metal1 12594 12635 12594 12635 7 dffrs_8.nand3_6.A
rlabel metal1 12594 12754 12594 12754 7 dffrs_8.nand3_6.B
rlabel metal1 12594 12870 12594 12870 7 dffrs_8.nand3_6.C
rlabel metal2 13198 11929 13198 11929 5 dffrs_8.nand3_6.VSS
rlabel metal2 14756 16084 14756 16084 1 dffrs_8.nand3_2.VDD
rlabel metal1 15166 14958 15166 14958 3 dffrs_8.nand3_2.Z
rlabel metal1 14080 14840 14080 14840 7 dffrs_8.nand3_2.A
rlabel metal1 14080 14959 14080 14959 7 dffrs_8.nand3_2.B
rlabel metal1 14080 15075 14080 15075 7 dffrs_8.nand3_2.C
rlabel metal2 14684 14134 14684 14134 5 dffrs_8.nand3_2.VSS
rlabel metal2 13270 16084 13270 16084 1 dffrs_8.nand3_1.VDD
rlabel metal1 13680 14958 13680 14958 3 dffrs_8.nand3_1.Z
rlabel metal1 12594 14840 12594 14840 7 dffrs_8.nand3_1.A
rlabel metal1 12594 14959 12594 14959 7 dffrs_8.nand3_1.B
rlabel metal1 12594 15075 12594 15075 7 dffrs_8.nand3_1.C
rlabel metal2 13198 14134 13198 14134 5 dffrs_8.nand3_1.VSS
rlabel metal2 13270 18289 13270 18289 1 dffrs_8.nand3_0.VDD
rlabel metal1 13680 17163 13680 17163 3 dffrs_8.nand3_0.Z
rlabel metal1 12594 17045 12594 17045 7 dffrs_8.nand3_0.A
rlabel metal1 12594 17164 12594 17164 7 dffrs_8.nand3_0.B
rlabel metal1 12594 17280 12594 17280 7 dffrs_8.nand3_0.C
rlabel metal2 13198 16339 13198 16339 5 dffrs_8.nand3_0.VSS
rlabel metal1 8064 17280 8064 17280 7 dffrs_7.setb
rlabel metal1 8064 14057 8064 14057 7 dffrs_7.clk
rlabel metal1 8064 10432 8064 10432 7 dffrs_7.d
rlabel metal1 8081 9645 8081 9645 7 dffrs_7.resetb
rlabel metal2 11532 14959 11532 14959 3 dffrs_7.Q
rlabel metal2 11532 12754 11532 12754 3 dffrs_7.Qb
rlabel metal5 10172 18385 10172 18385 1 dffrs_7.vdd
rlabel metal4 10280 9606 10280 9606 5 dffrs_7.vss
rlabel metal2 9228 11674 9228 11674 1 dffrs_7.nand3_8.VDD
rlabel metal1 9638 10548 9638 10548 3 dffrs_7.nand3_8.Z
rlabel metal1 8552 10430 8552 10430 7 dffrs_7.nand3_8.A
rlabel metal1 8552 10549 8552 10549 7 dffrs_7.nand3_8.B
rlabel metal1 8552 10665 8552 10665 7 dffrs_7.nand3_8.C
rlabel metal2 9156 9724 9156 9724 5 dffrs_7.nand3_8.VSS
rlabel metal2 10714 13880 10714 13880 1 dffrs_7.nand3_7.VDD
rlabel metal1 11124 12754 11124 12754 3 dffrs_7.nand3_7.Z
rlabel metal1 10038 12636 10038 12636 7 dffrs_7.nand3_7.A
rlabel metal1 10038 12755 10038 12755 7 dffrs_7.nand3_7.B
rlabel metal1 10038 12871 10038 12871 7 dffrs_7.nand3_7.C
rlabel metal2 10642 11930 10642 11930 5 dffrs_7.nand3_7.VSS
rlabel metal2 9228 13879 9228 13879 1 dffrs_7.nand3_6.VDD
rlabel metal1 9638 12753 9638 12753 3 dffrs_7.nand3_6.Z
rlabel metal1 8552 12635 8552 12635 7 dffrs_7.nand3_6.A
rlabel metal1 8552 12754 8552 12754 7 dffrs_7.nand3_6.B
rlabel metal1 8552 12870 8552 12870 7 dffrs_7.nand3_6.C
rlabel metal2 9156 11929 9156 11929 5 dffrs_7.nand3_6.VSS
rlabel metal2 10714 16084 10714 16084 1 dffrs_7.nand3_2.VDD
rlabel metal1 11124 14958 11124 14958 3 dffrs_7.nand3_2.Z
rlabel metal1 10038 14840 10038 14840 7 dffrs_7.nand3_2.A
rlabel metal1 10038 14959 10038 14959 7 dffrs_7.nand3_2.B
rlabel metal1 10038 15075 10038 15075 7 dffrs_7.nand3_2.C
rlabel metal2 10642 14134 10642 14134 5 dffrs_7.nand3_2.VSS
rlabel metal2 9228 16084 9228 16084 1 dffrs_7.nand3_1.VDD
rlabel metal1 9638 14958 9638 14958 3 dffrs_7.nand3_1.Z
rlabel metal1 8552 14840 8552 14840 7 dffrs_7.nand3_1.A
rlabel metal1 8552 14959 8552 14959 7 dffrs_7.nand3_1.B
rlabel metal1 8552 15075 8552 15075 7 dffrs_7.nand3_1.C
rlabel metal2 9156 14134 9156 14134 5 dffrs_7.nand3_1.VSS
rlabel metal2 9228 18289 9228 18289 1 dffrs_7.nand3_0.VDD
rlabel metal1 9638 17163 9638 17163 3 dffrs_7.nand3_0.Z
rlabel metal1 8552 17045 8552 17045 7 dffrs_7.nand3_0.A
rlabel metal1 8552 17164 8552 17164 7 dffrs_7.nand3_0.B
rlabel metal1 8552 17280 8552 17280 7 dffrs_7.nand3_0.C
rlabel metal2 9156 16339 9156 16339 5 dffrs_7.nand3_0.VSS
rlabel metal1 20190 17280 20190 17280 7 dffrs_10.setb
rlabel metal1 20190 14057 20190 14057 7 dffrs_10.clk
rlabel metal1 20190 10432 20190 10432 7 dffrs_10.d
rlabel metal1 20207 9645 20207 9645 7 dffrs_10.resetb
rlabel metal2 23658 14959 23658 14959 3 dffrs_10.Q
rlabel metal2 23658 12754 23658 12754 3 dffrs_10.Qb
rlabel metal5 22298 18385 22298 18385 1 dffrs_10.vdd
rlabel metal4 22406 9606 22406 9606 5 dffrs_10.vss
rlabel metal2 21354 11674 21354 11674 1 dffrs_10.nand3_8.VDD
rlabel metal1 21764 10548 21764 10548 3 dffrs_10.nand3_8.Z
rlabel metal1 20678 10430 20678 10430 7 dffrs_10.nand3_8.A
rlabel metal1 20678 10549 20678 10549 7 dffrs_10.nand3_8.B
rlabel metal1 20678 10665 20678 10665 7 dffrs_10.nand3_8.C
rlabel metal2 21282 9724 21282 9724 5 dffrs_10.nand3_8.VSS
rlabel metal2 22840 13880 22840 13880 1 dffrs_10.nand3_7.VDD
rlabel metal1 23250 12754 23250 12754 3 dffrs_10.nand3_7.Z
rlabel metal1 22164 12636 22164 12636 7 dffrs_10.nand3_7.A
rlabel metal1 22164 12755 22164 12755 7 dffrs_10.nand3_7.B
rlabel metal1 22164 12871 22164 12871 7 dffrs_10.nand3_7.C
rlabel metal2 22768 11930 22768 11930 5 dffrs_10.nand3_7.VSS
rlabel metal2 21354 13879 21354 13879 1 dffrs_10.nand3_6.VDD
rlabel metal1 21764 12753 21764 12753 3 dffrs_10.nand3_6.Z
rlabel metal1 20678 12635 20678 12635 7 dffrs_10.nand3_6.A
rlabel metal1 20678 12754 20678 12754 7 dffrs_10.nand3_6.B
rlabel metal1 20678 12870 20678 12870 7 dffrs_10.nand3_6.C
rlabel metal2 21282 11929 21282 11929 5 dffrs_10.nand3_6.VSS
rlabel metal2 22840 16084 22840 16084 1 dffrs_10.nand3_2.VDD
rlabel metal1 23250 14958 23250 14958 3 dffrs_10.nand3_2.Z
rlabel metal1 22164 14840 22164 14840 7 dffrs_10.nand3_2.A
rlabel metal1 22164 14959 22164 14959 7 dffrs_10.nand3_2.B
rlabel metal1 22164 15075 22164 15075 7 dffrs_10.nand3_2.C
rlabel metal2 22768 14134 22768 14134 5 dffrs_10.nand3_2.VSS
rlabel metal2 21354 16084 21354 16084 1 dffrs_10.nand3_1.VDD
rlabel metal1 21764 14958 21764 14958 3 dffrs_10.nand3_1.Z
rlabel metal1 20678 14840 20678 14840 7 dffrs_10.nand3_1.A
rlabel metal1 20678 14959 20678 14959 7 dffrs_10.nand3_1.B
rlabel metal1 20678 15075 20678 15075 7 dffrs_10.nand3_1.C
rlabel metal2 21282 14134 21282 14134 5 dffrs_10.nand3_1.VSS
rlabel metal2 21354 18289 21354 18289 1 dffrs_10.nand3_0.VDD
rlabel metal1 21764 17163 21764 17163 3 dffrs_10.nand3_0.Z
rlabel metal1 20678 17045 20678 17045 7 dffrs_10.nand3_0.A
rlabel metal1 20678 17164 20678 17164 7 dffrs_10.nand3_0.B
rlabel metal1 20678 17280 20678 17280 7 dffrs_10.nand3_0.C
rlabel metal2 21282 16339 21282 16339 5 dffrs_10.nand3_0.VSS
rlabel metal1 16148 17280 16148 17280 7 dffrs_9.setb
rlabel metal1 16148 14057 16148 14057 7 dffrs_9.clk
rlabel metal1 16148 10432 16148 10432 7 dffrs_9.d
rlabel metal1 16165 9645 16165 9645 7 dffrs_9.resetb
rlabel metal2 19616 14959 19616 14959 3 dffrs_9.Q
rlabel metal2 19616 12754 19616 12754 3 dffrs_9.Qb
rlabel metal5 18256 18385 18256 18385 1 dffrs_9.vdd
rlabel metal4 18364 9606 18364 9606 5 dffrs_9.vss
rlabel metal2 17312 11674 17312 11674 1 dffrs_9.nand3_8.VDD
rlabel metal1 17722 10548 17722 10548 3 dffrs_9.nand3_8.Z
rlabel metal1 16636 10430 16636 10430 7 dffrs_9.nand3_8.A
rlabel metal1 16636 10549 16636 10549 7 dffrs_9.nand3_8.B
rlabel metal1 16636 10665 16636 10665 7 dffrs_9.nand3_8.C
rlabel metal2 17240 9724 17240 9724 5 dffrs_9.nand3_8.VSS
rlabel metal2 18798 13880 18798 13880 1 dffrs_9.nand3_7.VDD
rlabel metal1 19208 12754 19208 12754 3 dffrs_9.nand3_7.Z
rlabel metal1 18122 12636 18122 12636 7 dffrs_9.nand3_7.A
rlabel metal1 18122 12755 18122 12755 7 dffrs_9.nand3_7.B
rlabel metal1 18122 12871 18122 12871 7 dffrs_9.nand3_7.C
rlabel metal2 18726 11930 18726 11930 5 dffrs_9.nand3_7.VSS
rlabel metal2 17312 13879 17312 13879 1 dffrs_9.nand3_6.VDD
rlabel metal1 17722 12753 17722 12753 3 dffrs_9.nand3_6.Z
rlabel metal1 16636 12635 16636 12635 7 dffrs_9.nand3_6.A
rlabel metal1 16636 12754 16636 12754 7 dffrs_9.nand3_6.B
rlabel metal1 16636 12870 16636 12870 7 dffrs_9.nand3_6.C
rlabel metal2 17240 11929 17240 11929 5 dffrs_9.nand3_6.VSS
rlabel metal2 18798 16084 18798 16084 1 dffrs_9.nand3_2.VDD
rlabel metal1 19208 14958 19208 14958 3 dffrs_9.nand3_2.Z
rlabel metal1 18122 14840 18122 14840 7 dffrs_9.nand3_2.A
rlabel metal1 18122 14959 18122 14959 7 dffrs_9.nand3_2.B
rlabel metal1 18122 15075 18122 15075 7 dffrs_9.nand3_2.C
rlabel metal2 18726 14134 18726 14134 5 dffrs_9.nand3_2.VSS
rlabel metal2 17312 16084 17312 16084 1 dffrs_9.nand3_1.VDD
rlabel metal1 17722 14958 17722 14958 3 dffrs_9.nand3_1.Z
rlabel metal1 16636 14840 16636 14840 7 dffrs_9.nand3_1.A
rlabel metal1 16636 14959 16636 14959 7 dffrs_9.nand3_1.B
rlabel metal1 16636 15075 16636 15075 7 dffrs_9.nand3_1.C
rlabel metal2 17240 14134 17240 14134 5 dffrs_9.nand3_1.VSS
rlabel metal2 17312 18289 17312 18289 1 dffrs_9.nand3_0.VDD
rlabel metal1 17722 17163 17722 17163 3 dffrs_9.nand3_0.Z
rlabel metal1 16636 17045 16636 17045 7 dffrs_9.nand3_0.A
rlabel metal1 16636 17164 16636 17164 7 dffrs_9.nand3_0.B
rlabel metal1 16636 17280 16636 17280 7 dffrs_9.nand3_0.C
rlabel metal2 17240 16339 17240 16339 5 dffrs_9.nand3_0.VSS
rlabel metal1 28274 17280 28274 17280 7 dffrs_12.setb
rlabel metal1 28274 14057 28274 14057 7 dffrs_12.clk
rlabel metal1 28274 10432 28274 10432 7 dffrs_12.d
rlabel metal1 28291 9645 28291 9645 7 dffrs_12.resetb
rlabel metal2 31742 14959 31742 14959 3 dffrs_12.Q
rlabel metal2 31742 12754 31742 12754 3 dffrs_12.Qb
rlabel metal5 30382 18385 30382 18385 1 dffrs_12.vdd
rlabel metal4 30490 9606 30490 9606 5 dffrs_12.vss
rlabel metal2 29438 11674 29438 11674 1 dffrs_12.nand3_8.VDD
rlabel metal1 29848 10548 29848 10548 3 dffrs_12.nand3_8.Z
rlabel metal1 28762 10430 28762 10430 7 dffrs_12.nand3_8.A
rlabel metal1 28762 10549 28762 10549 7 dffrs_12.nand3_8.B
rlabel metal1 28762 10665 28762 10665 7 dffrs_12.nand3_8.C
rlabel metal2 29366 9724 29366 9724 5 dffrs_12.nand3_8.VSS
rlabel metal2 30924 13880 30924 13880 1 dffrs_12.nand3_7.VDD
rlabel metal1 31334 12754 31334 12754 3 dffrs_12.nand3_7.Z
rlabel metal1 30248 12636 30248 12636 7 dffrs_12.nand3_7.A
rlabel metal1 30248 12755 30248 12755 7 dffrs_12.nand3_7.B
rlabel metal1 30248 12871 30248 12871 7 dffrs_12.nand3_7.C
rlabel metal2 30852 11930 30852 11930 5 dffrs_12.nand3_7.VSS
rlabel metal2 29438 13879 29438 13879 1 dffrs_12.nand3_6.VDD
rlabel metal1 29848 12753 29848 12753 3 dffrs_12.nand3_6.Z
rlabel metal1 28762 12635 28762 12635 7 dffrs_12.nand3_6.A
rlabel metal1 28762 12754 28762 12754 7 dffrs_12.nand3_6.B
rlabel metal1 28762 12870 28762 12870 7 dffrs_12.nand3_6.C
rlabel metal2 29366 11929 29366 11929 5 dffrs_12.nand3_6.VSS
rlabel metal2 30924 16084 30924 16084 1 dffrs_12.nand3_2.VDD
rlabel metal1 31334 14958 31334 14958 3 dffrs_12.nand3_2.Z
rlabel metal1 30248 14840 30248 14840 7 dffrs_12.nand3_2.A
rlabel metal1 30248 14959 30248 14959 7 dffrs_12.nand3_2.B
rlabel metal1 30248 15075 30248 15075 7 dffrs_12.nand3_2.C
rlabel metal2 30852 14134 30852 14134 5 dffrs_12.nand3_2.VSS
rlabel metal2 29438 16084 29438 16084 1 dffrs_12.nand3_1.VDD
rlabel metal1 29848 14958 29848 14958 3 dffrs_12.nand3_1.Z
rlabel metal1 28762 14840 28762 14840 7 dffrs_12.nand3_1.A
rlabel metal1 28762 14959 28762 14959 7 dffrs_12.nand3_1.B
rlabel metal1 28762 15075 28762 15075 7 dffrs_12.nand3_1.C
rlabel metal2 29366 14134 29366 14134 5 dffrs_12.nand3_1.VSS
rlabel metal2 29438 18289 29438 18289 1 dffrs_12.nand3_0.VDD
rlabel metal1 29848 17163 29848 17163 3 dffrs_12.nand3_0.Z
rlabel metal1 28762 17045 28762 17045 7 dffrs_12.nand3_0.A
rlabel metal1 28762 17164 28762 17164 7 dffrs_12.nand3_0.B
rlabel metal1 28762 17280 28762 17280 7 dffrs_12.nand3_0.C
rlabel metal2 29366 16339 29366 16339 5 dffrs_12.nand3_0.VSS
rlabel metal1 24232 17280 24232 17280 7 dffrs_11.setb
rlabel metal1 24232 14057 24232 14057 7 dffrs_11.clk
rlabel metal1 24232 10432 24232 10432 7 dffrs_11.d
rlabel metal1 24249 9645 24249 9645 7 dffrs_11.resetb
rlabel metal2 27700 14959 27700 14959 3 dffrs_11.Q
rlabel metal2 27700 12754 27700 12754 3 dffrs_11.Qb
rlabel metal5 26340 18385 26340 18385 1 dffrs_11.vdd
rlabel metal4 26448 9606 26448 9606 5 dffrs_11.vss
rlabel metal2 25396 11674 25396 11674 1 dffrs_11.nand3_8.VDD
rlabel metal1 25806 10548 25806 10548 3 dffrs_11.nand3_8.Z
rlabel metal1 24720 10430 24720 10430 7 dffrs_11.nand3_8.A
rlabel metal1 24720 10549 24720 10549 7 dffrs_11.nand3_8.B
rlabel metal1 24720 10665 24720 10665 7 dffrs_11.nand3_8.C
rlabel metal2 25324 9724 25324 9724 5 dffrs_11.nand3_8.VSS
rlabel metal2 26882 13880 26882 13880 1 dffrs_11.nand3_7.VDD
rlabel metal1 27292 12754 27292 12754 3 dffrs_11.nand3_7.Z
rlabel metal1 26206 12636 26206 12636 7 dffrs_11.nand3_7.A
rlabel metal1 26206 12755 26206 12755 7 dffrs_11.nand3_7.B
rlabel metal1 26206 12871 26206 12871 7 dffrs_11.nand3_7.C
rlabel metal2 26810 11930 26810 11930 5 dffrs_11.nand3_7.VSS
rlabel metal2 25396 13879 25396 13879 1 dffrs_11.nand3_6.VDD
rlabel metal1 25806 12753 25806 12753 3 dffrs_11.nand3_6.Z
rlabel metal1 24720 12635 24720 12635 7 dffrs_11.nand3_6.A
rlabel metal1 24720 12754 24720 12754 7 dffrs_11.nand3_6.B
rlabel metal1 24720 12870 24720 12870 7 dffrs_11.nand3_6.C
rlabel metal2 25324 11929 25324 11929 5 dffrs_11.nand3_6.VSS
rlabel metal2 26882 16084 26882 16084 1 dffrs_11.nand3_2.VDD
rlabel metal1 27292 14958 27292 14958 3 dffrs_11.nand3_2.Z
rlabel metal1 26206 14840 26206 14840 7 dffrs_11.nand3_2.A
rlabel metal1 26206 14959 26206 14959 7 dffrs_11.nand3_2.B
rlabel metal1 26206 15075 26206 15075 7 dffrs_11.nand3_2.C
rlabel metal2 26810 14134 26810 14134 5 dffrs_11.nand3_2.VSS
rlabel metal2 25396 16084 25396 16084 1 dffrs_11.nand3_1.VDD
rlabel metal1 25806 14958 25806 14958 3 dffrs_11.nand3_1.Z
rlabel metal1 24720 14840 24720 14840 7 dffrs_11.nand3_1.A
rlabel metal1 24720 14959 24720 14959 7 dffrs_11.nand3_1.B
rlabel metal1 24720 15075 24720 15075 7 dffrs_11.nand3_1.C
rlabel metal2 25324 14134 25324 14134 5 dffrs_11.nand3_1.VSS
rlabel metal2 25396 18289 25396 18289 1 dffrs_11.nand3_0.VDD
rlabel metal1 25806 17163 25806 17163 3 dffrs_11.nand3_0.Z
rlabel metal1 24720 17045 24720 17045 7 dffrs_11.nand3_0.A
rlabel metal1 24720 17164 24720 17164 7 dffrs_11.nand3_0.B
rlabel metal1 24720 17280 24720 17280 7 dffrs_11.nand3_0.C
rlabel metal2 25324 16339 25324 16339 5 dffrs_11.nand3_0.VSS
<< end >>
