* NGSPICE file created from comp_SAR_final.ext - technology: (null)

.subckt comp_SAR_final Clk_piso Vdd Vss Load Clk Piso_out Vin1 Vin2 Comp_out Reset SAR_in
X0 Vdd.t900 SARlogic_0.d3.t4 SARlogic_0.dffrs_7.nand3_8.C.t3 Vdd.t899 pfet_03v3
**devattr s=26000,604 d=26000,604
X1 a_5803_9634 SARlogic_0.dffrs_4.d.t4 Vss.t619 Vss.t618 nfet_03v3
**devattr s=17600,576 d=10400,304
X2 adc_PISO_0.dffrs_4.Qb Vdd.t730 Vdd.t732 Vdd.t731 pfet_03v3
**devattr s=26000,604 d=44000,1176
X3 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t4 Vdd.t928 Vdd.t927 pfet_03v3
**devattr s=26000,604 d=44000,1176
X4 a_37687_30440 inv2_0.out.t2 a_37499_31160.t2 Vss.t549 nfet_03v3
**devattr s=17600,576 d=10400,304
X5 a_n7937_n2793 a_n8017_n2885 a_n9429_n2007.t0 Vss.t116 nfet_03v3
**devattr s=8320,264 d=14080,496
X6 a_28027_28820.t2 SARlogic_0.d1.t4 Vdd.t804 Vdd.t803 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X7 Vss.t543 a_8377_29020 a_9271_28100 Vss.t542 nfet_03v3
**devattr s=10400,304 d=17600,576
X8 Vdd.t519 Reset.t0 SARlogic_0.dffrs_14.nand3_6.C.t1 Vdd.t518 pfet_03v3
**devattr s=26000,604 d=26000,604
X9 a_n7809_21417 SARlogic_0.dffrs_14.nand3_1.C Vss.t56 Vss.t55 nfet_03v3
**devattr s=17600,576 d=10400,304
X10 SARlogic_0.dffrs_2.nand3_1.C.t3 SARlogic_0.dffrs_2.nand3_6.C.t4 a_459_14043 Vss.t381 nfet_03v3
**devattr s=10400,304 d=17600,576
X11 SARlogic_0.d3.t3 SARlogic_0.dffrs_1.Qb.t4 Vdd.t491 Vdd.t490 pfet_03v3
**devattr s=44000,1176 d=26000,604
X12 SARlogic_0.dffrs_4.nand3_8.C.t0 SARlogic_0.dffrs_4.nand3_8.Z.t4 a_8543_9633 Vss.t334 nfet_03v3
**devattr s=10400,304 d=17600,576
X13 Vdd.t443 SARlogic_0.dffrs_1.nand3_8.C.t4 SARlogic_0.dffrs_1.Qb.t3 Vdd.t442 pfet_03v3
**devattr s=26000,604 d=26000,604
X14 adc_PISO_0.dffrs_0.Qb Vdd.t727 Vdd.t729 Vdd.t728 pfet_03v3
**devattr s=26000,604 d=44000,1176
X15 a_12401_7428 SARlogic_0.dffrs_5.nand3_8.C.t4 Vss.t404 Vss.t403 nfet_03v3
**devattr s=17600,576 d=10400,304
X16 SARlogic_0.dffrs_3.nand3_8.C.t1 SARlogic_0.dffrs_3.nand3_8.Z.t4 Vdd.t551 Vdd.t550 pfet_03v3
**devattr s=26000,604 d=44000,1176
X17 Vdd.t726 Vdd.t724 a_33257_31423.t0 Vdd.t725 pfet_03v3
**devattr s=26000,604 d=26000,604
X18 SARlogic_0.dffrs_5.nand3_8.C.t3 SARlogic_0.dffrs_5.nand3_6.C.t4 Vdd.t922 Vdd.t921 pfet_03v3
**devattr s=44000,1176 d=26000,604
X19 a_14071_9634 SARlogic_0.dffrs_5.nand3_8.C.t5 a_13887_9634 Vss.t405 nfet_03v3
**devattr s=10400,304 d=10400,304
X20 SARlogic_0.dffrs_1.Qb.t2 Reset.t1 Vdd.t449 Vdd.t448 pfet_03v3
**devattr s=26000,604 d=44000,1176
X21 a_18113_19210 SARlogic_0.dffrs_12.nand3_8.C.t4 a_17929_19210 Vss.t413 nfet_03v3
**devattr s=10400,304 d=10400,304
X22 Vdd.t391 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t8 Vdd.t390 pfet_03v3
**devattr s=10400,304 d=10400,304
X23 a_10029_9634 SARlogic_0.dffrs_4.nand3_8.C.t4 a_9845_9634 Vss.t396 nfet_03v3
**devattr s=10400,304 d=10400,304
X24 SARlogic_0.dffrs_1.nand3_6.C.t1 Clk.t0 a_n3583_11838 Vss.t48 nfet_03v3
**devattr s=10400,304 d=17600,576
X25 a_n4367_29309 Vdd.t945 a_n4551_29309 Vss.t523 nfet_03v3
**devattr s=10400,304 d=10400,304
X26 SARlogic_0.dffrs_9.Qb SARlogic_0.d2.t4 Vdd.t291 Vdd.t290 pfet_03v3
**devattr s=44000,1176 d=26000,604
X27 a_4841_33627.t3 a_4841_31422.t4 Vdd.t347 Vdd.t346 pfet_03v3
**devattr s=26000,604 d=44000,1176
X28 Vdd.t511 adc_PISO_0.2inmux_1.Bit.t4 a_37499_31160.t0 Vdd.t510 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X29 SARlogic_0.dffrs_5.nand3_6.C.t2 SARlogic_0.dffrs_5.nand3_1.C.t4 Vdd.t239 Vdd.t238 pfet_03v3
**devattr s=44000,1176 d=26000,604
X30 SARlogic_0.dffrs_4.d.t3 Vdd.t721 Vdd.t723 Vdd.t722 pfet_03v3
**devattr s=44000,1176 d=26000,604
X31 SARlogic_0.dffrs_3.nand3_6.C.t2 Clk.t1 Vdd.t65 Vdd.t64 pfet_03v3
**devattr s=26000,604 d=44000,1176
X32 Vdd.t451 Reset.t2 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t450 pfet_03v3
**devattr s=26000,604 d=26000,604
X33 Vdd.t822 a_33337_30170.t4 a_33257_33628.t2 Vdd.t821 pfet_03v3
**devattr s=26000,604 d=26000,604
X34 SARlogic_0.dffrs_13.Qb.t1 SARlogic_0.dffrs_0.d.t4 Vdd.t794 Vdd.t793 pfet_03v3
**devattr s=44000,1176 d=26000,604
X35 Vdd.t790 a_n10831_4320 Comp_out.t7 Vdd.t789 pfet_03v3
**devattr s=18700,450 d=18700,450
X36 a_10639_28100 a_9083_28820.t4 Vdd.t914 Vdd.t913 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X37 a_5987_21414 SARlogic_0.dffrs_9.nand3_6.C.t4 a_5803_21414 Vss.t656 nfet_03v3
**devattr s=10400,304 d=10400,304
X38 a_275_7428 SARlogic_0.dffrs_2.nand3_8.C.t4 Vss.t666 Vss.t665 nfet_03v3
**devattr s=17600,576 d=10400,304
X39 adc_PISO_0.2inmux_5.OUT.t0 a_30255_29264.t4 Vss.t201 Vss.t200 nfet_03v3
**devattr s=17600,576 d=17600,576
X40 SARlogic_0.dffrs_10.nand3_6.C.t3 SARlogic_0.d0.t4 Vdd.t259 Vdd.t258 pfet_03v3
**devattr s=26000,604 d=44000,1176
X41 SARlogic_0.d1.t1 SARlogic_0.dffrs_3.Qb.t4 Vdd.t395 Vdd.t394 pfet_03v3
**devattr s=44000,1176 d=26000,604
X42 a_12585_21414 Reset.t3 a_12401_21414 Vss.t348 nfet_03v3
**devattr s=10400,304 d=10400,304
X43 SARlogic_0.dffrs_3.Qb.t0 Reset.t4 a_5987_9634 Vss.t349 nfet_03v3
**devattr s=10400,304 d=17600,576
X44 SARlogic_0.dffrs_12.nand3_6.C.t0 SARlogic_0.dffrs_12.nand3_1.C Vdd.t103 Vdd.t102 pfet_03v3
**devattr s=44000,1176 d=26000,604
X45 SARlogic_0.dffrs_1.Qb.t1 Reset.t5 a_n2097_9634 Vss.t350 nfet_03v3
**devattr s=10400,304 d=17600,576
X46 a_n11637_11838 Vdd.t946 a_n11821_11838 Vss.t522 nfet_03v3
**devattr s=10400,304 d=10400,304
X47 a_n4551_35924 Vdd.t947 Vss.t521 Vss.t520 nfet_03v3
**devattr s=17600,576 d=10400,304
X48 SARlogic_0.dffrs_4.nand3_8.Z.t1 SARlogic_0.dffrs_4.nand3_8.C.t5 Vdd.t521 Vdd.t520 pfet_03v3
**devattr s=44000,1176 d=26000,604
X49 a_1761_19210 SARlogic_0.d3.t5 Vss.t643 Vss.t642 nfet_03v3
**devattr s=17600,576 d=10400,304
X50 a_14393_33720 a_14313_33628.t4 Vss.t267 Vss.t266 nfet_03v3
**devattr s=17600,576 d=10400,304
X51 a_9271_28100 SARlogic_0.d3.t6 a_9083_28820.t2 Vss.t641 nfet_03v3
**devattr s=17600,576 d=10400,304
X52 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t4 Vdd.t125 Vdd.t124 pfet_03v3
**devattr s=26000,604 d=44000,1176
X53 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_5.Qb.t4 Vdd.t427 Vdd.t426 pfet_03v3
**devattr s=44000,1176 d=26000,604
X54 a_12585_23619 SARlogic_0.dffrs_11.nand3_8.Z a_12401_23619 Vss.t135 nfet_03v3
**devattr s=10400,304 d=10400,304
X55 adc_PISO_0.dffrs_1.Qb adc_PISO_0.dffrs_1.Q.t4 Vdd.t267 Vdd.t266 pfet_03v3
**devattr s=44000,1176 d=26000,604
X56 Vdd.t483 SARlogic_0.dffrs_14.nand3_6.C.t4 SARlogic_0.d5.t0 Vdd.t482 pfet_03v3
**devattr s=26000,604 d=26000,604
X57 a_275_14043 Vdd.t948 Vss.t519 Vss.t518 nfet_03v3
**devattr s=17600,576 d=10400,304
X58 a_33257_29218.t2 a_33337_30170.t5 a_33521_31515 Vss.t589 nfet_03v3
**devattr s=10400,304 d=17600,576
X59 SARlogic_0.dffrs_0.Qb.t3 Reset.t6 a_n6139_9634 Vss.t351 nfet_03v3
**devattr s=10400,304 d=17600,576
X60 a_14393_35925 Vdd.t949 Vss.t517 Vss.t516 nfet_03v3
**devattr s=17600,576 d=10400,304
X61 SARlogic_0.dffrs_3.nand3_8.C.t2 SARlogic_0.dffrs_3.nand3_6.C.t4 Vdd.t433 Vdd.t432 pfet_03v3
**devattr s=44000,1176 d=26000,604
X62 a_9083_31160.t3 inv2_0.out.t3 a_9271_30440 Vss.t550 nfet_03v3
**devattr s=10400,304 d=17600,576
X63 a_23865_30170.t0 a_23785_29218.t4 Vdd.t181 Vdd.t180 pfet_03v3
**devattr s=44000,1176 d=26000,604
X64 a_18743_28100 a_17849_29020 Vss.t74 Vss.t73 nfet_03v3
**devattr s=17600,576 d=10400,304
X65 a_9845_19210 SARlogic_0.d1.t5 Vss.t583 Vss.t582 nfet_03v3
**devattr s=17600,576 d=10400,304
X66 SARlogic_0.dffrs_3.nand3_6.C.t3 SARlogic_0.dffrs_3.nand3_1.C.t4 Vdd.t189 Vdd.t188 pfet_03v3
**devattr s=44000,1176 d=26000,604
X67 a_42729_31423.t1 a_42729_33628.t4 Vdd.t131 Vdd.t130 pfet_03v3
**devattr s=44000,1176 d=26000,604
X68 a_29583_30440 a_28027_31160.t4 Vdd.t846 Vdd.t845 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X69 SARlogic_0.dffrs_13.Qb.t3 Vdd.t718 Vdd.t720 Vdd.t719 pfet_03v3
**devattr s=26000,604 d=44000,1176
X70 a_23785_29218.t2 a_23785_31423.t4 Vdd.t864 Vdd.t863 pfet_03v3
**devattr s=44000,1176 d=26000,604
X71 Vdd.t101 a_20111_30440 a_20971_29984 Vdd.t100 pfet_03v3
**devattr s=31200,704 d=52800,1376
X72 a_n9429_n2007.t16 Vin1.t0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t16 Vss.t181 nfet_03v3
**devattr s=15600,404 d=15600,404
X73 a_28027_31160.t2 inv2_0.out.t4 a_28215_30440 Vss.t551 nfet_03v3
**devattr s=10400,304 d=17600,576
X74 SARlogic_0.dffrs_10.nand3_6.C.t1 SARlogic_0.dffrs_10.nand3_1.C Vdd.t109 Vdd.t108 pfet_03v3
**devattr s=44000,1176 d=26000,604
X75 a_42729_33628.t1 Vdd.t715 Vdd.t717 Vdd.t716 pfet_03v3
**devattr s=44000,1176 d=26000,604
X76 a_n4631_33627.t0 a_n4631_31422.t4 a_n4367_35924 Vss.t524 nfet_03v3
**devattr s=10400,304 d=17600,576
X77 a_12401_17004 SARlogic_0.dffrs_11.nand3_8.C.t4 Vss.t167 Vss.t166 nfet_03v3
**devattr s=17600,576 d=10400,304
X78 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t0 a_4501_17004 Vss.t423 nfet_03v3
**devattr s=10400,304 d=17600,576
X79 a_n8305_30439 a_n9861_31159.t4 Vdd.t319 Vdd.t318 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X80 a_n6139_19213 SARlogic_0.dffrs_14.nand3_8.C.t4 a_n6323_19213 Vss.t532 nfet_03v3
**devattr s=10400,304 d=10400,304
X81 a_n201_28099 a_n1095_29019 Vss.t64 Vss.t63 nfet_03v3
**devattr s=17600,576 d=10400,304
X82 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_3.Qb.t5 Vdd.t397 Vdd.t396 pfet_03v3
**devattr s=44000,1176 d=26000,604
X83 SARlogic_0.d1.t3 SARlogic_0.dffrs_10.Qb Vdd.t750 Vdd.t749 pfet_03v3
**devattr s=26000,604 d=44000,1176
X84 Vdd.t714 Vdd.t712 SARlogic_0.dffrs_13.nand3_8.Z.t2 Vdd.t713 pfet_03v3
**devattr s=26000,604 d=26000,604
X85 SARlogic_0.dffrs_5.Qb.t1 Reset.t7 Vdd.t453 Vdd.t452 pfet_03v3
**devattr s=26000,604 d=44000,1176
X86 a_1167_30439 a_n389_31159.t4 Vdd.t201 Vdd.t200 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X87 SARlogic_0.dffrs_9.nand3_8.C.t1 SARlogic_0.dffrs_9.nand3_8.Z a_4501_19209 Vss.t127 nfet_03v3
**devattr s=10400,304 d=17600,576
X88 SARlogic_0.dffrs_0.nand3_8.C.t3 SARlogic_0.dffrs_0.nand3_6.C.t4 Vdd.t565 Vdd.t564 pfet_03v3
**devattr s=44000,1176 d=26000,604
X89 a_12401_19209 SARlogic_0.dffrs_11.nand3_6.C.t4 Vss.t428 Vss.t427 nfet_03v3
**devattr s=17600,576 d=10400,304
X90 a_33337_31515 a_33257_31423.t4 Vss.t529 Vss.t528 nfet_03v3
**devattr s=17600,576 d=10400,304
X91 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_13.Qb.t4 Vdd.t936 Vdd.t935 pfet_03v3
**devattr s=44000,1176 d=26000,604
X92 SARlogic_0.dffrs_3.nand3_8.C.t0 SARlogic_0.dffrs_3.nand3_8.Z.t5 a_4501_9633 Vss.t418 nfet_03v3
**devattr s=10400,304 d=17600,576
X93 a_10639_30440 a_9083_31160.t4 Vss.t608 Vss.t607 nfet_03v3
**devattr s=17600,576 d=17600,576
X94 Vdd.t529 SARlogic_0.dffrs_5.nand3_8.C.t6 SARlogic_0.dffrs_5.Qb.t3 Vdd.t528 pfet_03v3
**devattr s=26000,604 d=26000,604
X95 Vss.t131 a_29583_30440 a_30255_29264.t0 Vss.t130 nfet_03v3
**devattr s=17600,576 d=17600,576
X96 Vss.t389 adc_PISO_0.2inmux_1.Bit.t5 a_37687_30440 Vss.t388 nfet_03v3
**devattr s=10400,304 d=17600,576
X97 SARlogic_0.dffrs_8.nand3_6.C.t2 SARlogic_0.d2.t5 Vdd.t293 Vdd.t292 pfet_03v3
**devattr s=26000,604 d=44000,1176
X98 Vdd.t97 a_n1095_29019 a_n389_28819.t0 Vdd.t96 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X99 Vss.t636 a_1167_30439 a_1839_29263.t3 Vss.t635 nfet_03v3
**devattr s=17600,576 d=17600,576
X100 a_5987_9634 SARlogic_0.dffrs_3.nand3_8.C.t4 a_5803_9634 Vss.t77 nfet_03v3
**devattr s=10400,304 d=10400,304
X101 SARlogic_0.dffrs_0.nand3_6.C.t3 SARlogic_0.dffrs_0.nand3_1.C.t4 Vdd.t597 Vdd.t596 pfet_03v3
**devattr s=44000,1176 d=26000,604
X102 SARlogic_0.dffrs_5.nand3_1.C.t3 Vdd.t709 Vdd.t711 Vdd.t710 pfet_03v3
**devattr s=44000,1176 d=26000,604
X103 SARlogic_0.dffrs_3.nand3_1.C.t2 SARlogic_0.dffrs_3.nand3_6.C.t5 Vdd.t435 Vdd.t434 pfet_03v3
**devattr s=26000,604 d=44000,1176
X104 a_20971_29984 a_20111_28100 a_20783_29264.t2 Vdd.t135 pfet_03v3
**devattr s=52800,1376 d=31200,704
X105 a_n3065_31515 adc_PISO_0.2inmux_2.Bit.t4 Vss.t24 Vss.t23 nfet_03v3
**devattr s=17600,576 d=10400,304
X106 SARlogic_0.dffrs_12.Q.t3 SARlogic_0.dffrs_12.Qb Vdd.t507 Vdd.t506 pfet_03v3
**devattr s=26000,604 d=44000,1176
X107 SARlogic_0.dffrs_12.nand3_8.Z Vss.t677 Vdd.t5 Vdd.t4 pfet_03v3
**devattr s=26000,604 d=44000,1176
X108 a_4921_30169.t0 adc_PISO_0.2inmux_2.OUT.t2 a_5105_29309 Vss.t125 nfet_03v3
**devattr s=10400,304 d=17600,576
X109 Vdd.t331 a_27321_29020 a_28027_28820.t3 Vdd.t330 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X110 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t4 Vdd.t41 Vdd.t40 pfet_03v3
**devattr s=26000,604 d=44000,1176
X111 a_n2881_31515 a_n4631_29217.t4 a_n3065_31515 Vss.t673 nfet_03v3
**devattr s=10400,304 d=10400,304
X112 a_12585_7428 Reset.t8 a_12401_7428 Vss.t352 nfet_03v3
**devattr s=10400,304 d=10400,304
X113 SARlogic_0.dffrs_10.Qb Reset.t9 a_10029_19210 Vss.t353 nfet_03v3
**devattr s=10400,304 d=17600,576
X114 a_17849_29020 inv2_0.out.t5 Vdd.t766 Vdd.t765 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X115 SARlogic_0.dffrs_3.nand3_8.Z.t1 SARlogic_0.dffrs_3.nand3_8.C.t5 Vdd.t111 Vdd.t110 pfet_03v3
**devattr s=44000,1176 d=26000,604
X116 a_4317_17004 SARlogic_0.dffrs_9.nand3_8.C.t4 Vss.t34 Vss.t33 nfet_03v3
**devattr s=17600,576 d=10400,304
X117 Vdd.t455 Reset.t10 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t454 pfet_03v3
**devattr s=26000,604 d=26000,604
X118 SARlogic_0.dffrs_7.nand3_8.C.t2 SARlogic_0.dffrs_7.nand3_6.C.t4 Vdd.t798 Vdd.t797 pfet_03v3
**devattr s=44000,1176 d=26000,604
X119 SARlogic_0.d3.t1 SARlogic_0.dffrs_8.Qb Vdd.t241 Vdd.t240 pfet_03v3
**devattr s=26000,604 d=44000,1176
X120 Vdd.t279 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t2 Vdd.t278 pfet_03v3
**devattr s=10400,304 d=10400,304
X121 a_14393_30170.t1 adc_PISO_0.2inmux_3.OUT.t2 Vdd.t884 Vdd.t883 pfet_03v3
**devattr s=26000,604 d=44000,1176
X122 Vdd.t43 SARlogic_0.dffrs_8.nand3_6.C.t5 SARlogic_0.d3.t0 Vdd.t42 pfet_03v3
**devattr s=26000,604 d=26000,604
X123 a_4317_19209 SARlogic_0.dffrs_9.nand3_6.C.t5 Vss.t658 Vss.t657 nfet_03v3
**devattr s=17600,576 d=10400,304
X124 a_459_7428 Reset.t11 a_275_7428 Vss.t354 nfet_03v3
**devattr s=10400,304 d=10400,304
X125 a_n9429_n2007.t1 Vin2.t0 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t178 nfet_03v3
**devattr s=15600,404 d=15600,404
X126 Vdd.t67 Clk.t2 SARlogic_0.dffrs_5.nand3_8.C.t0 Vdd.t66 pfet_03v3
**devattr s=26000,604 d=26000,604
X127 a_33257_31423.t2 Clk_piso.t0 Vdd.t852 Vdd.t851 pfet_03v3
**devattr s=26000,604 d=44000,1176
X128 adc_PISO_0.2inmux_1.Bit.t1 Vdd.t706 Vdd.t708 Vdd.t707 pfet_03v3
**devattr s=44000,1176 d=26000,604
X129 SARlogic_0.dffrs_8.nand3_6.C.t3 SARlogic_0.dffrs_8.nand3_1.C Vdd.t329 Vdd.t328 pfet_03v3
**devattr s=44000,1176 d=26000,604
X130 SARlogic_0.dffrs_12.Qb Reset.t12 a_18113_19210 Vss.t355 nfet_03v3
**devattr s=10400,304 d=17600,576
X131 a_14313_29218.t1 a_14393_30170.t4 Vdd.t854 Vdd.t853 pfet_03v3
**devattr s=26000,604 d=44000,1176
X132 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t0 a_n7971_249 a_n8059_341 Vss.t303 nfet_03v3
**devattr s=35200,976 d=20800,504
X133 SARlogic_0.dffrs_3.nand3_1.C.t3 Vdd.t703 Vdd.t705 Vdd.t704 pfet_03v3
**devattr s=44000,1176 d=26000,604
X134 Vdd.t45 SARlogic_0.dffrs_9.nand3_8.C.t5 SARlogic_0.dffrs_9.Qb Vdd.t44 pfet_03v3
**devattr s=26000,604 d=26000,604
X135 SARlogic_0.dffrs_5.nand3_6.C.t0 Clk.t3 a_12585_11838 Vss.t49 nfet_03v3
**devattr s=10400,304 d=17600,576
X136 Vdd.t457 Reset.t13 SARlogic_0.dffrs_5.nand3_6.C.t1 Vdd.t456 pfet_03v3
**devattr s=26000,604 d=26000,604
X137 Vdd.t437 SARlogic_0.dffrs_3.nand3_6.C.t6 SARlogic_0.dffrs_4.d.t2 Vdd.t436 pfet_03v3
**devattr s=26000,604 d=26000,604
X138 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_8.C.t5 Vdd.t509 Vdd.t508 pfet_03v3
**devattr s=44000,1176 d=26000,604
X139 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t1 Vdd.t557 Vdd.t556 pfet_03v3
**devattr s=26000,604 d=44000,1176
X140 a_33257_33628.t1 a_33257_31423.t5 Vdd.t740 Vdd.t739 pfet_03v3
**devattr s=26000,604 d=44000,1176
X141 a_6591_31515 a_4841_29217.t4 a_6407_31515 Vss.t176 nfet_03v3
**devattr s=10400,304 d=10400,304
X142 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_1.Qb.t5 Vdd.t493 Vdd.t492 pfet_03v3
**devattr s=44000,1176 d=26000,604
X143 SARlogic_0.dffrs_14.nand3_6.C.t3 SARlogic_0.d4.t4 a_n7625_21417 Vss.t616 nfet_03v3
**devattr s=10400,304 d=17600,576
X144 a_n6323_21417 SARlogic_0.dffrs_13.Qb.t5 Vss.t669 Vss.t668 nfet_03v3
**devattr s=17600,576 d=10400,304
X145 a_13887_21414 SARlogic_0.dffrs_4.Qb.t4 Vss.t247 Vss.t246 nfet_03v3
**devattr s=17600,576 d=10400,304
X146 Vdd.t127 SARlogic_0.dffrs_10.nand3_6.C.t5 SARlogic_0.d1.t0 Vdd.t126 pfet_03v3
**devattr s=26000,604 d=26000,604
X147 Vdd.t459 Reset.t14 SARlogic_0.dffrs_12.nand3_6.C.t3 Vdd.t458 pfet_03v3
**devattr s=26000,604 d=26000,604
X148 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t1 a_n9429_n2007.t2 Vss.t179 nfet_03v3
**devattr s=15600,404 d=15600,404
X149 a_n3583_9633 Clk.t4 a_n3767_9633 Vss.t50 nfet_03v3
**devattr s=10400,304 d=10400,304
X150 a_n6139_9634 SARlogic_0.dffrs_0.nand3_8.C.t4 a_n6323_9634 Vss.t10 nfet_03v3
**devattr s=10400,304 d=10400,304
X151 SARlogic_0.dffrs_8.Qb Reset.t15 a_1945_19210 Vss.t356 nfet_03v3
**devattr s=10400,304 d=17600,576
X152 a_44295_33720 Vdd.t950 Vss.t515 Vss.t514 nfet_03v3
**devattr s=17600,576 d=10400,304
X153 a_n7445_29983 a_n8305_30439 Vdd.t165 Vdd.t164 pfet_03v3
**devattr s=52800,1376 d=31200,704
X154 a_23785_29218.t0 a_23865_30170.t4 a_24049_31515 Vss.t120 nfet_03v3
**devattr s=10400,304 d=17600,576
X155 a_1945_19210 SARlogic_0.dffrs_8.nand3_8.C.t4 a_1761_19210 Vss.t249 nfet_03v3
**devattr s=10400,304 d=10400,304
X156 a_5105_35924 a_4921_30169.t4 a_4921_35924 Vss.t216 nfet_03v3
**devattr s=10400,304 d=10400,304
X157 a_n201_30439 adc_PISO_0.2inmux_2.Bit.t5 Vss.t26 Vss.t25 nfet_03v3
**devattr s=17600,576 d=10400,304
X158 Vdd.t760 SARlogic_0.dffrs_12.nand3_8.Z SARlogic_0.dffrs_12.nand3_1.C Vdd.t759 pfet_03v3
**devattr s=26000,604 d=26000,604
X159 SARlogic_0.dffrs_7.nand3_8.C.t0 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t211 Vdd.t210 pfet_03v3
**devattr s=26000,604 d=44000,1176
X160 a_4501_11838 Reset.t16 a_4317_11838 Vss.t357 nfet_03v3
**devattr s=10400,304 d=10400,304
X161 a_42993_33720 Vdd.t951 a_42809_33720 Vss.t513 nfet_03v3
**devattr s=10400,304 d=10400,304
X162 a_4921_35924 Vdd.t952 Vss.t512 Vss.t511 nfet_03v3
**devattr s=17600,576 d=10400,304
X163 adc_PISO_0.dffrs_4.Qb adc_PISO_0.2inmux_1.Bit.t6 Vdd.t513 Vdd.t512 pfet_03v3
**devattr s=44000,1176 d=26000,604
X164 a_459_14043 SARlogic_0.dffrs_2.nand3_8.Z.t4 a_275_14043 Vss.t164 nfet_03v3
**devattr s=10400,304 d=10400,304
X165 a_28215_30440 adc_PISO_0.dffrs_3.Q.t4 Vss.t187 Vss.t186 nfet_03v3
**devattr s=17600,576 d=10400,304
X166 a_39727_29264.t2 a_39055_28100 a_39915_29984 Vdd.t389 pfet_03v3
**devattr s=31200,704 d=52800,1376
X167 a_8543_21414 Reset.t17 a_8359_21414 Vss.t358 nfet_03v3
**devattr s=10400,304 d=10400,304
X168 a_n7809_9633 SARlogic_0.dffrs_0.nand3_6.C.t5 Vss.t42 Vss.t41 nfet_03v3
**devattr s=17600,576 d=10400,304
X169 comparator_no_offsetcal_0.no_offsetLatch_0.Vq a_n9933_n2099 a_n10021_n2007 Vss.t368 nfet_03v3
**devattr s=26400,776 d=15600,404
X170 SARlogic_0.dffrs_0.nand3_1.C.t1 Vdd.t700 Vdd.t702 Vdd.t701 pfet_03v3
**devattr s=44000,1176 d=26000,604
X171 a_n7809_17007 SARlogic_0.dffrs_14.nand3_8.C.t5 Vss.t534 Vss.t533 nfet_03v3
**devattr s=17600,576 d=10400,304
X172 a_42993_35925 a_42809_30170.t4 a_42809_35925 Vss.t258 nfet_03v3
**devattr s=10400,304 d=10400,304
X173 a_33257_31423.t1 a_33257_33628.t4 Vdd.t796 Vdd.t795 pfet_03v3
**devattr s=44000,1176 d=26000,604
X174 a_28215_28100 SARlogic_0.d1.t6 a_28027_28820.t1 Vss.t584 nfet_03v3
**devattr s=17600,576 d=10400,304
X175 Vdd.t699 Vdd.t697 a_23865_30170.t2 Vdd.t698 pfet_03v3
**devattr s=26000,604 d=26000,604
X176 a_8543_23619 SARlogic_0.dffrs_10.nand3_8.Z a_8359_23619 Vss.t9 nfet_03v3
**devattr s=10400,304 d=10400,304
X177 a_10029_19210 SARlogic_0.dffrs_10.nand3_8.C.t4 a_9845_19210 Vss.t189 nfet_03v3
**devattr s=10400,304 d=10400,304
X178 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_8.C.t5 Vdd.t245 Vdd.t244 pfet_03v3
**devattr s=44000,1176 d=26000,604
X179 a_33257_33628.t3 Vdd.t694 Vdd.t696 Vdd.t695 pfet_03v3
**devattr s=44000,1176 d=26000,604
X180 Vdd.t872 Clk_piso.t1 a_23785_29218.t3 Vdd.t871 pfet_03v3
**devattr s=26000,604 d=26000,604
X181 SARlogic_0.d5.t1 SARlogic_0.dffrs_14.Qb a_n6139_21417 Vss.t157 nfet_03v3
**devattr s=10400,304 d=17600,576
X182 a_44295_31516 Piso_out.t4 Vss.t15 Vss.t14 nfet_03v3
**devattr s=17600,576 d=10400,304
X183 a_n4367_35924 a_n4551_30169.t4 a_n4551_35924 Vss.t648 nfet_03v3
**devattr s=10400,304 d=10400,304
X184 a_n4551_30169.t0 a_n4631_29217.t5 Vdd.t942 Vdd.t941 pfet_03v3
**devattr s=44000,1176 d=26000,604
X185 a_12585_17004 Reset.t18 a_12401_17004 Vss.t359 nfet_03v3
**devattr s=10400,304 d=10400,304
X186 a_8377_29020 inv2_0.out.t6 Vss.t553 Vss.t552 nfet_03v3
**devattr s=17600,576 d=17600,576
X187 SARlogic_0.dffrs_0.nand3_8.Z.t3 SARlogic_0.dffrs_0.d.t5 Vdd.t824 Vdd.t823 pfet_03v3
**devattr s=26000,604 d=44000,1176
X188 a_14393_29310 a_14313_29218.t4 Vss.t675 Vss.t674 nfet_03v3
**devattr s=17600,576 d=10400,304
X189 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t2 Vdd.t559 Vdd.t558 pfet_03v3
**devattr s=26000,604 d=44000,1176
X190 a_12585_19209 SARlogic_0.dffrs_12.Q.t4 a_12401_19209 Vss.t406 nfet_03v3
**devattr s=10400,304 d=10400,304
X191 a_39727_29264.t0 a_39055_28100 Vss.t302 Vss.t301 nfet_03v3
**devattr s=17600,576 d=17600,576
X192 a_11499_29984 a_10639_28100 a_11311_29264.t2 Vdd.t595 pfet_03v3
**devattr s=52800,1376 d=31200,704
X193 a_n6555_341 a_n6755_249 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t177 nfet_03v3
**devattr s=20800,504 d=35200,976
X194 Vdd.t147 SARlogic_0.dffrs_5.nand3_8.Z.t4 SARlogic_0.dffrs_5.nand3_1.C.t2 Vdd.t146 pfet_03v3
**devattr s=26000,604 d=26000,604
X195 a_n10151_9634 SARlogic_0.dffrs_13.nand3_8.C.t4 a_n10335_9634 Vss.t634 nfet_03v3
**devattr s=10400,304 d=10400,304
X196 SARlogic_0.d2.t1 SARlogic_0.dffrs_9.Qb Vdd.t89 Vdd.t88 pfet_03v3
**devattr s=26000,604 d=44000,1176
X197 adc_PISO_0.2inmux_1.Bit.t2 adc_PISO_0.dffrs_4.Qb a_35007_33720 Vss.t660 nfet_03v3
**devattr s=10400,304 d=17600,576
X198 adc_PISO_0.2inmux_0.OUT.t1 a_n7633_29263.t4 Vdd.t171 Vdd.t170 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X199 SARlogic_0.d4.t3 SARlogic_0.dffrs_0.Qb.t4 Vdd.t195 Vdd.t194 pfet_03v3
**devattr s=44000,1176 d=26000,604
X200 SARlogic_0.dffrs_0.nand3_8.C.t1 SARlogic_0.dffrs_0.nand3_8.Z.t4 Vdd.t149 Vdd.t148 pfet_03v3
**devattr s=26000,604 d=44000,1176
X201 a_36793_29020 inv2_0.out.t7 Vdd.t768 Vdd.t767 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X202 Vdd.t393 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t7 Vdd.t392 pfet_03v3
**devattr s=10400,304 d=10400,304
X203 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t5 Vdd.t485 Vdd.t484 pfet_03v3
**devattr s=26000,604 d=44000,1176
X204 SARlogic_0.dffrs_5.nand3_8.Z.t1 SARlogic_0.dffrs_4.Q.t4 Vdd.t137 Vdd.t136 pfet_03v3
**devattr s=26000,604 d=44000,1176
X205 a_n9429_n2007.t3 Vin2.t2 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t180 nfet_03v3
**devattr s=15600,404 d=15600,404
X206 SARlogic_0.dffrs_0.nand3_6.C.t2 Clk.t5 Vdd.t69 Vdd.t68 pfet_03v3
**devattr s=26000,604 d=44000,1176
X207 a_n4551_30169.t1 adc_PISO_0.2inmux_0.OUT.t2 Vdd.t141 Vdd.t140 pfet_03v3
**devattr s=26000,604 d=44000,1176
X208 SARlogic_0.dffrs_0.Q.t0 Vdd.t691 Vdd.t693 Vdd.t692 pfet_03v3
**devattr s=44000,1176 d=26000,604
X209 adc_PISO_0.dffrs_3.Q.t2 Vdd.t688 Vdd.t690 Vdd.t689 pfet_03v3
**devattr s=44000,1176 d=26000,604
X210 a_18555_28820.t1 SARlogic_0.d2.t6 Vdd.t295 Vdd.t294 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X211 a_18113_21414 SARlogic_0.dffrs_12.nand3_6.C.t5 a_17929_21414 Vss.t661 nfet_03v3
**devattr s=10400,304 d=10400,304
X212 a_23785_31423.t3 Clk_piso.t2 Vdd.t874 Vdd.t873 pfet_03v3
**devattr s=26000,604 d=44000,1176
X213 SARlogic_0.dffrs_13.nand3_8.Z.t1 Vss.t109 a_n11637_7428 Vss.t110 nfet_03v3
**devattr s=10400,304 d=17600,576
X214 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t243 Vdd.t242 pfet_03v3
**devattr s=17600,576 d=17600,576
X215 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_8.C.t5 Vdd.t311 Vdd.t310 pfet_03v3
**devattr s=44000,1176 d=26000,604
X216 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x3.out Vss.t163 Vss.t162 nfet_03v3
**devattr s=17600,576 d=17600,576
X217 SARlogic_0.dffrs_12.nand3_6.C.t1 Vss.t107 a_16627_21414 Vss.t108 nfet_03v3
**devattr s=10400,304 d=17600,576
X218 a_n3767_9633 SARlogic_0.dffrs_1.nand3_6.C.t4 Vss.t218 Vss.t217 nfet_03v3
**devattr s=17600,576 d=10400,304
X219 Vdd.t742 a_33257_31423.t6 adc_PISO_0.2inmux_1.Bit.t0 Vdd.t741 pfet_03v3
**devattr s=26000,604 d=26000,604
X220 SARlogic_0.dffrs_9.Qb Reset.t19 a_5987_19210 Vss.t360 nfet_03v3
**devattr s=10400,304 d=17600,576
X221 a_23785_33628.t3 a_23785_31423.t5 Vdd.t866 Vdd.t865 pfet_03v3
**devattr s=26000,604 d=44000,1176
X222 Vdd.t461 Reset.t20 SARlogic_0.dffrs_8.nand3_6.C.t0 Vdd.t460 pfet_03v3
**devattr s=26000,604 d=26000,604
X223 SARlogic_0.dffrs_14.Qb SARlogic_0.d5.t4 Vdd.t121 Vdd.t120 pfet_03v3
**devattr s=44000,1176 d=26000,604
X224 a_n2281_19210 SARlogic_0.d4.t5 Vss.t172 Vss.t171 nfet_03v3
**devattr s=17600,576 d=10400,304
X225 a_n3583_14043 SARlogic_0.dffrs_1.nand3_8.Z.t4 a_n3767_14043 Vss.t13 nfet_03v3
**devattr s=10400,304 d=10400,304
X226 a_n7633_29263.t3 a_n8305_28099 a_n7445_29983 Vdd.t303 pfet_03v3
**devattr s=31200,704 d=52800,1376
X227 SARlogic_0.dffrs_2.nand3_8.Z.t0 SARlogic_0.dffrs_2.d.t4 Vdd.t31 Vdd.t30 pfet_03v3
**devattr s=26000,604 d=44000,1176
X228 SARlogic_0.dffrs_12.nand3_1.C SARlogic_0.dffrs_12.nand3_6.C.t6 a_16627_23619 Vss.t662 nfet_03v3
**devattr s=10400,304 d=17600,576
X229 SARlogic_0.dffrs_11.Qb SARlogic_0.d0.t5 Vdd.t261 Vdd.t260 pfet_03v3
**devattr s=44000,1176 d=26000,604
X230 adc_PISO_0.dffrs_4.Qb Vdd.t953 a_35007_31516 Vss.t510 nfet_03v3
**devattr s=10400,304 d=17600,576
X231 SARlogic_0.dffrs_5.Q.t3 Vdd.t685 Vdd.t687 Vdd.t686 pfet_03v3
**devattr s=44000,1176 d=26000,604
X232 Vdd.t463 Reset.t21 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t462 pfet_03v3
**devattr s=26000,604 d=26000,604
X233 a_n389_31159.t3 inv2_0.out.t8 Vdd.t770 Vdd.t769 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X234 a_n7625_21417 Reset.t22 a_n7809_21417 Vss.t361 nfet_03v3
**devattr s=10400,304 d=10400,304
X235 Vdd.t317 SARlogic_0.dffrs_8.nand3_8.Z SARlogic_0.dffrs_8.nand3_1.C Vdd.t316 pfet_03v3
**devattr s=26000,604 d=26000,604
X236 adc_PISO_0.dffrs_0.Qb Vdd.t954 a_n2881_31515 Vss.t509 nfet_03v3
**devattr s=10400,304 d=17600,576
X237 a_1761_21414 SARlogic_0.dffrs_1.Qb.t6 Vss.t376 Vss.t375 nfet_03v3
**devattr s=17600,576 d=10400,304
X238 a_n10567_29019 inv2_0.out.t9 Vss.t555 Vss.t554 nfet_03v3
**devattr s=17600,576 d=17600,576
X239 a_n201_28099 SARlogic_0.d4.t6 a_n389_28819.t1 Vss.t173 nfet_03v3
**devattr s=17600,576 d=10400,304
X240 SARlogic_0.dffrs_12.Q.t1 SARlogic_0.dffrs_5.Qb.t5 Vdd.t429 Vdd.t428 pfet_03v3
**devattr s=44000,1176 d=26000,604
X241 a_n11821_14043 Reset.t23 Vss.t363 Vss.t362 nfet_03v3
**devattr s=17600,576 d=10400,304
X242 a_33521_33720 Vdd.t955 a_33337_33720 Vss.t508 nfet_03v3
**devattr s=10400,304 d=10400,304
X243 Vdd.t71 Clk.t6 SARlogic_0.dffrs_4.nand3_8.C.t2 Vdd.t70 pfet_03v3
**devattr s=26000,604 d=26000,604
X244 SARlogic_0.dffrs_1.nand3_8.Z.t2 SARlogic_0.dffrs_0.Q.t4 Vdd.t944 Vdd.t943 pfet_03v3
**devattr s=26000,604 d=44000,1176
X245 SARlogic_0.dffrs_0.Q.t2 SARlogic_0.dffrs_0.Qb.t5 Vdd.t197 Vdd.t196 pfet_03v3
**devattr s=26000,604 d=44000,1176
X246 adc_PISO_0.dffrs_3.Qb adc_PISO_0.dffrs_3.Q.t5 Vdd.t253 Vdd.t252 pfet_03v3
**devattr s=44000,1176 d=26000,604
X247 a_30255_29264.t3 a_29583_28100 a_30443_29984 Vdd.t301 pfet_03v3
**devattr s=31200,704 d=52800,1376
X248 a_5803_11838 Vdd.t956 Vss.t507 Vss.t506 nfet_03v3
**devattr s=17600,576 d=10400,304
X249 a_4841_33627.t2 a_4841_31422.t5 a_5105_35924 Vss.t275 nfet_03v3
**devattr s=10400,304 d=17600,576
X250 a_1839_29263.t2 a_1167_28099 a_2027_29983 Vdd.t299 pfet_03v3
**devattr s=31200,704 d=52800,1376
X251 a_12401_11838 SARlogic_0.dffrs_5.nand3_1.C.t5 Vss.t387 Vss.t386 nfet_03v3
**devattr s=17600,576 d=10400,304
X252 SARlogic_0.dffrs_3.nand3_6.C.t1 Clk.t7 a_4501_11838 Vss.t51 nfet_03v3
**devattr s=10400,304 d=17600,576
X253 Vdd.t465 Reset.t24 SARlogic_0.dffrs_4.nand3_6.C.t0 Vdd.t464 pfet_03v3
**devattr s=26000,604 d=26000,604
X254 a_33521_35925 a_33337_30170.t6 a_33337_35925 Vss.t590 nfet_03v3
**devattr s=10400,304 d=10400,304
X255 a_42809_30170.t2 adc_PISO_0.2inmux_1.OUT.t2 Vdd.t838 Vdd.t837 pfet_03v3
**devattr s=26000,604 d=44000,1176
X256 inv2_0.out.t0 Load.t0 Vss.t1 Vss.t0 nfet_03v3
**devattr s=17600,576 d=17600,576
X257 Vdd.t684 Vdd.t682 a_14393_30170.t3 Vdd.t683 pfet_03v3
**devattr s=26000,604 d=26000,604
X258 Comp_out.t3 a_n10831_4320 Vss.t572 Vss.t571 nfet_03v3
**devattr s=17000,540 d=9350,280
X259 Vdd.t185 a_33257_29218.t4 adc_PISO_0.dffrs_4.Qb Vdd.t184 pfet_03v3
**devattr s=26000,604 d=26000,604
X260 SARlogic_0.dffrs_11.nand3_8.C.t1 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t175 Vdd.t174 pfet_03v3
**devattr s=26000,604 d=44000,1176
X261 SARlogic_0.dffrs_10.nand3_6.C.t2 SARlogic_0.d0.t6 a_8543_21414 Vss.t202 nfet_03v3
**devattr s=10400,304 d=17600,576
X262 a_9845_21414 SARlogic_0.dffrs_3.Qb.t6 Vss.t308 Vss.t307 nfet_03v3
**devattr s=17600,576 d=10400,304
X263 a_16443_21414 SARlogic_0.dffrs_12.nand3_1.C Vss.t68 Vss.t67 nfet_03v3
**devattr s=17600,576 d=10400,304
X264 a_42729_29218.t2 a_42809_30170.t5 Vdd.t325 Vdd.t324 pfet_03v3
**devattr s=26000,604 d=44000,1176
X265 a_8359_7428 SARlogic_0.dffrs_4.nand3_8.C.t6 Vss.t398 Vss.t397 nfet_03v3
**devattr s=17600,576 d=10400,304
X266 Vdd.t876 Clk_piso.t3 a_14313_29218.t3 Vdd.t875 pfet_03v3
**devattr s=26000,604 d=26000,604
X267 SARlogic_0.dffrs_14.Qb Reset.t25 Vdd.t467 Vdd.t466 pfet_03v3
**devattr s=26000,604 d=44000,1176
X268 inv2_0.out.t1 Load.t1 Vdd.t850 Vdd.t849 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X269 SARlogic_0.dffrs_10.nand3_1.C SARlogic_0.dffrs_10.nand3_6.C.t6 a_8543_23619 Vss.t88 nfet_03v3
**devattr s=10400,304 d=17600,576
X270 a_16443_23619 SARlogic_0.dffrs_5.Qb.t6 Vss.t326 Vss.t325 nfet_03v3
**devattr s=17600,576 d=10400,304
X271 a_17929_19210 SARlogic_0.dffrs_12.Q.t5 Vss.t408 Vss.t407 nfet_03v3
**devattr s=17600,576 d=10400,304
X272 a_n9429_n2007.t4 Vin2.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t181 nfet_03v3
**devattr s=15600,404 d=15600,404
X273 a_6407_31515 adc_PISO_0.dffrs_1.Q.t5 Vss.t209 Vss.t208 nfet_03v3
**devattr s=17600,576 d=10400,304
X274 a_18555_31160.t2 inv2_0.out.t10 a_18743_30440 Vss.t556 nfet_03v3
**devattr s=10400,304 d=17600,576
X275 Vdd.t806 SARlogic_0.d1.t7 SARlogic_0.dffrs_9.nand3_8.C.t0 Vdd.t805 pfet_03v3
**devattr s=26000,604 d=26000,604
X276 Vdd.t469 Reset.t26 SARlogic_0.dffrs_0.nand3_8.Z.t0 Vdd.t468 pfet_03v3
**devattr s=26000,604 d=26000,604
X277 a_n6139_21417 SARlogic_0.dffrs_14.nand3_6.C.t6 a_n6323_21417 Vss.t370 nfet_03v3
**devattr s=10400,304 d=10400,304
X278 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t11 Vss.t305 Vss.t304 nfet_03v3
**devattr s=35200,976 d=35200,976
X279 SARlogic_0.dffrs_13.nand3_1.C.t2 SARlogic_0.dffrs_13.nand3_6.C.t4 a_n11637_14043 Vss.t597 nfet_03v3
**devattr s=10400,304 d=17600,576
X280 SARlogic_0.dffrs_0.nand3_1.C.t3 SARlogic_0.dffrs_0.nand3_6.C.t6 Vdd.t57 Vdd.t56 pfet_03v3
**devattr s=26000,604 d=44000,1176
X281 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t3 a_n7625_17007 Vss.t424 nfet_03v3
**devattr s=10400,304 d=17600,576
X282 adc_PISO_0.2inmux_5.OUT.t1 a_30255_29264.t5 Vdd.t257 Vdd.t256 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X283 a_n10335_9634 SARlogic_0.dffrs_0.d.t6 Vss.t592 Vss.t591 nfet_03v3
**devattr s=17600,576 d=10400,304
X284 a_42809_33720 a_42729_33628.t5 Vss.t93 Vss.t92 nfet_03v3
**devattr s=17600,576 d=10400,304
X285 Vdd.t681 Vdd.t679 a_4921_30169.t3 Vdd.t680 pfet_03v3
**devattr s=26000,604 d=26000,604
X286 a_4317_11838 SARlogic_0.dffrs_3.nand3_1.C.t5 Vss.t148 Vss.t147 nfet_03v3
**devattr s=17600,576 d=10400,304
X287 a_23865_31515 a_23785_31423.t6 Vss.t621 Vss.t620 nfet_03v3
**devattr s=17600,576 d=10400,304
X288 a_4921_30169.t2 a_4841_29217.t5 Vdd.t225 Vdd.t224 pfet_03v3
**devattr s=44000,1176 d=26000,604
X289 a_42993_29310 Vdd.t957 a_42809_29310 Vss.t505 nfet_03v3
**devattr s=10400,304 d=10400,304
X290 Vss.t66 a_20111_30440 a_20783_29264.t0 Vss.t65 nfet_03v3
**devattr s=17600,576 d=17600,576
X291 a_8359_21414 SARlogic_0.dffrs_10.nand3_1.C Vss.t76 Vss.t75 nfet_03v3
**devattr s=17600,576 d=10400,304
X292 a_42809_35925 Vdd.t958 Vss.t504 Vss.t503 nfet_03v3
**devattr s=17600,576 d=10400,304
X293 a_n9673_28099 a_n10567_29019 Vss.t653 Vss.t652 nfet_03v3
**devattr s=17600,576 d=10400,304
X294 a_8543_17004 Reset.t27 a_8359_17004 Vss.t364 nfet_03v3
**devattr s=10400,304 d=10400,304
X295 SARlogic_0.d1.t2 SARlogic_0.dffrs_10.Qb a_10029_21414 Vss.t535 nfet_03v3
**devattr s=10400,304 d=17600,576
X296 a_8359_23619 SARlogic_0.dffrs_3.Qb.t7 Vss.t310 Vss.t309 nfet_03v3
**devattr s=17600,576 d=10400,304
X297 a_n11637_7428 Vdd.t959 a_n11821_7428 Vss.t502 nfet_03v3
**devattr s=10400,304 d=10400,304
X298 Vdd.t107 a_17849_29020 a_18555_28820.t0 Vdd.t106 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X299 Vdd.t471 Reset.t28 SARlogic_0.dffrs_7.nand3_6.C.t0 Vdd.t470 pfet_03v3
**devattr s=26000,604 d=26000,604
X300 Vdd.t73 Clk.t8 SARlogic_0.dffrs_0.nand3_8.C.t0 Vdd.t72 pfet_03v3
**devattr s=26000,604 d=26000,604
X301 a_n201_30439 inv2_0.out.t11 a_n389_31159.t2 Vss.t557 nfet_03v3
**devattr s=17600,576 d=10400,304
X302 a_20111_28100 a_18555_28820.t4 Vss.t575 Vss.t574 nfet_03v3
**devattr s=17600,576 d=17600,576
X303 a_8543_19209 SARlogic_0.d0.t7 a_8359_19209 Vss.t203 nfet_03v3
**devattr s=10400,304 d=10400,304
X304 Vdd.t912 a_n10567_29019 a_n9861_28819.t3 Vdd.t911 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X305 Vdd.t207 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_1.C Vdd.t206 pfet_03v3
**devattr s=26000,604 d=26000,604
X306 a_n7809_23622 SARlogic_0.dffrs_13.Qb.t6 Vss.t671 Vss.t670 nfet_03v3
**devattr s=17600,576 d=10400,304
X307 Vss.t211 adc_PISO_0.dffrs_1.Q.t6 a_9271_30440 Vss.t210 nfet_03v3
**devattr s=10400,304 d=17600,576
X308 a_37499_28820.t2 SARlogic_0.d0.t8 a_37687_28100 Vss.t204 nfet_03v3
**devattr s=10400,304 d=17600,576
X309 Vdd.t209 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_1.C Vdd.t208 pfet_03v3
**devattr s=26000,604 d=26000,604
X310 SARlogic_0.dffrs_8.nand3_6.C.t1 SARlogic_0.d2.t7 a_459_21414 Vss.t230 nfet_03v3
**devattr s=10400,304 d=17600,576
X311 Vdd.t3 SARlogic_0.dffrs_12.nand3_8.C.t6 SARlogic_0.dffrs_12.Qb Vdd.t2 pfet_03v3
**devattr s=26000,604 d=26000,604
X312 Vdd.t678 Vdd.t676 a_n4551_30169.t2 Vdd.t677 pfet_03v3
**devattr s=26000,604 d=26000,604
X313 a_12401_9633 SARlogic_0.dffrs_5.nand3_6.C.t5 Vss.t537 Vss.t536 nfet_03v3
**devattr s=17600,576 d=10400,304
X314 a_n7809_11838 SARlogic_0.dffrs_0.nand3_1.C.t5 Vss.t452 Vss.t451 nfet_03v3
**devattr s=17600,576 d=10400,304
X315 Vdd.t473 Reset.t29 SARlogic_0.dffrs_0.nand3_6.C.t0 Vdd.t472 pfet_03v3
**devattr s=26000,604 d=26000,604
X316 Vdd.t439 SARlogic_0.dffrs_4.nand3_8.Z.t5 SARlogic_0.dffrs_4.nand3_1.C.t0 Vdd.t438 pfet_03v3
**devattr s=26000,604 d=26000,604
X317 a_1761_9634 SARlogic_0.dffrs_2.Q.t4 Vss.t270 Vss.t269 nfet_03v3
**devattr s=17600,576 d=10400,304
X318 Vdd.t868 a_23785_31423.t7 adc_PISO_0.dffrs_3.Q.t3 Vdd.t867 pfet_03v3
**devattr s=26000,604 d=26000,604
X319 SARlogic_0.dffrs_12.Q.t2 SARlogic_0.dffrs_12.Qb a_18113_21414 Vss.t385 nfet_03v3
**devattr s=10400,304 d=17600,576
X320 SARlogic_0.dffrs_8.nand3_1.C SARlogic_0.dffrs_8.nand3_6.C.t6 a_459_23619 Vss.t29 nfet_03v3
**devattr s=10400,304 d=17600,576
X321 Vdd.t475 Reset.t30 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t474 pfet_03v3
**devattr s=26000,604 d=26000,604
X322 Vdd.t75 Clk.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vdd.t74 pfet_03v3
**devattr s=14080,496 d=14080,496
X323 a_275_9633 SARlogic_0.dffrs_2.nand3_6.C.t5 Vss.t383 Vss.t382 nfet_03v3
**devattr s=17600,576 d=10400,304
X324 adc_PISO_0.dffrs_1.Q.t1 adc_PISO_0.dffrs_1.Qb Vdd.t35 Vdd.t34 pfet_03v3
**devattr s=26000,604 d=44000,1176
X325 a_4317_7428 SARlogic_0.dffrs_3.nand3_8.C.t6 Vss.t79 Vss.t78 nfet_03v3
**devattr s=17600,576 d=10400,304
X326 a_n3767_14043 Vdd.t960 Vss.t501 Vss.t500 nfet_03v3
**devattr s=17600,576 d=10400,304
X327 SARlogic_0.dffrs_8.Qb SARlogic_0.d3.t7 Vdd.t898 Vdd.t897 pfet_03v3
**devattr s=44000,1176 d=26000,604
X328 a_30443_29984 a_29583_30440 Vdd.t169 Vdd.t168 pfet_03v3
**devattr s=52800,1376 d=31200,704
X329 SARlogic_0.dffrs_2.Q.t0 Vdd.t673 Vdd.t675 Vdd.t674 pfet_03v3
**devattr s=44000,1176 d=26000,604
X330 SARlogic_0.d3.t2 SARlogic_0.dffrs_8.Qb a_1945_21414 Vss.t188 nfet_03v3
**devattr s=10400,304 d=17600,576
X331 a_2027_29983 a_1167_30439 Vdd.t890 Vdd.t889 pfet_03v3
**devattr s=52800,1376 d=31200,704
X332 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t15 Vin1.t1 a_n9429_n2007.t17 Vss.t179 nfet_03v3
**devattr s=15600,404 d=15600,404
X333 a_9271_30440 inv2_0.out.t12 a_9083_31160.t2 Vss.t558 nfet_03v3
**devattr s=17600,576 d=10400,304
X334 a_39055_28100 a_37499_28820.t4 Vss.t612 Vss.t611 nfet_03v3
**devattr s=17600,576 d=17600,576
X335 Vdd.t800 SARlogic_0.dffrs_7.nand3_6.C.t5 SARlogic_0.d4.t0 Vdd.t799 pfet_03v3
**devattr s=26000,604 d=26000,604
X336 comparator_no_offsetcal_0.no_offsetLatch_0.Vq comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t4 Vss.t306 nfet_03v3
**devattr s=20800,504 d=20800,504
X337 a_n7633_29263.t1 a_n8305_28099 Vss.t241 Vss.t240 nfet_03v3
**devattr s=17600,576 d=17600,576
X338 a_1945_21414 SARlogic_0.dffrs_8.nand3_6.C.t7 a_1761_21414 Vss.t30 nfet_03v3
**devattr s=10400,304 d=10400,304
X339 SARlogic_0.dffrs_3.Qb.t2 SARlogic_0.dffrs_4.d.t5 Vdd.t814 Vdd.t813 pfet_03v3
**devattr s=44000,1176 d=26000,604
X340 a_33257_31423.t3 Clk_piso.t4 a_33521_33720 Vss.t629 nfet_03v3
**devattr s=10400,304 d=17600,576
X341 a_34823_33720 Vdd.t961 Vss.t499 Vss.t498 nfet_03v3
**devattr s=17600,576 d=10400,304
X342 SARlogic_0.d4.t2 SARlogic_0.dffrs_7.Qb Vdd.t541 Vdd.t540 pfet_03v3
**devattr s=26000,604 d=44000,1176
X343 SARlogic_0.dffrs_4.nand3_8.C.t1 SARlogic_0.dffrs_4.nand3_8.Z.t6 Vdd.t441 Vdd.t440 pfet_03v3
**devattr s=26000,604 d=44000,1176
X344 a_14313_29218.t0 a_14393_30170.t5 a_14577_31515 Vss.t609 nfet_03v3
**devattr s=10400,304 d=17600,576
X345 a_275_21414 SARlogic_0.dffrs_8.nand3_1.C Vss.t261 Vss.t260 nfet_03v3
**devattr s=17600,576 d=10400,304
X346 a_9083_31160.t1 inv2_0.out.t13 Vdd.t772 Vdd.t771 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X347 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t10 Vdd.t281 Vdd.t280 pfet_03v3
**devattr s=10400,304 d=10400,304
X348 Vdd.t59 SARlogic_0.dffrs_0.nand3_6.C.t7 SARlogic_0.dffrs_0.Q.t3 Vdd.t58 pfet_03v3
**devattr s=26000,604 d=26000,604
X349 Vdd.t183 a_23785_29218.t5 adc_PISO_0.dffrs_3.Qb Vdd.t182 pfet_03v3
**devattr s=26000,604 d=26000,604
X350 SARlogic_0.dffrs_10.Qb SARlogic_0.d1.t8 Vdd.t808 Vdd.t807 pfet_03v3
**devattr s=44000,1176 d=26000,604
X351 a_5987_11838 SARlogic_0.dffrs_3.nand3_6.C.t7 a_5803_11838 Vss.t330 nfet_03v3
**devattr s=10400,304 d=10400,304
X352 a_n1095_29019 inv2_0.out.t14 Vss.t560 Vss.t559 nfet_03v3
**devattr s=17600,576 d=17600,576
X353 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vss.t257 Vss.t256 nfet_03v3
**devattr s=9350,280 d=17000,540
X354 a_12585_11838 Reset.t31 a_12401_11838 Vss.t365 nfet_03v3
**devattr s=10400,304 d=10400,304
X355 SARlogic_0.dffrs_4.Q.t2 Vdd.t670 Vdd.t672 Vdd.t671 pfet_03v3
**devattr s=44000,1176 d=26000,604
X356 SARlogic_0.dffrs_4.nand3_6.C.t3 Clk.t10 Vdd.t77 Vdd.t76 pfet_03v3
**devattr s=26000,604 d=44000,1176
X357 a_33257_33628.t0 a_33257_31423.t7 a_33521_35925 Vss.t530 nfet_03v3
**devattr s=10400,304 d=17600,576
X358 a_18743_30440 adc_PISO_0.dffrs_2.Q.t4 Vss.t286 Vss.t285 nfet_03v3
**devattr s=17600,576 d=10400,304
X359 a_275_23619 SARlogic_0.dffrs_1.Qb.t7 Vss.t378 Vss.t377 nfet_03v3
**devattr s=17600,576 d=10400,304
X360 a_n6389_n1044 a_n6589_n1136 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t156 nfet_03v3
**devattr s=15600,404 d=26400,776
X361 a_23785_31423.t0 a_23785_33628.t4 Vdd.t95 Vdd.t94 pfet_03v3
**devattr s=44000,1176 d=26000,604
X362 a_28027_31160.t3 inv2_0.out.t15 Vdd.t774 Vdd.t773 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X363 a_10029_21414 SARlogic_0.dffrs_10.nand3_6.C.t7 a_9845_21414 Vss.t89 nfet_03v3
**devattr s=10400,304 d=10400,304
X364 a_16627_21414 Reset.t32 a_16443_21414 Vss.t366 nfet_03v3
**devattr s=10400,304 d=10400,304
X365 a_n9673_30439 Vss.t104 Vss.t106 Vss.t105 nfet_03v3
**devattr s=17600,576 d=10400,304
X366 Vdd.t746 SARlogic_0.dffrs_14.nand3_8.C.t6 SARlogic_0.dffrs_14.Qb Vdd.t745 pfet_03v3
**devattr s=26000,604 d=26000,604
X367 a_n2097_19210 SARlogic_0.dffrs_7.nand3_8.C.t4 a_n2281_19210 Vss.t60 nfet_03v3
**devattr s=10400,304 d=10400,304
X368 SARlogic_0.dffrs_1.nand3_1.C.t0 SARlogic_0.dffrs_1.nand3_6.C.t5 a_n3583_14043 Vss.t219 nfet_03v3
**devattr s=10400,304 d=17600,576
X369 SARlogic_0.dffrs_12.nand3_8.Z Vss.t102 a_16627_17004 Vss.t103 nfet_03v3
**devattr s=10400,304 d=17600,576
X370 a_23785_33628.t0 Vdd.t667 Vdd.t669 Vdd.t668 pfet_03v3
**devattr s=44000,1176 d=26000,604
X371 a_1839_29263.t0 a_1167_28099 Vss.t237 Vss.t236 nfet_03v3
**devattr s=17600,576 d=17600,576
X372 adc_PISO_0.2inmux_4.OUT.t0 a_20783_29264.t4 Vss.t150 Vss.t149 nfet_03v3
**devattr s=17600,576 d=17600,576
X373 a_16627_23619 SARlogic_0.dffrs_12.nand3_8.Z a_16443_23619 Vss.t546 nfet_03v3
**devattr s=10400,304 d=10400,304
X374 SARlogic_0.dffrs_7.Qb Reset.t33 a_n2097_19210 Vss.t367 nfet_03v3
**devattr s=10400,304 d=17600,576
X375 SARlogic_0.dffrs_9.nand3_8.C.t2 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t161 Vdd.t160 pfet_03v3
**devattr s=26000,604 d=44000,1176
X376 SARlogic_0.dffrs_11.nand3_8.C.t3 SARlogic_0.dffrs_11.nand3_6.C.t5 Vdd.t569 Vdd.t568 pfet_03v3
**devattr s=44000,1176 d=26000,604
X377 Vdd.t359 Reset.t34 SARlogic_0.dffrs_4.nand3_8.Z.t0 Vdd.t358 pfet_03v3
**devattr s=26000,604 d=26000,604
X378 a_34823_31516 adc_PISO_0.2inmux_1.Bit.t7 Vss.t391 Vss.t390 nfet_03v3
**devattr s=17600,576 d=10400,304
X379 a_9271_28100 a_8377_29020 Vss.t541 Vss.t540 nfet_03v3
**devattr s=17600,576 d=10400,304
X380 SARlogic_0.dffrs_12.nand3_8.C.t2 SARlogic_0.dffrs_12.nand3_8.Z a_16627_19209 Vss.t545 nfet_03v3
**devattr s=10400,304 d=17600,576
X381 Vdd.t151 SARlogic_0.dffrs_0.nand3_8.Z.t5 SARlogic_0.dffrs_0.nand3_1.C.t0 Vdd.t150 pfet_03v3
**devattr s=26000,604 d=26000,604
X382 a_10639_30440 a_9083_31160.t5 Vdd.t848 Vdd.t847 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X383 a_27321_29020 inv2_0.out.t16 Vss.t562 Vss.t561 nfet_03v3
**devattr s=17600,576 d=17600,576
X384 SARlogic_0.dffrs_4.nand3_8.C.t3 SARlogic_0.dffrs_4.nand3_6.C.t4 Vdd.t832 Vdd.t831 pfet_03v3
**devattr s=44000,1176 d=26000,604
X385 a_n11637_14043 SARlogic_0.dffrs_13.nand3_8.Z.t4 a_n11821_14043 Vss.t547 nfet_03v3
**devattr s=10400,304 d=10400,304
X386 a_n7625_17007 Reset.t35 a_n7809_17007 Vss.t287 nfet_03v3
**devattr s=10400,304 d=10400,304
X387 a_33337_33720 a_33257_33628.t5 Vss.t579 Vss.t578 nfet_03v3
**devattr s=17600,576 d=10400,304
X388 a_n9861_28819.t2 SARlogic_0.d5.t5 a_n9673_28099 Vss.t84 nfet_03v3
**devattr s=10400,304 d=17600,576
X389 a_33521_29310 Vdd.t962 a_33337_29310 Vss.t497 nfet_03v3
**devattr s=10400,304 d=10400,304
X390 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t0 Clk.t11 Vdd.t79 Vdd.t78 pfet_03v3
**devattr s=14080,496 d=14080,496
X391 a_4921_30169.t1 adc_PISO_0.2inmux_2.OUT.t3 Vdd.t157 Vdd.t156 pfet_03v3
**devattr s=26000,604 d=44000,1176
X392 SARlogic_0.dffrs_4.nand3_6.C.t1 SARlogic_0.dffrs_4.nand3_1.C.t4 Vdd.t105 Vdd.t104 pfet_03v3
**devattr s=44000,1176 d=26000,604
X393 a_33337_35925 Vdd.t963 Vss.t496 Vss.t495 nfet_03v3
**devattr s=17600,576 d=10400,304
X394 a_24049_31515 Clk_piso.t5 a_23865_31515 Vss.t630 nfet_03v3
**devattr s=10400,304 d=10400,304
X395 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t0 Clk.t12 Vdd.t81 Vdd.t80 pfet_03v3
**devattr s=14080,496 d=14080,496
X396 a_n9861_28819.t0 SARlogic_0.d5.t6 Vdd.t123 Vdd.t122 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X397 a_37687_28100 a_36793_29020 Vss.t83 Vss.t82 nfet_03v3
**devattr s=17600,576 d=10400,304
X398 SARlogic_0.dffrs_10.Qb Reset.t36 Vdd.t361 Vdd.t360 pfet_03v3
**devattr s=26000,604 d=44000,1176
X399 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t3 Vss.t221 nfet_03v3
**devattr s=20800,504 d=20800,504
X400 a_12585_9633 Clk.t13 a_12401_9633 Vss.t52 nfet_03v3
**devattr s=10400,304 d=10400,304
X401 SARlogic_0.dffrs_4.Q.t1 SARlogic_0.dffrs_4.Qb.t5 Vdd.t305 Vdd.t304 pfet_03v3
**devattr s=26000,604 d=44000,1176
X402 Vdd.t363 Reset.t37 SARlogic_0.dffrs_7.nand3_8.Z Vdd.t362 pfet_03v3
**devattr s=26000,604 d=26000,604
X403 SARlogic_0.dffrs_2.nand3_8.C.t1 SARlogic_0.dffrs_2.nand3_8.Z.t5 Vdd.t213 Vdd.t212 pfet_03v3
**devattr s=26000,604 d=44000,1176
X404 SARlogic_0.dffrs_10.nand3_8.Z SAR_in.t4 a_8543_17004 Vss.t425 nfet_03v3
**devattr s=10400,304 d=17600,576
X405 a_16443_17004 SARlogic_0.dffrs_12.nand3_8.C.t7 Vss.t5 Vss.t4 nfet_03v3
**devattr s=17600,576 d=10400,304
X406 a_1945_9634 SARlogic_0.dffrs_2.nand3_8.C.t5 a_1761_9634 Vss.t667 nfet_03v3
**devattr s=10400,304 d=10400,304
X407 SARlogic_0.d0.t1 SARlogic_0.dffrs_11.Qb Vdd.t133 Vdd.t132 pfet_03v3
**devattr s=26000,604 d=44000,1176
X408 a_13887_9634 SARlogic_0.dffrs_5.Q.t4 Vss.t410 Vss.t409 nfet_03v3
**devattr s=17600,576 d=10400,304
X409 SARlogic_0.dffrs_7.nand3_6.C.t1 SARlogic_0.dffrs_7.nand3_1.C Vdd.t425 Vdd.t424 pfet_03v3
**devattr s=44000,1176 d=26000,604
X410 SARlogic_0.dffrs_0.nand3_8.Z.t2 SARlogic_0.dffrs_0.d.t7 a_n7625_7428 Vss.t593 nfet_03v3
**devattr s=10400,304 d=17600,576
X411 SARlogic_0.dffrs_9.nand3_8.C.t3 SARlogic_0.dffrs_9.nand3_6.C.t6 Vdd.t916 Vdd.t915 pfet_03v3
**devattr s=44000,1176 d=26000,604
X412 SARlogic_0.dffrs_2.nand3_6.C.t0 Clk.t14 Vdd.t83 Vdd.t82 pfet_03v3
**devattr s=26000,604 d=44000,1176
X413 a_16443_19209 SARlogic_0.dffrs_12.nand3_6.C.t7 Vss.t664 Vss.t663 nfet_03v3
**devattr s=17600,576 d=10400,304
X414 SARlogic_0.dffrs_10.nand3_8.C.t1 SARlogic_0.dffrs_10.nand3_8.Z a_8543_19209 Vss.t8 nfet_03v3
**devattr s=10400,304 d=17600,576
X415 Vdd.t571 SARlogic_0.dffrs_11.nand3_6.C.t6 SARlogic_0.d0.t2 Vdd.t570 pfet_03v3
**devattr s=26000,604 d=26000,604
X416 a_n9429_n2007.t18 Vin1.t2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t14 Vss.t180 nfet_03v3
**devattr s=15600,404 d=15600,404
X417 SARlogic_0.dffrs_12.Qb Reset.t38 Vdd.t365 Vdd.t364 pfet_03v3
**devattr s=26000,604 d=44000,1176
X418 a_459_9633 Clk.t15 a_275_9633 Vss.t53 nfet_03v3
**devattr s=10400,304 d=10400,304
X419 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_0.Qb.t6 Vdd.t199 Vdd.t198 pfet_03v3
**devattr s=44000,1176 d=26000,604
X420 SARlogic_0.dffrs_13.nand3_8.Z.t3 SARlogic_0.dffrs_13.nand3_8.C.t5 Vdd.t886 Vdd.t885 pfet_03v3
**devattr s=44000,1176 d=26000,604
X421 SARlogic_0.dffrs_4.nand3_1.C.t1 SARlogic_0.dffrs_4.nand3_6.C.t5 Vdd.t834 Vdd.t833 pfet_03v3
**devattr s=26000,604 d=44000,1176
X422 a_14313_31423.t2 Clk_piso.t6 Vdd.t878 Vdd.t877 pfet_03v3
**devattr s=26000,604 d=44000,1176
X423 Vss.t223 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t12 comparator_no_offsetcal_0.x5.out Vss.t222 nfet_03v3
**devattr s=35200,976 d=35200,976
X424 adc_PISO_0.dffrs_3.Q.t1 adc_PISO_0.dffrs_3.Qb Vdd.t517 Vdd.t516 pfet_03v3
**devattr s=26000,604 d=44000,1176
X425 SARlogic_0.d2.t0 SARlogic_0.dffrs_9.Qb a_5987_21414 Vss.t57 nfet_03v3
**devattr s=10400,304 d=17600,576
X426 a_8377_29020 inv2_0.out.t17 Vdd.t776 Vdd.t775 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X427 a_n2281_21414 SARlogic_0.dffrs_0.Qb.t7 Vss.t152 Vss.t151 nfet_03v3
**devattr s=17600,576 d=10400,304
X428 Comp_out.t2 a_n10831_4320 Vss.t570 Vss.t569 nfet_03v3
**devattr s=9350,280 d=9350,280
X429 Comp_out.t6 a_n10831_4320 Vdd.t788 Vdd.t787 pfet_03v3
**devattr s=34000,880 d=18700,450
X430 SARlogic_0.dffrs_14.nand3_1.C SARlogic_0.dffrs_14.nand3_6.C.t7 a_n7625_23622 Vss.t371 nfet_03v3
**devattr s=10400,304 d=17600,576
X431 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t13 Vin1.t3 a_n9429_n2007.t19 Vss.t193 nfet_03v3
**devattr s=15600,404 d=15600,404
X432 a_14313_33628.t2 a_14313_31423.t4 Vdd.t816 Vdd.t815 pfet_03v3
**devattr s=26000,604 d=44000,1176
X433 a_42809_29310 a_42729_29218.t4 Vss.t39 Vss.t38 nfet_03v3
**devattr s=17600,576 d=10400,304
X434 SARlogic_0.dffrs_8.Qb Reset.t39 Vdd.t367 Vdd.t366 pfet_03v3
**devattr s=26000,604 d=44000,1176
X435 SARlogic_0.dffrs_5.nand3_8.Z.t2 SARlogic_0.dffrs_4.Q.t5 a_12585_7428 Vss.t113 nfet_03v3
**devattr s=10400,304 d=17600,576
X436 SARlogic_0.dffrs_5.Qb.t0 Reset.t40 a_14071_9634 Vss.t288 nfet_03v3
**devattr s=10400,304 d=17600,576
X437 SARlogic_0.dffrs_2.Q.t1 SARlogic_0.dffrs_2.Qb.t4 Vdd.t870 Vdd.t869 pfet_03v3
**devattr s=26000,604 d=44000,1176
X438 SARlogic_0.dffrs_11.Qb Reset.t41 a_14071_19210 Vss.t289 nfet_03v3
**devattr s=10400,304 d=17600,576
X439 a_39915_29984 a_39055_28100 a_39727_29264.t1 Vdd.t388 pfet_03v3
**devattr s=52800,1376 d=31200,704
X440 a_n6323_11838 Vdd.t964 Vss.t494 Vss.t493 nfet_03v3
**devattr s=17600,576 d=10400,304
X441 SARlogic_0.dffrs_0.nand3_6.C.t1 Clk.t16 a_n7625_11838 Vss.t54 nfet_03v3
**devattr s=10400,304 d=17600,576
X442 a_29583_28100 a_28027_28820.t4 Vss.t595 Vss.t594 nfet_03v3
**devattr s=17600,576 d=17600,576
X443 Vdd.t313 SARlogic_0.dffrs_8.nand3_8.C.t6 SARlogic_0.dffrs_8.Qb Vdd.t312 pfet_03v3
**devattr s=26000,604 d=26000,604
X444 SARlogic_0.dffrs_2.nand3_8.C.t3 SARlogic_0.dffrs_2.nand3_6.C.t6 Vdd.t501 Vdd.t500 pfet_03v3
**devattr s=44000,1176 d=26000,604
X445 a_8359_17004 SARlogic_0.dffrs_10.nand3_8.C.t6 Vss.t191 Vss.t190 nfet_03v3
**devattr s=17600,576 d=10400,304
X446 Vdd.t37 adc_PISO_0.2inmux_2.Bit.t6 a_n389_31159.t0 Vdd.t36 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X447 Vdd.t503 SARlogic_0.dffrs_2.nand3_6.C.t7 SARlogic_0.dffrs_2.Q.t3 Vdd.t502 pfet_03v3
**devattr s=26000,604 d=26000,604
X448 a_14071_19210 SARlogic_0.dffrs_11.nand3_8.C.t5 a_13887_19210 Vss.t168 nfet_03v3
**devattr s=10400,304 d=10400,304
X449 a_23785_31423.t1 Clk_piso.t7 a_24049_33720 Vss.t184 nfet_03v3
**devattr s=10400,304 d=17600,576
X450 a_25351_33720 Vdd.t965 Vss.t492 Vss.t491 nfet_03v3
**devattr s=17600,576 d=10400,304
X451 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t13 Vdd.t339 Vdd.t338 pfet_03v3
**devattr s=10400,304 d=10400,304
X452 SARlogic_0.dffrs_7.nand3_6.C.t2 SARlogic_0.d3.t8 Vdd.t896 Vdd.t895 pfet_03v3
**devattr s=26000,604 d=44000,1176
X453 Vdd.t369 Reset.t42 SARlogic_0.dffrs_3.nand3_8.Z.t0 Vdd.t368 pfet_03v3
**devattr s=26000,604 d=26000,604
X454 SARlogic_0.dffrs_2.nand3_6.C.t2 SARlogic_0.dffrs_2.nand3_1.C.t4 Vdd.t477 Vdd.t476 pfet_03v3
**devattr s=44000,1176 d=26000,604
X455 a_8359_19209 SARlogic_0.dffrs_10.nand3_6.C.t8 Vss.t91 Vss.t90 nfet_03v3
**devattr s=17600,576 d=10400,304
X456 a_35007_33720 a_33257_31423.t8 a_34823_33720 Vss.t531 nfet_03v3
**devattr s=10400,304 d=10400,304
X457 Vdd.t255 adc_PISO_0.dffrs_3.Q.t6 a_28027_31160.t0 Vdd.t254 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X458 a_n2097_9634 SARlogic_0.dffrs_1.nand3_8.C.t5 a_n2281_9634 Vss.t341 nfet_03v3
**devattr s=10400,304 d=10400,304
X459 Vdd.t113 SARlogic_0.dffrs_3.nand3_8.C.t7 SARlogic_0.dffrs_3.Qb.t3 Vdd.t112 pfet_03v3
**devattr s=26000,604 d=26000,604
X460 a_23785_33628.t2 a_23785_31423.t8 a_24049_35925 Vss.t622 nfet_03v3
**devattr s=10400,304 d=17600,576
X461 a_n9861_31159.t3 inv2_0.out.t18 a_n9673_30439 Vss.t563 nfet_03v3
**devattr s=10400,304 d=17600,576
X462 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t6 Vdd.t802 Vdd.t801 pfet_03v3
**devattr s=26000,604 d=44000,1176
X463 a_459_21414 Reset.t43 a_275_21414 Vss.t290 nfet_03v3
**devattr s=10400,304 d=10400,304
X464 a_n7809_19212 SARlogic_0.dffrs_14.nand3_6.C.t8 Vss.t373 Vss.t372 nfet_03v3
**devattr s=17600,576 d=10400,304
X465 Vss.t265 a_27321_29020 a_28215_28100 Vss.t264 nfet_03v3
**devattr s=10400,304 d=17600,576
X466 SARlogic_0.dffrs_2.nand3_8.Z.t1 SARlogic_0.dffrs_2.d.t5 a_459_7428 Vss.t16 nfet_03v3
**devattr s=10400,304 d=17600,576
X467 SARlogic_0.dffrs_4.nand3_1.C.t3 Vdd.t664 Vdd.t666 Vdd.t665 pfet_03v3
**devattr s=44000,1176 d=26000,604
X468 adc_PISO_0.dffrs_3.Qb Vdd.t661 Vdd.t663 Vdd.t662 pfet_03v3
**devattr s=26000,604 d=44000,1176
X469 Vdd.t247 SARlogic_0.dffrs_10.nand3_8.C.t7 SARlogic_0.dffrs_10.Qb Vdd.t246 pfet_03v3
**devattr s=26000,604 d=26000,604
X470 a_13887_11838 Vdd.t966 Vss.t490 Vss.t489 nfet_03v3
**devattr s=17600,576 d=10400,304
X471 a_28215_30440 inv2_0.out.t19 a_28027_31160.t1 Vss.t564 nfet_03v3
**devattr s=17600,576 d=10400,304
X472 Vdd.t836 SARlogic_0.dffrs_4.nand3_6.C.t6 SARlogic_0.dffrs_4.Q.t3 Vdd.t835 pfet_03v3
**devattr s=26000,604 d=26000,604
X473 SARlogic_0.dffrs_8.nand3_8.Z SAR_in.t5 a_459_17004 Vss.t426 nfet_03v3
**devattr s=10400,304 d=17600,576
X474 SARlogic_0.dffrs_4.nand3_8.Z.t3 SARlogic_0.dffrs_4.d.t6 Vdd.t812 Vdd.t811 pfet_03v3
**devattr s=26000,604 d=44000,1176
X475 a_459_23619 SARlogic_0.dffrs_8.nand3_8.Z a_275_23619 Vss.t253 nfet_03v3
**devattr s=10400,304 d=10400,304
X476 Vdd.t660 Vdd.t658 a_23785_31423.t2 Vdd.t659 pfet_03v3
**devattr s=26000,604 d=26000,604
X477 a_17929_21414 SARlogic_0.dffrs_5.Qb.t7 Vss.t328 Vss.t327 nfet_03v3
**devattr s=17600,576 d=10400,304
X478 adc_PISO_0.2inmux_1.OUT.t0 a_39727_29264.t4 Vss.t645 Vss.t644 nfet_03v3
**devattr s=17600,576 d=17600,576
X479 SARlogic_0.dffrs_8.nand3_8.C.t1 SARlogic_0.dffrs_8.nand3_8.Z a_459_19209 Vss.t252 nfet_03v3
**devattr s=10400,304 d=17600,576
X480 SARlogic_0.dffrs_1.nand3_8.Z.t1 SARlogic_0.dffrs_0.Q.t5 a_n3583_7428 Vss.t676 nfet_03v3
**devattr s=10400,304 d=17600,576
X481 a_25351_31516 adc_PISO_0.dffrs_3.Q.t7 Vss.t197 Vss.t196 nfet_03v3
**devattr s=17600,576 d=10400,304
X482 SARlogic_0.dffrs_0.Q.t1 SARlogic_0.dffrs_0.Qb.t8 a_n6139_11838 Vss.t153 nfet_03v3
**devattr s=10400,304 d=17600,576
X483 a_n4631_29217.t0 a_n4631_31422.t5 Vdd.t734 Vdd.t733 pfet_03v3
**devattr s=44000,1176 d=26000,604
X484 a_n6323_9634 SARlogic_0.dffrs_0.Q.t6 Vss.t3 Vss.t2 nfet_03v3
**devattr s=17600,576 d=10400,304
X485 Vdd.t153 a_23865_30170.t5 a_23785_33628.t1 Vdd.t152 pfet_03v3
**devattr s=26000,604 d=26000,604
X486 a_8543_11838 Reset.t44 a_8359_11838 Vss.t291 nfet_03v3
**devattr s=10400,304 d=10400,304
X487 SARlogic_0.dffrs_5.nand3_1.C.t0 SARlogic_0.dffrs_5.nand3_6.C.t6 a_12585_14043 Vss.t538 nfet_03v3
**devattr s=10400,304 d=17600,576
X488 SARlogic_0.dffrs_2.nand3_1.C.t2 SARlogic_0.dffrs_2.nand3_6.C.t8 Vdd.t505 Vdd.t504 pfet_03v3
**devattr s=26000,604 d=44000,1176
X489 a_14393_30170.t2 a_14313_29218.t5 Vdd.t307 Vdd.t306 pfet_03v3
**devattr s=44000,1176 d=26000,604
X490 Vdd.t533 SARlogic_0.dffrs_12.Q.t6 SARlogic_0.dffrs_11.nand3_8.C.t2 Vdd.t532 pfet_03v3
**devattr s=26000,604 d=26000,604
X491 a_35007_31516 a_33257_29218.t5 a_34823_31516 Vss.t143 nfet_03v3
**devattr s=10400,304 d=10400,304
X492 a_n4631_31422.t2 a_n4631_33627.t4 Vdd.t555 Vdd.t554 pfet_03v3
**devattr s=44000,1176 d=26000,604
X493 a_42729_29218.t1 a_42809_30170.t6 a_42993_31515 Vss.t259 nfet_03v3
**devattr s=10400,304 d=17600,576
X494 a_14313_29218.t2 a_14313_31423.t5 Vdd.t547 Vdd.t546 pfet_03v3
**devattr s=44000,1176 d=26000,604
X495 a_14577_31515 Clk_piso.t8 a_14393_31515 Vss.t185 nfet_03v3
**devattr s=10400,304 d=10400,304
X496 a_n10567_29019 inv2_0.out.t20 Vdd.t778 Vdd.t777 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X497 a_33337_30170.t2 adc_PISO_0.2inmux_5.OUT.t2 a_33521_29310 Vss.t369 nfet_03v3
**devattr s=10400,304 d=17600,576
X498 a_4501_14043 SARlogic_0.dffrs_3.nand3_8.Z.t6 a_4317_14043 Vss.t419 nfet_03v3
**devattr s=10400,304 d=10400,304
X499 a_275_17004 SARlogic_0.dffrs_8.nand3_8.C.t7 Vss.t251 Vss.t250 nfet_03v3
**devattr s=17600,576 d=10400,304
X500 a_n7625_7428 Reset.t45 a_n7809_7428 Vss.t292 nfet_03v3
**devattr s=10400,304 d=10400,304
X501 a_275_19209 SARlogic_0.dffrs_8.nand3_6.C.t8 Vss.t32 Vss.t31 nfet_03v3
**devattr s=17600,576 d=10400,304
X502 Vdd.t283 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t5 Vdd.t282 pfet_03v3
**devattr s=10400,304 d=10400,304
X503 SARlogic_0.dffrs_4.Qb.t0 Reset.t46 a_10029_9634 Vss.t293 nfet_03v3
**devattr s=10400,304 d=17600,576
X504 SARlogic_0.dffrs_7.nand3_8.Z SARlogic_0.dffrs_7.nand3_8.C.t5 Vdd.t93 Vdd.t92 pfet_03v3
**devattr s=44000,1176 d=26000,604
X505 a_16627_17004 Reset.t47 a_16443_17004 Vss.t294 nfet_03v3
**devattr s=10400,304 d=10400,304
X506 a_n4631_29217.t2 a_n4551_30169.t5 Vdd.t908 Vdd.t907 pfet_03v3
**devattr s=26000,604 d=44000,1176
X507 Vdd.t163 a_n8305_30439 a_n7445_29983 Vdd.t162 pfet_03v3
**devattr s=31200,704 d=52800,1376
X508 SARlogic_0.dffrs_2.nand3_1.C.t1 Vdd.t655 Vdd.t657 Vdd.t656 pfet_03v3
**devattr s=44000,1176 d=26000,604
X509 SARlogic_0.dffrs_13.nand3_8.C.t1 SARlogic_0.dffrs_13.nand3_8.Z.t5 a_n11637_9633 Vss.t548 nfet_03v3
**devattr s=10400,304 d=17600,576
X510 a_16627_19209 Vss.t100 a_16443_19209 Vss.t101 nfet_03v3
**devattr s=10400,304 d=10400,304
X511 a_n4631_31422.t1 Clk_piso.t9 Vdd.t231 Vdd.t230 pfet_03v3
**devattr s=26000,604 d=44000,1176
X512 adc_PISO_0.2inmux_2.Bit.t1 Vdd.t652 Vdd.t654 Vdd.t653 pfet_03v3
**devattr s=44000,1176 d=26000,604
X513 adc_PISO_0.dffrs_2.Q.t1 adc_PISO_0.dffrs_2.Qb Vdd.t515 Vdd.t514 pfet_03v3
**devattr s=26000,604 d=44000,1176
X514 SARlogic_0.dffrs_9.Qb Reset.t48 Vdd.t371 Vdd.t370 pfet_03v3
**devattr s=26000,604 d=44000,1176
X515 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t14 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t271 nfet_03v3
**devattr s=20800,504 d=20800,504
X516 SARlogic_0.dffrs_7.Qb SARlogic_0.d4.t7 Vdd.t221 Vdd.t220 pfet_03v3
**devattr s=44000,1176 d=26000,604
X517 SARlogic_0.dffrs_4.d.t0 SARlogic_0.dffrs_3.Qb.t8 Vdd.t399 Vdd.t398 pfet_03v3
**devattr s=26000,604 d=44000,1176
X518 Piso_out.t2 adc_PISO_0.dffrs_5.Qb Vdd.t487 Vdd.t486 pfet_03v3
**devattr s=26000,604 d=44000,1176
X519 SARlogic_0.dffrs_2.d.t3 Vdd.t649 Vdd.t651 Vdd.t650 pfet_03v3
**devattr s=44000,1176 d=26000,604
X520 Vdd.t736 a_n4631_31422.t6 adc_PISO_0.2inmux_2.Bit.t0 Vdd.t735 pfet_03v3
**devattr s=26000,604 d=26000,604
X521 Vdd.t549 a_14313_31423.t6 adc_PISO_0.dffrs_2.Q.t2 Vdd.t548 pfet_03v3
**devattr s=26000,604 d=26000,604
X522 a_33337_29310 a_33257_29218.t6 Vss.t145 Vss.t144 nfet_03v3
**devattr s=17600,576 d=10400,304
X523 a_n10831_4320 comparator_no_offsetcal_0.x4.A Vdd.t323 Vdd.t322 pfet_03v3
**devattr s=18700,450 d=34000,880
X524 a_n3583_21414 Reset.t49 a_n3767_21414 Vss.t295 nfet_03v3
**devattr s=10400,304 d=10400,304
X525 SARlogic_0.dffrs_3.nand3_8.Z.t3 SARlogic_0.dffrs_2.Q.t5 Vdd.t335 Vdd.t334 pfet_03v3
**devattr s=26000,604 d=44000,1176
X526 SARlogic_0.dffrs_0.Qb.t0 SARlogic_0.dffrs_0.Q.t7 Vdd.t1 Vdd.t0 pfet_03v3
**devattr s=44000,1176 d=26000,604
X527 a_n7625_23622 SARlogic_0.dffrs_14.nand3_8.Z a_n7809_23622 Vss.t159 nfet_03v3
**devattr s=10400,304 d=10400,304
X528 a_n3583_23619 SARlogic_0.dffrs_7.nand3_8.Z a_n3767_23619 Vss.t161 nfet_03v3
**devattr s=10400,304 d=10400,304
X529 a_20971_29984 a_20111_30440 Vdd.t99 Vdd.t98 pfet_03v3
**devattr s=52800,1376 d=31200,704
X530 Vdd.t85 Clk.t17 SARlogic_0.dffrs_2.nand3_8.C.t0 Vdd.t84 pfet_03v3
**devattr s=26000,604 d=26000,604
X531 a_n7625_11838 Reset.t50 a_n7809_11838 Vss.t296 nfet_03v3
**devattr s=10400,304 d=10400,304
X532 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t6 Vdd.t561 Vdd.t560 pfet_03v3
**devattr s=26000,604 d=44000,1176
X533 a_25535_33720 a_23785_31423.t9 a_25351_33720 Vss.t623 nfet_03v3
**devattr s=10400,304 d=10400,304
X534 Vss.t402 a_39055_30440 a_39727_29264.t3 Vss.t401 nfet_03v3
**devattr s=17600,576 d=17600,576
X535 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t4 a_n9767_249 a_n9855_341 Vss.t336 nfet_03v3
**devattr s=35200,976 d=20800,504
X536 Vdd.t373 Reset.t51 SARlogic_0.dffrs_2.nand3_6.C.t1 Vdd.t372 pfet_03v3
**devattr s=26000,604 d=26000,604
X537 adc_PISO_0.dffrs_2.Qb Vdd.t646 Vdd.t648 Vdd.t647 pfet_03v3
**devattr s=26000,604 d=44000,1176
X538 adc_PISO_0.dffrs_5.Qb Vdd.t643 Vdd.t645 Vdd.t644 pfet_03v3
**devattr s=26000,604 d=44000,1176
X539 a_20111_28100 a_18555_28820.t5 Vdd.t792 Vdd.t791 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X540 SARlogic_0.dffrs_11.nand3_6.C.t3 SARlogic_0.dffrs_12.Q.t7 Vdd.t535 Vdd.t534 pfet_03v3
**devattr s=26000,604 d=44000,1176
X541 SARlogic_0.dffrs_5.Qb.t2 SARlogic_0.dffrs_5.Q.t5 Vdd.t537 Vdd.t536 pfet_03v3
**devattr s=44000,1176 d=26000,604
X542 Vdd.t349 a_4841_31422.t6 adc_PISO_0.dffrs_1.Q.t3 Vdd.t348 pfet_03v3
**devattr s=26000,604 d=26000,604
X543 adc_PISO_0.dffrs_1.Q.t0 adc_PISO_0.dffrs_1.Qb a_6591_33719 Vss.t22 nfet_03v3
**devattr s=10400,304 d=17600,576
X544 Vdd.t309 a_14313_29218.t6 adc_PISO_0.dffrs_2.Qb Vdd.t308 pfet_03v3
**devattr s=26000,604 d=26000,604
X545 a_37499_28820.t3 SARlogic_0.d0.t9 Vdd.t263 Vdd.t262 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X546 a_42729_31423.t2 Clk_piso.t10 Vdd.t233 Vdd.t232 pfet_03v3
**devattr s=26000,604 d=44000,1176
X547 a_8359_9633 SARlogic_0.dffrs_4.nand3_6.C.t7 Vss.t599 Vss.t598 nfet_03v3
**devattr s=17600,576 d=10400,304
X548 Vdd.t642 Vdd.t640 a_14313_31423.t0 Vdd.t641 pfet_03v3
**devattr s=26000,604 d=26000,604
X549 SARlogic_0.dffrs_12.Qb SARlogic_0.dffrs_12.Q.t8 Vdd.t499 Vdd.t498 pfet_03v3
**devattr s=44000,1176 d=26000,604
X550 a_1761_11838 Vdd.t967 Vss.t488 Vss.t487 nfet_03v3
**devattr s=17600,576 d=10400,304
X551 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t7 Vdd.t573 Vdd.t572 pfet_03v3
**devattr s=26000,604 d=44000,1176
X552 a_n6389_n2007 a_n6589_n2099 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t6 Vss.t156 nfet_03v3
**devattr s=15600,404 d=26400,776
X553 a_18555_31160.t3 inv2_0.out.t21 Vdd.t780 Vdd.t779 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X554 adc_PISO_0.2inmux_2.OUT.t0 a_1839_29263.t4 Vss.t274 Vss.t273 nfet_03v3
**devattr s=17600,576 d=17600,576
X555 a_n2097_21414 SARlogic_0.dffrs_7.nand3_6.C.t7 a_n2281_21414 Vss.t624 nfet_03v3
**devattr s=10400,304 d=10400,304
X556 SARlogic_0.dffrs_0.Qb.t2 Reset.t52 Vdd.t375 Vdd.t374 pfet_03v3
**devattr s=26000,604 d=44000,1176
X557 a_42729_33628.t2 a_42729_31423.t4 Vdd.t840 Vdd.t839 pfet_03v3
**devattr s=26000,604 d=44000,1176
X558 Vdd.t377 Reset.t53 SARlogic_0.dffrs_9.nand3_6.C.t2 Vdd.t376 pfet_03v3
**devattr s=26000,604 d=26000,604
X559 Vdd.t856 a_14393_30170.t6 a_14313_33628.t3 Vdd.t855 pfet_03v3
**devattr s=26000,604 d=26000,604
X560 SARlogic_0.d4.t1 SARlogic_0.dffrs_7.Qb a_n2097_21414 Vss.t414 nfet_03v3
**devattr s=10400,304 d=17600,576
X561 Vdd.t830 SARlogic_0.dffrs_13.nand3_6.C.t5 SARlogic_0.dffrs_0.d.t1 Vdd.t829 pfet_03v3
**devattr s=26000,604 d=26000,604
X562 SARlogic_0.dffrs_14.nand3_8.C.t1 SARlogic_0.dffrs_14.nand3_8.Z a_n7625_19212 Vss.t158 nfet_03v3
**devattr s=10400,304 d=17600,576
X563 a_n6139_11838 SARlogic_0.dffrs_0.nand3_6.C.t8 a_n6323_11838 Vss.t43 nfet_03v3
**devattr s=10400,304 d=10400,304
X564 a_n8351_341 a_n8551_249 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t1 Vss.t139 nfet_03v3
**devattr s=20800,504 d=35200,976
X565 adc_PISO_0.2inmux_3.OUT.t0 a_11311_29264.t4 Vss.t138 Vss.t137 nfet_03v3
**devattr s=17600,576 d=17600,576
X566 a_25535_31516 a_23785_29218.t6 a_25351_31516 Vss.t142 nfet_03v3
**devattr s=10400,304 d=10400,304
X567 Vdd.t159 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_1.C Vdd.t158 pfet_03v3
**devattr s=26000,604 d=26000,604
X568 SARlogic_0.dffrs_4.nand3_6.C.t2 Clk.t18 a_8543_11838 Vss.t431 nfet_03v3
**devattr s=10400,304 d=17600,576
X569 a_9845_11838 Vdd.t968 Vss.t486 Vss.t485 nfet_03v3
**devattr s=17600,576 d=10400,304
X570 a_18743_28100 SARlogic_0.d2.t8 a_18555_28820.t3 Vss.t231 nfet_03v3
**devattr s=17600,576 d=10400,304
X571 Vdd.t379 Reset.t54 SARlogic_0.dffrs_1.nand3_8.Z.t0 Vdd.t378 pfet_03v3
**devattr s=26000,604 d=26000,604
X572 Vdd.t235 Clk_piso.t11 a_4841_29217.t3 Vdd.t234 pfet_03v3
**devattr s=26000,604 d=26000,604
X573 Vdd.t639 Vdd.t637 a_42809_30170.t1 Vdd.t638 pfet_03v3
**devattr s=26000,604 d=26000,604
X574 a_39055_28100 a_37499_28820.t5 Vdd.t858 Vdd.t857 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X575 a_23865_30170.t1 adc_PISO_0.2inmux_4.OUT.t2 a_24049_29310 Vss.t422 nfet_03v3
**devattr s=10400,304 d=17600,576
X576 Vdd.t888 a_1167_30439 a_2027_29983 Vdd.t887 pfet_03v3
**devattr s=31200,704 d=52800,1376
X577 a_23865_33720 a_23785_33628.t5 Vss.t577 Vss.t576 nfet_03v3
**devattr s=17600,576 d=10400,304
X578 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 Vdd.t341 Vdd.t340 pfet_03v3
**devattr s=10400,304 d=10400,304
X579 a_n7445_29983 a_n8305_28099 a_n7633_29263.t2 Vdd.t302 pfet_03v3
**devattr s=52800,1376 d=31200,704
X580 a_4841_29217.t2 a_4841_31422.t7 Vdd.t351 Vdd.t350 pfet_03v3
**devattr s=44000,1176 d=26000,604
X581 a_n9429_n2007.t5 Vin2.t4 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t182 nfet_03v3
**devattr s=15600,404 d=15600,404
X582 Vdd.t636 Vdd.t634 a_4841_31422.t3 Vdd.t635 pfet_03v3
**devattr s=26000,604 d=26000,604
X583 Vdd.t237 Clk_piso.t12 a_42729_29218.t3 Vdd.t236 pfet_03v3
**devattr s=26000,604 d=26000,604
X584 a_459_17004 Reset.t55 a_275_17004 Vss.t297 nfet_03v3
**devattr s=10400,304 d=10400,304
X585 SARlogic_0.dffrs_3.nand3_1.C.t1 SARlogic_0.dffrs_3.nand3_6.C.t8 a_4501_14043 Vss.t331 nfet_03v3
**devattr s=10400,304 d=17600,576
X586 a_12401_14043 Vdd.t970 Vss.t482 Vss.t481 nfet_03v3
**devattr s=17600,576 d=10400,304
X587 Vdd.t906 a_10639_30440 a_11499_29984 Vdd.t905 pfet_03v3
**devattr s=31200,704 d=52800,1376
X588 a_23865_35925 Vdd.t969 Vss.t484 Vss.t483 nfet_03v3
**devattr s=17600,576 d=10400,304
X589 Comp_out.t5 a_n10831_4320 Vdd.t786 Vdd.t785 pfet_03v3
**devattr s=18700,450 d=18700,450
X590 a_8543_7428 Reset.t56 a_8359_7428 Vss.t298 nfet_03v3
**devattr s=10400,304 d=10400,304
X591 a_4841_31422.t1 a_4841_33627.t4 Vdd.t229 Vdd.t228 pfet_03v3
**devattr s=44000,1176 d=26000,604
X592 SARlogic_0.dffrs_0.nand3_8.Z.t1 SARlogic_0.dffrs_0.nand3_8.C.t5 Vdd.t21 Vdd.t20 pfet_03v3
**devattr s=44000,1176 d=26000,604
X593 Vdd.t265 SARlogic_0.d0.t10 SARlogic_0.dffrs_10.nand3_8.C.t2 Vdd.t264 pfet_03v3
**devattr s=26000,604 d=26000,604
X594 a_n1095_29019 inv2_0.out.t22 Vdd.t782 Vdd.t781 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X595 a_n11637_9633 Clk.t19 a_n11821_9633 Vss.t432 nfet_03v3
**devattr s=10400,304 d=10400,304
X596 a_459_19209 SARlogic_0.d2.t9 a_275_19209 Vss.t232 nfet_03v3
**devattr s=10400,304 d=10400,304
X597 a_20111_30440 a_18555_31160.t4 Vss.t21 Vss.t20 nfet_03v3
**devattr s=17600,576 d=17600,576
X598 a_37499_31160.t1 inv2_0.out.t23 a_37687_30440 Vss.t441 nfet_03v3
**devattr s=10400,304 d=17600,576
X599 a_30255_29264.t1 a_29583_28100 Vss.t239 Vss.t238 nfet_03v3
**devattr s=17600,576 d=17600,576
X600 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t5 a_n9429_n2007.t6 Vss.t183 nfet_03v3
**devattr s=15600,404 d=15600,404
X601 Vdd.t47 Clk_piso.t13 a_n4631_29217.t1 Vdd.t46 pfet_03v3
**devattr s=26000,604 d=26000,604
X602 Vdd.t215 SARlogic_0.dffrs_2.nand3_8.Z.t6 SARlogic_0.dffrs_2.nand3_1.C.t0 Vdd.t214 pfet_03v3
**devattr s=26000,604 d=26000,604
X603 a_8359_11838 SARlogic_0.dffrs_4.nand3_1.C.t5 Vss.t70 Vss.t69 nfet_03v3
**devattr s=17600,576 d=10400,304
X604 Vss.t400 a_n8385_n2885 a_n8473_n2793 Vss.t399 nfet_03v3
**devattr s=14080,496 d=8320,264
X605 Vdd.t575 Clk.t20 SARlogic_0.dffrs_1.nand3_8.C.t3 Vdd.t574 pfet_03v3
**devattr s=26000,604 d=26000,604
X606 adc_PISO_0.2inmux_4.OUT.t1 a_20783_29264.t5 Vdd.t191 Vdd.t190 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X607 a_2027_29983 a_1167_28099 a_1839_29263.t1 Vdd.t298 pfet_03v3
**devattr s=52800,1376 d=31200,704
X608 SARlogic_0.dffrs_4.Q.t0 SARlogic_0.dffrs_4.Qb.t6 a_10029_11838 Vss.t613 nfet_03v3
**devattr s=10400,304 d=17600,576
X609 Vdd.t633 Vdd.t631 a_n4631_31422.t3 Vdd.t632 pfet_03v3
**devattr s=26000,604 d=26000,604
X610 Vdd.t756 a_8377_29020 a_9083_28820.t0 Vdd.t755 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X611 Vdd.t381 Reset.t57 SARlogic_0.dffrs_1.nand3_6.C.t0 Vdd.t380 pfet_03v3
**devattr s=26000,604 d=26000,604
X612 a_27321_29020 inv2_0.out.t24 Vdd.t589 Vdd.t588 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X613 a_4317_9633 SARlogic_0.dffrs_3.nand3_6.C.t9 Vss.t333 Vss.t332 nfet_03v3
**devattr s=17600,576 d=10400,304
X614 a_4317_14043 Vdd.t971 Vss.t480 Vss.t479 nfet_03v3
**devattr s=17600,576 d=10400,304
X615 SARlogic_0.dffrs_13.nand3_8.C.t3 SARlogic_0.dffrs_13.nand3_6.C.t6 Vdd.t826 Vdd.t825 pfet_03v3
**devattr s=44000,1176 d=26000,604
X616 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t6 a_n9429_n2007.t7 Vss.t192 nfet_03v3
**devattr s=15600,404 d=15600,404
X617 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t7 a_n9429_n2007.t8 Vss.t193 nfet_03v3
**devattr s=15600,404 d=15600,404
X618 SARlogic_0.d0.t0 SARlogic_0.dffrs_11.Qb a_14071_21414 Vss.t94 nfet_03v3
**devattr s=10400,304 d=17600,576
X619 a_n3767_21414 SARlogic_0.dffrs_7.nand3_1.C Vss.t324 Vss.t323 nfet_03v3
**devattr s=17600,576 d=10400,304
X620 Vss.t62 a_n1095_29019 a_n201_28099 Vss.t61 nfet_03v3
**devattr s=10400,304 d=17600,576
X621 Vss.t647 a_10639_30440 a_11311_29264.t3 Vss.t646 nfet_03v3
**devattr s=17600,576 d=17600,576
X622 SARlogic_0.dffrs_2.nand3_6.C.t3 Clk.t21 a_459_11838 Vss.t433 nfet_03v3
**devattr s=10400,304 d=17600,576
X623 a_14071_21414 SARlogic_0.dffrs_11.nand3_6.C.t8 a_13887_21414 Vss.t429 nfet_03v3
**devattr s=10400,304 d=10400,304
X624 SARlogic_0.dffrs_13.nand3_6.C.t3 SARlogic_0.dffrs_13.nand3_1.C.t4 Vdd.t924 Vdd.t923 pfet_03v3
**devattr s=44000,1176 d=26000,604
X625 a_n11821_7428 SARlogic_0.dffrs_13.nand3_8.C.t6 Vss.t7 Vss.t6 nfet_03v3
**devattr s=17600,576 d=10400,304
X626 a_n3767_23619 SARlogic_0.dffrs_0.Qb.t9 Vss.t155 Vss.t154 nfet_03v3
**devattr s=17600,576 d=10400,304
X627 a_39055_30440 a_37499_31160.t4 Vss.t581 Vss.t580 nfet_03v3
**devattr s=17600,576 d=17600,576
X628 Vdd.t119 a_36793_29020 a_37499_28820.t0 Vdd.t118 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X629 a_14313_31423.t1 Clk_piso.t14 a_14577_33720 Vss.t35 nfet_03v3
**devattr s=10400,304 d=17600,576
X630 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t7 Vdd.t563 Vdd.t562 pfet_03v3
**devattr s=26000,604 d=44000,1176
X631 a_n9429_n2007.t20 Vin1.t4 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t12 Vss.t194 nfet_03v3
**devattr s=15600,404 d=15600,404
X632 adc_PISO_0.dffrs_3.Q.t0 adc_PISO_0.dffrs_3.Qb a_25535_33720 Vss.t395 nfet_03v3
**devattr s=10400,304 d=17600,576
X633 adc_PISO_0.dffrs_1.Qb Vdd.t628 Vdd.t630 Vdd.t629 pfet_03v3
**devattr s=26000,604 d=44000,1176
X634 Vdd.t353 adc_PISO_0.dffrs_2.Q.t5 a_18555_31160.t0 Vdd.t352 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X635 SARlogic_0.dffrs_2.Qb.t3 SARlogic_0.dffrs_2.Q.t6 Vdd.t337 Vdd.t336 pfet_03v3
**devattr s=44000,1176 d=26000,604
X636 a_14313_33628.t0 a_14313_31423.t7 a_14577_35925 Vss.t417 nfet_03v3
**devattr s=10400,304 d=17600,576
X637 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t16 Vdd.t343 Vdd.t342 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X638 SARlogic_0.dffrs_2.Q.t2 SARlogic_0.dffrs_2.Qb.t5 a_1945_11838 Vss.t628 nfet_03v3
**devattr s=10400,304 d=17600,576
X639 Vdd.t7 Vss.t678 a_n9861_31159.t0 Vdd.t6 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X640 a_n7809_14043 Vdd.t972 Vss.t478 Vss.t477 nfet_03v3
**devattr s=17600,576 d=10400,304
X641 Vdd.t91 SARlogic_0.dffrs_7.nand3_8.C.t6 SARlogic_0.dffrs_7.Qb Vdd.t90 pfet_03v3
**devattr s=26000,604 d=26000,604
X642 Vss.t72 a_17849_29020 a_18743_28100 Vss.t71 nfet_03v3
**devattr s=10400,304 d=17600,576
X643 Vdd.t842 a_42729_31423.t5 Piso_out.t0 Vdd.t841 pfet_03v3
**devattr s=26000,604 d=26000,604
X644 Vdd.t273 SARlogic_0.dffrs_1.nand3_6.C.t6 SARlogic_0.dffrs_2.d.t0 Vdd.t272 pfet_03v3
**devattr s=26000,604 d=26000,604
X645 Vdd.t383 Reset.t58 SARlogic_0.dffrs_9.nand3_8.Z Vdd.t382 pfet_03v3
**devattr s=26000,604 d=26000,604
X646 a_1945_11838 SARlogic_0.dffrs_2.nand3_6.C.t9 a_1761_11838 Vss.t384 nfet_03v3
**devattr s=10400,304 d=10400,304
X647 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t11 Vin1.t5 a_n9429_n2007.t11 Vss.t195 nfet_03v3
**devattr s=15600,404 d=15600,404
X648 Vdd.t577 Clk.t22 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t1 Vdd.t576 pfet_03v3
**devattr s=14080,496 d=14080,496
X649 adc_PISO_0.dffrs_2.Q.t3 Vdd.t625 Vdd.t627 Vdd.t626 pfet_03v3
**devattr s=44000,1176 d=26000,604
X650 adc_PISO_0.2inmux_2.Bit.t3 adc_PISO_0.dffrs_0.Qb Vdd.t892 Vdd.t891 pfet_03v3
**devattr s=26000,604 d=44000,1176
X651 SARlogic_0.dffrs_13.nand3_8.C.t2 SARlogic_0.dffrs_13.nand3_8.Z.t6 Vdd.t762 Vdd.t761 pfet_03v3
**devattr s=26000,604 d=44000,1176
X652 SARlogic_0.dffrs_7.Qb Reset.t59 Vdd.t385 Vdd.t384 pfet_03v3
**devattr s=26000,604 d=44000,1176
X653 SARlogic_0.dffrs_2.d.t2 SARlogic_0.dffrs_1.Qb.t8 Vdd.t495 Vdd.t494 pfet_03v3
**devattr s=26000,604 d=44000,1176
X654 a_4501_7428 Reset.t60 a_4317_7428 Vss.t299 nfet_03v3
**devattr s=10400,304 d=10400,304
X655 SARlogic_0.dffrs_7.nand3_6.C.t3 SARlogic_0.d3.t9 a_n3583_21414 Vss.t640 nfet_03v3
**devattr s=10400,304 d=17600,576
X656 a_275_11838 SARlogic_0.dffrs_2.nand3_1.C.t5 Vss.t340 Vss.t339 nfet_03v3
**devattr s=17600,576 d=10400,304
X657 Vdd.t23 SARlogic_0.dffrs_0.nand3_8.C.t6 SARlogic_0.dffrs_0.Qb.t1 Vdd.t22 pfet_03v3
**devattr s=26000,604 d=26000,604
X658 SARlogic_0.dffrs_1.nand3_8.Z.t3 SARlogic_0.dffrs_1.nand3_8.C.t6 Vdd.t445 Vdd.t444 pfet_03v3
**devattr s=44000,1176 d=26000,604
X659 SARlogic_0.dffrs_12.nand3_8.C.t3 SARlogic_0.dffrs_12.nand3_8.Z Vdd.t758 Vdd.t757 pfet_03v3
**devattr s=26000,604 d=44000,1176
X660 SARlogic_0.dffrs_11.nand3_6.C.t1 SARlogic_0.dffrs_11.nand3_1.C Vdd.t447 Vdd.t446 pfet_03v3
**devattr s=44000,1176 d=26000,604
X661 SARlogic_0.d2.t2 SARlogic_0.dffrs_2.Qb.t6 Vdd.t880 Vdd.t879 pfet_03v3
**devattr s=44000,1176 d=26000,604
X662 SARlogic_0.dffrs_9.nand3_6.C.t1 SARlogic_0.d1.t9 Vdd.t810 Vdd.t809 pfet_03v3
**devattr s=26000,604 d=44000,1176
X663 a_n3583_17004 Reset.t61 a_n3767_17004 Vss.t300 nfet_03v3
**devattr s=10400,304 d=10400,304
X664 SARlogic_0.dffrs_13.nand3_6.C.t1 Clk.t23 Vdd.t579 Vdd.t578 pfet_03v3
**devattr s=26000,604 d=44000,1176
X665 SARlogic_0.dffrs_4.Qb.t2 SARlogic_0.dffrs_4.Q.t6 Vdd.t139 Vdd.t138 pfet_03v3
**devattr s=44000,1176 d=26000,604
X666 SARlogic_0.dffrs_0.d.t0 Reset.t62 Vdd.t387 Vdd.t386 pfet_03v3
**devattr s=44000,1176 d=26000,604
X667 a_n7625_19212 SARlogic_0.d4.t8 a_n7809_19212 Vss.t174 nfet_03v3
**devattr s=10400,304 d=10400,304
X668 SARlogic_0.dffrs_7.nand3_1.C SARlogic_0.dffrs_7.nand3_6.C.t8 a_n3583_23619 Vss.t625 nfet_03v3
**devattr s=10400,304 d=17600,576
X669 a_37687_28100 SARlogic_0.d0.t11 a_37499_28820.t1 Vss.t205 nfet_03v3
**devattr s=17600,576 d=10400,304
X670 a_9271_30440 adc_PISO_0.dffrs_1.Q.t7 Vss.t213 Vss.t212 nfet_03v3
**devattr s=17600,576 d=10400,304
X671 Vdd.t624 Vdd.t622 a_33337_30170.t3 Vdd.t623 pfet_03v3
**devattr s=26000,604 d=26000,604
X672 adc_PISO_0.dffrs_3.Qb Vdd.t973 a_25535_31516 Vss.t476 nfet_03v3
**devattr s=10400,304 d=17600,576
X673 a_10029_11838 SARlogic_0.dffrs_4.nand3_6.C.t8 a_9845_11838 Vss.t600 nfet_03v3
**devattr s=10400,304 d=10400,304
X674 Vdd.t489 a_n9629_1405 a_n9717_1497 Vdd.t488 pfet_03v3
**devattr s=17600,576 d=10400,304
X675 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_4.Qb.t7 Vdd.t860 Vdd.t859 pfet_03v3
**devattr s=44000,1176 d=26000,604
X676 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t7 Vdd.t918 Vdd.t917 pfet_03v3
**devattr s=26000,604 d=44000,1176
X677 a_n8305_28099 a_n9861_28819.t4 Vss.t412 Vss.t411 nfet_03v3
**devattr s=17600,576 d=17600,576
X678 a_n3583_19209 SARlogic_0.d3.t10 a_n3767_19209 Vss.t639 nfet_03v3
**devattr s=10400,304 d=10400,304
X679 a_29583_28100 a_28027_28820.t5 Vdd.t357 Vdd.t356 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X680 SARlogic_0.dffrs_4.nand3_8.Z.t2 SARlogic_0.dffrs_4.d.t7 a_8543_7428 Vss.t617 nfet_03v3
**devattr s=10400,304 d=17600,576
X681 a_4841_29217.t0 a_4921_30169.t5 Vdd.t143 Vdd.t142 pfet_03v3
**devattr s=26000,604 d=44000,1176
X682 a_1167_28099 a_n389_28819.t4 Vss.t47 Vss.t46 nfet_03v3
**devattr s=17600,576 d=17600,576
X683 Vdd.t49 Clk_piso.t15 a_33257_29218.t0 Vdd.t48 pfet_03v3
**devattr s=26000,604 d=26000,604
X684 Vdd.t25 SARlogic_0.dffrs_1.nand3_8.Z.t5 SARlogic_0.dffrs_1.nand3_1.C.t2 Vdd.t24 pfet_03v3
**devattr s=26000,604 d=26000,604
X685 a_24049_33720 Vdd.t974 a_23865_33720 Vss.t475 nfet_03v3
**devattr s=10400,304 d=10400,304
X686 Vdd.t53 a_42729_29218.t5 adc_PISO_0.dffrs_5.Qb Vdd.t52 pfet_03v3
**devattr s=26000,604 d=26000,604
X687 a_n8305_28099 a_n9861_28819.t5 Vdd.t539 Vdd.t538 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X688 adc_PISO_0.dffrs_2.Qb adc_PISO_0.dffrs_2.Q.t6 Vdd.t355 Vdd.t354 pfet_03v3
**devattr s=44000,1176 d=26000,604
X689 adc_PISO_0.dffrs_1.Q.t2 Vdd.t619 Vdd.t621 Vdd.t620 pfet_03v3
**devattr s=44000,1176 d=26000,604
X690 a_20783_29264.t1 a_20111_28100 a_20971_29984 Vdd.t134 pfet_03v3
**devattr s=31200,704 d=52800,1376
X691 a_4841_31422.t0 Clk_piso.t16 Vdd.t51 Vdd.t50 pfet_03v3
**devattr s=26000,604 d=44000,1176
X692 a_5803_19210 SARlogic_0.d2.t10 Vss.t234 Vss.t233 nfet_03v3
**devattr s=17600,576 d=10400,304
X693 a_37687_30440 adc_PISO_0.2inmux_1.Bit.t8 Vss.t393 Vss.t392 nfet_03v3
**devattr s=17600,576 d=10400,304
X694 a_n4551_31514 a_n4631_31422.t7 Vss.t526 Vss.t525 nfet_03v3
**devattr s=17600,576 d=10400,304
X695 a_12585_14043 SARlogic_0.dffrs_5.nand3_8.Z.t5 a_12401_14043 Vss.t118 nfet_03v3
**devattr s=10400,304 d=10400,304
X696 Vss.t28 adc_PISO_0.2inmux_2.Bit.t7 a_n201_30439 Vss.t27 nfet_03v3
**devattr s=10400,304 d=17600,576
X697 a_24049_35925 a_23865_30170.t6 a_23865_35925 Vss.t121 nfet_03v3
**devattr s=10400,304 d=10400,304
X698 a_1167_28099 a_n389_28819.t5 Vdd.t63 Vdd.t62 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X699 SARlogic_0.dffrs_13.nand3_1.C.t0 Reset.t63 Vdd.t401 Vdd.t400 pfet_03v3
**devattr s=44000,1176 d=26000,604
X700 SARlogic_0.dffrs_12.nand3_8.C.t0 SARlogic_0.dffrs_12.nand3_6.C.t8 Vdd.t930 Vdd.t929 pfet_03v3
**devattr s=44000,1176 d=26000,604
X701 SARlogic_0.dffrs_10.nand3_8.C.t0 SARlogic_0.dffrs_10.nand3_8.Z Vdd.t19 Vdd.t18 pfet_03v3
**devattr s=26000,604 d=44000,1176
X702 SARlogic_0.dffrs_0.nand3_8.C.t2 SARlogic_0.dffrs_0.nand3_8.Z.t6 a_n7625_9633 Vss.t119 nfet_03v3
**devattr s=10400,304 d=17600,576
X703 SARlogic_0.dffrs_9.nand3_6.C.t3 SARlogic_0.dffrs_9.nand3_1.C Vdd.t285 Vdd.t284 pfet_03v3
**devattr s=44000,1176 d=26000,604
X704 a_n4551_33719 a_n4631_33627.t5 Vss.t421 Vss.t420 nfet_03v3
**devattr s=17600,576 d=10400,304
X705 SARlogic_0.dffrs_0.d.t2 SARlogic_0.dffrs_13.Qb.t7 Vdd.t938 Vdd.t937 pfet_03v3
**devattr s=26000,604 d=44000,1176
X706 a_14393_31515 a_14313_31423.t8 Vss.t587 Vss.t586 nfet_03v3
**devattr s=17600,576 d=10400,304
X707 adc_PISO_0.2inmux_1.OUT.t1 a_39727_29264.t5 Vdd.t902 Vdd.t901 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X708 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_2.Qb.t7 Vdd.t882 Vdd.t881 pfet_03v3
**devattr s=44000,1176 d=26000,604
X709 SARlogic_0.dffrs_4.Qb.t1 Reset.t64 Vdd.t403 Vdd.t402 pfet_03v3
**devattr s=26000,604 d=44000,1176
X710 SARlogic_0.dffrs_1.nand3_8.C.t2 SARlogic_0.dffrs_1.nand3_6.C.t7 Vdd.t275 Vdd.t274 pfet_03v3
**devattr s=44000,1176 d=26000,604
X711 a_9083_28820.t1 SARlogic_0.d3.t11 a_9271_28100 Vss.t638 nfet_03v3
**devattr s=10400,304 d=17600,576
X712 a_42809_30170.t0 a_42729_29218.t6 Vdd.t55 Vdd.t54 pfet_03v3
**devattr s=44000,1176 d=26000,604
X713 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t2 Vss.t224 nfet_03v3
**devattr s=20800,504 d=20800,504
X714 SARlogic_0.dffrs_11.Qb Reset.t65 Vdd.t405 Vdd.t404 pfet_03v3
**devattr s=26000,604 d=44000,1176
X715 SARlogic_0.dffrs_5.Q.t2 SARlogic_0.dffrs_5.Qb.t8 Vdd.t431 Vdd.t430 pfet_03v3
**devattr s=26000,604 d=44000,1176
X716 SARlogic_0.dffrs_5.nand3_8.C.t1 SARlogic_0.dffrs_5.nand3_8.Z.t6 a_12585_9633 Vss.t136 nfet_03v3
**devattr s=10400,304 d=17600,576
X717 SARlogic_0.dffrs_1.nand3_6.C.t3 SARlogic_0.dffrs_1.nand3_1.C.t4 Vdd.t423 Vdd.t422 pfet_03v3
**devattr s=44000,1176 d=26000,604
X718 a_23865_29310 a_23785_29218.t7 Vss.t141 Vss.t140 nfet_03v3
**devattr s=17600,576 d=10400,304
X719 Vdd.t217 SARlogic_0.dffrs_11.nand3_8.C.t6 SARlogic_0.dffrs_11.Qb Vdd.t216 pfet_03v3
**devattr s=26000,604 d=26000,604
X720 Vdd.t527 a_39055_30440 a_39915_29984 Vdd.t526 pfet_03v3
**devattr s=31200,704 d=52800,1376
X721 a_42729_29218.t0 a_42729_31423.t6 Vdd.t844 Vdd.t843 pfet_03v3
**devattr s=44000,1176 d=26000,604
X722 Vdd.t752 SARlogic_0.dffrs_5.nand3_6.C.t7 SARlogic_0.dffrs_5.Q.t0 Vdd.t751 pfet_03v3
**devattr s=26000,604 d=26000,604
X723 a_28027_28820.t0 SARlogic_0.d1.t10 a_28215_28100 Vss.t585 nfet_03v3
**devattr s=10400,304 d=17600,576
X724 a_n4631_29217.t3 a_n4551_30169.t6 a_n4367_31514 Vss.t649 nfet_03v3
**devattr s=10400,304 d=17600,576
X725 comparator_no_offsetcal_0.no_offsetLatch_0.Vq comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t17 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t2 Vss.t272 nfet_03v3
**devattr s=20800,504 d=20800,504
X726 a_29583_30440 a_28027_31160.t5 Vss.t606 Vss.t605 nfet_03v3
**devattr s=17600,576 d=17600,576
X727 SARlogic_0.dffrs_13.nand3_1.C.t3 SARlogic_0.dffrs_13.nand3_6.C.t7 Vdd.t828 Vdd.t827 pfet_03v3
**devattr s=26000,604 d=44000,1176
X728 SARlogic_0.dffrs_10.nand3_8.C.t3 SARlogic_0.dffrs_10.nand3_6.C.t9 Vdd.t129 Vdd.t128 pfet_03v3
**devattr s=44000,1176 d=26000,604
X729 a_n4631_31422.t0 Clk_piso.t17 a_n4367_33719 Vss.t36 nfet_03v3
**devattr s=10400,304 d=17600,576
X730 SARlogic_0.dffrs_4.d.t1 SARlogic_0.dffrs_3.Qb.t9 a_5987_11838 Vss.t311 nfet_03v3
**devattr s=10400,304 d=17600,576
X731 adc_PISO_0.dffrs_2.Q.t0 adc_PISO_0.dffrs_2.Qb a_16063_33720 Vss.t394 nfet_03v3
**devattr s=10400,304 d=17600,576
X732 a_n3065_33719 Vdd.t975 Vss.t474 Vss.t473 nfet_03v3
**devattr s=17600,576 d=10400,304
X733 SARlogic_0.dffrs_14.nand3_8.C.t0 SARlogic_0.dffrs_14.nand3_6.C.t9 Vdd.t481 Vdd.t480 pfet_03v3
**devattr s=44000,1176 d=26000,604
X734 a_n9861_31159.t1 inv2_0.out.t25 Vdd.t591 Vdd.t590 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X735 Piso_out.t1 adc_PISO_0.dffrs_5.Qb a_44479_33720 Vss.t374 nfet_03v3
**devattr s=10400,304 d=17600,576
X736 a_n2281_11838 Vdd.t976 Vss.t458 Vss.t457 nfet_03v3
**devattr s=17600,576 d=10400,304
X737 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t15 Vdd.t287 Vdd.t286 pfet_03v3
**devattr s=10400,304 d=10400,304
X738 a_n8305_30439 a_n9861_31159.t5 Vss.t255 Vss.t254 nfet_03v3
**devattr s=17600,576 d=17600,576
X739 a_16063_33720 a_14313_31423.t9 a_15879_33720 Vss.t588 nfet_03v3
**devattr s=10400,304 d=10400,304
X740 a_n2881_33719 a_n4631_31422.t8 a_n3065_33719 Vss.t527 nfet_03v3
**devattr s=10400,304 d=10400,304
X741 SARlogic_0.dffrs_2.nand3_8.C.t2 SARlogic_0.dffrs_2.nand3_8.Z.t7 a_459_9633 Vss.t165 nfet_03v3
**devattr s=10400,304 d=17600,576
X742 SARlogic_0.dffrs_2.Qb.t1 Reset.t66 Vdd.t407 Vdd.t406 pfet_03v3
**devattr s=26000,604 d=44000,1176
X743 Vss.t568 a_n10831_4320 Comp_out.t1 Vss.t567 nfet_03v3
**devattr s=9350,280 d=9350,280
X744 a_10639_28100 a_9083_28820.t5 Vss.t655 Vss.t654 nfet_03v3
**devattr s=17600,576 d=17600,576
X745 SARlogic_0.dffrs_1.nand3_8.C.t0 SARlogic_0.dffrs_1.nand3_8.Z.t6 Vdd.t27 Vdd.t26 pfet_03v3
**devattr s=26000,604 d=44000,1176
X746 SARlogic_0.dffrs_3.nand3_8.Z.t2 SARlogic_0.dffrs_2.Q.t7 a_4501_7428 Vss.t268 nfet_03v3
**devattr s=10400,304 d=17600,576
X747 SARlogic_0.dffrs_14.nand3_6.C.t0 SARlogic_0.dffrs_14.nand3_1.C Vdd.t87 Vdd.t86 pfet_03v3
**devattr s=44000,1176 d=26000,604
X748 Vss.t199 adc_PISO_0.dffrs_3.Q.t8 a_28215_30440 Vss.t198 nfet_03v3
**devattr s=10400,304 d=17600,576
X749 Vss.t81 a_36793_29020 a_37687_28100 Vss.t80 nfet_03v3
**devattr s=10400,304 d=17600,576
X750 a_1167_30439 a_n389_31159.t5 Vss.t338 Vss.t337 nfet_03v3
**devattr s=17600,576 d=17600,576
X751 Vdd.t932 SARlogic_0.dffrs_2.nand3_8.C.t6 SARlogic_0.dffrs_2.Qb.t2 Vdd.t931 pfet_03v3
**devattr s=26000,604 d=26000,604
X752 SARlogic_0.dffrs_5.nand3_8.Z.t3 SARlogic_0.dffrs_5.nand3_8.C.t7 Vdd.t531 Vdd.t530 pfet_03v3
**devattr s=44000,1176 d=26000,604
X753 SARlogic_0.dffrs_8.nand3_8.C.t2 SARlogic_0.dffrs_8.nand3_8.Z Vdd.t315 Vdd.t314 pfet_03v3
**devattr s=26000,604 d=44000,1176
X754 SARlogic_0.dffrs_1.nand3_6.C.t2 Clk.t24 Vdd.t581 Vdd.t580 pfet_03v3
**devattr s=26000,604 d=44000,1176
X755 SARlogic_0.dffrs_9.nand3_8.Z SAR_in.t8 Vdd.t543 Vdd.t542 pfet_03v3
**devattr s=26000,604 d=44000,1176
X756 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_8.C.t7 Vdd.t219 Vdd.t218 pfet_03v3
**devattr s=44000,1176 d=26000,604
X757 Vdd.t583 Clk.t25 SARlogic_0.dffrs_13.nand3_8.C.t0 Vdd.t582 pfet_03v3
**devattr s=26000,604 d=26000,604
X758 SARlogic_0.dffrs_1.nand3_8.C.t1 SARlogic_0.dffrs_1.nand3_8.Z.t7 a_n3583_9633 Vss.t146 nfet_03v3
**devattr s=10400,304 d=17600,576
X759 a_459_11838 Reset.t67 a_275_11838 Vss.t312 nfet_03v3
**devattr s=10400,304 d=10400,304
X760 SARlogic_0.dffrs_2.nand3_8.Z.t3 SARlogic_0.dffrs_2.nand3_8.C.t7 Vdd.t934 Vdd.t933 pfet_03v3
**devattr s=44000,1176 d=26000,604
X761 SARlogic_0.dffrs_11.nand3_6.C.t2 SARlogic_0.dffrs_12.Q.t9 a_12585_21414 Vss.t380 nfet_03v3
**devattr s=10400,304 d=17600,576
X762 Vdd.t409 Reset.t68 SARlogic_0.dffrs_11.nand3_6.C.t0 Vdd.t408 pfet_03v3
**devattr s=26000,604 d=26000,604
X763 Vdd.t920 SARlogic_0.dffrs_9.nand3_6.C.t8 SARlogic_0.d2.t3 Vdd.t919 pfet_03v3
**devattr s=26000,604 d=26000,604
X764 adc_PISO_0.dffrs_2.Qb Vdd.t977 a_16063_31516 Vss.t472 nfet_03v3
**devattr s=10400,304 d=17600,576
X765 a_n3767_17004 SARlogic_0.dffrs_7.nand3_8.C.t7 Vss.t59 Vss.t58 nfet_03v3
**devattr s=17600,576 d=10400,304
X766 Vdd.t618 Vdd.t616 SARlogic_0.dffrs_13.nand3_6.C.t2 Vdd.t617 pfet_03v3
**devattr s=26000,604 d=26000,604
X767 Vdd.t523 SARlogic_0.dffrs_4.nand3_8.C.t7 SARlogic_0.dffrs_4.Qb.t3 Vdd.t522 pfet_03v3
**devattr s=26000,604 d=26000,604
X768 adc_PISO_0.dffrs_5.Qb Vdd.t978 a_44479_31516 Vss.t471 nfet_03v3
**devattr s=10400,304 d=17600,576
X769 a_16063_31516 a_14313_29218.t7 a_15879_31516 Vss.t248 nfet_03v3
**devattr s=10400,304 d=10400,304
X770 a_6591_33719 a_4841_31422.t8 a_6407_33719 Vss.t276 nfet_03v3
**devattr s=10400,304 d=10400,304
X771 a_n4631_33627.t2 Vdd.t613 Vdd.t615 Vdd.t614 pfet_03v3
**devattr s=44000,1176 d=26000,604
X772 SARlogic_0.dffrs_0.nand3_1.C.t2 SARlogic_0.dffrs_0.nand3_6.C.t9 a_n7625_14043 Vss.t44 nfet_03v3
**devattr s=10400,304 d=17600,576
X773 a_42729_31423.t0 Clk_piso.t18 a_42993_33720 Vss.t37 nfet_03v3
**devattr s=10400,304 d=17600,576
X774 a_33337_30170.t0 adc_PISO_0.2inmux_5.OUT.t3 Vdd.t115 Vdd.t114 pfet_03v3
**devattr s=26000,604 d=44000,1176
X775 a_n3767_19209 SARlogic_0.dffrs_7.nand3_6.C.t9 Vss.t627 Vss.t626 nfet_03v3
**devattr s=17600,576 d=10400,304
X776 SARlogic_0.dffrs_11.nand3_1.C SARlogic_0.dffrs_11.nand3_6.C.t9 a_12585_23619 Vss.t430 nfet_03v3
**devattr s=10400,304 d=17600,576
X777 Vdd.t173 SARlogic_0.dffrs_11.nand3_8.Z SARlogic_0.dffrs_11.nand3_1.C Vdd.t172 pfet_03v3
**devattr s=26000,604 d=26000,604
X778 a_14577_33720 Vdd.t979 a_14393_33720 Vss.t470 nfet_03v3
**devattr s=10400,304 d=10400,304
X779 a_14313_31423.t3 a_14313_33628.t5 Vdd.t333 Vdd.t332 pfet_03v3
**devattr s=44000,1176 d=26000,604
X780 a_n2281_9634 SARlogic_0.dffrs_2.d.t6 Vss.t18 Vss.t17 nfet_03v3
**devattr s=17600,576 d=10400,304
X781 a_n7625_9633 Clk.t26 a_n7809_9633 Vss.t434 nfet_03v3
**devattr s=10400,304 d=10400,304
X782 a_14393_30170.t0 adc_PISO_0.2inmux_3.OUT.t3 a_14577_29310 Vss.t633 nfet_03v3
**devattr s=10400,304 d=17600,576
X783 a_11311_29264.t1 a_10639_28100 a_11499_29984 Vdd.t594 pfet_03v3
**devattr s=31200,704 d=52800,1376
X784 a_42729_33628.t3 a_42729_31423.t7 a_42993_35925 Vss.t604 nfet_03v3
**devattr s=10400,304 d=17600,576
X785 a_4501_21414 Reset.t69 a_4317_21414 Vss.t313 nfet_03v3
**devattr s=10400,304 d=10400,304
X786 a_33257_29218.t3 a_33337_30170.t7 Vdd.t818 Vdd.t817 pfet_03v3
**devattr s=26000,604 d=44000,1176
X787 SARlogic_0.dffrs_1.nand3_1.C.t3 Vdd.t607 Vdd.t609 Vdd.t608 pfet_03v3
**devattr s=44000,1176 d=26000,604
X788 a_n9429_n2007.t12 Vin1.t6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t10 Vss.t182 nfet_03v3
**devattr s=15600,404 d=15600,404
X789 SARlogic_0.dffrs_8.nand3_8.C.t3 SARlogic_0.dffrs_8.nand3_6.C.t9 Vdd.t193 Vdd.t192 pfet_03v3
**devattr s=44000,1176 d=26000,604
X790 a_39915_29984 a_39055_30440 Vdd.t525 Vdd.t524 pfet_03v3
**devattr s=52800,1376 d=31200,704
X791 a_14577_35925 a_14393_30170.t7 a_14393_35925 Vss.t610 nfet_03v3
**devattr s=10400,304 d=10400,304
X792 a_14313_33628.t1 Vdd.t610 Vdd.t612 Vdd.t611 pfet_03v3
**devattr s=44000,1176 d=26000,604
X793 a_n10151_11838 SARlogic_0.dffrs_13.nand3_6.C.t8 a_n10335_11838 Vss.t596 nfet_03v3
**devattr s=10400,304 d=10400,304
X794 a_5987_19210 SARlogic_0.dffrs_9.nand3_8.C.t6 a_5803_19210 Vss.t45 nfet_03v3
**devattr s=10400,304 d=10400,304
X795 a_4501_23619 SARlogic_0.dffrs_9.nand3_8.Z a_4317_23619 Vss.t126 nfet_03v3
**devattr s=10400,304 d=10400,304
X796 SARlogic_0.dffrs_9.nand3_8.Z SARlogic_0.dffrs_9.nand3_8.C.t7 Vdd.t61 Vdd.t60 pfet_03v3
**devattr s=44000,1176 d=26000,604
X797 Vdd.t289 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t16 comparator_no_offsetcal_0.x5.out Vdd.t288 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X798 a_n3583_7428 Reset.t70 a_n3767_7428 Vss.t314 nfet_03v3
**devattr s=10400,304 d=10400,304
X799 Vdd.t9 Vss.t679 SARlogic_0.dffrs_12.nand3_8.C.t1 Vdd.t8 pfet_03v3
**devattr s=26000,604 d=26000,604
X800 a_5105_31514 Clk_piso.t19 a_4921_31514 Vss.t242 nfet_03v3
**devattr s=10400,304 d=10400,304
X801 SARlogic_0.dffrs_7.nand3_8.Z SAR_in.t9 a_n3583_17004 Vss.t415 nfet_03v3
**devattr s=10400,304 d=17600,576
X802 adc_PISO_0.2inmux_2.OUT.t1 a_1839_29263.t5 Vdd.t345 Vdd.t344 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X803 a_4921_31514 a_4841_31422.t9 Vss.t278 Vss.t277 nfet_03v3
**devattr s=17600,576 d=10400,304
X804 a_20783_29264.t3 a_20111_28100 Vss.t112 Vss.t111 nfet_03v3
**devattr s=17600,576 d=17600,576
X805 a_5105_33719 Vdd.t980 a_4921_33719 Vss.t469 nfet_03v3
**devattr s=10400,304 d=10400,304
X806 a_n4631_33627.t1 a_n4631_31422.t9 Vdd.t738 Vdd.t737 pfet_03v3
**devattr s=26000,604 d=44000,1176
X807 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t9 Vin1.t7 a_n9429_n2007.t13 Vss.t183 nfet_03v3
**devattr s=15600,404 d=15600,404
X808 SARlogic_0.dffrs_2.Qb.t0 Reset.t71 a_1945_9634 Vss.t315 nfet_03v3
**devattr s=10400,304 d=17600,576
X809 a_33337_30170.t1 a_33257_29218.t7 Vdd.t187 Vdd.t186 pfet_03v3
**devattr s=44000,1176 d=26000,604
X810 a_42993_31515 Clk_piso.t20 a_42809_31515 Vss.t243 nfet_03v3
**devattr s=10400,304 d=10400,304
X811 a_8543_14043 SARlogic_0.dffrs_4.nand3_8.Z.t7 a_8359_14043 Vss.t335 nfet_03v3
**devattr s=10400,304 d=10400,304
X812 SARlogic_0.dffrs_7.nand3_8.C.t1 SARlogic_0.dffrs_7.nand3_8.Z a_n3583_19209 Vss.t160 nfet_03v3
**devattr s=10400,304 d=17600,576
X813 a_28215_28100 a_27321_29020 Vss.t263 Vss.t262 nfet_03v3
**devattr s=17600,576 d=10400,304
X814 adc_PISO_0.2inmux_3.OUT.t1 a_11311_29264.t5 Vdd.t179 Vdd.t178 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X815 a_4921_33719 a_4841_33627.t5 Vss.t280 Vss.t279 nfet_03v3
**devattr s=17600,576 d=10400,304
X816 a_n7809_7428 SARlogic_0.dffrs_0.nand3_8.C.t7 Vss.t12 Vss.t11 nfet_03v3
**devattr s=17600,576 d=10400,304
X817 Vss.t566 a_n10831_4320 Comp_out.t0 Vss.t565 nfet_03v3
**devattr s=9350,280 d=9350,280
X818 SARlogic_0.dffrs_13.Qb.t2 Vdd.t981 a_n10151_9634 Vss.t468 nfet_03v3
**devattr s=10400,304 d=17600,576
X819 SARlogic_0.dffrs_1.nand3_1.C.t1 SARlogic_0.dffrs_1.nand3_6.C.t8 Vdd.t277 Vdd.t276 pfet_03v3
**devattr s=26000,604 d=44000,1176
X820 a_17849_29020 inv2_0.out.t26 Vss.t443 Vss.t442 nfet_03v3
**devattr s=17600,576 d=17600,576
X821 a_33257_29218.t1 a_33257_31423.t9 Vdd.t744 Vdd.t743 pfet_03v3
**devattr s=44000,1176 d=26000,604
X822 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t8 Vin1.t8 a_n9429_n2007.t14 Vss.t192 nfet_03v3
**devattr s=15600,404 d=15600,404
X823 a_24049_29310 Vdd.t982 a_23865_29310 Vss.t467 nfet_03v3
**devattr s=10400,304 d=10400,304
X824 a_n4367_31514 Clk_piso.t21 a_n4551_31514 Vss.t244 nfet_03v3
**devattr s=10400,304 d=10400,304
X825 adc_PISO_0.dffrs_0.Qb adc_PISO_0.2inmux_2.Bit.t8 Vdd.t39 Vdd.t38 pfet_03v3
**devattr s=44000,1176 d=26000,604
X826 SARlogic_0.dffrs_3.Qb.t1 Reset.t72 Vdd.t411 Vdd.t410 pfet_03v3
**devattr s=26000,604 d=44000,1176
X827 a_n9429_n2007.t21 Clk.t27 Vss.t436 Vss.t435 nfet_03v3
**devattr s=8320,264 d=8320,264
X828 SARlogic_0.dffrs_1.Qb.t0 SARlogic_0.dffrs_2.d.t7 Vdd.t33 Vdd.t32 pfet_03v3
**devattr s=44000,1176 d=26000,604
X829 a_n389_28819.t2 SARlogic_0.d4.t9 a_n201_28099 Vss.t175 nfet_03v3
**devattr s=10400,304 d=17600,576
X830 Vdd.t764 SARlogic_0.dffrs_13.nand3_8.Z.t7 SARlogic_0.dffrs_13.nand3_1.C.t1 Vdd.t763 pfet_03v3
**devattr s=26000,604 d=26000,604
X831 Vdd.t271 a_n4631_29217.t6 adc_PISO_0.dffrs_0.Qb Vdd.t270 pfet_03v3
**devattr s=26000,604 d=26000,604
X832 Vdd.t413 Reset.t73 SARlogic_0.dffrs_5.nand3_8.Z.t0 Vdd.t412 pfet_03v3
**devattr s=26000,604 d=26000,604
X833 a_n4367_33719 Vdd.t983 a_n4551_33719 Vss.t466 nfet_03v3
**devattr s=10400,304 d=10400,304
X834 a_n3583_11838 Reset.t74 a_n3767_11838 Vss.t316 nfet_03v3
**devattr s=10400,304 d=10400,304
X835 SARlogic_0.dffrs_14.nand3_8.Z SARlogic_0.dffrs_14.nand3_8.C.t7 Vdd.t748 Vdd.t747 pfet_03v3
**devattr s=44000,1176 d=26000,604
X836 a_n4551_29309 a_n4631_29217.t7 Vss.t215 Vss.t214 nfet_03v3
**devattr s=17600,576 d=10400,304
X837 a_n9429_n2007.t9 Vin2.t8 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vss.t194 nfet_03v3
**devattr s=15600,404 d=15600,404
X838 a_n389_28819.t3 SARlogic_0.d4.t10 Vdd.t223 Vdd.t222 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X839 a_30443_29984 a_29583_28100 a_30255_29264.t2 Vdd.t300 pfet_03v3
**devattr s=52800,1376 d=31200,704
X840 Vdd.t415 Reset.t75 SARlogic_0.dffrs_2.nand3_8.Z.t2 Vdd.t414 pfet_03v3
**devattr s=26000,604 d=26000,604
X841 a_n11821_11838 SARlogic_0.dffrs_13.nand3_1.C.t5 Vss.t228 Vss.t227 nfet_03v3
**devattr s=17600,576 d=10400,304
X842 SARlogic_0.dffrs_5.nand3_8.C.t2 SARlogic_0.dffrs_5.nand3_8.Z.t7 Vdd.t177 Vdd.t176 pfet_03v3
**devattr s=26000,604 d=44000,1176
X843 Vss.t129 a_n8305_30439 a_n7633_29263.t0 Vss.t128 nfet_03v3
**devattr s=17600,576 d=17600,576
X844 SARlogic_0.dffrs_14.nand3_8.C.t2 SARlogic_0.dffrs_14.nand3_8.Z Vdd.t205 Vdd.t204 pfet_03v3
**devattr s=26000,604 d=44000,1176
X845 comparator_no_offsetcal_0.no_offsetLatch_0.Vq Vin2.t9 a_n9429_n2007.t10 Vss.t195 nfet_03v3
**devattr s=15600,404 d=15600,404
X846 Vdd.t417 Reset.t76 SARlogic_0.dffrs_11.nand3_8.Z Vdd.t416 pfet_03v3
**devattr s=26000,604 d=26000,604
X847 SARlogic_0.dffrs_5.nand3_6.C.t3 Clk.t28 Vdd.t585 Vdd.t584 pfet_03v3
**devattr s=26000,604 d=44000,1176
X848 SARlogic_0.dffrs_14.nand3_6.C.t2 SARlogic_0.d4.t11 Vdd.t249 Vdd.t248 pfet_03v3
**devattr s=26000,604 d=44000,1176
X849 SARlogic_0.d5.t3 SARlogic_0.dffrs_13.Qb.t8 Vdd.t940 Vdd.t939 pfet_03v3
**devattr s=44000,1176 d=26000,604
X850 Vdd.t321 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t320 pfet_03v3
**devattr s=17600,576 d=17600,576
X851 a_n9673_28099 SARlogic_0.d5.t7 a_n9861_28819.t1 Vss.t85 nfet_03v3
**devattr s=17600,576 d=10400,304
X852 adc_PISO_0.dffrs_1.Qb Vdd.t984 a_6591_31515 Vss.t465 nfet_03v3
**devattr s=10400,304 d=17600,576
X853 Vdd.t227 a_4841_29217.t6 adc_PISO_0.dffrs_1.Qb Vdd.t226 pfet_03v3
**devattr s=26000,604 d=26000,604
X854 a_11499_29984 a_10639_30440 Vdd.t904 Vdd.t903 pfet_03v3
**devattr s=52800,1376 d=31200,704
X855 a_23865_30170.t3 adc_PISO_0.2inmux_4.OUT.t3 Vdd.t820 Vdd.t819 pfet_03v3
**devattr s=26000,604 d=44000,1176
X856 SARlogic_0.d0.t3 SARlogic_0.dffrs_4.Qb.t8 Vdd.t862 Vdd.t861 pfet_03v3
**devattr s=44000,1176 d=26000,604
X857 Vss.t345 comparator_no_offsetcal_0.x5.out comparator_no_offsetcal_0.x2.Vout2 Vss.t344 nfet_03v3
**devattr s=17600,576 d=17600,576
X858 a_18743_30440 inv2_0.out.t27 a_18555_31160.t1 Vss.t444 nfet_03v3
**devattr s=17600,576 d=10400,304
X859 Vdd.t587 Clk.t29 SARlogic_0.dffrs_3.nand3_8.C.t3 Vdd.t586 pfet_03v3
**devattr s=26000,604 d=26000,604
X860 a_n9429_n2007.t15 Vin1.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t7 Vss.t178 nfet_03v3
**devattr s=15600,404 d=15600,404
X861 Piso_out.t3 Vdd.t604 Vdd.t606 Vdd.t605 pfet_03v3
**devattr s=44000,1176 d=26000,604
X862 a_44479_33720 a_42729_31423.t8 a_44295_33720 Vss.t122 nfet_03v3
**devattr s=10400,304 d=10400,304
X863 a_n2097_11838 SARlogic_0.dffrs_1.nand3_6.C.t9 a_n2281_11838 Vss.t220 nfet_03v3
**devattr s=10400,304 d=10400,304
X864 a_n7625_14043 SARlogic_0.dffrs_0.nand3_8.Z.t7 a_n7809_14043 Vss.t573 nfet_03v3
**devattr s=10400,304 d=10400,304
X865 adc_PISO_0.2inmux_2.Bit.t2 adc_PISO_0.dffrs_0.Qb a_n2881_33719 Vss.t637 nfet_03v3
**devattr s=10400,304 d=17600,576
X866 a_15879_33720 Vdd.t985 Vss.t464 Vss.t463 nfet_03v3
**devattr s=17600,576 d=10400,304
X867 a_23785_29218.t1 a_23865_30170.t7 Vdd.t155 Vdd.t154 pfet_03v3
**devattr s=26000,604 d=44000,1176
X868 a_n4551_30169.t3 adc_PISO_0.2inmux_0.OUT.t3 a_n4367_29309 Vss.t544 nfet_03v3
**devattr s=10400,304 d=17600,576
X869 Vdd.t145 a_4921_30169.t6 a_4841_33627.t0 Vdd.t144 pfet_03v3
**devattr s=26000,604 d=26000,604
X870 Vdd.t419 Reset.t77 SARlogic_0.dffrs_3.nand3_6.C.t0 Vdd.t418 pfet_03v3
**devattr s=26000,604 d=26000,604
X871 Vdd.t603 Vdd.t601 a_42729_31423.t3 Vdd.t602 pfet_03v3
**devattr s=26000,604 d=26000,604
X872 Vdd.t15 SARlogic_0.dffrs_13.nand3_8.C.t7 SARlogic_0.dffrs_13.Qb.t0 Vdd.t14 pfet_03v3
**devattr s=26000,604 d=26000,604
X873 SARlogic_0.dffrs_2.d.t1 SARlogic_0.dffrs_1.Qb.t9 a_n2097_11838 Vss.t379 nfet_03v3
**devattr s=10400,304 d=17600,576
X874 a_n3767_7428 SARlogic_0.dffrs_1.nand3_8.C.t7 Vss.t343 Vss.t342 nfet_03v3
**devattr s=17600,576 d=10400,304
X875 a_4841_33627.t1 Vdd.t598 Vdd.t600 Vdd.t599 pfet_03v3
**devattr s=44000,1176 d=26000,604
X876 SARlogic_0.dffrs_9.nand3_6.C.t0 SARlogic_0.d1.t11 a_4501_21414 Vss.t453 nfet_03v3
**devattr s=10400,304 d=17600,576
X877 a_5803_21414 SARlogic_0.dffrs_2.Qb.t8 Vss.t632 Vss.t631 nfet_03v3
**devattr s=17600,576 d=10400,304
X878 a_12401_21414 SARlogic_0.dffrs_11.nand3_1.C Vss.t347 Vss.t346 nfet_03v3
**devattr s=17600,576 d=10400,304
X879 a_8543_9633 Clk.t30 a_8359_9633 Vss.t437 nfet_03v3
**devattr s=10400,304 d=10400,304
X880 Vdd.t421 Reset.t78 SARlogic_0.dffrs_10.nand3_6.C.t0 Vdd.t420 pfet_03v3
**devattr s=26000,604 d=26000,604
X881 Vdd.t297 SARlogic_0.d2.t11 SARlogic_0.dffrs_8.nand3_8.C.t0 Vdd.t296 pfet_03v3
**devattr s=26000,604 d=26000,604
X882 SARlogic_0.dffrs_13.nand3_6.C.t0 Clk.t31 a_n11637_11838 Vss.t438 nfet_03v3
**devattr s=10400,304 d=17600,576
X883 Vdd.t327 a_42809_30170.t7 a_42729_33628.t0 Vdd.t326 pfet_03v3
**devattr s=26000,604 d=26000,604
X884 a_20111_30440 a_18555_31160.t5 Vdd.t117 Vdd.t116 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X885 a_n10335_11838 Reset.t79 Vss.t318 Vss.t317 nfet_03v3
**devattr s=17600,576 d=10400,304
X886 a_n6693_1497 a_n6893_1405 Vdd.t497 Vdd.t496 pfet_03v3
**devattr s=10400,304 d=17600,576
X887 a_n6323_19213 SARlogic_0.d5.t8 Vss.t87 Vss.t86 nfet_03v3
**devattr s=17600,576 d=10400,304
X888 a_9845_9634 SARlogic_0.dffrs_4.Q.t7 Vss.t115 Vss.t114 nfet_03v3
**devattr s=17600,576 d=10400,304
X889 a_37499_31160.t3 inv2_0.out.t28 Vdd.t593 Vdd.t592 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X890 Vss.t651 a_n10567_29019 a_n9673_28099 Vss.t650 nfet_03v3
**devattr s=10400,304 d=17600,576
X891 Vdd.t17 SARlogic_0.dffrs_10.nand3_8.Z SARlogic_0.dffrs_10.nand3_1.C Vdd.t16 pfet_03v3
**devattr s=26000,604 d=26000,604
X892 SARlogic_0.dffrs_9.nand3_1.C SARlogic_0.dffrs_9.nand3_6.C.t9 a_4501_23619 Vss.t659 nfet_03v3
**devattr s=10400,304 d=17600,576
X893 a_12401_23619 SARlogic_0.dffrs_4.Qb.t9 Vss.t615 Vss.t614 nfet_03v3
**devattr s=17600,576 d=10400,304
X894 a_13887_19210 SARlogic_0.d0.t12 Vss.t207 Vss.t206 nfet_03v3
**devattr s=17600,576 d=10400,304
X895 a_n389_31159.t1 inv2_0.out.t29 a_n201_30439 Vss.t445 nfet_03v3
**devattr s=10400,304 d=17600,576
X896 a_4841_29217.t1 a_4921_30169.t7 a_5105_31514 Vss.t117 nfet_03v3
**devattr s=10400,304 d=17600,576
X897 a_11311_29264.t0 a_10639_28100 Vss.t450 Vss.t449 nfet_03v3
**devattr s=17600,576 d=17600,576
X898 SARlogic_0.d5.t2 SARlogic_0.dffrs_14.Qb Vdd.t203 Vdd.t202 pfet_03v3
**devattr s=26000,604 d=44000,1176
X899 a_33521_31515 Clk_piso.t22 a_33337_31515 Vss.t245 nfet_03v3
**devattr s=10400,304 d=10400,304
X900 adc_PISO_0.dffrs_5.Qb Piso_out.t5 Vdd.t29 Vdd.t28 pfet_03v3
**devattr s=44000,1176 d=26000,604
X901 a_44479_31516 a_42729_29218.t7 a_44295_31516 Vss.t19 nfet_03v3
**devattr s=10400,304 d=10400,304
X902 Vdd.t910 a_n4551_30169.t7 a_n4631_33627.t3 Vdd.t909 pfet_03v3
**devattr s=26000,604 d=26000,604
X903 a_4841_31422.t2 Clk_piso.t23 a_5105_33719 Vss.t440 nfet_03v3
**devattr s=10400,304 d=17600,576
X904 a_6407_33719 Vdd.t986 Vss.t462 Vss.t461 nfet_03v3
**devattr s=17600,576 d=10400,304
X905 a_15879_31516 adc_PISO_0.dffrs_2.Q.t7 Vss.t284 Vss.t283 nfet_03v3
**devattr s=17600,576 d=10400,304
X906 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t5 a_n9933_n1136 a_n10021_n1044 Vss.t368 nfet_03v3
**devattr s=26400,776 d=15600,404
X907 adc_PISO_0.2inmux_0.OUT.t0 a_n7633_29263.t5 Vss.t133 Vss.t132 nfet_03v3
**devattr s=17600,576 d=17600,576
X908 SARlogic_0.dffrs_11.nand3_8.Z SAR_in.t10 a_12585_17004 Vss.t416 nfet_03v3
**devattr s=10400,304 d=17600,576
X909 a_36793_29020 inv2_0.out.t30 Vss.t447 Vss.t446 nfet_03v3
**devattr s=17600,576 d=17600,576
X910 Vdd.t784 a_n10831_4320 Comp_out.t4 Vdd.t783 pfet_03v3
**devattr s=18700,450 d=18700,450
X911 SARlogic_0.dffrs_4.nand3_1.C.t2 SARlogic_0.dffrs_4.nand3_6.C.t9 a_8543_14043 Vss.t40 nfet_03v3
**devattr s=10400,304 d=17600,576
X912 a_42809_30170.t3 adc_PISO_0.2inmux_1.OUT.t3 a_42993_29310 Vss.t603 nfet_03v3
**devattr s=10400,304 d=17600,576
X913 a_14577_29310 Vdd.t987 a_14393_29310 Vss.t460 nfet_03v3
**devattr s=10400,304 d=10400,304
X914 SARlogic_0.dffrs_11.nand3_8.C.t0 SARlogic_0.dffrs_11.nand3_8.Z a_12585_19209 Vss.t134 nfet_03v3
**devattr s=10400,304 d=17600,576
X915 a_4317_21414 SARlogic_0.dffrs_9.nand3_1.C Vss.t226 Vss.t225 nfet_03v3
**devattr s=17600,576 d=10400,304
X916 SARlogic_0.dffrs_0.d.t3 SARlogic_0.dffrs_13.Qb.t9 a_n10151_11838 Vss.t672 nfet_03v3
**devattr s=10400,304 d=17600,576
X917 a_39055_30440 a_37499_31160.t5 Vdd.t567 Vdd.t566 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X918 Vdd.t167 a_29583_30440 a_30443_29984 Vdd.t166 pfet_03v3
**devattr s=31200,704 d=52800,1376
X919 a_4501_17004 Reset.t80 a_4317_17004 Vss.t319 nfet_03v3
**devattr s=10400,304 d=10400,304
X920 a_18555_28820.t2 SARlogic_0.d2.t12 a_18743_28100 Vss.t235 nfet_03v3
**devattr s=10400,304 d=17600,576
X921 SARlogic_0.dffrs_14.Qb Reset.t81 a_n6139_19213 Vss.t320 nfet_03v3
**devattr s=10400,304 d=17600,576
X922 a_n11821_9633 SARlogic_0.dffrs_13.nand3_6.C.t9 Vss.t602 Vss.t601 nfet_03v3
**devattr s=17600,576 d=10400,304
X923 SARlogic_0.dffrs_5.nand3_1.C.t1 SARlogic_0.dffrs_5.nand3_6.C.t8 Vdd.t754 Vdd.t753 pfet_03v3
**devattr s=26000,604 d=44000,1176
X924 a_4317_23619 SARlogic_0.dffrs_2.Qb.t9 Vss.t96 Vss.t95 nfet_03v3
**devattr s=17600,576 d=10400,304
X925 adc_PISO_0.2inmux_1.Bit.t3 adc_PISO_0.dffrs_4.Qb Vdd.t926 Vdd.t925 pfet_03v3
**devattr s=26000,604 d=44000,1176
X926 a_n9673_30439 inv2_0.out.t31 a_n9861_31159.t2 Vss.t448 nfet_03v3
**devattr s=17600,576 d=10400,304
X927 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t17 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t8 Vss.t229 nfet_03v3
**devattr s=20800,504 d=20800,504
X928 a_4501_19209 SARlogic_0.d1.t12 a_4317_19209 Vss.t454 nfet_03v3
**devattr s=10400,304 d=10400,304
X929 SARlogic_0.dffrs_5.Q.t1 SARlogic_0.dffrs_5.Qb.t9 a_14071_11838 Vss.t329 nfet_03v3
**devattr s=10400,304 d=17600,576
X930 a_n3767_11838 SARlogic_0.dffrs_1.nand3_1.C.t5 Vss.t322 Vss.t321 nfet_03v3
**devattr s=17600,576 d=10400,304
X931 Vdd.t553 SARlogic_0.dffrs_3.nand3_8.Z.t7 SARlogic_0.dffrs_3.nand3_1.C.t0 Vdd.t552 pfet_03v3
**devattr s=26000,604 d=26000,604
X932 a_42809_31515 a_42729_31423.t9 Vss.t124 Vss.t123 nfet_03v3
**devattr s=17600,576 d=10400,304
X933 a_14071_11838 SARlogic_0.dffrs_5.nand3_6.C.t9 a_13887_11838 Vss.t539 nfet_03v3
**devattr s=10400,304 d=10400,304
X934 Vss.t282 adc_PISO_0.dffrs_2.Q.t8 a_18743_30440 Vss.t281 nfet_03v3
**devattr s=10400,304 d=17600,576
X935 a_5105_29309 Vdd.t988 a_4921_29309 Vss.t459 nfet_03v3
**devattr s=10400,304 d=10400,304
X936 Vdd.t479 SARlogic_0.dffrs_12.nand3_6.C.t9 SARlogic_0.dffrs_12.Q.t0 Vdd.t478 pfet_03v3
**devattr s=26000,604 d=26000,604
X937 SARlogic_0.dffrs_13.nand3_8.Z.t0 Vss.t680 Vdd.t11 Vdd.t10 pfet_03v3
**devattr s=26000,604 d=44000,1176
X938 a_8359_14043 Vdd.t989 Vss.t456 Vss.t455 nfet_03v3
**devattr s=17600,576 d=10400,304
X939 a_4921_29309 a_4841_29217.t7 Vss.t170 Vss.t169 nfet_03v3
**devattr s=17600,576 d=10400,304
X940 SARlogic_0.dffrs_12.nand3_6.C.t2 Vss.t681 Vdd.t13 Vdd.t12 pfet_03v3
**devattr s=26000,604 d=44000,1176
X941 a_4501_9633 Clk.t32 a_4317_9633 Vss.t439 nfet_03v3
**devattr s=10400,304 d=10400,304
X942 a_9083_28820.t3 SARlogic_0.d3.t12 Vdd.t894 Vdd.t893 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X943 Vdd.t251 SARlogic_0.d4.t12 SARlogic_0.dffrs_14.nand3_8.C.t3 Vdd.t250 pfet_03v3
**devattr s=26000,604 d=26000,604
X944 Vdd.t269 adc_PISO_0.dffrs_1.Q.t8 a_9083_31160.t0 Vdd.t268 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X945 Vss.t99 Vss.t97 a_n9673_30439 Vss.t98 nfet_03v3
**devattr s=10400,304 d=17600,576
X946 SARlogic_0.dffrs_14.nand3_8.Z SAR_in.t11 Vdd.t545 Vdd.t544 pfet_03v3
**devattr s=26000,604 d=44000,1176
R0 SARlogic_0.d3.n3 SARlogic_0.d3.t8 41.0041
R1 SARlogic_0.d3.n4 SARlogic_0.d3.t4 40.8177
R2 SARlogic_0.d3.n7 SARlogic_0.d3.t7 40.6313
R3 SARlogic_0.d3.n1 SARlogic_0.d3.t12 34.2529
R4 SARlogic_0.d3.n6 SARlogic_0.dffrs_7.clk 33.3108
R5 SARlogic_0.d3.n7 SARlogic_0.d3.t5 27.3166
R6 SARlogic_0.d3.n4 SARlogic_0.d3.t10 27.1302
R7 SARlogic_0.d3.n3 SARlogic_0.d3.t9 26.9438
R8 SARlogic_0.d3.n0 SARlogic_0.d3.t6 19.673
R9 SARlogic_0.d3.n0 SARlogic_0.d3.t11 19.4007
R10 SARlogic_0.d3.n9 SARlogic_0.d3.n8 14.0582
R11 SARlogic_0.d3.n9 SARlogic_0.d3.n6 11.1633
R12 SARlogic_0.d3 SARlogic_0.d3.n2 10.6816
R13 SARlogic_0.d3.n12 SARlogic_0.d3.t2 10.0473
R14 SARlogic_0.d3.n2 SARlogic_0.d3.n1 8.05164
R15 SARlogic_0.d3.n11 SARlogic_0.d3.t1 6.51042
R16 SARlogic_0.d3.n11 SARlogic_0.d3.n10 6.04952
R17 SARlogic_0.dffrs_7.nand3_1.A SARlogic_0.d3.n3 5.7755
R18 SARlogic_0.dffrs_7.nand3_6.B SARlogic_0.d3.n4 5.47979
R19 SARlogic_0.d3.n8 SARlogic_0.d3.n7 5.13907
R20 SARlogic_0.dffrs_8.nand3_2.Z SARlogic_0.d3.n12 4.72925
R21 SARlogic_0.d3.n5 SARlogic_0.dffrs_7.nand3_6.B 2.17818
R22 SARlogic_0.d3.n6 SARlogic_0.d3 1.54657
R23 SARlogic_0.d3.n5 SARlogic_0.dffrs_7.nand3_1.A 1.34729
R24 SARlogic_0.d3.n12 SARlogic_0.d3.n11 0.732092
R25 SARlogic_0.d3.n10 SARlogic_0.d3.t0 0.7285
R26 SARlogic_0.d3.n10 SARlogic_0.d3.t3 0.7285
R27 SARlogic_0.dffrs_7.clk SARlogic_0.d3.n5 0.610571
R28 SARlogic_0.dffrs_8.nand3_2.Z SARlogic_0.d3.n9 0.166901
R29 SARlogic_0.d3.n1 SARlogic_0.d3.n0 0.106438
R30 SARlogic_0.d3.n8 SARlogic_0.dffrs_8.nand3_7.C 0.0455
R31 SARlogic_0.d3.n2 adc_PISO_0.2inmux_3.In 0.0455
R32 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t6 40.8177
R33 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t5 40.6313
R34 SARlogic_0.dffrs_7.nand3_8.C.n1 SARlogic_0.dffrs_7.nand3_8.C.t7 27.3166
R35 SARlogic_0.dffrs_7.nand3_8.C.n0 SARlogic_0.dffrs_7.nand3_8.C.t4 27.1302
R36 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_8.C.n2 14.119
R37 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.t1 10.0473
R38 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.t0 6.51042
R39 SARlogic_0.dffrs_7.nand3_8.C.n5 SARlogic_0.dffrs_7.nand3_8.C.n4 6.04952
R40 SARlogic_0.dffrs_7.nand3_7.B SARlogic_0.dffrs_7.nand3_8.C.n0 5.47979
R41 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C.n1 5.13907
R42 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n6 4.72925
R43 SARlogic_0.dffrs_7.nand3_8.C.n6 SARlogic_0.dffrs_7.nand3_8.C.n5 0.732092
R44 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t3 0.7285
R45 SARlogic_0.dffrs_7.nand3_8.C.n4 SARlogic_0.dffrs_7.nand3_8.C.t2 0.7285
R46 SARlogic_0.dffrs_7.nand3_8.C.n3 SARlogic_0.dffrs_7.nand3_7.B 0.438233
R47 SARlogic_0.dffrs_7.nand3_6.Z SARlogic_0.dffrs_7.nand3_8.C.n3 0.166901
R48 SARlogic_0.dffrs_7.nand3_8.C.n2 SARlogic_0.dffrs_7.nand3_8.C 0.0455
R49 Vdd.n1020 Vdd.t342 869.717
R50 Vdd.n1009 Vdd.t288 869.717
R51 Vdd.t282 Vdd.t496 490.324
R52 Vdd.t286 Vdd.t282 490.324
R53 Vdd.t390 Vdd.t286 490.324
R54 Vdd.t340 Vdd.t390 490.324
R55 Vdd.t278 Vdd.t340 490.324
R56 Vdd.t280 Vdd.t278 490.324
R57 Vdd.t392 Vdd.t280 490.324
R58 Vdd.t338 Vdd.t392 490.324
R59 Vdd.t488 Vdd.t338 490.324
R60 Vdd.t496 Vdd.n1056 467.743
R61 Vdd.n1058 Vdd.t488 467.743
R62 Vdd.n1059 Vdd.t78 398.652
R63 Vdd.n1041 Vdd.t576 398.652
R64 Vdd.t78 Vdd.n1058 389.878
R65 Vdd.n1056 Vdd.t576 389.878
R66 Vdd.t320 Vdd.n1013 372.543
R67 Vdd.n1016 Vdd.t242 372.543
R68 Vdd.n1015 Vdd.t320 370.969
R69 Vdd.t242 Vdd.n1015 370.969
R70 Vdd.n1036 Vdd.n1034 287.351
R71 Vdd.n1037 Vdd.n1035 287.351
R72 Vdd.t785 Vdd.t783 265.625
R73 Vdd.t865 Vdd.n4 250.9
R74 Vdd.n5 Vdd.t668 250.9
R75 Vdd.t873 Vdd.n1095 250.9
R76 Vdd.n1096 Vdd.t94 250.9
R77 Vdd.t516 Vdd.n9 250.9
R78 Vdd.n10 Vdd.t689 250.9
R79 Vdd.t154 Vdd.n1083 250.9
R80 Vdd.n1084 Vdd.t863 250.9
R81 Vdd.t662 Vdd.n1089 250.9
R82 Vdd.n1090 Vdd.t252 250.9
R83 Vdd.t819 Vdd.n1076 250.9
R84 Vdd.n1077 Vdd.t180 250.9
R85 Vdd.t839 Vdd.n51 250.9
R86 Vdd.n52 Vdd.t716 250.9
R87 Vdd.t232 Vdd.n62 250.9
R88 Vdd.n63 Vdd.t130 250.9
R89 Vdd.t486 Vdd.n57 250.9
R90 Vdd.n58 Vdd.t605 250.9
R91 Vdd.t324 Vdd.n74 250.9
R92 Vdd.n75 Vdd.t843 250.9
R93 Vdd.t644 Vdd.n68 250.9
R94 Vdd.n69 Vdd.t28 250.9
R95 Vdd.t837 Vdd.n85 250.9
R96 Vdd.n86 Vdd.t54 250.9
R97 Vdd.t739 Vdd.n124 250.9
R98 Vdd.n125 Vdd.t695 250.9
R99 Vdd.t851 Vdd.n135 250.9
R100 Vdd.n136 Vdd.t795 250.9
R101 Vdd.t925 Vdd.n130 250.9
R102 Vdd.n131 Vdd.t707 250.9
R103 Vdd.t817 Vdd.n147 250.9
R104 Vdd.n148 Vdd.t743 250.9
R105 Vdd.t731 Vdd.n141 250.9
R106 Vdd.n142 Vdd.t512 250.9
R107 Vdd.t114 Vdd.n158 250.9
R108 Vdd.n159 Vdd.t186 250.9
R109 Vdd.t514 Vdd.n204 250.9
R110 Vdd.n205 Vdd.t626 250.9
R111 Vdd.t647 Vdd.n209 250.9
R112 Vdd.n210 Vdd.t354 250.9
R113 Vdd.t927 Vdd.n198 250.9
R114 Vdd.n199 Vdd.t426 250.9
R115 Vdd.t12 Vdd.n1001 250.9
R116 Vdd.n1002 Vdd.t102 250.9
R117 Vdd.t506 Vdd.n984 250.9
R118 Vdd.n985 Vdd.t428 250.9
R119 Vdd.t757 Vdd.n989 250.9
R120 Vdd.n990 Vdd.t929 250.9
R121 Vdd.t364 Vdd.n995 250.9
R122 Vdd.n996 Vdd.t498 250.9
R123 Vdd.t4 Vdd.n977 250.9
R124 Vdd.n978 Vdd.t508 250.9
R125 Vdd.t815 Vdd.n505 250.9
R126 Vdd.n506 Vdd.t611 250.9
R127 Vdd.t877 Vdd.n511 250.9
R128 Vdd.n512 Vdd.t332 250.9
R129 Vdd.t853 Vdd.n517 250.9
R130 Vdd.n518 Vdd.t546 250.9
R131 Vdd.t883 Vdd.n968 250.9
R132 Vdd.n969 Vdd.t306 250.9
R133 Vdd.t484 Vdd.n754 250.9
R134 Vdd.n755 Vdd.t935 250.9
R135 Vdd.t801 Vdd.n793 250.9
R136 Vdd.n794 Vdd.t198 250.9
R137 Vdd.t40 Vdd.n831 250.9
R138 Vdd.n832 Vdd.t492 250.9
R139 Vdd.t917 Vdd.n869 250.9
R140 Vdd.n870 Vdd.t881 250.9
R141 Vdd.t124 Vdd.n908 250.9
R142 Vdd.n909 Vdd.t396 250.9
R143 Vdd.t572 Vdd.n946 250.9
R144 Vdd.n947 Vdd.t859 250.9
R145 Vdd.t248 Vdd.n672 250.9
R146 Vdd.n673 Vdd.t86 250.9
R147 Vdd.t202 Vdd.n765 250.9
R148 Vdd.n766 Vdd.t939 250.9
R149 Vdd.t895 Vdd.n398 250.9
R150 Vdd.n399 Vdd.t424 250.9
R151 Vdd.t540 Vdd.n804 250.9
R152 Vdd.n805 Vdd.t194 250.9
R153 Vdd.t292 Vdd.n368 250.9
R154 Vdd.n369 Vdd.t328 250.9
R155 Vdd.t240 Vdd.n842 250.9
R156 Vdd.n843 Vdd.t490 250.9
R157 Vdd.t809 Vdd.n338 250.9
R158 Vdd.n339 Vdd.t284 250.9
R159 Vdd.t88 Vdd.n881 250.9
R160 Vdd.n882 Vdd.t879 250.9
R161 Vdd.t258 Vdd.n302 250.9
R162 Vdd.n303 Vdd.t108 250.9
R163 Vdd.t749 Vdd.n919 250.9
R164 Vdd.n920 Vdd.t394 250.9
R165 Vdd.t534 Vdd.n272 250.9
R166 Vdd.n273 Vdd.t446 250.9
R167 Vdd.t132 Vdd.n957 250.9
R168 Vdd.n958 Vdd.t861 250.9
R169 Vdd.t204 Vdd.n749 250.9
R170 Vdd.n750 Vdd.t480 250.9
R171 Vdd.t466 Vdd.n662 250.9
R172 Vdd.n663 Vdd.t120 250.9
R173 Vdd.t210 Vdd.n788 250.9
R174 Vdd.n789 Vdd.t797 250.9
R175 Vdd.t384 Vdd.n388 250.9
R176 Vdd.n389 Vdd.t220 250.9
R177 Vdd.t314 Vdd.n826 250.9
R178 Vdd.n827 Vdd.t192 250.9
R179 Vdd.t366 Vdd.n358 250.9
R180 Vdd.n359 Vdd.t897 250.9
R181 Vdd.t160 Vdd.n864 250.9
R182 Vdd.n865 Vdd.t915 250.9
R183 Vdd.t370 Vdd.n322 250.9
R184 Vdd.n323 Vdd.t290 250.9
R185 Vdd.t18 Vdd.n903 250.9
R186 Vdd.n904 Vdd.t128 250.9
R187 Vdd.t360 Vdd.n292 250.9
R188 Vdd.n293 Vdd.t807 250.9
R189 Vdd.t174 Vdd.n941 250.9
R190 Vdd.n942 Vdd.t568 250.9
R191 Vdd.t404 Vdd.n262 250.9
R192 Vdd.n263 Vdd.t260 250.9
R193 Vdd.t544 Vdd.n677 250.9
R194 Vdd.n678 Vdd.t747 250.9
R195 Vdd.t560 Vdd.n403 250.9
R196 Vdd.n404 Vdd.t92 250.9
R197 Vdd.t558 Vdd.n373 250.9
R198 Vdd.n374 Vdd.t310 250.9
R199 Vdd.t542 Vdd.n343 250.9
R200 Vdd.n344 Vdd.t60 250.9
R201 Vdd.t556 Vdd.n307 250.9
R202 Vdd.n308 Vdd.t244 250.9
R203 Vdd.t562 Vdd.n277 250.9
R204 Vdd.n278 Vdd.t218 250.9
R205 Vdd.t56 Vdd.n744 250.9
R206 Vdd.n745 Vdd.t701 250.9
R207 Vdd.t68 Vdd.n682 250.9
R208 Vdd.n683 Vdd.t596 250.9
R209 Vdd.t276 Vdd.n783 250.9
R210 Vdd.n784 Vdd.t608 250.9
R211 Vdd.t196 Vdd.n760 250.9
R212 Vdd.n761 Vdd.t692 250.9
R213 Vdd.t580 Vdd.n408 250.9
R214 Vdd.n409 Vdd.t422 250.9
R215 Vdd.t504 Vdd.n821 250.9
R216 Vdd.n822 Vdd.t656 250.9
R217 Vdd.t494 Vdd.n799 250.9
R218 Vdd.n800 Vdd.t650 250.9
R219 Vdd.t82 Vdd.n378 250.9
R220 Vdd.n379 Vdd.t476 250.9
R221 Vdd.t434 Vdd.n859 250.9
R222 Vdd.n860 Vdd.t704 250.9
R223 Vdd.t869 Vdd.n837 250.9
R224 Vdd.n838 Vdd.t674 250.9
R225 Vdd.t64 Vdd.n348 250.9
R226 Vdd.n349 Vdd.t188 250.9
R227 Vdd.t833 Vdd.n898 250.9
R228 Vdd.n899 Vdd.t665 250.9
R229 Vdd.t398 Vdd.n876 250.9
R230 Vdd.n877 Vdd.t722 250.9
R231 Vdd.t76 Vdd.n312 250.9
R232 Vdd.n313 Vdd.t104 250.9
R233 Vdd.t753 Vdd.n936 250.9
R234 Vdd.n937 Vdd.t710 250.9
R235 Vdd.t304 Vdd.n914 250.9
R236 Vdd.n915 Vdd.t671 250.9
R237 Vdd.t584 Vdd.n282 250.9
R238 Vdd.n283 Vdd.t238 250.9
R239 Vdd.t430 Vdd.n952 250.9
R240 Vdd.n953 Vdd.t686 250.9
R241 Vdd.t148 Vdd.n739 250.9
R242 Vdd.n740 Vdd.t564 250.9
R243 Vdd.t374 Vdd.n667 250.9
R244 Vdd.n668 Vdd.t0 250.9
R245 Vdd.t26 Vdd.n778 250.9
R246 Vdd.n779 Vdd.t274 250.9
R247 Vdd.t448 Vdd.n393 250.9
R248 Vdd.n394 Vdd.t32 250.9
R249 Vdd.t212 Vdd.n816 250.9
R250 Vdd.n817 Vdd.t500 250.9
R251 Vdd.t406 Vdd.n363 250.9
R252 Vdd.n364 Vdd.t336 250.9
R253 Vdd.t550 Vdd.n854 250.9
R254 Vdd.n855 Vdd.t432 250.9
R255 Vdd.t410 Vdd.n327 250.9
R256 Vdd.n328 Vdd.t813 250.9
R257 Vdd.t440 Vdd.n893 250.9
R258 Vdd.n894 Vdd.t831 250.9
R259 Vdd.t402 Vdd.n297 250.9
R260 Vdd.n298 Vdd.t138 250.9
R261 Vdd.t176 Vdd.n931 250.9
R262 Vdd.n932 Vdd.t921 250.9
R263 Vdd.t452 Vdd.n267 250.9
R264 Vdd.n268 Vdd.t536 250.9
R265 Vdd.t823 Vdd.n687 250.9
R266 Vdd.n688 Vdd.t20 250.9
R267 Vdd.t943 Vdd.n413 250.9
R268 Vdd.n414 Vdd.t444 250.9
R269 Vdd.t30 Vdd.n383 250.9
R270 Vdd.n384 Vdd.t933 250.9
R271 Vdd.t334 Vdd.n353 250.9
R272 Vdd.n354 Vdd.t110 250.9
R273 Vdd.t811 Vdd.n317 250.9
R274 Vdd.n318 Vdd.t520 250.9
R275 Vdd.t136 Vdd.n287 250.9
R276 Vdd.n288 Vdd.t530 250.9
R277 Vdd.t827 Vdd.n692 250.9
R278 Vdd.n693 Vdd.t400 250.9
R279 Vdd.t578 Vdd.n708 250.9
R280 Vdd.n709 Vdd.t923 250.9
R281 Vdd.t937 Vdd.n703 250.9
R282 Vdd.n704 Vdd.t386 250.9
R283 Vdd.t761 Vdd.n726 250.9
R284 Vdd.n727 Vdd.t825 250.9
R285 Vdd.t719 Vdd.n732 250.9
R286 Vdd.n733 Vdd.t793 250.9
R287 Vdd.t10 Vdd.n720 250.9
R288 Vdd.n721 Vdd.t885 250.9
R289 Vdd.t737 Vdd.n625 250.9
R290 Vdd.n626 Vdd.t614 250.9
R291 Vdd.t230 Vdd.n636 250.9
R292 Vdd.n637 Vdd.t554 250.9
R293 Vdd.t891 Vdd.n631 250.9
R294 Vdd.n632 Vdd.t653 250.9
R295 Vdd.t907 Vdd.n648 250.9
R296 Vdd.n649 Vdd.t733 250.9
R297 Vdd.t728 Vdd.n642 250.9
R298 Vdd.n643 Vdd.t38 250.9
R299 Vdd.t140 Vdd.n655 250.9
R300 Vdd.n656 Vdd.t941 250.9
R301 Vdd.t346 Vdd.n556 250.9
R302 Vdd.n557 Vdd.t599 250.9
R303 Vdd.t50 Vdd.n567 250.9
R304 Vdd.n568 Vdd.t228 250.9
R305 Vdd.t34 Vdd.n562 250.9
R306 Vdd.n563 Vdd.t620 250.9
R307 Vdd.t142 Vdd.n579 250.9
R308 Vdd.n580 Vdd.t350 250.9
R309 Vdd.t629 Vdd.n573 250.9
R310 Vdd.n574 Vdd.t266 250.9
R311 Vdd.t156 Vdd.n586 250.9
R312 Vdd.n587 Vdd.t224 250.9
R313 Vdd.n1027 Vdd.t322 242.189
R314 Vdd.n186 Vdd.t845 236.083
R315 Vdd.t773 Vdd.n183 236.083
R316 Vdd.t356 Vdd.n166 236.083
R317 Vdd.n172 Vdd.t803 236.083
R318 Vdd.n113 Vdd.t566 236.083
R319 Vdd.t592 Vdd.n110 236.083
R320 Vdd.t857 Vdd.n93 236.083
R321 Vdd.n99 Vdd.t262 236.083
R322 Vdd.n45 Vdd.t901 236.083
R323 Vdd.n39 Vdd.t524 236.083
R324 Vdd.n29 Vdd.t256 236.083
R325 Vdd.n23 Vdd.t168 236.083
R326 Vdd.t791 Vdd.n231 236.083
R327 Vdd.n237 Vdd.t294 236.083
R328 Vdd.n614 Vdd.t200 236.083
R329 Vdd.t769 Vdd.n611 236.083
R330 Vdd.t62 Vdd.n594 236.083
R331 Vdd.n600 Vdd.t222 236.083
R332 Vdd.n545 Vdd.t847 236.083
R333 Vdd.t771 Vdd.n542 236.083
R334 Vdd.t913 Vdd.n525 236.083
R335 Vdd.n531 Vdd.t893 236.083
R336 Vdd.n499 Vdd.t178 236.083
R337 Vdd.n493 Vdd.t903 236.083
R338 Vdd.n483 Vdd.t344 236.083
R339 Vdd.n477 Vdd.t889 236.083
R340 Vdd.t538 Vdd.n453 236.083
R341 Vdd.n459 Vdd.t122 236.083
R342 Vdd.t318 Vdd.n435 236.083
R343 Vdd.n445 Vdd.t590 236.083
R344 Vdd.t170 Vdd.n422 236.083
R345 Vdd.n433 Vdd.t164 236.083
R346 Vdd.t116 Vdd.n247 236.083
R347 Vdd.n251 Vdd.t779 236.083
R348 Vdd.t190 Vdd.n221 236.083
R349 Vdd.n223 Vdd.t98 236.083
R350 Vdd.t845 Vdd.n185 235.294
R351 Vdd.n185 Vdd.t773 235.294
R352 Vdd.n171 Vdd.t356 235.294
R353 Vdd.t803 Vdd.n171 235.294
R354 Vdd.t566 Vdd.n112 235.294
R355 Vdd.n112 Vdd.t592 235.294
R356 Vdd.n98 Vdd.t857 235.294
R357 Vdd.t262 Vdd.n98 235.294
R358 Vdd.t901 Vdd.n44 235.294
R359 Vdd.n44 Vdd.t389 235.294
R360 Vdd.t388 Vdd.n42 235.294
R361 Vdd.n42 Vdd.t526 235.294
R362 Vdd.t256 Vdd.n28 235.294
R363 Vdd.n28 Vdd.t301 235.294
R364 Vdd.t300 Vdd.n26 235.294
R365 Vdd.n26 Vdd.t166 235.294
R366 Vdd.n236 Vdd.t791 235.294
R367 Vdd.t294 Vdd.n236 235.294
R368 Vdd.t200 Vdd.n613 235.294
R369 Vdd.n613 Vdd.t769 235.294
R370 Vdd.n599 Vdd.t62 235.294
R371 Vdd.t222 Vdd.n599 235.294
R372 Vdd.t847 Vdd.n544 235.294
R373 Vdd.n544 Vdd.t771 235.294
R374 Vdd.n530 Vdd.t913 235.294
R375 Vdd.t893 Vdd.n530 235.294
R376 Vdd.t178 Vdd.n498 235.294
R377 Vdd.n498 Vdd.t594 235.294
R378 Vdd.t595 Vdd.n496 235.294
R379 Vdd.n496 Vdd.t905 235.294
R380 Vdd.t344 Vdd.n482 235.294
R381 Vdd.n482 Vdd.t299 235.294
R382 Vdd.t298 Vdd.n480 235.294
R383 Vdd.n480 Vdd.t887 235.294
R384 Vdd.n458 Vdd.t538 235.294
R385 Vdd.t122 Vdd.n458 235.294
R386 Vdd.n444 Vdd.t318 235.294
R387 Vdd.t590 Vdd.n444 235.294
R388 Vdd.n430 Vdd.t170 235.294
R389 Vdd.t303 Vdd.n430 235.294
R390 Vdd.n432 Vdd.t302 235.294
R391 Vdd.t162 Vdd.n432 235.294
R392 Vdd.n250 Vdd.t116 235.294
R393 Vdd.t779 Vdd.n250 235.294
R394 Vdd.n227 Vdd.t190 235.294
R395 Vdd.n227 Vdd.t134 235.294
R396 Vdd.t135 Vdd.n226 235.294
R397 Vdd.n226 Vdd.t100 235.294
R398 Vdd.t152 Vdd.t865 200
R399 Vdd.t668 Vdd.t152 200
R400 Vdd.t659 Vdd.t873 200
R401 Vdd.t94 Vdd.t659 200
R402 Vdd.t867 Vdd.t516 200
R403 Vdd.t689 Vdd.t867 200
R404 Vdd.t871 Vdd.t154 200
R405 Vdd.t863 Vdd.t871 200
R406 Vdd.t182 Vdd.t662 200
R407 Vdd.t252 Vdd.t182 200
R408 Vdd.t698 Vdd.t819 200
R409 Vdd.t180 Vdd.t698 200
R410 Vdd.t326 Vdd.t839 200
R411 Vdd.t716 Vdd.t326 200
R412 Vdd.t602 Vdd.t232 200
R413 Vdd.t130 Vdd.t602 200
R414 Vdd.t841 Vdd.t486 200
R415 Vdd.t605 Vdd.t841 200
R416 Vdd.t236 Vdd.t324 200
R417 Vdd.t843 Vdd.t236 200
R418 Vdd.t52 Vdd.t644 200
R419 Vdd.t28 Vdd.t52 200
R420 Vdd.t638 Vdd.t837 200
R421 Vdd.t54 Vdd.t638 200
R422 Vdd.t389 Vdd.t388 200
R423 Vdd.t524 Vdd.t526 200
R424 Vdd.t821 Vdd.t739 200
R425 Vdd.t695 Vdd.t821 200
R426 Vdd.t725 Vdd.t851 200
R427 Vdd.t795 Vdd.t725 200
R428 Vdd.t741 Vdd.t925 200
R429 Vdd.t707 Vdd.t741 200
R430 Vdd.t48 Vdd.t817 200
R431 Vdd.t743 Vdd.t48 200
R432 Vdd.t184 Vdd.t731 200
R433 Vdd.t512 Vdd.t184 200
R434 Vdd.t623 Vdd.t114 200
R435 Vdd.t186 Vdd.t623 200
R436 Vdd.t301 Vdd.t300 200
R437 Vdd.t168 Vdd.t166 200
R438 Vdd.t548 Vdd.t514 200
R439 Vdd.t626 Vdd.t548 200
R440 Vdd.t308 Vdd.t647 200
R441 Vdd.t354 Vdd.t308 200
R442 Vdd.t759 Vdd.t927 200
R443 Vdd.t426 Vdd.t759 200
R444 Vdd.t458 Vdd.t12 200
R445 Vdd.t102 Vdd.t458 200
R446 Vdd.t478 Vdd.t506 200
R447 Vdd.t428 Vdd.t478 200
R448 Vdd.t8 Vdd.t757 200
R449 Vdd.t929 Vdd.t8 200
R450 Vdd.t2 Vdd.t364 200
R451 Vdd.t498 Vdd.t2 200
R452 Vdd.t462 Vdd.t4 200
R453 Vdd.t508 Vdd.t462 200
R454 Vdd.t855 Vdd.t815 200
R455 Vdd.t611 Vdd.t855 200
R456 Vdd.t641 Vdd.t877 200
R457 Vdd.t332 Vdd.t641 200
R458 Vdd.t875 Vdd.t853 200
R459 Vdd.t546 Vdd.t875 200
R460 Vdd.t683 Vdd.t883 200
R461 Vdd.t306 Vdd.t683 200
R462 Vdd.t206 Vdd.t484 200
R463 Vdd.t935 Vdd.t206 200
R464 Vdd.t208 Vdd.t801 200
R465 Vdd.t198 Vdd.t208 200
R466 Vdd.t316 Vdd.t40 200
R467 Vdd.t492 Vdd.t316 200
R468 Vdd.t158 Vdd.t917 200
R469 Vdd.t881 Vdd.t158 200
R470 Vdd.t16 Vdd.t124 200
R471 Vdd.t396 Vdd.t16 200
R472 Vdd.t172 Vdd.t572 200
R473 Vdd.t859 Vdd.t172 200
R474 Vdd.t518 Vdd.t248 200
R475 Vdd.t86 Vdd.t518 200
R476 Vdd.t482 Vdd.t202 200
R477 Vdd.t939 Vdd.t482 200
R478 Vdd.t470 Vdd.t895 200
R479 Vdd.t424 Vdd.t470 200
R480 Vdd.t799 Vdd.t540 200
R481 Vdd.t194 Vdd.t799 200
R482 Vdd.t460 Vdd.t292 200
R483 Vdd.t328 Vdd.t460 200
R484 Vdd.t42 Vdd.t240 200
R485 Vdd.t490 Vdd.t42 200
R486 Vdd.t376 Vdd.t809 200
R487 Vdd.t284 Vdd.t376 200
R488 Vdd.t919 Vdd.t88 200
R489 Vdd.t879 Vdd.t919 200
R490 Vdd.t420 Vdd.t258 200
R491 Vdd.t108 Vdd.t420 200
R492 Vdd.t126 Vdd.t749 200
R493 Vdd.t394 Vdd.t126 200
R494 Vdd.t408 Vdd.t534 200
R495 Vdd.t446 Vdd.t408 200
R496 Vdd.t570 Vdd.t132 200
R497 Vdd.t861 Vdd.t570 200
R498 Vdd.t250 Vdd.t204 200
R499 Vdd.t480 Vdd.t250 200
R500 Vdd.t745 Vdd.t466 200
R501 Vdd.t120 Vdd.t745 200
R502 Vdd.t899 Vdd.t210 200
R503 Vdd.t797 Vdd.t899 200
R504 Vdd.t90 Vdd.t384 200
R505 Vdd.t220 Vdd.t90 200
R506 Vdd.t296 Vdd.t314 200
R507 Vdd.t192 Vdd.t296 200
R508 Vdd.t312 Vdd.t366 200
R509 Vdd.t897 Vdd.t312 200
R510 Vdd.t805 Vdd.t160 200
R511 Vdd.t915 Vdd.t805 200
R512 Vdd.t44 Vdd.t370 200
R513 Vdd.t290 Vdd.t44 200
R514 Vdd.t264 Vdd.t18 200
R515 Vdd.t128 Vdd.t264 200
R516 Vdd.t246 Vdd.t360 200
R517 Vdd.t807 Vdd.t246 200
R518 Vdd.t532 Vdd.t174 200
R519 Vdd.t568 Vdd.t532 200
R520 Vdd.t216 Vdd.t404 200
R521 Vdd.t260 Vdd.t216 200
R522 Vdd.t454 Vdd.t544 200
R523 Vdd.t747 Vdd.t454 200
R524 Vdd.t362 Vdd.t560 200
R525 Vdd.t92 Vdd.t362 200
R526 Vdd.t474 Vdd.t558 200
R527 Vdd.t310 Vdd.t474 200
R528 Vdd.t382 Vdd.t542 200
R529 Vdd.t60 Vdd.t382 200
R530 Vdd.t450 Vdd.t556 200
R531 Vdd.t244 Vdd.t450 200
R532 Vdd.t416 Vdd.t562 200
R533 Vdd.t218 Vdd.t416 200
R534 Vdd.t150 Vdd.t56 200
R535 Vdd.t701 Vdd.t150 200
R536 Vdd.t472 Vdd.t68 200
R537 Vdd.t596 Vdd.t472 200
R538 Vdd.t24 Vdd.t276 200
R539 Vdd.t608 Vdd.t24 200
R540 Vdd.t58 Vdd.t196 200
R541 Vdd.t692 Vdd.t58 200
R542 Vdd.t380 Vdd.t580 200
R543 Vdd.t422 Vdd.t380 200
R544 Vdd.t214 Vdd.t504 200
R545 Vdd.t656 Vdd.t214 200
R546 Vdd.t272 Vdd.t494 200
R547 Vdd.t650 Vdd.t272 200
R548 Vdd.t372 Vdd.t82 200
R549 Vdd.t476 Vdd.t372 200
R550 Vdd.t552 Vdd.t434 200
R551 Vdd.t704 Vdd.t552 200
R552 Vdd.t502 Vdd.t869 200
R553 Vdd.t674 Vdd.t502 200
R554 Vdd.t418 Vdd.t64 200
R555 Vdd.t188 Vdd.t418 200
R556 Vdd.t438 Vdd.t833 200
R557 Vdd.t665 Vdd.t438 200
R558 Vdd.t436 Vdd.t398 200
R559 Vdd.t722 Vdd.t436 200
R560 Vdd.t464 Vdd.t76 200
R561 Vdd.t104 Vdd.t464 200
R562 Vdd.t146 Vdd.t753 200
R563 Vdd.t710 Vdd.t146 200
R564 Vdd.t835 Vdd.t304 200
R565 Vdd.t671 Vdd.t835 200
R566 Vdd.t456 Vdd.t584 200
R567 Vdd.t238 Vdd.t456 200
R568 Vdd.t751 Vdd.t430 200
R569 Vdd.t686 Vdd.t751 200
R570 Vdd.t72 Vdd.t148 200
R571 Vdd.t564 Vdd.t72 200
R572 Vdd.t22 Vdd.t374 200
R573 Vdd.t0 Vdd.t22 200
R574 Vdd.t574 Vdd.t26 200
R575 Vdd.t274 Vdd.t574 200
R576 Vdd.t442 Vdd.t448 200
R577 Vdd.t32 Vdd.t442 200
R578 Vdd.t84 Vdd.t212 200
R579 Vdd.t500 Vdd.t84 200
R580 Vdd.t931 Vdd.t406 200
R581 Vdd.t336 Vdd.t931 200
R582 Vdd.t586 Vdd.t550 200
R583 Vdd.t432 Vdd.t586 200
R584 Vdd.t112 Vdd.t410 200
R585 Vdd.t813 Vdd.t112 200
R586 Vdd.t70 Vdd.t440 200
R587 Vdd.t831 Vdd.t70 200
R588 Vdd.t522 Vdd.t402 200
R589 Vdd.t138 Vdd.t522 200
R590 Vdd.t66 Vdd.t176 200
R591 Vdd.t921 Vdd.t66 200
R592 Vdd.t528 Vdd.t452 200
R593 Vdd.t536 Vdd.t528 200
R594 Vdd.t468 Vdd.t823 200
R595 Vdd.t20 Vdd.t468 200
R596 Vdd.t378 Vdd.t943 200
R597 Vdd.t444 Vdd.t378 200
R598 Vdd.t414 Vdd.t30 200
R599 Vdd.t933 Vdd.t414 200
R600 Vdd.t368 Vdd.t334 200
R601 Vdd.t110 Vdd.t368 200
R602 Vdd.t358 Vdd.t811 200
R603 Vdd.t520 Vdd.t358 200
R604 Vdd.t412 Vdd.t136 200
R605 Vdd.t530 Vdd.t412 200
R606 Vdd.t763 Vdd.t827 200
R607 Vdd.t400 Vdd.t763 200
R608 Vdd.t617 Vdd.t578 200
R609 Vdd.t923 Vdd.t617 200
R610 Vdd.t829 Vdd.t937 200
R611 Vdd.t386 Vdd.t829 200
R612 Vdd.t582 Vdd.t761 200
R613 Vdd.t825 Vdd.t582 200
R614 Vdd.t14 Vdd.t719 200
R615 Vdd.t793 Vdd.t14 200
R616 Vdd.t713 Vdd.t10 200
R617 Vdd.t885 Vdd.t713 200
R618 Vdd.t909 Vdd.t737 200
R619 Vdd.t614 Vdd.t909 200
R620 Vdd.t632 Vdd.t230 200
R621 Vdd.t554 Vdd.t632 200
R622 Vdd.t735 Vdd.t891 200
R623 Vdd.t653 Vdd.t735 200
R624 Vdd.t46 Vdd.t907 200
R625 Vdd.t733 Vdd.t46 200
R626 Vdd.t270 Vdd.t728 200
R627 Vdd.t38 Vdd.t270 200
R628 Vdd.t677 Vdd.t140 200
R629 Vdd.t941 Vdd.t677 200
R630 Vdd.t144 Vdd.t346 200
R631 Vdd.t599 Vdd.t144 200
R632 Vdd.t635 Vdd.t50 200
R633 Vdd.t228 Vdd.t635 200
R634 Vdd.t348 Vdd.t34 200
R635 Vdd.t620 Vdd.t348 200
R636 Vdd.t234 Vdd.t142 200
R637 Vdd.t350 Vdd.t234 200
R638 Vdd.t226 Vdd.t629 200
R639 Vdd.t266 Vdd.t226 200
R640 Vdd.t680 Vdd.t156 200
R641 Vdd.t224 Vdd.t680 200
R642 Vdd.t594 Vdd.t595 200
R643 Vdd.t903 Vdd.t905 200
R644 Vdd.t299 Vdd.t298 200
R645 Vdd.t889 Vdd.t887 200
R646 Vdd.t302 Vdd.t303 200
R647 Vdd.t164 Vdd.t162 200
R648 Vdd.t134 Vdd.t135 200
R649 Vdd.t98 Vdd.t100 200
R650 Vdd.t789 Vdd.n1029 195.312
R651 Vdd.n1063 Vdd.t80 190.464
R652 Vdd.n1039 Vdd.t74 190.464
R653 Vdd.n1030 Vdd.t789 179.689
R654 Vdd.t322 Vdd.n1026 145.413
R655 Vdd.n15 Vdd.t254 131.589
R656 Vdd.n174 Vdd.t330 131.589
R657 Vdd.n31 Vdd.t510 131.589
R658 Vdd.n101 Vdd.t118 131.589
R659 Vdd.n239 Vdd.t106 131.589
R660 Vdd.n253 Vdd.t352 131.589
R661 Vdd.n469 Vdd.t36 131.589
R662 Vdd.n602 Vdd.t96 131.589
R663 Vdd.n485 Vdd.t268 131.589
R664 Vdd.n533 Vdd.t755 131.589
R665 Vdd.n461 Vdd.t911 131.589
R666 Vdd.n447 Vdd.t6 131.589
R667 Vdd.n1006 Vdd.n259 130.231
R668 Vdd.n1006 Vdd.n982 121.085
R669 Vdd.n117 Vdd.t767 118.543
R670 Vdd.n190 Vdd.t588 118.543
R671 Vdd.n549 Vdd.t775 118.543
R672 Vdd.n618 Vdd.t781 118.543
R673 Vdd.n438 Vdd.t777 118.543
R674 Vdd.n255 Vdd.t765 118.543
R675 Vdd.n437 Vdd.t849 118.519
R676 Vdd.n259 Vdd.n258 117.481
R677 Vdd.n39 Vdd.n38 96.0755
R678 Vdd.n40 Vdd.n39 96.0755
R679 Vdd.n23 Vdd.n22 96.0755
R680 Vdd.n24 Vdd.n23 96.0755
R681 Vdd.n493 Vdd.n492 96.0755
R682 Vdd.n494 Vdd.n493 96.0755
R683 Vdd.n477 Vdd.n476 96.0755
R684 Vdd.n478 Vdd.n477 96.0755
R685 Vdd.n433 Vdd.n425 96.0755
R686 Vdd.n433 Vdd.n426 96.0755
R687 Vdd.n223 Vdd.n222 96.0755
R688 Vdd.n224 Vdd.n223 96.0755
R689 Vdd.n1030 Vdd.t785 85.938
R690 Vdd.n168 Vdd.n166 78.2255
R691 Vdd.n172 Vdd.n168 78.2255
R692 Vdd.n172 Vdd.n169 78.2255
R693 Vdd.n169 Vdd.n166 78.2255
R694 Vdd.n95 Vdd.n93 78.2255
R695 Vdd.n99 Vdd.n95 78.2255
R696 Vdd.n99 Vdd.n96 78.2255
R697 Vdd.n96 Vdd.n93 78.2255
R698 Vdd.n45 Vdd.n36 78.2255
R699 Vdd.n45 Vdd.n37 78.2255
R700 Vdd.n113 Vdd.n108 78.2255
R701 Vdd.n113 Vdd.n109 78.2255
R702 Vdd.n110 Vdd.n108 78.2255
R703 Vdd.n110 Vdd.n109 78.2255
R704 Vdd.n29 Vdd.n20 78.2255
R705 Vdd.n29 Vdd.n21 78.2255
R706 Vdd.n186 Vdd.n181 78.2255
R707 Vdd.n186 Vdd.n182 78.2255
R708 Vdd.n183 Vdd.n181 78.2255
R709 Vdd.n183 Vdd.n182 78.2255
R710 Vdd.n233 Vdd.n231 78.2255
R711 Vdd.n237 Vdd.n233 78.2255
R712 Vdd.n237 Vdd.n234 78.2255
R713 Vdd.n234 Vdd.n231 78.2255
R714 Vdd.n596 Vdd.n594 78.2255
R715 Vdd.n600 Vdd.n596 78.2255
R716 Vdd.n600 Vdd.n597 78.2255
R717 Vdd.n597 Vdd.n594 78.2255
R718 Vdd.n527 Vdd.n525 78.2255
R719 Vdd.n531 Vdd.n527 78.2255
R720 Vdd.n531 Vdd.n528 78.2255
R721 Vdd.n528 Vdd.n525 78.2255
R722 Vdd.n499 Vdd.n490 78.2255
R723 Vdd.n499 Vdd.n491 78.2255
R724 Vdd.n545 Vdd.n540 78.2255
R725 Vdd.n545 Vdd.n541 78.2255
R726 Vdd.n542 Vdd.n540 78.2255
R727 Vdd.n542 Vdd.n541 78.2255
R728 Vdd.n483 Vdd.n474 78.2255
R729 Vdd.n483 Vdd.n475 78.2255
R730 Vdd.n614 Vdd.n609 78.2255
R731 Vdd.n614 Vdd.n610 78.2255
R732 Vdd.n611 Vdd.n609 78.2255
R733 Vdd.n611 Vdd.n610 78.2255
R734 Vdd.n455 Vdd.n453 78.2255
R735 Vdd.n459 Vdd.n455 78.2255
R736 Vdd.n459 Vdd.n456 78.2255
R737 Vdd.n456 Vdd.n453 78.2255
R738 Vdd.n441 Vdd.n435 78.2255
R739 Vdd.n445 Vdd.n441 78.2255
R740 Vdd.n445 Vdd.n442 78.2255
R741 Vdd.n442 Vdd.n435 78.2255
R742 Vdd.n427 Vdd.n422 78.2255
R743 Vdd.n428 Vdd.n422 78.2255
R744 Vdd.n247 Vdd.n215 78.2255
R745 Vdd.n251 Vdd.n215 78.2255
R746 Vdd.n251 Vdd.n216 78.2255
R747 Vdd.n247 Vdd.n216 78.2255
R748 Vdd.n221 Vdd.n219 78.2255
R749 Vdd.n221 Vdd.n220 78.2255
R750 Vdd.n1029 Vdd.t787 70.313
R751 Vdd.n5 Vdd.n4 68.0765
R752 Vdd.n1096 Vdd.n1095 68.0765
R753 Vdd.n10 Vdd.n9 68.0765
R754 Vdd.n1084 Vdd.n1083 68.0765
R755 Vdd.n1090 Vdd.n1089 68.0765
R756 Vdd.n1077 Vdd.n1076 68.0765
R757 Vdd.n52 Vdd.n51 68.0765
R758 Vdd.n63 Vdd.n62 68.0765
R759 Vdd.n58 Vdd.n57 68.0765
R760 Vdd.n75 Vdd.n74 68.0765
R761 Vdd.n69 Vdd.n68 68.0765
R762 Vdd.n86 Vdd.n85 68.0765
R763 Vdd.n125 Vdd.n124 68.0765
R764 Vdd.n136 Vdd.n135 68.0765
R765 Vdd.n131 Vdd.n130 68.0765
R766 Vdd.n148 Vdd.n147 68.0765
R767 Vdd.n142 Vdd.n141 68.0765
R768 Vdd.n159 Vdd.n158 68.0765
R769 Vdd.n205 Vdd.n204 68.0765
R770 Vdd.n210 Vdd.n209 68.0765
R771 Vdd.n199 Vdd.n198 68.0765
R772 Vdd.n1002 Vdd.n1001 68.0765
R773 Vdd.n985 Vdd.n984 68.0765
R774 Vdd.n990 Vdd.n989 68.0765
R775 Vdd.n996 Vdd.n995 68.0765
R776 Vdd.n978 Vdd.n977 68.0765
R777 Vdd.n506 Vdd.n505 68.0765
R778 Vdd.n512 Vdd.n511 68.0765
R779 Vdd.n518 Vdd.n517 68.0765
R780 Vdd.n969 Vdd.n968 68.0765
R781 Vdd.n755 Vdd.n754 68.0765
R782 Vdd.n794 Vdd.n793 68.0765
R783 Vdd.n832 Vdd.n831 68.0765
R784 Vdd.n870 Vdd.n869 68.0765
R785 Vdd.n909 Vdd.n908 68.0765
R786 Vdd.n947 Vdd.n946 68.0765
R787 Vdd.n673 Vdd.n672 68.0765
R788 Vdd.n766 Vdd.n765 68.0765
R789 Vdd.n399 Vdd.n398 68.0765
R790 Vdd.n805 Vdd.n804 68.0765
R791 Vdd.n369 Vdd.n368 68.0765
R792 Vdd.n843 Vdd.n842 68.0765
R793 Vdd.n339 Vdd.n338 68.0765
R794 Vdd.n882 Vdd.n881 68.0765
R795 Vdd.n303 Vdd.n302 68.0765
R796 Vdd.n920 Vdd.n919 68.0765
R797 Vdd.n273 Vdd.n272 68.0765
R798 Vdd.n958 Vdd.n957 68.0765
R799 Vdd.n750 Vdd.n749 68.0765
R800 Vdd.n663 Vdd.n662 68.0765
R801 Vdd.n789 Vdd.n788 68.0765
R802 Vdd.n389 Vdd.n388 68.0765
R803 Vdd.n827 Vdd.n826 68.0765
R804 Vdd.n359 Vdd.n358 68.0765
R805 Vdd.n865 Vdd.n864 68.0765
R806 Vdd.n323 Vdd.n322 68.0765
R807 Vdd.n904 Vdd.n903 68.0765
R808 Vdd.n293 Vdd.n292 68.0765
R809 Vdd.n942 Vdd.n941 68.0765
R810 Vdd.n263 Vdd.n262 68.0765
R811 Vdd.n678 Vdd.n677 68.0765
R812 Vdd.n404 Vdd.n403 68.0765
R813 Vdd.n374 Vdd.n373 68.0765
R814 Vdd.n344 Vdd.n343 68.0765
R815 Vdd.n308 Vdd.n307 68.0765
R816 Vdd.n278 Vdd.n277 68.0765
R817 Vdd.n745 Vdd.n744 68.0765
R818 Vdd.n683 Vdd.n682 68.0765
R819 Vdd.n784 Vdd.n783 68.0765
R820 Vdd.n761 Vdd.n760 68.0765
R821 Vdd.n409 Vdd.n408 68.0765
R822 Vdd.n822 Vdd.n821 68.0765
R823 Vdd.n800 Vdd.n799 68.0765
R824 Vdd.n379 Vdd.n378 68.0765
R825 Vdd.n860 Vdd.n859 68.0765
R826 Vdd.n838 Vdd.n837 68.0765
R827 Vdd.n349 Vdd.n348 68.0765
R828 Vdd.n899 Vdd.n898 68.0765
R829 Vdd.n877 Vdd.n876 68.0765
R830 Vdd.n313 Vdd.n312 68.0765
R831 Vdd.n937 Vdd.n936 68.0765
R832 Vdd.n915 Vdd.n914 68.0765
R833 Vdd.n283 Vdd.n282 68.0765
R834 Vdd.n953 Vdd.n952 68.0765
R835 Vdd.n740 Vdd.n739 68.0765
R836 Vdd.n668 Vdd.n667 68.0765
R837 Vdd.n779 Vdd.n778 68.0765
R838 Vdd.n394 Vdd.n393 68.0765
R839 Vdd.n817 Vdd.n816 68.0765
R840 Vdd.n364 Vdd.n363 68.0765
R841 Vdd.n855 Vdd.n854 68.0765
R842 Vdd.n328 Vdd.n327 68.0765
R843 Vdd.n894 Vdd.n893 68.0765
R844 Vdd.n298 Vdd.n297 68.0765
R845 Vdd.n932 Vdd.n931 68.0765
R846 Vdd.n268 Vdd.n267 68.0765
R847 Vdd.n688 Vdd.n687 68.0765
R848 Vdd.n414 Vdd.n413 68.0765
R849 Vdd.n384 Vdd.n383 68.0765
R850 Vdd.n354 Vdd.n353 68.0765
R851 Vdd.n318 Vdd.n317 68.0765
R852 Vdd.n288 Vdd.n287 68.0765
R853 Vdd.n693 Vdd.n692 68.0765
R854 Vdd.n709 Vdd.n708 68.0765
R855 Vdd.n704 Vdd.n703 68.0765
R856 Vdd.n727 Vdd.n726 68.0765
R857 Vdd.n733 Vdd.n732 68.0765
R858 Vdd.n721 Vdd.n720 68.0765
R859 Vdd.n626 Vdd.n625 68.0765
R860 Vdd.n637 Vdd.n636 68.0765
R861 Vdd.n632 Vdd.n631 68.0765
R862 Vdd.n649 Vdd.n648 68.0765
R863 Vdd.n643 Vdd.n642 68.0765
R864 Vdd.n656 Vdd.n655 68.0765
R865 Vdd.n557 Vdd.n556 68.0765
R866 Vdd.n568 Vdd.n567 68.0765
R867 Vdd.n563 Vdd.n562 68.0765
R868 Vdd.n580 Vdd.n579 68.0765
R869 Vdd.n574 Vdd.n573 68.0765
R870 Vdd.n587 Vdd.n586 68.0765
R871 Vdd.n38 Vdd.n36 59.8505
R872 Vdd.n40 Vdd.n37 59.8505
R873 Vdd.n22 Vdd.n20 59.8505
R874 Vdd.n24 Vdd.n21 59.8505
R875 Vdd.n492 Vdd.n490 59.8505
R876 Vdd.n494 Vdd.n491 59.8505
R877 Vdd.n476 Vdd.n474 59.8505
R878 Vdd.n478 Vdd.n475 59.8505
R879 Vdd.n427 Vdd.n425 59.8505
R880 Vdd.n428 Vdd.n426 59.8505
R881 Vdd.n222 Vdd.n219 59.8505
R882 Vdd.n224 Vdd.n220 59.8505
R883 Vdd.n1013 Vdd.n1011 58.9755
R884 Vdd.n1016 Vdd.n1011 58.9755
R885 Vdd.n1016 Vdd.n1012 58.9755
R886 Vdd.n1013 Vdd.n1012 58.9755
R887 Vdd.n1059 Vdd.n1034 54.0755
R888 Vdd.n1041 Vdd.n1036 54.0755
R889 Vdd.n1041 Vdd.n1037 54.0755
R890 Vdd.n1059 Vdd.n1035 54.0755
R891 Vdd.n192 Vdd.t661 41.0041
R892 Vdd.n79 Vdd.t643 41.0041
R893 Vdd.n152 Vdd.t730 41.0041
R894 Vdd.n962 Vdd.t646 41.0041
R895 Vdd.n713 Vdd.t718 41.0041
R896 Vdd.n417 Vdd.t727 41.0041
R897 Vdd.n331 Vdd.t628 41.0041
R898 Vdd.n194 Vdd.t697 40.8177
R899 Vdd.n193 Vdd.t658 40.8177
R900 Vdd.n81 Vdd.t637 40.8177
R901 Vdd.n80 Vdd.t601 40.8177
R902 Vdd.n154 Vdd.t622 40.8177
R903 Vdd.n153 Vdd.t724 40.8177
R904 Vdd.n964 Vdd.t682 40.8177
R905 Vdd.n963 Vdd.t640 40.8177
R906 Vdd.n716 Vdd.t712 40.8177
R907 Vdd.n715 Vdd.t616 40.8177
R908 Vdd.n419 Vdd.t676 40.8177
R909 Vdd.n418 Vdd.t631 40.8177
R910 Vdd.n333 Vdd.t679 40.8177
R911 Vdd.n332 Vdd.t634 40.8177
R912 Vdd.n47 Vdd.t715 40.6313
R913 Vdd.n46 Vdd.t604 40.6313
R914 Vdd.n120 Vdd.t694 40.6313
R915 Vdd.n119 Vdd.t706 40.6313
R916 Vdd.n501 Vdd.t610 40.6313
R917 Vdd.n500 Vdd.t625 40.6313
R918 Vdd.n773 Vdd.t607 40.6313
R919 Vdd.n771 Vdd.t649 40.6313
R920 Vdd.n811 Vdd.t655 40.6313
R921 Vdd.n809 Vdd.t673 40.6313
R922 Vdd.n849 Vdd.t703 40.6313
R923 Vdd.n847 Vdd.t721 40.6313
R924 Vdd.n888 Vdd.t664 40.6313
R925 Vdd.n886 Vdd.t670 40.6313
R926 Vdd.n926 Vdd.t709 40.6313
R927 Vdd.n924 Vdd.t685 40.6313
R928 Vdd.n698 Vdd.t700 40.6313
R929 Vdd.n696 Vdd.t691 40.6313
R930 Vdd.n552 Vdd.t598 40.6313
R931 Vdd.n551 Vdd.t619 40.6313
R932 Vdd.n621 Vdd.t613 40.6313
R933 Vdd.n620 Vdd.t652 40.6313
R934 Vdd.n1 Vdd.t667 40.6313
R935 Vdd.n0 Vdd.t688 40.6313
R936 Vdd.n170 Vdd.n168 36.2255
R937 Vdd.n170 Vdd.n169 36.2255
R938 Vdd.n97 Vdd.n95 36.2255
R939 Vdd.n97 Vdd.n96 36.2255
R940 Vdd.n41 Vdd.n38 36.2255
R941 Vdd.n41 Vdd.n40 36.2255
R942 Vdd.n43 Vdd.n36 36.2255
R943 Vdd.n43 Vdd.n37 36.2255
R944 Vdd.n111 Vdd.n108 36.2255
R945 Vdd.n111 Vdd.n109 36.2255
R946 Vdd.n25 Vdd.n22 36.2255
R947 Vdd.n25 Vdd.n24 36.2255
R948 Vdd.n27 Vdd.n20 36.2255
R949 Vdd.n27 Vdd.n21 36.2255
R950 Vdd.n184 Vdd.n181 36.2255
R951 Vdd.n184 Vdd.n182 36.2255
R952 Vdd.n235 Vdd.n233 36.2255
R953 Vdd.n235 Vdd.n234 36.2255
R954 Vdd.n598 Vdd.n596 36.2255
R955 Vdd.n598 Vdd.n597 36.2255
R956 Vdd.n529 Vdd.n527 36.2255
R957 Vdd.n529 Vdd.n528 36.2255
R958 Vdd.n495 Vdd.n492 36.2255
R959 Vdd.n495 Vdd.n494 36.2255
R960 Vdd.n497 Vdd.n490 36.2255
R961 Vdd.n497 Vdd.n491 36.2255
R962 Vdd.n543 Vdd.n540 36.2255
R963 Vdd.n543 Vdd.n541 36.2255
R964 Vdd.n479 Vdd.n476 36.2255
R965 Vdd.n479 Vdd.n478 36.2255
R966 Vdd.n481 Vdd.n474 36.2255
R967 Vdd.n481 Vdd.n475 36.2255
R968 Vdd.n612 Vdd.n609 36.2255
R969 Vdd.n612 Vdd.n610 36.2255
R970 Vdd.n457 Vdd.n455 36.2255
R971 Vdd.n457 Vdd.n456 36.2255
R972 Vdd.n443 Vdd.n441 36.2255
R973 Vdd.n443 Vdd.n442 36.2255
R974 Vdd.n431 Vdd.n425 36.2255
R975 Vdd.n431 Vdd.n426 36.2255
R976 Vdd.n429 Vdd.n427 36.2255
R977 Vdd.n429 Vdd.n428 36.2255
R978 Vdd.n249 Vdd.n215 36.2255
R979 Vdd.n249 Vdd.n216 36.2255
R980 Vdd.n225 Vdd.n222 36.2255
R981 Vdd.n225 Vdd.n224 36.2255
R982 Vdd.n228 Vdd.n219 36.2255
R983 Vdd.n228 Vdd.n220 36.2255
R984 Vdd.n770 Vdd.n660 32.646
R985 Vdd.n1063 Vdd.n1062 29.3622
R986 Vdd.n1040 Vdd.n1039 29.3622
R987 Vdd.n47 Vdd.t958 27.3166
R988 Vdd.n46 Vdd.t950 27.3166
R989 Vdd.n120 Vdd.t963 27.3166
R990 Vdd.n119 Vdd.t961 27.3166
R991 Vdd.n501 Vdd.t949 27.3166
R992 Vdd.n500 Vdd.t985 27.3166
R993 Vdd.n773 Vdd.t960 27.3166
R994 Vdd.n771 Vdd.t976 27.3166
R995 Vdd.n811 Vdd.t948 27.3166
R996 Vdd.n809 Vdd.t967 27.3166
R997 Vdd.n849 Vdd.t971 27.3166
R998 Vdd.n847 Vdd.t956 27.3166
R999 Vdd.n888 Vdd.t989 27.3166
R1000 Vdd.n886 Vdd.t968 27.3166
R1001 Vdd.n926 Vdd.t970 27.3166
R1002 Vdd.n924 Vdd.t966 27.3166
R1003 Vdd.n698 Vdd.t972 27.3166
R1004 Vdd.n696 Vdd.t964 27.3166
R1005 Vdd.n552 Vdd.t952 27.3166
R1006 Vdd.n551 Vdd.t986 27.3166
R1007 Vdd.n621 Vdd.t947 27.3166
R1008 Vdd.n620 Vdd.t975 27.3166
R1009 Vdd.n1 Vdd.t969 27.3166
R1010 Vdd.n0 Vdd.t965 27.3166
R1011 Vdd.n194 Vdd.t982 27.1302
R1012 Vdd.n193 Vdd.t974 27.1302
R1013 Vdd.n81 Vdd.t957 27.1302
R1014 Vdd.n80 Vdd.t951 27.1302
R1015 Vdd.n154 Vdd.t962 27.1302
R1016 Vdd.n153 Vdd.t955 27.1302
R1017 Vdd.n964 Vdd.t987 27.1302
R1018 Vdd.n963 Vdd.t979 27.1302
R1019 Vdd.n716 Vdd.t959 27.1302
R1020 Vdd.n715 Vdd.t946 27.1302
R1021 Vdd.n419 Vdd.t945 27.1302
R1022 Vdd.n418 Vdd.t983 27.1302
R1023 Vdd.n333 Vdd.t988 27.1302
R1024 Vdd.n332 Vdd.t980 27.1302
R1025 Vdd.n192 Vdd.t973 26.9438
R1026 Vdd.n79 Vdd.t978 26.9438
R1027 Vdd.n152 Vdd.t953 26.9438
R1028 Vdd.n962 Vdd.t977 26.9438
R1029 Vdd.n713 Vdd.t981 26.9438
R1030 Vdd.n417 Vdd.t954 26.9438
R1031 Vdd.n331 Vdd.t984 26.9438
R1032 Vdd.t783 Vdd.n1027 23.438
R1033 Vdd.n1055 Vdd.n1036 20.1255
R1034 Vdd.n1055 Vdd.n1037 20.1255
R1035 Vdd.n1057 Vdd.n1034 20.1255
R1036 Vdd.n1057 Vdd.n1035 20.1255
R1037 Vdd.n1064 Vdd.n1063 19.9167
R1038 Vdd.n1039 Vdd.n1038 19.9167
R1039 Vdd.n1014 Vdd.n1011 18.7255
R1040 Vdd.n1014 Vdd.n1012 18.7255
R1041 Vdd.n724 SARlogic_0.dffrs_13.resetb 18.2673
R1042 Vdd.n89 adc_PISO_0.dffrs_5.resetb 18.2415
R1043 Vdd.n162 adc_PISO_0.dffrs_4.resetb 18.2415
R1044 Vdd.n1074 adc_PISO_0.dffrs_3.resetb 18.2061
R1045 Vdd.n973 adc_PISO_0.dffrs_2.resetb 18.2061
R1046 Vdd.n660 adc_PISO_0.dffrs_0.resetb 18.2061
R1047 Vdd.n336 adc_PISO_0.dffrs_1.resetb 18.2061
R1048 Vdd.n55 Vdd.n49 18.0418
R1049 Vdd.n128 Vdd.n122 18.0418
R1050 Vdd.n509 Vdd.n503 18.0418
R1051 Vdd.n560 Vdd.n554 18.0418
R1052 Vdd.n629 Vdd.n623 18.0418
R1053 Vdd.n1101 Vdd.n1100 18.0418
R1054 Vdd.n776 Vdd.n775 18.0005
R1055 Vdd.n814 Vdd.n813 18.0005
R1056 Vdd.n852 Vdd.n851 18.0005
R1057 Vdd.n891 Vdd.n890 18.0005
R1058 Vdd.n929 Vdd.n928 18.0005
R1059 Vdd.n701 Vdd.n700 18.0005
R1060 Vdd.n195 Vdd.n193 17.6364
R1061 Vdd.n82 Vdd.n80 17.6364
R1062 Vdd.n155 Vdd.n153 17.6364
R1063 Vdd.n965 Vdd.n963 17.6364
R1064 Vdd.n420 Vdd.n418 17.6364
R1065 Vdd.n334 Vdd.n332 17.6364
R1066 Vdd.n1066 Vdd.n1065 14.6602
R1067 Vdd.n48 Vdd.n46 14.3609
R1068 Vdd.n121 Vdd.n119 14.3609
R1069 Vdd.n502 Vdd.n500 14.3609
R1070 Vdd.n553 Vdd.n551 14.3609
R1071 Vdd.n622 Vdd.n620 14.3609
R1072 Vdd.n2 Vdd.n0 14.3609
R1073 Vdd.n213 Vdd.n207 13.5842
R1074 Vdd.n509 Vdd.n508 13.5431
R1075 Vdd.n1100 Vdd.n7 13.5174
R1076 Vdd.n55 Vdd.n54 13.5174
R1077 Vdd.n128 Vdd.n127 13.5174
R1078 Vdd.n629 Vdd.n628 13.5174
R1079 Vdd.n560 Vdd.n559 13.5174
R1080 Vdd.n701 Vdd.n695 13.5152
R1081 Vdd.n1099 Vdd.n1098 13.5005
R1082 Vdd.n1099 Vdd.n12 13.5005
R1083 Vdd.n1087 Vdd.n1086 13.5005
R1084 Vdd.n1093 Vdd.n1092 13.5005
R1085 Vdd.n1080 Vdd.n1079 13.5005
R1086 Vdd.n66 Vdd.n65 13.5005
R1087 Vdd.n66 Vdd.n60 13.5005
R1088 Vdd.n78 Vdd.n77 13.5005
R1089 Vdd.n72 Vdd.n71 13.5005
R1090 Vdd.n89 Vdd.n88 13.5005
R1091 Vdd.n139 Vdd.n138 13.5005
R1092 Vdd.n139 Vdd.n133 13.5005
R1093 Vdd.n151 Vdd.n150 13.5005
R1094 Vdd.n145 Vdd.n144 13.5005
R1095 Vdd.n162 Vdd.n161 13.5005
R1096 Vdd.n213 Vdd.n212 13.5005
R1097 Vdd.n202 Vdd.n201 13.5005
R1098 Vdd.n1005 Vdd.n1004 13.5005
R1099 Vdd.n1005 Vdd.n987 13.5005
R1100 Vdd.n993 Vdd.n992 13.5005
R1101 Vdd.n999 Vdd.n998 13.5005
R1102 Vdd.n981 Vdd.n980 13.5005
R1103 Vdd.n515 Vdd.n514 13.5005
R1104 Vdd.n521 Vdd.n520 13.5005
R1105 Vdd.n972 Vdd.n971 13.5005
R1106 Vdd.n758 Vdd.n757 13.5005
R1107 Vdd.n797 Vdd.n796 13.5005
R1108 Vdd.n835 Vdd.n834 13.5005
R1109 Vdd.n873 Vdd.n872 13.5005
R1110 Vdd.n912 Vdd.n911 13.5005
R1111 Vdd.n950 Vdd.n949 13.5005
R1112 Vdd.n758 Vdd.n675 13.5005
R1113 Vdd.n769 Vdd.n768 13.5005
R1114 Vdd.n797 Vdd.n401 13.5005
R1115 Vdd.n808 Vdd.n807 13.5005
R1116 Vdd.n835 Vdd.n371 13.5005
R1117 Vdd.n846 Vdd.n845 13.5005
R1118 Vdd.n873 Vdd.n341 13.5005
R1119 Vdd.n885 Vdd.n884 13.5005
R1120 Vdd.n912 Vdd.n305 13.5005
R1121 Vdd.n923 Vdd.n922 13.5005
R1122 Vdd.n950 Vdd.n275 13.5005
R1123 Vdd.n961 Vdd.n960 13.5005
R1124 Vdd.n758 Vdd.n752 13.5005
R1125 Vdd.n769 Vdd.n665 13.5005
R1126 Vdd.n797 Vdd.n791 13.5005
R1127 Vdd.n808 Vdd.n391 13.5005
R1128 Vdd.n835 Vdd.n829 13.5005
R1129 Vdd.n846 Vdd.n361 13.5005
R1130 Vdd.n873 Vdd.n867 13.5005
R1131 Vdd.n885 Vdd.n325 13.5005
R1132 Vdd.n912 Vdd.n906 13.5005
R1133 Vdd.n923 Vdd.n295 13.5005
R1134 Vdd.n950 Vdd.n944 13.5005
R1135 Vdd.n961 Vdd.n265 13.5005
R1136 Vdd.n758 Vdd.n680 13.5005
R1137 Vdd.n797 Vdd.n406 13.5005
R1138 Vdd.n835 Vdd.n376 13.5005
R1139 Vdd.n873 Vdd.n346 13.5005
R1140 Vdd.n912 Vdd.n310 13.5005
R1141 Vdd.n950 Vdd.n280 13.5005
R1142 Vdd.n758 Vdd.n747 13.5005
R1143 Vdd.n758 Vdd.n685 13.5005
R1144 Vdd.n797 Vdd.n786 13.5005
R1145 Vdd.n769 Vdd.n763 13.5005
R1146 Vdd.n797 Vdd.n411 13.5005
R1147 Vdd.n835 Vdd.n824 13.5005
R1148 Vdd.n808 Vdd.n802 13.5005
R1149 Vdd.n835 Vdd.n381 13.5005
R1150 Vdd.n873 Vdd.n862 13.5005
R1151 Vdd.n846 Vdd.n840 13.5005
R1152 Vdd.n873 Vdd.n351 13.5005
R1153 Vdd.n912 Vdd.n901 13.5005
R1154 Vdd.n885 Vdd.n879 13.5005
R1155 Vdd.n912 Vdd.n315 13.5005
R1156 Vdd.n950 Vdd.n939 13.5005
R1157 Vdd.n923 Vdd.n917 13.5005
R1158 Vdd.n950 Vdd.n285 13.5005
R1159 Vdd.n961 Vdd.n955 13.5005
R1160 Vdd.n758 Vdd.n742 13.5005
R1161 Vdd.n769 Vdd.n670 13.5005
R1162 Vdd.n797 Vdd.n781 13.5005
R1163 Vdd.n808 Vdd.n396 13.5005
R1164 Vdd.n835 Vdd.n819 13.5005
R1165 Vdd.n846 Vdd.n366 13.5005
R1166 Vdd.n873 Vdd.n857 13.5005
R1167 Vdd.n885 Vdd.n330 13.5005
R1168 Vdd.n912 Vdd.n896 13.5005
R1169 Vdd.n923 Vdd.n300 13.5005
R1170 Vdd.n950 Vdd.n934 13.5005
R1171 Vdd.n961 Vdd.n270 13.5005
R1172 Vdd.n758 Vdd.n690 13.5005
R1173 Vdd.n797 Vdd.n416 13.5005
R1174 Vdd.n835 Vdd.n386 13.5005
R1175 Vdd.n873 Vdd.n356 13.5005
R1176 Vdd.n912 Vdd.n320 13.5005
R1177 Vdd.n950 Vdd.n290 13.5005
R1178 Vdd.n712 Vdd.n711 13.5005
R1179 Vdd.n712 Vdd.n706 13.5005
R1180 Vdd.n730 Vdd.n729 13.5005
R1181 Vdd.n736 Vdd.n735 13.5005
R1182 Vdd.n724 Vdd.n723 13.5005
R1183 Vdd.n640 Vdd.n639 13.5005
R1184 Vdd.n640 Vdd.n634 13.5005
R1185 Vdd.n652 Vdd.n651 13.5005
R1186 Vdd.n646 Vdd.n645 13.5005
R1187 Vdd.n659 Vdd.n658 13.5005
R1188 Vdd.n571 Vdd.n570 13.5005
R1189 Vdd.n571 Vdd.n565 13.5005
R1190 Vdd.n583 Vdd.n582 13.5005
R1191 Vdd.n577 Vdd.n576 13.5005
R1192 Vdd.n590 Vdd.n589 13.5005
R1193 Vdd.n1071 Vdd.n1008 13.4987
R1194 Vdd.n196 Vdd.n192 13.4839
R1195 Vdd.n83 Vdd.n79 13.4839
R1196 Vdd.n156 Vdd.n152 13.4839
R1197 Vdd.n966 Vdd.n962 13.4839
R1198 Vdd.n421 Vdd.n417 13.4839
R1199 Vdd.n335 Vdd.n331 13.4839
R1200 Vdd.n1027 Vdd.n1021 12.6005
R1201 Vdd.n1031 Vdd.n1030 12.6005
R1202 Vdd.n1029 Vdd.n1028 12.6005
R1203 Vdd.n717 SARlogic_0.dffrs_13.nand3_1.B 12.1571
R1204 Vdd.n1053 Vdd.n1052 12.136
R1205 Vdd.n1051 Vdd.n1050 12.136
R1206 Vdd.n1049 Vdd.n1048 12.136
R1207 Vdd.n1047 Vdd.n1046 12.136
R1208 Vdd.n1045 Vdd.n1044 12.136
R1209 Vdd.n1057 Vdd.n1033 11.111
R1210 Vdd.n1055 Vdd.n1054 11.111
R1211 Vdd.n195 Vdd.n194 10.5752
R1212 Vdd.n82 Vdd.n81 10.5752
R1213 Vdd.n155 Vdd.n154 10.5752
R1214 Vdd.n965 Vdd.n964 10.5752
R1215 Vdd.n420 Vdd.n419 10.5752
R1216 Vdd.n334 Vdd.n333 10.5752
R1217 Vdd.n1038 Vdd.n1008 9.86945
R1218 Vdd.n1043 Vdd.n1042 9.536
R1219 Vdd.n1061 Vdd.n1060 9.536
R1220 Vdd.n1065 Vdd.n1064 9.536
R1221 Vdd.n774 Vdd.n772 9.22229
R1222 Vdd.n812 Vdd.n810 9.22229
R1223 Vdd.n850 Vdd.n848 9.22229
R1224 Vdd.n889 Vdd.n887 9.22229
R1225 Vdd.n927 Vdd.n925 9.22229
R1226 Vdd.n699 Vdd.n697 9.22229
R1227 Vdd.n718 Vdd.n714 7.75389
R1228 Vdd.n1042 Vdd.t577 7.4755
R1229 Vdd.n1060 Vdd.t79 7.4755
R1230 Vdd.n1064 Vdd.t81 7.4755
R1231 Vdd.n1038 Vdd.t75 7.4755
R1232 Vdd.n975 Vdd.n974 6.55364
R1233 Vdd.n7 Vdd.n4 6.4802
R1234 Vdd.n1098 Vdd.n1095 6.4802
R1235 Vdd.n12 Vdd.n9 6.4802
R1236 Vdd.n1086 Vdd.n1083 6.4802
R1237 Vdd.n1092 Vdd.n1089 6.4802
R1238 Vdd.n1079 Vdd.n1076 6.4802
R1239 Vdd.n54 Vdd.n51 6.4802
R1240 Vdd.n65 Vdd.n62 6.4802
R1241 Vdd.n60 Vdd.n57 6.4802
R1242 Vdd.n77 Vdd.n74 6.4802
R1243 Vdd.n71 Vdd.n68 6.4802
R1244 Vdd.n88 Vdd.n85 6.4802
R1245 Vdd.n127 Vdd.n124 6.4802
R1246 Vdd.n138 Vdd.n135 6.4802
R1247 Vdd.n133 Vdd.n130 6.4802
R1248 Vdd.n150 Vdd.n147 6.4802
R1249 Vdd.n144 Vdd.n141 6.4802
R1250 Vdd.n161 Vdd.n158 6.4802
R1251 Vdd.n207 Vdd.n204 6.4802
R1252 Vdd.n212 Vdd.n209 6.4802
R1253 Vdd.n201 Vdd.n198 6.4802
R1254 Vdd.n1004 Vdd.n1001 6.4802
R1255 Vdd.n987 Vdd.n984 6.4802
R1256 Vdd.n992 Vdd.n989 6.4802
R1257 Vdd.n998 Vdd.n995 6.4802
R1258 Vdd.n980 Vdd.n977 6.4802
R1259 Vdd.n508 Vdd.n505 6.4802
R1260 Vdd.n514 Vdd.n511 6.4802
R1261 Vdd.n520 Vdd.n517 6.4802
R1262 Vdd.n971 Vdd.n968 6.4802
R1263 Vdd.n757 Vdd.n754 6.4802
R1264 Vdd.n796 Vdd.n793 6.4802
R1265 Vdd.n834 Vdd.n831 6.4802
R1266 Vdd.n872 Vdd.n869 6.4802
R1267 Vdd.n911 Vdd.n908 6.4802
R1268 Vdd.n949 Vdd.n946 6.4802
R1269 Vdd.n675 Vdd.n672 6.4802
R1270 Vdd.n768 Vdd.n765 6.4802
R1271 Vdd.n401 Vdd.n398 6.4802
R1272 Vdd.n807 Vdd.n804 6.4802
R1273 Vdd.n371 Vdd.n368 6.4802
R1274 Vdd.n845 Vdd.n842 6.4802
R1275 Vdd.n341 Vdd.n338 6.4802
R1276 Vdd.n884 Vdd.n881 6.4802
R1277 Vdd.n305 Vdd.n302 6.4802
R1278 Vdd.n922 Vdd.n919 6.4802
R1279 Vdd.n275 Vdd.n272 6.4802
R1280 Vdd.n960 Vdd.n957 6.4802
R1281 Vdd.n752 Vdd.n749 6.4802
R1282 Vdd.n665 Vdd.n662 6.4802
R1283 Vdd.n791 Vdd.n788 6.4802
R1284 Vdd.n391 Vdd.n388 6.4802
R1285 Vdd.n829 Vdd.n826 6.4802
R1286 Vdd.n361 Vdd.n358 6.4802
R1287 Vdd.n867 Vdd.n864 6.4802
R1288 Vdd.n325 Vdd.n322 6.4802
R1289 Vdd.n906 Vdd.n903 6.4802
R1290 Vdd.n295 Vdd.n292 6.4802
R1291 Vdd.n944 Vdd.n941 6.4802
R1292 Vdd.n265 Vdd.n262 6.4802
R1293 Vdd.n680 Vdd.n677 6.4802
R1294 Vdd.n406 Vdd.n403 6.4802
R1295 Vdd.n376 Vdd.n373 6.4802
R1296 Vdd.n346 Vdd.n343 6.4802
R1297 Vdd.n310 Vdd.n307 6.4802
R1298 Vdd.n280 Vdd.n277 6.4802
R1299 Vdd.n747 Vdd.n744 6.4802
R1300 Vdd.n685 Vdd.n682 6.4802
R1301 Vdd.n786 Vdd.n783 6.4802
R1302 Vdd.n763 Vdd.n760 6.4802
R1303 Vdd.n411 Vdd.n408 6.4802
R1304 Vdd.n824 Vdd.n821 6.4802
R1305 Vdd.n802 Vdd.n799 6.4802
R1306 Vdd.n381 Vdd.n378 6.4802
R1307 Vdd.n862 Vdd.n859 6.4802
R1308 Vdd.n840 Vdd.n837 6.4802
R1309 Vdd.n351 Vdd.n348 6.4802
R1310 Vdd.n901 Vdd.n898 6.4802
R1311 Vdd.n879 Vdd.n876 6.4802
R1312 Vdd.n315 Vdd.n312 6.4802
R1313 Vdd.n939 Vdd.n936 6.4802
R1314 Vdd.n917 Vdd.n914 6.4802
R1315 Vdd.n285 Vdd.n282 6.4802
R1316 Vdd.n955 Vdd.n952 6.4802
R1317 Vdd.n742 Vdd.n739 6.4802
R1318 Vdd.n670 Vdd.n667 6.4802
R1319 Vdd.n781 Vdd.n778 6.4802
R1320 Vdd.n396 Vdd.n393 6.4802
R1321 Vdd.n819 Vdd.n816 6.4802
R1322 Vdd.n366 Vdd.n363 6.4802
R1323 Vdd.n857 Vdd.n854 6.4802
R1324 Vdd.n330 Vdd.n327 6.4802
R1325 Vdd.n896 Vdd.n893 6.4802
R1326 Vdd.n300 Vdd.n297 6.4802
R1327 Vdd.n934 Vdd.n931 6.4802
R1328 Vdd.n270 Vdd.n267 6.4802
R1329 Vdd.n690 Vdd.n687 6.4802
R1330 Vdd.n416 Vdd.n413 6.4802
R1331 Vdd.n386 Vdd.n383 6.4802
R1332 Vdd.n356 Vdd.n353 6.4802
R1333 Vdd.n320 Vdd.n317 6.4802
R1334 Vdd.n290 Vdd.n287 6.4802
R1335 Vdd.n695 Vdd.n692 6.4802
R1336 Vdd.n711 Vdd.n708 6.4802
R1337 Vdd.n706 Vdd.n703 6.4802
R1338 Vdd.n729 Vdd.n726 6.4802
R1339 Vdd.n735 Vdd.n732 6.4802
R1340 Vdd.n723 Vdd.n720 6.4802
R1341 Vdd.n628 Vdd.n625 6.4802
R1342 Vdd.n639 Vdd.n636 6.4802
R1343 Vdd.n634 Vdd.n631 6.4802
R1344 Vdd.n651 Vdd.n648 6.4802
R1345 Vdd.n645 Vdd.n642 6.4802
R1346 Vdd.n658 Vdd.n655 6.4802
R1347 Vdd.n559 Vdd.n556 6.4802
R1348 Vdd.n570 Vdd.n567 6.4802
R1349 Vdd.n565 Vdd.n562 6.4802
R1350 Vdd.n582 Vdd.n579 6.4802
R1351 Vdd.n576 Vdd.n573 6.4802
R1352 Vdd.n589 Vdd.n586 6.4802
R1353 Vdd.n7 Vdd.n3 6.25878
R1354 Vdd.n1098 Vdd.n1094 6.25878
R1355 Vdd.n12 Vdd.n8 6.25878
R1356 Vdd.n1086 Vdd.n1082 6.25878
R1357 Vdd.n1092 Vdd.n1088 6.25878
R1358 Vdd.n1079 Vdd.n1075 6.25878
R1359 Vdd.n54 Vdd.n50 6.25878
R1360 Vdd.n65 Vdd.n61 6.25878
R1361 Vdd.n60 Vdd.n56 6.25878
R1362 Vdd.n77 Vdd.n73 6.25878
R1363 Vdd.n71 Vdd.n67 6.25878
R1364 Vdd.n88 Vdd.n84 6.25878
R1365 Vdd.n127 Vdd.n123 6.25878
R1366 Vdd.n138 Vdd.n134 6.25878
R1367 Vdd.n133 Vdd.n129 6.25878
R1368 Vdd.n150 Vdd.n146 6.25878
R1369 Vdd.n144 Vdd.n140 6.25878
R1370 Vdd.n161 Vdd.n157 6.25878
R1371 Vdd.n207 Vdd.n203 6.25878
R1372 Vdd.n212 Vdd.n208 6.25878
R1373 Vdd.n201 Vdd.n197 6.25878
R1374 Vdd.n1004 Vdd.n1000 6.25878
R1375 Vdd.n987 Vdd.n983 6.25878
R1376 Vdd.n992 Vdd.n988 6.25878
R1377 Vdd.n998 Vdd.n994 6.25878
R1378 Vdd.n980 Vdd.n976 6.25878
R1379 Vdd.n508 Vdd.n504 6.25878
R1380 Vdd.n514 Vdd.n510 6.25878
R1381 Vdd.n520 Vdd.n516 6.25878
R1382 Vdd.n971 Vdd.n967 6.25878
R1383 Vdd.n757 Vdd.n753 6.25878
R1384 Vdd.n796 Vdd.n792 6.25878
R1385 Vdd.n834 Vdd.n830 6.25878
R1386 Vdd.n872 Vdd.n868 6.25878
R1387 Vdd.n911 Vdd.n907 6.25878
R1388 Vdd.n949 Vdd.n945 6.25878
R1389 Vdd.n675 Vdd.n671 6.25878
R1390 Vdd.n768 Vdd.n764 6.25878
R1391 Vdd.n401 Vdd.n397 6.25878
R1392 Vdd.n807 Vdd.n803 6.25878
R1393 Vdd.n371 Vdd.n367 6.25878
R1394 Vdd.n845 Vdd.n841 6.25878
R1395 Vdd.n341 Vdd.n337 6.25878
R1396 Vdd.n884 Vdd.n880 6.25878
R1397 Vdd.n305 Vdd.n301 6.25878
R1398 Vdd.n922 Vdd.n918 6.25878
R1399 Vdd.n275 Vdd.n271 6.25878
R1400 Vdd.n960 Vdd.n956 6.25878
R1401 Vdd.n752 Vdd.n748 6.25878
R1402 Vdd.n665 Vdd.n661 6.25878
R1403 Vdd.n791 Vdd.n787 6.25878
R1404 Vdd.n391 Vdd.n387 6.25878
R1405 Vdd.n829 Vdd.n825 6.25878
R1406 Vdd.n361 Vdd.n357 6.25878
R1407 Vdd.n867 Vdd.n863 6.25878
R1408 Vdd.n325 Vdd.n321 6.25878
R1409 Vdd.n906 Vdd.n902 6.25878
R1410 Vdd.n295 Vdd.n291 6.25878
R1411 Vdd.n944 Vdd.n940 6.25878
R1412 Vdd.n265 Vdd.n261 6.25878
R1413 Vdd.n680 Vdd.n676 6.25878
R1414 Vdd.n406 Vdd.n402 6.25878
R1415 Vdd.n376 Vdd.n372 6.25878
R1416 Vdd.n346 Vdd.n342 6.25878
R1417 Vdd.n310 Vdd.n306 6.25878
R1418 Vdd.n280 Vdd.n276 6.25878
R1419 Vdd.n747 Vdd.n743 6.25878
R1420 Vdd.n685 Vdd.n681 6.25878
R1421 Vdd.n786 Vdd.n782 6.25878
R1422 Vdd.n763 Vdd.n759 6.25878
R1423 Vdd.n411 Vdd.n407 6.25878
R1424 Vdd.n824 Vdd.n820 6.25878
R1425 Vdd.n802 Vdd.n798 6.25878
R1426 Vdd.n381 Vdd.n377 6.25878
R1427 Vdd.n862 Vdd.n858 6.25878
R1428 Vdd.n840 Vdd.n836 6.25878
R1429 Vdd.n351 Vdd.n347 6.25878
R1430 Vdd.n901 Vdd.n897 6.25878
R1431 Vdd.n879 Vdd.n875 6.25878
R1432 Vdd.n315 Vdd.n311 6.25878
R1433 Vdd.n939 Vdd.n935 6.25878
R1434 Vdd.n917 Vdd.n913 6.25878
R1435 Vdd.n285 Vdd.n281 6.25878
R1436 Vdd.n955 Vdd.n951 6.25878
R1437 Vdd.n742 Vdd.n738 6.25878
R1438 Vdd.n670 Vdd.n666 6.25878
R1439 Vdd.n781 Vdd.n777 6.25878
R1440 Vdd.n396 Vdd.n392 6.25878
R1441 Vdd.n819 Vdd.n815 6.25878
R1442 Vdd.n366 Vdd.n362 6.25878
R1443 Vdd.n857 Vdd.n853 6.25878
R1444 Vdd.n330 Vdd.n326 6.25878
R1445 Vdd.n896 Vdd.n892 6.25878
R1446 Vdd.n300 Vdd.n296 6.25878
R1447 Vdd.n934 Vdd.n930 6.25878
R1448 Vdd.n270 Vdd.n266 6.25878
R1449 Vdd.n690 Vdd.n686 6.25878
R1450 Vdd.n416 Vdd.n412 6.25878
R1451 Vdd.n386 Vdd.n382 6.25878
R1452 Vdd.n356 Vdd.n352 6.25878
R1453 Vdd.n320 Vdd.n316 6.25878
R1454 Vdd.n290 Vdd.n286 6.25878
R1455 Vdd.n695 Vdd.n691 6.25878
R1456 Vdd.n711 Vdd.n707 6.25878
R1457 Vdd.n706 Vdd.n702 6.25878
R1458 Vdd.n729 Vdd.n725 6.25878
R1459 Vdd.n735 Vdd.n731 6.25878
R1460 Vdd.n723 Vdd.n719 6.25878
R1461 Vdd.n628 Vdd.n624 6.25878
R1462 Vdd.n639 Vdd.n635 6.25878
R1463 Vdd.n634 Vdd.n630 6.25878
R1464 Vdd.n651 Vdd.n647 6.25878
R1465 Vdd.n645 Vdd.n641 6.25878
R1466 Vdd.n658 Vdd.n654 6.25878
R1467 Vdd.n559 Vdd.n555 6.25878
R1468 Vdd.n570 Vdd.n566 6.25878
R1469 Vdd.n565 Vdd.n561 6.25878
R1470 Vdd.n582 Vdd.n578 6.25878
R1471 Vdd.n576 Vdd.n572 6.25878
R1472 Vdd.n589 Vdd.n585 6.25878
R1473 Vdd.n196 Vdd.n195 5.93546
R1474 Vdd.n83 Vdd.n82 5.93546
R1475 Vdd.n156 Vdd.n155 5.93546
R1476 Vdd.n966 Vdd.n965 5.93546
R1477 Vdd.n718 Vdd.n717 5.93546
R1478 Vdd.n421 Vdd.n420 5.93546
R1479 Vdd.n335 Vdd.n334 5.93546
R1480 Vdd.n714 Vdd.n713 5.7305
R1481 SARlogic_0.dffrs_13.nand3_8.B Vdd.n716 5.47979
R1482 SARlogic_0.dffrs_13.nand3_1.B Vdd.n715 5.47979
R1483 Vdd.n7 Vdd.n6 5.44497
R1484 Vdd.n1098 Vdd.n1097 5.44497
R1485 Vdd.n12 Vdd.n11 5.44497
R1486 Vdd.n1086 Vdd.n1085 5.44497
R1487 Vdd.n1092 Vdd.n1091 5.44497
R1488 Vdd.n1079 Vdd.n1078 5.44497
R1489 Vdd.n54 Vdd.n53 5.44497
R1490 Vdd.n65 Vdd.n64 5.44497
R1491 Vdd.n60 Vdd.n59 5.44497
R1492 Vdd.n77 Vdd.n76 5.44497
R1493 Vdd.n71 Vdd.n70 5.44497
R1494 Vdd.n88 Vdd.n87 5.44497
R1495 Vdd.n127 Vdd.n126 5.44497
R1496 Vdd.n138 Vdd.n137 5.44497
R1497 Vdd.n133 Vdd.n132 5.44497
R1498 Vdd.n150 Vdd.n149 5.44497
R1499 Vdd.n144 Vdd.n143 5.44497
R1500 Vdd.n161 Vdd.n160 5.44497
R1501 Vdd.n207 Vdd.n206 5.44497
R1502 Vdd.n212 Vdd.n211 5.44497
R1503 Vdd.n201 Vdd.n200 5.44497
R1504 Vdd.n1004 Vdd.n1003 5.44497
R1505 Vdd.n987 Vdd.n986 5.44497
R1506 Vdd.n992 Vdd.n991 5.44497
R1507 Vdd.n998 Vdd.n997 5.44497
R1508 Vdd.n980 Vdd.n979 5.44497
R1509 Vdd.n508 Vdd.n507 5.44497
R1510 Vdd.n514 Vdd.n513 5.44497
R1511 Vdd.n520 Vdd.n519 5.44497
R1512 Vdd.n971 Vdd.n970 5.44497
R1513 Vdd.n757 Vdd.n756 5.44497
R1514 Vdd.n796 Vdd.n795 5.44497
R1515 Vdd.n834 Vdd.n833 5.44497
R1516 Vdd.n872 Vdd.n871 5.44497
R1517 Vdd.n911 Vdd.n910 5.44497
R1518 Vdd.n949 Vdd.n948 5.44497
R1519 Vdd.n675 Vdd.n674 5.44497
R1520 Vdd.n768 Vdd.n767 5.44497
R1521 Vdd.n401 Vdd.n400 5.44497
R1522 Vdd.n807 Vdd.n806 5.44497
R1523 Vdd.n371 Vdd.n370 5.44497
R1524 Vdd.n845 Vdd.n844 5.44497
R1525 Vdd.n341 Vdd.n340 5.44497
R1526 Vdd.n884 Vdd.n883 5.44497
R1527 Vdd.n305 Vdd.n304 5.44497
R1528 Vdd.n922 Vdd.n921 5.44497
R1529 Vdd.n275 Vdd.n274 5.44497
R1530 Vdd.n960 Vdd.n959 5.44497
R1531 Vdd.n752 Vdd.n751 5.44497
R1532 Vdd.n665 Vdd.n664 5.44497
R1533 Vdd.n791 Vdd.n790 5.44497
R1534 Vdd.n391 Vdd.n390 5.44497
R1535 Vdd.n829 Vdd.n828 5.44497
R1536 Vdd.n361 Vdd.n360 5.44497
R1537 Vdd.n867 Vdd.n866 5.44497
R1538 Vdd.n325 Vdd.n324 5.44497
R1539 Vdd.n906 Vdd.n905 5.44497
R1540 Vdd.n295 Vdd.n294 5.44497
R1541 Vdd.n944 Vdd.n943 5.44497
R1542 Vdd.n265 Vdd.n264 5.44497
R1543 Vdd.n680 Vdd.n679 5.44497
R1544 Vdd.n406 Vdd.n405 5.44497
R1545 Vdd.n376 Vdd.n375 5.44497
R1546 Vdd.n346 Vdd.n345 5.44497
R1547 Vdd.n310 Vdd.n309 5.44497
R1548 Vdd.n280 Vdd.n279 5.44497
R1549 Vdd.n747 Vdd.n746 5.44497
R1550 Vdd.n685 Vdd.n684 5.44497
R1551 Vdd.n786 Vdd.n785 5.44497
R1552 Vdd.n763 Vdd.n762 5.44497
R1553 Vdd.n411 Vdd.n410 5.44497
R1554 Vdd.n824 Vdd.n823 5.44497
R1555 Vdd.n802 Vdd.n801 5.44497
R1556 Vdd.n381 Vdd.n380 5.44497
R1557 Vdd.n862 Vdd.n861 5.44497
R1558 Vdd.n840 Vdd.n839 5.44497
R1559 Vdd.n351 Vdd.n350 5.44497
R1560 Vdd.n901 Vdd.n900 5.44497
R1561 Vdd.n879 Vdd.n878 5.44497
R1562 Vdd.n315 Vdd.n314 5.44497
R1563 Vdd.n939 Vdd.n938 5.44497
R1564 Vdd.n917 Vdd.n916 5.44497
R1565 Vdd.n285 Vdd.n284 5.44497
R1566 Vdd.n955 Vdd.n954 5.44497
R1567 Vdd.n742 Vdd.n741 5.44497
R1568 Vdd.n670 Vdd.n669 5.44497
R1569 Vdd.n781 Vdd.n780 5.44497
R1570 Vdd.n396 Vdd.n395 5.44497
R1571 Vdd.n819 Vdd.n818 5.44497
R1572 Vdd.n366 Vdd.n365 5.44497
R1573 Vdd.n857 Vdd.n856 5.44497
R1574 Vdd.n330 Vdd.n329 5.44497
R1575 Vdd.n896 Vdd.n895 5.44497
R1576 Vdd.n300 Vdd.n299 5.44497
R1577 Vdd.n934 Vdd.n933 5.44497
R1578 Vdd.n270 Vdd.n269 5.44497
R1579 Vdd.n690 Vdd.n689 5.44497
R1580 Vdd.n416 Vdd.n415 5.44497
R1581 Vdd.n386 Vdd.n385 5.44497
R1582 Vdd.n356 Vdd.n355 5.44497
R1583 Vdd.n320 Vdd.n319 5.44497
R1584 Vdd.n290 Vdd.n289 5.44497
R1585 Vdd.n695 Vdd.n694 5.44497
R1586 Vdd.n711 Vdd.n710 5.44497
R1587 Vdd.n706 Vdd.n705 5.44497
R1588 Vdd.n729 Vdd.n728 5.44497
R1589 Vdd.n735 Vdd.n734 5.44497
R1590 Vdd.n723 Vdd.n722 5.44497
R1591 Vdd.n628 Vdd.n627 5.44497
R1592 Vdd.n639 Vdd.n638 5.44497
R1593 Vdd.n634 Vdd.n633 5.44497
R1594 Vdd.n651 Vdd.n650 5.44497
R1595 Vdd.n645 Vdd.n644 5.44497
R1596 Vdd.n658 Vdd.n657 5.44497
R1597 Vdd.n559 Vdd.n558 5.44497
R1598 Vdd.n570 Vdd.n569 5.44497
R1599 Vdd.n565 Vdd.n564 5.44497
R1600 Vdd.n582 Vdd.n581 5.44497
R1601 Vdd.n576 Vdd.n575 5.44497
R1602 Vdd.n589 Vdd.n588 5.44497
R1603 Vdd.n48 Vdd.n47 5.14711
R1604 Vdd.n121 Vdd.n120 5.14711
R1605 Vdd.n502 Vdd.n501 5.14711
R1606 Vdd.n774 Vdd.n773 5.14711
R1607 Vdd.n812 Vdd.n811 5.14711
R1608 Vdd.n850 Vdd.n849 5.14711
R1609 Vdd.n889 Vdd.n888 5.14711
R1610 Vdd.n927 Vdd.n926 5.14711
R1611 Vdd.n699 Vdd.n698 5.14711
R1612 Vdd.n553 Vdd.n552 5.14711
R1613 Vdd.n622 Vdd.n621 5.14711
R1614 Vdd.n2 Vdd.n1 5.14711
R1615 Vdd.n772 Vdd.n771 5.13907
R1616 Vdd.n810 Vdd.n809 5.13907
R1617 Vdd.n848 Vdd.n847 5.13907
R1618 Vdd.n887 Vdd.n886 5.13907
R1619 Vdd.n925 Vdd.n924 5.13907
R1620 Vdd.n697 Vdd.n696 5.13907
R1621 Vdd.n717 SARlogic_0.dffrs_13.nand3_8.B 5.09593
R1622 Vdd.n1072 Vdd.n1071 4.98176
R1623 Vdd.n1017 Vdd.t243 4.4205
R1624 Vdd.n1010 Vdd.t321 4.4205
R1625 Vdd.n975 Vdd.n260 4.3905
R1626 Vdd.n1028 Vdd.t788 3.38176
R1627 Vdd.n178 Vdd.n177 2.49936
R1628 Vdd.n105 Vdd.n104 2.49936
R1629 Vdd.n243 Vdd.n242 2.49936
R1630 Vdd.n606 Vdd.n605 2.49936
R1631 Vdd.n537 Vdd.n536 2.49936
R1632 Vdd.n465 Vdd.n464 2.49936
R1633 Vdd.n1042 Vdd.n1041 2.1905
R1634 Vdd.n1060 Vdd.n1059 2.1905
R1635 Vdd.n1023 Vdd.n1022 2.16583
R1636 Vdd.n1025 Vdd.n1024 2.16583
R1637 Vdd.n1009 Vdd.t289 1.99236
R1638 Vdd.n177 Vdd.n166 1.93883
R1639 Vdd.n104 Vdd.n93 1.93883
R1640 Vdd.n242 Vdd.n231 1.93883
R1641 Vdd.n605 Vdd.n594 1.93883
R1642 Vdd.n536 Vdd.n525 1.93883
R1643 Vdd.n464 Vdd.n453 1.93883
R1644 Vdd.n1019 Vdd.t343 1.91107
R1645 Vdd.n981 Vdd.n975 1.89424
R1646 Vdd.n6 Vdd.t669 1.85637
R1647 Vdd.n1097 Vdd.t95 1.85637
R1648 Vdd.n11 Vdd.t690 1.85637
R1649 Vdd.n1085 Vdd.t864 1.85637
R1650 Vdd.n1091 Vdd.t253 1.85637
R1651 Vdd.n1078 Vdd.t181 1.85637
R1652 Vdd.n53 Vdd.t717 1.85637
R1653 Vdd.n64 Vdd.t131 1.85637
R1654 Vdd.n59 Vdd.t606 1.85637
R1655 Vdd.n76 Vdd.t844 1.85637
R1656 Vdd.n70 Vdd.t29 1.85637
R1657 Vdd.n87 Vdd.t55 1.85637
R1658 Vdd.n126 Vdd.t696 1.85637
R1659 Vdd.n137 Vdd.t796 1.85637
R1660 Vdd.n132 Vdd.t708 1.85637
R1661 Vdd.n149 Vdd.t744 1.85637
R1662 Vdd.n143 Vdd.t513 1.85637
R1663 Vdd.n160 Vdd.t187 1.85637
R1664 Vdd.n206 Vdd.t627 1.85637
R1665 Vdd.n211 Vdd.t355 1.85637
R1666 Vdd.n200 Vdd.t427 1.85637
R1667 Vdd.n1003 Vdd.t103 1.85637
R1668 Vdd.n986 Vdd.t429 1.85637
R1669 Vdd.n991 Vdd.t930 1.85637
R1670 Vdd.n997 Vdd.t499 1.85637
R1671 Vdd.n979 Vdd.t509 1.85637
R1672 Vdd.n507 Vdd.t612 1.85637
R1673 Vdd.n513 Vdd.t333 1.85637
R1674 Vdd.n519 Vdd.t547 1.85637
R1675 Vdd.n970 Vdd.t307 1.85637
R1676 Vdd.n756 Vdd.t936 1.85637
R1677 Vdd.n795 Vdd.t199 1.85637
R1678 Vdd.n833 Vdd.t493 1.85637
R1679 Vdd.n871 Vdd.t882 1.85637
R1680 Vdd.n910 Vdd.t397 1.85637
R1681 Vdd.n948 Vdd.t860 1.85637
R1682 Vdd.n674 Vdd.t87 1.85637
R1683 Vdd.n767 Vdd.t940 1.85637
R1684 Vdd.n400 Vdd.t425 1.85637
R1685 Vdd.n806 Vdd.t195 1.85637
R1686 Vdd.n370 Vdd.t329 1.85637
R1687 Vdd.n844 Vdd.t491 1.85637
R1688 Vdd.n340 Vdd.t285 1.85637
R1689 Vdd.n883 Vdd.t880 1.85637
R1690 Vdd.n304 Vdd.t109 1.85637
R1691 Vdd.n921 Vdd.t395 1.85637
R1692 Vdd.n274 Vdd.t447 1.85637
R1693 Vdd.n959 Vdd.t862 1.85637
R1694 Vdd.n751 Vdd.t481 1.85637
R1695 Vdd.n664 Vdd.t121 1.85637
R1696 Vdd.n790 Vdd.t798 1.85637
R1697 Vdd.n390 Vdd.t221 1.85637
R1698 Vdd.n828 Vdd.t193 1.85637
R1699 Vdd.n360 Vdd.t898 1.85637
R1700 Vdd.n866 Vdd.t916 1.85637
R1701 Vdd.n324 Vdd.t291 1.85637
R1702 Vdd.n905 Vdd.t129 1.85637
R1703 Vdd.n294 Vdd.t808 1.85637
R1704 Vdd.n943 Vdd.t569 1.85637
R1705 Vdd.n264 Vdd.t261 1.85637
R1706 Vdd.n679 Vdd.t748 1.85637
R1707 Vdd.n405 Vdd.t93 1.85637
R1708 Vdd.n375 Vdd.t311 1.85637
R1709 Vdd.n345 Vdd.t61 1.85637
R1710 Vdd.n309 Vdd.t245 1.85637
R1711 Vdd.n279 Vdd.t219 1.85637
R1712 Vdd.n746 Vdd.t702 1.85637
R1713 Vdd.n684 Vdd.t597 1.85637
R1714 Vdd.n785 Vdd.t609 1.85637
R1715 Vdd.n762 Vdd.t693 1.85637
R1716 Vdd.n410 Vdd.t423 1.85637
R1717 Vdd.n823 Vdd.t657 1.85637
R1718 Vdd.n801 Vdd.t651 1.85637
R1719 Vdd.n380 Vdd.t477 1.85637
R1720 Vdd.n861 Vdd.t705 1.85637
R1721 Vdd.n839 Vdd.t675 1.85637
R1722 Vdd.n350 Vdd.t189 1.85637
R1723 Vdd.n900 Vdd.t666 1.85637
R1724 Vdd.n878 Vdd.t723 1.85637
R1725 Vdd.n314 Vdd.t105 1.85637
R1726 Vdd.n938 Vdd.t711 1.85637
R1727 Vdd.n916 Vdd.t672 1.85637
R1728 Vdd.n284 Vdd.t239 1.85637
R1729 Vdd.n954 Vdd.t687 1.85637
R1730 Vdd.n741 Vdd.t565 1.85637
R1731 Vdd.n669 Vdd.t1 1.85637
R1732 Vdd.n780 Vdd.t275 1.85637
R1733 Vdd.n395 Vdd.t33 1.85637
R1734 Vdd.n818 Vdd.t501 1.85637
R1735 Vdd.n365 Vdd.t337 1.85637
R1736 Vdd.n856 Vdd.t433 1.85637
R1737 Vdd.n329 Vdd.t814 1.85637
R1738 Vdd.n895 Vdd.t832 1.85637
R1739 Vdd.n299 Vdd.t139 1.85637
R1740 Vdd.n933 Vdd.t922 1.85637
R1741 Vdd.n269 Vdd.t537 1.85637
R1742 Vdd.n689 Vdd.t21 1.85637
R1743 Vdd.n415 Vdd.t445 1.85637
R1744 Vdd.n385 Vdd.t934 1.85637
R1745 Vdd.n355 Vdd.t111 1.85637
R1746 Vdd.n319 Vdd.t521 1.85637
R1747 Vdd.n289 Vdd.t531 1.85637
R1748 Vdd.n694 Vdd.t401 1.85637
R1749 Vdd.n710 Vdd.t924 1.85637
R1750 Vdd.n705 Vdd.t387 1.85637
R1751 Vdd.n728 Vdd.t826 1.85637
R1752 Vdd.n734 Vdd.t794 1.85637
R1753 Vdd.n722 Vdd.t886 1.85637
R1754 Vdd.n627 Vdd.t615 1.85637
R1755 Vdd.n638 Vdd.t555 1.85637
R1756 Vdd.n633 Vdd.t654 1.85637
R1757 Vdd.n650 Vdd.t734 1.85637
R1758 Vdd.n644 Vdd.t39 1.85637
R1759 Vdd.n657 Vdd.t942 1.85637
R1760 Vdd.n558 Vdd.t600 1.85637
R1761 Vdd.n569 Vdd.t229 1.85637
R1762 Vdd.n564 Vdd.t621 1.85637
R1763 Vdd.n581 Vdd.t351 1.85637
R1764 Vdd.n575 Vdd.t267 1.85637
R1765 Vdd.n588 Vdd.t225 1.85637
R1766 Vdd.n1068 Vdd.n1020 1.83762
R1767 Vdd.n1070 Vdd.n1009 1.83762
R1768 Vdd.n1052 Vdd.t497 1.8205
R1769 Vdd.n1052 Vdd.t283 1.8205
R1770 Vdd.n1050 Vdd.t287 1.8205
R1771 Vdd.n1050 Vdd.t391 1.8205
R1772 Vdd.n1048 Vdd.t341 1.8205
R1773 Vdd.n1048 Vdd.t279 1.8205
R1774 Vdd.n1046 Vdd.t281 1.8205
R1775 Vdd.n1046 Vdd.t393 1.8205
R1776 Vdd.n1044 Vdd.t339 1.8205
R1777 Vdd.n1044 Vdd.t489 1.8205
R1778 Vdd.n437 Vdd.t850 1.80717
R1779 Vdd.n91 Vdd.n45 1.80479
R1780 Vdd.n164 Vdd.n29 1.80479
R1781 Vdd.n523 Vdd.n499 1.80479
R1782 Vdd.n592 Vdd.n483 1.80479
R1783 Vdd.n467 Vdd.n422 1.80479
R1784 Vdd.n221 Vdd.n13 1.80479
R1785 Vdd.n114 Vdd.n113 1.78583
R1786 Vdd.n187 Vdd.n186 1.78583
R1787 Vdd.n546 Vdd.n545 1.78583
R1788 Vdd.n615 Vdd.n614 1.78583
R1789 Vdd.n450 Vdd.n435 1.78583
R1790 Vdd.n247 Vdd.n246 1.78583
R1791 Vdd.n117 Vdd.t768 1.74654
R1792 Vdd.n190 Vdd.t589 1.74654
R1793 Vdd.n549 Vdd.t776 1.74654
R1794 Vdd.n618 Vdd.t782 1.74654
R1795 Vdd.n438 Vdd.t778 1.74654
R1796 Vdd.n255 Vdd.t766 1.74654
R1797 Vdd.n439 Vdd.n437 1.62809
R1798 Vdd.n1015 Vdd.n1014 1.5755
R1799 Vdd.n1017 Vdd.n1016 1.5755
R1800 Vdd.n1013 Vdd.n1010 1.5755
R1801 Vdd.n1056 Vdd.n1055 1.5755
R1802 Vdd.n1058 Vdd.n1057 1.5755
R1803 Vdd.n15 Vdd.t255 1.49467
R1804 Vdd.n174 Vdd.t331 1.49467
R1805 Vdd.n173 Vdd.t804 1.49467
R1806 Vdd.n31 Vdd.t511 1.49467
R1807 Vdd.n101 Vdd.t119 1.49467
R1808 Vdd.n100 Vdd.t263 1.49467
R1809 Vdd.n30 Vdd.t593 1.49467
R1810 Vdd.n14 Vdd.t774 1.49467
R1811 Vdd.n239 Vdd.t107 1.49467
R1812 Vdd.n238 Vdd.t295 1.49467
R1813 Vdd.n253 Vdd.t353 1.49467
R1814 Vdd.n252 Vdd.t780 1.49467
R1815 Vdd.n469 Vdd.t37 1.49467
R1816 Vdd.n602 Vdd.t97 1.49467
R1817 Vdd.n601 Vdd.t223 1.49467
R1818 Vdd.n485 Vdd.t269 1.49467
R1819 Vdd.n533 Vdd.t756 1.49467
R1820 Vdd.n532 Vdd.t894 1.49467
R1821 Vdd.n484 Vdd.t772 1.49467
R1822 Vdd.n468 Vdd.t770 1.49467
R1823 Vdd.n461 Vdd.t912 1.49467
R1824 Vdd.n460 Vdd.t123 1.49467
R1825 Vdd.n447 Vdd.t7 1.49467
R1826 Vdd.n446 Vdd.t591 1.49467
R1827 Vdd.n167 Vdd.t357 1.47383
R1828 Vdd.n94 Vdd.t858 1.47383
R1829 Vdd.n33 Vdd.t525 1.47383
R1830 Vdd.n34 Vdd.t527 1.47383
R1831 Vdd.n35 Vdd.t902 1.47383
R1832 Vdd.n32 Vdd.t567 1.47383
R1833 Vdd.n17 Vdd.t169 1.47383
R1834 Vdd.n18 Vdd.t167 1.47383
R1835 Vdd.n19 Vdd.t257 1.47383
R1836 Vdd.n16 Vdd.t846 1.47383
R1837 Vdd.n232 Vdd.t792 1.47383
R1838 Vdd.n595 Vdd.t63 1.47383
R1839 Vdd.n526 Vdd.t914 1.47383
R1840 Vdd.n487 Vdd.t904 1.47383
R1841 Vdd.n488 Vdd.t906 1.47383
R1842 Vdd.n489 Vdd.t179 1.47383
R1843 Vdd.n486 Vdd.t848 1.47383
R1844 Vdd.n471 Vdd.t890 1.47383
R1845 Vdd.n472 Vdd.t888 1.47383
R1846 Vdd.n473 Vdd.t345 1.47383
R1847 Vdd.n470 Vdd.t201 1.47383
R1848 Vdd.n454 Vdd.t539 1.47383
R1849 Vdd.n436 Vdd.t319 1.47383
R1850 Vdd.n434 Vdd.t165 1.47383
R1851 Vdd.n424 Vdd.t163 1.47383
R1852 Vdd.n423 Vdd.t171 1.47383
R1853 Vdd.n248 Vdd.t117 1.47383
R1854 Vdd.n217 Vdd.t99 1.47383
R1855 Vdd.n218 Vdd.t101 1.47383
R1856 Vdd.n229 Vdd.t191 1.47383
R1857 Vdd.n163 Vdd.n118 1.19311
R1858 Vdd.n1081 Vdd.n191 1.19311
R1859 Vdd.n584 Vdd.n550 1.19311
R1860 Vdd.n653 Vdd.n619 1.19311
R1861 Vdd.n257 Vdd.n256 1.19311
R1862 Vdd.n1022 Vdd.t786 1.13285
R1863 Vdd.n1022 Vdd.t790 1.13285
R1864 Vdd.n1024 Vdd.t323 1.13285
R1865 Vdd.n1024 Vdd.t784 1.13285
R1866 Vdd.n1069 Vdd.n1018 1.058
R1867 Vdd.n6 Vdd.n5 1.04105
R1868 Vdd.n1097 Vdd.n1096 1.04105
R1869 Vdd.n11 Vdd.n10 1.04105
R1870 Vdd.n1085 Vdd.n1084 1.04105
R1871 Vdd.n1091 Vdd.n1090 1.04105
R1872 Vdd.n1078 Vdd.n1077 1.04105
R1873 Vdd.n53 Vdd.n52 1.04105
R1874 Vdd.n64 Vdd.n63 1.04105
R1875 Vdd.n59 Vdd.n58 1.04105
R1876 Vdd.n76 Vdd.n75 1.04105
R1877 Vdd.n70 Vdd.n69 1.04105
R1878 Vdd.n87 Vdd.n86 1.04105
R1879 Vdd.n126 Vdd.n125 1.04105
R1880 Vdd.n137 Vdd.n136 1.04105
R1881 Vdd.n132 Vdd.n131 1.04105
R1882 Vdd.n149 Vdd.n148 1.04105
R1883 Vdd.n143 Vdd.n142 1.04105
R1884 Vdd.n160 Vdd.n159 1.04105
R1885 Vdd.n206 Vdd.n205 1.04105
R1886 Vdd.n211 Vdd.n210 1.04105
R1887 Vdd.n200 Vdd.n199 1.04105
R1888 Vdd.n1003 Vdd.n1002 1.04105
R1889 Vdd.n986 Vdd.n985 1.04105
R1890 Vdd.n991 Vdd.n990 1.04105
R1891 Vdd.n997 Vdd.n996 1.04105
R1892 Vdd.n979 Vdd.n978 1.04105
R1893 Vdd.n507 Vdd.n506 1.04105
R1894 Vdd.n513 Vdd.n512 1.04105
R1895 Vdd.n519 Vdd.n518 1.04105
R1896 Vdd.n970 Vdd.n969 1.04105
R1897 Vdd.n756 Vdd.n755 1.04105
R1898 Vdd.n795 Vdd.n794 1.04105
R1899 Vdd.n833 Vdd.n832 1.04105
R1900 Vdd.n871 Vdd.n870 1.04105
R1901 Vdd.n910 Vdd.n909 1.04105
R1902 Vdd.n948 Vdd.n947 1.04105
R1903 Vdd.n674 Vdd.n673 1.04105
R1904 Vdd.n767 Vdd.n766 1.04105
R1905 Vdd.n400 Vdd.n399 1.04105
R1906 Vdd.n806 Vdd.n805 1.04105
R1907 Vdd.n370 Vdd.n369 1.04105
R1908 Vdd.n844 Vdd.n843 1.04105
R1909 Vdd.n340 Vdd.n339 1.04105
R1910 Vdd.n883 Vdd.n882 1.04105
R1911 Vdd.n304 Vdd.n303 1.04105
R1912 Vdd.n921 Vdd.n920 1.04105
R1913 Vdd.n274 Vdd.n273 1.04105
R1914 Vdd.n959 Vdd.n958 1.04105
R1915 Vdd.n751 Vdd.n750 1.04105
R1916 Vdd.n664 Vdd.n663 1.04105
R1917 Vdd.n790 Vdd.n789 1.04105
R1918 Vdd.n390 Vdd.n389 1.04105
R1919 Vdd.n828 Vdd.n827 1.04105
R1920 Vdd.n360 Vdd.n359 1.04105
R1921 Vdd.n866 Vdd.n865 1.04105
R1922 Vdd.n324 Vdd.n323 1.04105
R1923 Vdd.n905 Vdd.n904 1.04105
R1924 Vdd.n294 Vdd.n293 1.04105
R1925 Vdd.n943 Vdd.n942 1.04105
R1926 Vdd.n264 Vdd.n263 1.04105
R1927 Vdd.n679 Vdd.n678 1.04105
R1928 Vdd.n405 Vdd.n404 1.04105
R1929 Vdd.n375 Vdd.n374 1.04105
R1930 Vdd.n345 Vdd.n344 1.04105
R1931 Vdd.n309 Vdd.n308 1.04105
R1932 Vdd.n279 Vdd.n278 1.04105
R1933 Vdd.n746 Vdd.n745 1.04105
R1934 Vdd.n684 Vdd.n683 1.04105
R1935 Vdd.n785 Vdd.n784 1.04105
R1936 Vdd.n762 Vdd.n761 1.04105
R1937 Vdd.n410 Vdd.n409 1.04105
R1938 Vdd.n823 Vdd.n822 1.04105
R1939 Vdd.n801 Vdd.n800 1.04105
R1940 Vdd.n380 Vdd.n379 1.04105
R1941 Vdd.n861 Vdd.n860 1.04105
R1942 Vdd.n839 Vdd.n838 1.04105
R1943 Vdd.n350 Vdd.n349 1.04105
R1944 Vdd.n900 Vdd.n899 1.04105
R1945 Vdd.n878 Vdd.n877 1.04105
R1946 Vdd.n314 Vdd.n313 1.04105
R1947 Vdd.n938 Vdd.n937 1.04105
R1948 Vdd.n916 Vdd.n915 1.04105
R1949 Vdd.n284 Vdd.n283 1.04105
R1950 Vdd.n954 Vdd.n953 1.04105
R1951 Vdd.n741 Vdd.n740 1.04105
R1952 Vdd.n669 Vdd.n668 1.04105
R1953 Vdd.n780 Vdd.n779 1.04105
R1954 Vdd.n395 Vdd.n394 1.04105
R1955 Vdd.n818 Vdd.n817 1.04105
R1956 Vdd.n365 Vdd.n364 1.04105
R1957 Vdd.n856 Vdd.n855 1.04105
R1958 Vdd.n329 Vdd.n328 1.04105
R1959 Vdd.n895 Vdd.n894 1.04105
R1960 Vdd.n299 Vdd.n298 1.04105
R1961 Vdd.n933 Vdd.n932 1.04105
R1962 Vdd.n269 Vdd.n268 1.04105
R1963 Vdd.n689 Vdd.n688 1.04105
R1964 Vdd.n415 Vdd.n414 1.04105
R1965 Vdd.n385 Vdd.n384 1.04105
R1966 Vdd.n355 Vdd.n354 1.04105
R1967 Vdd.n319 Vdd.n318 1.04105
R1968 Vdd.n289 Vdd.n288 1.04105
R1969 Vdd.n694 Vdd.n693 1.04105
R1970 Vdd.n710 Vdd.n709 1.04105
R1971 Vdd.n705 Vdd.n704 1.04105
R1972 Vdd.n728 Vdd.n727 1.04105
R1973 Vdd.n734 Vdd.n733 1.04105
R1974 Vdd.n722 Vdd.n721 1.04105
R1975 Vdd.n627 Vdd.n626 1.04105
R1976 Vdd.n638 Vdd.n637 1.04105
R1977 Vdd.n633 Vdd.n632 1.04105
R1978 Vdd.n650 Vdd.n649 1.04105
R1979 Vdd.n644 Vdd.n643 1.04105
R1980 Vdd.n657 Vdd.n656 1.04105
R1981 Vdd.n558 Vdd.n557 1.04105
R1982 Vdd.n569 Vdd.n568 1.04105
R1983 Vdd.n564 Vdd.n563 1.04105
R1984 Vdd.n581 Vdd.n580 1.04105
R1985 Vdd.n575 Vdd.n574 1.04105
R1986 Vdd.n588 Vdd.n587 1.04105
R1987 Vdd.n1018 Vdd.n1010 1.01373
R1988 Vdd.n1018 Vdd.n1017 0.979984
R1989 Vdd.n91 Vdd.n90 0.809622
R1990 Vdd.n164 Vdd.n163 0.809622
R1991 Vdd.n523 Vdd.n522 0.809622
R1992 Vdd.n592 Vdd.n591 0.809622
R1993 Vdd.n653 Vdd.n467 0.809622
R1994 Vdd.n1081 Vdd.n13 0.809622
R1995 Vdd.n170 Vdd.n167 0.788
R1996 Vdd.n171 Vdd.n170 0.788
R1997 Vdd.n173 Vdd.n172 0.788
R1998 Vdd.n97 Vdd.n94 0.788
R1999 Vdd.n98 Vdd.n97 0.788
R2000 Vdd.n100 Vdd.n99 0.788
R2001 Vdd.n41 Vdd.n34 0.788
R2002 Vdd.n42 Vdd.n41 0.788
R2003 Vdd.n43 Vdd.n35 0.788
R2004 Vdd.n44 Vdd.n43 0.788
R2005 Vdd.n39 Vdd.n33 0.788
R2006 Vdd.n111 Vdd.n32 0.788
R2007 Vdd.n112 Vdd.n111 0.788
R2008 Vdd.n110 Vdd.n30 0.788
R2009 Vdd.n25 Vdd.n18 0.788
R2010 Vdd.n26 Vdd.n25 0.788
R2011 Vdd.n27 Vdd.n19 0.788
R2012 Vdd.n28 Vdd.n27 0.788
R2013 Vdd.n23 Vdd.n17 0.788
R2014 Vdd.n184 Vdd.n16 0.788
R2015 Vdd.n185 Vdd.n184 0.788
R2016 Vdd.n183 Vdd.n14 0.788
R2017 Vdd.n235 Vdd.n232 0.788
R2018 Vdd.n236 Vdd.n235 0.788
R2019 Vdd.n238 Vdd.n237 0.788
R2020 Vdd.n598 Vdd.n595 0.788
R2021 Vdd.n599 Vdd.n598 0.788
R2022 Vdd.n601 Vdd.n600 0.788
R2023 Vdd.n529 Vdd.n526 0.788
R2024 Vdd.n530 Vdd.n529 0.788
R2025 Vdd.n532 Vdd.n531 0.788
R2026 Vdd.n495 Vdd.n488 0.788
R2027 Vdd.n496 Vdd.n495 0.788
R2028 Vdd.n497 Vdd.n489 0.788
R2029 Vdd.n498 Vdd.n497 0.788
R2030 Vdd.n493 Vdd.n487 0.788
R2031 Vdd.n543 Vdd.n486 0.788
R2032 Vdd.n544 Vdd.n543 0.788
R2033 Vdd.n542 Vdd.n484 0.788
R2034 Vdd.n479 Vdd.n472 0.788
R2035 Vdd.n480 Vdd.n479 0.788
R2036 Vdd.n481 Vdd.n473 0.788
R2037 Vdd.n482 Vdd.n481 0.788
R2038 Vdd.n477 Vdd.n471 0.788
R2039 Vdd.n612 Vdd.n470 0.788
R2040 Vdd.n613 Vdd.n612 0.788
R2041 Vdd.n611 Vdd.n468 0.788
R2042 Vdd.n457 Vdd.n454 0.788
R2043 Vdd.n458 Vdd.n457 0.788
R2044 Vdd.n460 Vdd.n459 0.788
R2045 Vdd.n443 Vdd.n436 0.788
R2046 Vdd.n444 Vdd.n443 0.788
R2047 Vdd.n446 Vdd.n445 0.788
R2048 Vdd.n431 Vdd.n424 0.788
R2049 Vdd.n432 Vdd.n431 0.788
R2050 Vdd.n429 Vdd.n423 0.788
R2051 Vdd.n430 Vdd.n429 0.788
R2052 Vdd.n434 Vdd.n433 0.788
R2053 Vdd.n249 Vdd.n248 0.788
R2054 Vdd.n250 Vdd.n249 0.788
R2055 Vdd.n252 Vdd.n251 0.788
R2056 Vdd.n225 Vdd.n218 0.788
R2057 Vdd.n226 Vdd.n225 0.788
R2058 Vdd.n229 Vdd.n228 0.788
R2059 Vdd.n228 Vdd.n227 0.788
R2060 Vdd.n223 Vdd.n217 0.788
R2061 Vdd.n49 Vdd.n48 0.754571
R2062 Vdd.n122 Vdd.n121 0.754571
R2063 Vdd.n503 Vdd.n502 0.754571
R2064 Vdd.n554 Vdd.n553 0.754571
R2065 Vdd.n623 Vdd.n622 0.754571
R2066 Vdd.n1101 Vdd.n2 0.754571
R2067 Vdd.n1067 Vdd.n1032 0.750875
R2068 Vdd.n3 Vdd.t866 0.7285
R2069 Vdd.n3 Vdd.t153 0.7285
R2070 Vdd.n1094 Vdd.t874 0.7285
R2071 Vdd.n1094 Vdd.t660 0.7285
R2072 Vdd.n8 Vdd.t517 0.7285
R2073 Vdd.n8 Vdd.t868 0.7285
R2074 Vdd.n1082 Vdd.t155 0.7285
R2075 Vdd.n1082 Vdd.t872 0.7285
R2076 Vdd.n1088 Vdd.t663 0.7285
R2077 Vdd.n1088 Vdd.t183 0.7285
R2078 Vdd.n1075 Vdd.t820 0.7285
R2079 Vdd.n1075 Vdd.t699 0.7285
R2080 Vdd.n50 Vdd.t840 0.7285
R2081 Vdd.n50 Vdd.t327 0.7285
R2082 Vdd.n61 Vdd.t233 0.7285
R2083 Vdd.n61 Vdd.t603 0.7285
R2084 Vdd.n56 Vdd.t487 0.7285
R2085 Vdd.n56 Vdd.t842 0.7285
R2086 Vdd.n73 Vdd.t325 0.7285
R2087 Vdd.n73 Vdd.t237 0.7285
R2088 Vdd.n67 Vdd.t645 0.7285
R2089 Vdd.n67 Vdd.t53 0.7285
R2090 Vdd.n84 Vdd.t838 0.7285
R2091 Vdd.n84 Vdd.t639 0.7285
R2092 Vdd.n123 Vdd.t740 0.7285
R2093 Vdd.n123 Vdd.t822 0.7285
R2094 Vdd.n134 Vdd.t852 0.7285
R2095 Vdd.n134 Vdd.t726 0.7285
R2096 Vdd.n129 Vdd.t926 0.7285
R2097 Vdd.n129 Vdd.t742 0.7285
R2098 Vdd.n146 Vdd.t818 0.7285
R2099 Vdd.n146 Vdd.t49 0.7285
R2100 Vdd.n140 Vdd.t732 0.7285
R2101 Vdd.n140 Vdd.t185 0.7285
R2102 Vdd.n157 Vdd.t115 0.7285
R2103 Vdd.n157 Vdd.t624 0.7285
R2104 Vdd.n203 Vdd.t515 0.7285
R2105 Vdd.n203 Vdd.t549 0.7285
R2106 Vdd.n208 Vdd.t648 0.7285
R2107 Vdd.n208 Vdd.t309 0.7285
R2108 Vdd.n197 Vdd.t928 0.7285
R2109 Vdd.n197 Vdd.t760 0.7285
R2110 Vdd.n1000 Vdd.t13 0.7285
R2111 Vdd.n1000 Vdd.t459 0.7285
R2112 Vdd.n983 Vdd.t507 0.7285
R2113 Vdd.n983 Vdd.t479 0.7285
R2114 Vdd.n988 Vdd.t758 0.7285
R2115 Vdd.n988 Vdd.t9 0.7285
R2116 Vdd.n994 Vdd.t365 0.7285
R2117 Vdd.n994 Vdd.t3 0.7285
R2118 Vdd.n976 Vdd.t5 0.7285
R2119 Vdd.n976 Vdd.t463 0.7285
R2120 Vdd.n504 Vdd.t816 0.7285
R2121 Vdd.n504 Vdd.t856 0.7285
R2122 Vdd.n510 Vdd.t878 0.7285
R2123 Vdd.n510 Vdd.t642 0.7285
R2124 Vdd.n516 Vdd.t854 0.7285
R2125 Vdd.n516 Vdd.t876 0.7285
R2126 Vdd.n967 Vdd.t884 0.7285
R2127 Vdd.n967 Vdd.t684 0.7285
R2128 Vdd.n753 Vdd.t485 0.7285
R2129 Vdd.n753 Vdd.t207 0.7285
R2130 Vdd.n792 Vdd.t802 0.7285
R2131 Vdd.n792 Vdd.t209 0.7285
R2132 Vdd.n830 Vdd.t41 0.7285
R2133 Vdd.n830 Vdd.t317 0.7285
R2134 Vdd.n868 Vdd.t918 0.7285
R2135 Vdd.n868 Vdd.t159 0.7285
R2136 Vdd.n907 Vdd.t125 0.7285
R2137 Vdd.n907 Vdd.t17 0.7285
R2138 Vdd.n945 Vdd.t573 0.7285
R2139 Vdd.n945 Vdd.t173 0.7285
R2140 Vdd.n671 Vdd.t249 0.7285
R2141 Vdd.n671 Vdd.t519 0.7285
R2142 Vdd.n764 Vdd.t203 0.7285
R2143 Vdd.n764 Vdd.t483 0.7285
R2144 Vdd.n397 Vdd.t896 0.7285
R2145 Vdd.n397 Vdd.t471 0.7285
R2146 Vdd.n803 Vdd.t541 0.7285
R2147 Vdd.n803 Vdd.t800 0.7285
R2148 Vdd.n367 Vdd.t293 0.7285
R2149 Vdd.n367 Vdd.t461 0.7285
R2150 Vdd.n841 Vdd.t241 0.7285
R2151 Vdd.n841 Vdd.t43 0.7285
R2152 Vdd.n337 Vdd.t810 0.7285
R2153 Vdd.n337 Vdd.t377 0.7285
R2154 Vdd.n880 Vdd.t89 0.7285
R2155 Vdd.n880 Vdd.t920 0.7285
R2156 Vdd.n301 Vdd.t259 0.7285
R2157 Vdd.n301 Vdd.t421 0.7285
R2158 Vdd.n918 Vdd.t750 0.7285
R2159 Vdd.n918 Vdd.t127 0.7285
R2160 Vdd.n271 Vdd.t535 0.7285
R2161 Vdd.n271 Vdd.t409 0.7285
R2162 Vdd.n956 Vdd.t133 0.7285
R2163 Vdd.n956 Vdd.t571 0.7285
R2164 Vdd.n748 Vdd.t205 0.7285
R2165 Vdd.n748 Vdd.t251 0.7285
R2166 Vdd.n661 Vdd.t467 0.7285
R2167 Vdd.n661 Vdd.t746 0.7285
R2168 Vdd.n787 Vdd.t211 0.7285
R2169 Vdd.n787 Vdd.t900 0.7285
R2170 Vdd.n387 Vdd.t385 0.7285
R2171 Vdd.n387 Vdd.t91 0.7285
R2172 Vdd.n825 Vdd.t315 0.7285
R2173 Vdd.n825 Vdd.t297 0.7285
R2174 Vdd.n357 Vdd.t367 0.7285
R2175 Vdd.n357 Vdd.t313 0.7285
R2176 Vdd.n863 Vdd.t161 0.7285
R2177 Vdd.n863 Vdd.t806 0.7285
R2178 Vdd.n321 Vdd.t371 0.7285
R2179 Vdd.n321 Vdd.t45 0.7285
R2180 Vdd.n902 Vdd.t19 0.7285
R2181 Vdd.n902 Vdd.t265 0.7285
R2182 Vdd.n291 Vdd.t361 0.7285
R2183 Vdd.n291 Vdd.t247 0.7285
R2184 Vdd.n940 Vdd.t175 0.7285
R2185 Vdd.n940 Vdd.t533 0.7285
R2186 Vdd.n261 Vdd.t405 0.7285
R2187 Vdd.n261 Vdd.t217 0.7285
R2188 Vdd.n676 Vdd.t545 0.7285
R2189 Vdd.n676 Vdd.t455 0.7285
R2190 Vdd.n402 Vdd.t561 0.7285
R2191 Vdd.n402 Vdd.t363 0.7285
R2192 Vdd.n372 Vdd.t559 0.7285
R2193 Vdd.n372 Vdd.t475 0.7285
R2194 Vdd.n342 Vdd.t543 0.7285
R2195 Vdd.n342 Vdd.t383 0.7285
R2196 Vdd.n306 Vdd.t557 0.7285
R2197 Vdd.n306 Vdd.t451 0.7285
R2198 Vdd.n276 Vdd.t563 0.7285
R2199 Vdd.n276 Vdd.t417 0.7285
R2200 Vdd.n743 Vdd.t57 0.7285
R2201 Vdd.n743 Vdd.t151 0.7285
R2202 Vdd.n681 Vdd.t69 0.7285
R2203 Vdd.n681 Vdd.t473 0.7285
R2204 Vdd.n782 Vdd.t277 0.7285
R2205 Vdd.n782 Vdd.t25 0.7285
R2206 Vdd.n759 Vdd.t197 0.7285
R2207 Vdd.n759 Vdd.t59 0.7285
R2208 Vdd.n407 Vdd.t581 0.7285
R2209 Vdd.n407 Vdd.t381 0.7285
R2210 Vdd.n820 Vdd.t505 0.7285
R2211 Vdd.n820 Vdd.t215 0.7285
R2212 Vdd.n798 Vdd.t495 0.7285
R2213 Vdd.n798 Vdd.t273 0.7285
R2214 Vdd.n377 Vdd.t83 0.7285
R2215 Vdd.n377 Vdd.t373 0.7285
R2216 Vdd.n858 Vdd.t435 0.7285
R2217 Vdd.n858 Vdd.t553 0.7285
R2218 Vdd.n836 Vdd.t870 0.7285
R2219 Vdd.n836 Vdd.t503 0.7285
R2220 Vdd.n347 Vdd.t65 0.7285
R2221 Vdd.n347 Vdd.t419 0.7285
R2222 Vdd.n897 Vdd.t834 0.7285
R2223 Vdd.n897 Vdd.t439 0.7285
R2224 Vdd.n875 Vdd.t399 0.7285
R2225 Vdd.n875 Vdd.t437 0.7285
R2226 Vdd.n311 Vdd.t77 0.7285
R2227 Vdd.n311 Vdd.t465 0.7285
R2228 Vdd.n935 Vdd.t754 0.7285
R2229 Vdd.n935 Vdd.t147 0.7285
R2230 Vdd.n913 Vdd.t305 0.7285
R2231 Vdd.n913 Vdd.t836 0.7285
R2232 Vdd.n281 Vdd.t585 0.7285
R2233 Vdd.n281 Vdd.t457 0.7285
R2234 Vdd.n951 Vdd.t431 0.7285
R2235 Vdd.n951 Vdd.t752 0.7285
R2236 Vdd.n738 Vdd.t149 0.7285
R2237 Vdd.n738 Vdd.t73 0.7285
R2238 Vdd.n666 Vdd.t375 0.7285
R2239 Vdd.n666 Vdd.t23 0.7285
R2240 Vdd.n777 Vdd.t27 0.7285
R2241 Vdd.n777 Vdd.t575 0.7285
R2242 Vdd.n392 Vdd.t449 0.7285
R2243 Vdd.n392 Vdd.t443 0.7285
R2244 Vdd.n815 Vdd.t213 0.7285
R2245 Vdd.n815 Vdd.t85 0.7285
R2246 Vdd.n362 Vdd.t407 0.7285
R2247 Vdd.n362 Vdd.t932 0.7285
R2248 Vdd.n853 Vdd.t551 0.7285
R2249 Vdd.n853 Vdd.t587 0.7285
R2250 Vdd.n326 Vdd.t411 0.7285
R2251 Vdd.n326 Vdd.t113 0.7285
R2252 Vdd.n892 Vdd.t441 0.7285
R2253 Vdd.n892 Vdd.t71 0.7285
R2254 Vdd.n296 Vdd.t403 0.7285
R2255 Vdd.n296 Vdd.t523 0.7285
R2256 Vdd.n930 Vdd.t177 0.7285
R2257 Vdd.n930 Vdd.t67 0.7285
R2258 Vdd.n266 Vdd.t453 0.7285
R2259 Vdd.n266 Vdd.t529 0.7285
R2260 Vdd.n686 Vdd.t824 0.7285
R2261 Vdd.n686 Vdd.t469 0.7285
R2262 Vdd.n412 Vdd.t944 0.7285
R2263 Vdd.n412 Vdd.t379 0.7285
R2264 Vdd.n382 Vdd.t31 0.7285
R2265 Vdd.n382 Vdd.t415 0.7285
R2266 Vdd.n352 Vdd.t335 0.7285
R2267 Vdd.n352 Vdd.t369 0.7285
R2268 Vdd.n316 Vdd.t812 0.7285
R2269 Vdd.n316 Vdd.t359 0.7285
R2270 Vdd.n286 Vdd.t137 0.7285
R2271 Vdd.n286 Vdd.t413 0.7285
R2272 Vdd.n691 Vdd.t828 0.7285
R2273 Vdd.n691 Vdd.t764 0.7285
R2274 Vdd.n707 Vdd.t579 0.7285
R2275 Vdd.n707 Vdd.t618 0.7285
R2276 Vdd.n702 Vdd.t938 0.7285
R2277 Vdd.n702 Vdd.t830 0.7285
R2278 Vdd.n725 Vdd.t762 0.7285
R2279 Vdd.n725 Vdd.t583 0.7285
R2280 Vdd.n731 Vdd.t720 0.7285
R2281 Vdd.n731 Vdd.t15 0.7285
R2282 Vdd.n719 Vdd.t11 0.7285
R2283 Vdd.n719 Vdd.t714 0.7285
R2284 Vdd.n624 Vdd.t738 0.7285
R2285 Vdd.n624 Vdd.t910 0.7285
R2286 Vdd.n635 Vdd.t231 0.7285
R2287 Vdd.n635 Vdd.t633 0.7285
R2288 Vdd.n630 Vdd.t892 0.7285
R2289 Vdd.n630 Vdd.t736 0.7285
R2290 Vdd.n647 Vdd.t908 0.7285
R2291 Vdd.n647 Vdd.t47 0.7285
R2292 Vdd.n641 Vdd.t729 0.7285
R2293 Vdd.n641 Vdd.t271 0.7285
R2294 Vdd.n654 Vdd.t141 0.7285
R2295 Vdd.n654 Vdd.t678 0.7285
R2296 Vdd.n555 Vdd.t347 0.7285
R2297 Vdd.n555 Vdd.t145 0.7285
R2298 Vdd.n566 Vdd.t51 0.7285
R2299 Vdd.n566 Vdd.t636 0.7285
R2300 Vdd.n561 Vdd.t35 0.7285
R2301 Vdd.n561 Vdd.t349 0.7285
R2302 Vdd.n578 Vdd.t143 0.7285
R2303 Vdd.n578 Vdd.t235 0.7285
R2304 Vdd.n572 Vdd.t630 0.7285
R2305 Vdd.n572 Vdd.t227 0.7285
R2306 Vdd.n585 Vdd.t157 0.7285
R2307 Vdd.n585 Vdd.t681 0.7285
R2308 Vdd.n775 SARlogic_0.dffrs_1.nand3_0.C 0.717607
R2309 Vdd.n813 SARlogic_0.dffrs_2.nand3_0.C 0.717607
R2310 Vdd.n851 SARlogic_0.dffrs_3.nand3_0.C 0.717607
R2311 Vdd.n890 SARlogic_0.dffrs_4.nand3_0.C 0.717607
R2312 Vdd.n928 SARlogic_0.dffrs_5.nand3_0.C 0.717607
R2313 Vdd.n700 SARlogic_0.dffrs_0.nand3_0.C 0.717607
R2314 Vdd.n1047 Vdd.n1045 0.667
R2315 Vdd.n1053 Vdd.n1051 0.662
R2316 Vdd.n1049 Vdd.n1047 0.643429
R2317 Vdd.n1051 Vdd.n1049 0.638429
R2318 Vdd.n1062 Vdd.n1061 0.58325
R2319 Vdd.n1043 Vdd.n1040 0.58325
R2320 Vdd.n176 Vdd.n167 0.561043
R2321 Vdd.n103 Vdd.n94 0.561043
R2322 Vdd.n107 Vdd.n33 0.561043
R2323 Vdd.n106 Vdd.n34 0.561043
R2324 Vdd.n92 Vdd.n35 0.561043
R2325 Vdd.n115 Vdd.n32 0.561043
R2326 Vdd.n180 Vdd.n17 0.561043
R2327 Vdd.n179 Vdd.n18 0.561043
R2328 Vdd.n165 Vdd.n19 0.561043
R2329 Vdd.n188 Vdd.n16 0.561043
R2330 Vdd.n241 Vdd.n232 0.561043
R2331 Vdd.n604 Vdd.n595 0.561043
R2332 Vdd.n535 Vdd.n526 0.561043
R2333 Vdd.n539 Vdd.n487 0.561043
R2334 Vdd.n538 Vdd.n488 0.561043
R2335 Vdd.n524 Vdd.n489 0.561043
R2336 Vdd.n547 Vdd.n486 0.561043
R2337 Vdd.n608 Vdd.n471 0.561043
R2338 Vdd.n607 Vdd.n472 0.561043
R2339 Vdd.n593 Vdd.n473 0.561043
R2340 Vdd.n616 Vdd.n470 0.561043
R2341 Vdd.n463 Vdd.n454 0.561043
R2342 Vdd.n449 Vdd.n436 0.561043
R2343 Vdd.n451 Vdd.n434 0.561043
R2344 Vdd.n452 Vdd.n424 0.561043
R2345 Vdd.n466 Vdd.n423 0.561043
R2346 Vdd.n248 Vdd.n214 0.561043
R2347 Vdd.n245 Vdd.n217 0.561043
R2348 Vdd.n244 Vdd.n218 0.561043
R2349 Vdd.n230 Vdd.n229 0.561043
R2350 Vdd.n118 Vdd.n116 0.490037
R2351 Vdd.n191 Vdd.n189 0.490037
R2352 Vdd.n550 Vdd.n548 0.490037
R2353 Vdd.n619 Vdd.n617 0.490037
R2354 Vdd.n256 Vdd.n254 0.490037
R2355 Vdd.n1045 Vdd.n1033 0.47525
R2356 Vdd.n1054 Vdd.n1053 0.47525
R2357 Vdd.n118 Vdd.n117 0.436534
R2358 Vdd.n191 Vdd.n190 0.436534
R2359 Vdd.n550 Vdd.n549 0.436534
R2360 Vdd.n619 Vdd.n618 0.436534
R2361 Vdd.n256 Vdd.n255 0.436534
R2362 Vdd.n448 Vdd.n440 0.415037
R2363 Vdd.n758 Vdd.n737 0.403945
R2364 Vdd.n439 Vdd.n438 0.3862
R2365 Vdd.n1067 Vdd.n1066 0.381816
R2366 Vdd.n1065 Vdd.n1062 0.34025
R2367 Vdd.n1061 Vdd.n1033 0.34025
R2368 Vdd.n1054 Vdd.n1043 0.34025
R2369 Vdd.n1071 Vdd.n1070 0.313132
R2370 Vdd.n1070 Vdd.n1069 0.289447
R2371 Vdd.n1069 Vdd.n1068 0.279974
R2372 Vdd.n1073 Vdd.n1072 0.265225
R2373 Vdd.n1068 Vdd.n1067 0.256289
R2374 Vdd.n176 Vdd.n175 0.255737
R2375 Vdd.n103 Vdd.n102 0.255737
R2376 Vdd.n116 Vdd.n115 0.255737
R2377 Vdd.n189 Vdd.n188 0.255737
R2378 Vdd.n241 Vdd.n240 0.255737
R2379 Vdd.n604 Vdd.n603 0.255737
R2380 Vdd.n535 Vdd.n534 0.255737
R2381 Vdd.n548 Vdd.n547 0.255737
R2382 Vdd.n617 Vdd.n616 0.255737
R2383 Vdd.n463 Vdd.n462 0.255737
R2384 Vdd.n449 Vdd.n448 0.255737
R2385 Vdd.n254 Vdd.n214 0.255737
R2386 Vdd.n258 Vdd.n202 0.236406
R2387 Vdd.n115 Vdd.n114 0.2165
R2388 Vdd.n188 Vdd.n187 0.2165
R2389 Vdd.n547 Vdd.n546 0.2165
R2390 Vdd.n616 Vdd.n615 0.2165
R2391 Vdd.n450 Vdd.n449 0.2165
R2392 Vdd.n246 Vdd.n214 0.2165
R2393 Vdd.n1019 comparator_no_offsetcal_0.x3.avdd 0.207699
R2394 Vdd.n1066 comparator_no_offsetcal_0.VDD 0.193526
R2395 Vdd.n974 Vdd.n973 0.165959
R2396 Vdd.n1072 Vdd 0.162037
R2397 Vdd.n114 Vdd.n107 0.148424
R2398 Vdd.n187 Vdd.n180 0.148424
R2399 Vdd.n546 Vdd.n539 0.148424
R2400 Vdd.n615 Vdd.n608 0.148424
R2401 Vdd.n451 Vdd.n450 0.148424
R2402 Vdd.n246 Vdd.n245 0.148424
R2403 adc_PISO_0.dffrs_3.resetb Vdd.n196 0.136036
R2404 adc_PISO_0.dffrs_5.resetb Vdd.n83 0.136036
R2405 adc_PISO_0.dffrs_4.resetb Vdd.n156 0.136036
R2406 adc_PISO_0.dffrs_2.resetb Vdd.n966 0.136036
R2407 SARlogic_0.dffrs_13.resetb Vdd.n718 0.136036
R2408 adc_PISO_0.dffrs_0.resetb Vdd.n421 0.136036
R2409 adc_PISO_0.dffrs_1.resetb Vdd.n335 0.136036
R2410 Vdd.n1028 Vdd.n1023 0.1355
R2411 Vdd.n440 Vdd.n439 0.124324
R2412 Vdd.n1026 Vdd.n1025 0.109786
R2413 Vdd.n1032 Vdd.n1021 0.103357
R2414 Vdd.n521 Vdd.n515 0.101647
R2415 Vdd.n1073 Vdd.n1007 0.0967961
R2416 Vdd.n1020 Vdd.n1019 0.0965492
R2417 Vdd.n973 Vdd.n972 0.0898578
R2418 Vdd.n975 Vdd.n259 0.0817571
R2419 Vdd.n522 Vdd.n521 0.0720596
R2420 Vdd.n1074 Vdd.n1073 0.0680047
R2421 Vdd.n874 Vdd.n336 0.0660636
R2422 Vdd.n177 Vdd.n176 0.0635
R2423 Vdd.n104 Vdd.n103 0.0635
R2424 Vdd.n242 Vdd.n241 0.0635
R2425 Vdd.n605 Vdd.n604 0.0635
R2426 Vdd.n536 Vdd.n535 0.0635
R2427 Vdd.n464 Vdd.n463 0.0635
R2428 Vdd.n257 Vdd.n213 0.0597785
R2429 Vdd.n515 Vdd.n509 0.0590321
R2430 Vdd.n1032 Vdd.n1031 0.0519286
R2431 Vdd.n1025 Vdd.n1021 0.0455
R2432 Vdd.n772 SARlogic_0.dffrs_1.nand3_2.C 0.0455
R2433 Vdd.n810 SARlogic_0.dffrs_2.nand3_2.C 0.0455
R2434 Vdd.n848 SARlogic_0.dffrs_3.nand3_2.C 0.0455
R2435 Vdd.n887 SARlogic_0.dffrs_4.nand3_2.C 0.0455
R2436 Vdd.n925 SARlogic_0.dffrs_5.nand3_2.C 0.0455
R2437 Vdd.n697 SARlogic_0.dffrs_0.nand3_2.C 0.0455
R2438 Vdd.n714 SARlogic_0.dffrs_13.nand3_7.A 0.0455
R2439 Vdd.n107 Vdd.n106 0.0452384
R2440 Vdd.n180 Vdd.n179 0.0452384
R2441 Vdd.n539 Vdd.n538 0.0452384
R2442 Vdd.n608 Vdd.n607 0.0452384
R2443 Vdd.n452 Vdd.n451 0.0452384
R2444 Vdd.n245 Vdd.n244 0.0452384
R2445 Vdd.n72 Vdd.n66 0.0405727
R2446 Vdd.n145 Vdd.n139 0.0405727
R2447 Vdd.n577 Vdd.n571 0.0405727
R2448 Vdd.n646 Vdd.n640 0.0405727
R2449 Vdd.n1099 Vdd.n1093 0.0405727
R2450 SARlogic_0.dffrs_1.nand3_0.C Vdd.n774 0.0374643
R2451 SARlogic_0.dffrs_2.nand3_0.C Vdd.n812 0.0374643
R2452 SARlogic_0.dffrs_3.nand3_0.C Vdd.n850 0.0374643
R2453 SARlogic_0.dffrs_4.nand3_0.C Vdd.n889 0.0374643
R2454 SARlogic_0.dffrs_5.nand3_0.C Vdd.n927 0.0374643
R2455 SARlogic_0.dffrs_0.nand3_0.C Vdd.n699 0.0374643
R2456 Vdd.n1005 Vdd.n999 0.0373206
R2457 Vdd.n590 Vdd.n336 0.0359182
R2458 Vdd.n660 Vdd.n659 0.0359182
R2459 Vdd.n1080 Vdd.n1074 0.0359182
R2460 Vdd.n730 Vdd.n724 0.0339767
R2461 Vdd.n49 adc_PISO_0.dffrs_5.setb 0.032
R2462 Vdd.n122 adc_PISO_0.dffrs_4.setb 0.032
R2463 Vdd.n503 adc_PISO_0.dffrs_2.setb 0.032
R2464 Vdd.n775 SARlogic_0.dffrs_1.setb 0.032
R2465 Vdd.n813 SARlogic_0.dffrs_2.setb 0.032
R2466 Vdd.n851 SARlogic_0.dffrs_3.setb 0.032
R2467 Vdd.n890 SARlogic_0.dffrs_4.setb 0.032
R2468 Vdd.n928 SARlogic_0.dffrs_5.setb 0.032
R2469 Vdd.n700 SARlogic_0.dffrs_0.setb 0.032
R2470 Vdd.n554 adc_PISO_0.dffrs_1.setb 0.032
R2471 Vdd.n623 adc_PISO_0.dffrs_0.setb 0.032
R2472 adc_PISO_0.dffrs_3.setb Vdd.n1101 0.032
R2473 Vdd.n737 Vdd.n712 0.0316083
R2474 Vdd.n175 Vdd.n173 0.0313054
R2475 Vdd.n175 Vdd.n174 0.0313054
R2476 Vdd.n102 Vdd.n100 0.0313054
R2477 Vdd.n102 Vdd.n101 0.0313054
R2478 Vdd.n116 Vdd.n30 0.0313054
R2479 Vdd.n116 Vdd.n31 0.0313054
R2480 Vdd.n189 Vdd.n14 0.0313054
R2481 Vdd.n189 Vdd.n15 0.0313054
R2482 Vdd.n240 Vdd.n238 0.0313054
R2483 Vdd.n240 Vdd.n239 0.0313054
R2484 Vdd.n603 Vdd.n601 0.0313054
R2485 Vdd.n603 Vdd.n602 0.0313054
R2486 Vdd.n534 Vdd.n532 0.0313054
R2487 Vdd.n534 Vdd.n533 0.0313054
R2488 Vdd.n548 Vdd.n484 0.0313054
R2489 Vdd.n548 Vdd.n485 0.0313054
R2490 Vdd.n617 Vdd.n468 0.0313054
R2491 Vdd.n617 Vdd.n469 0.0313054
R2492 Vdd.n462 Vdd.n460 0.0313054
R2493 Vdd.n462 Vdd.n461 0.0313054
R2494 Vdd.n448 Vdd.n446 0.0313054
R2495 Vdd.n448 Vdd.n447 0.0313054
R2496 Vdd.n254 Vdd.n252 0.0313054
R2497 Vdd.n254 Vdd.n253 0.0313054
R2498 Vdd.n105 Vdd.n92 0.0295407
R2499 Vdd.n178 Vdd.n165 0.0295407
R2500 Vdd.n537 Vdd.n524 0.0295407
R2501 Vdd.n606 Vdd.n593 0.0295407
R2502 Vdd.n466 Vdd.n465 0.0295407
R2503 Vdd.n243 Vdd.n230 0.0295407
R2504 Vdd.n90 Vdd.n78 0.0288636
R2505 Vdd.n163 Vdd.n151 0.0288636
R2506 Vdd.n653 Vdd.n652 0.0288636
R2507 Vdd.n1087 Vdd.n1081 0.0288636
R2508 Vdd.n584 Vdd.n583 0.0288455
R2509 Vdd.n993 Vdd.n982 0.0286958
R2510 Vdd.n972 Vdd.n260 0.0279312
R2511 Vdd.n1007 Vdd.n202 0.0273926
R2512 Vdd.n66 Vdd.n55 0.0237
R2513 Vdd.n139 Vdd.n128 0.0237
R2514 Vdd.n571 Vdd.n560 0.0237
R2515 Vdd.n640 Vdd.n629 0.0237
R2516 Vdd.n1100 Vdd.n1099 0.0237
R2517 Vdd.n1031 Vdd.n1023 0.0197857
R2518 Vdd.n712 Vdd.n701 0.0192652
R2519 Vdd.n106 Vdd.n105 0.0161977
R2520 Vdd.n179 Vdd.n178 0.0161977
R2521 Vdd.n538 Vdd.n537 0.0161977
R2522 Vdd.n607 Vdd.n606 0.0161977
R2523 Vdd.n465 Vdd.n452 0.0161977
R2524 Vdd.n244 Vdd.n243 0.0161977
R2525 Vdd.n92 Vdd.n91 0.0129273
R2526 Vdd.n165 Vdd.n164 0.0129273
R2527 Vdd.n524 Vdd.n523 0.0129273
R2528 Vdd.n593 Vdd.n592 0.0129273
R2529 Vdd.n467 Vdd.n466 0.0129273
R2530 Vdd.n230 Vdd.n13 0.0129273
R2531 Vdd.n440 adc_PISO_0.avdd 0.0128676
R2532 Vdd.n90 Vdd.n89 0.0122273
R2533 Vdd.n163 Vdd.n162 0.0122273
R2534 Vdd.n591 Vdd.n590 0.0122273
R2535 Vdd.n659 Vdd.n653 0.0122273
R2536 Vdd.n1081 Vdd.n1080 0.0122273
R2537 Vdd.n982 Vdd.n981 0.0113078
R2538 Vdd.n1040 Vdd.n1008 0.0068
R2539 Vdd.n1007 Vdd.n1006 0.00613636
R2540 Vdd.n929 Vdd.n923 0.00505026
R2541 Vdd.n891 Vdd.n885 0.00505026
R2542 Vdd.n852 Vdd.n846 0.00505026
R2543 Vdd.n814 Vdd.n808 0.00505026
R2544 Vdd.n1006 Vdd.n1005 0.00441736
R2545 Vdd.n950 Vdd.n929 0.00430496
R2546 Vdd.n912 Vdd.n891 0.00430496
R2547 Vdd.n873 Vdd.n852 0.00430496
R2548 Vdd.n835 Vdd.n814 0.00430496
R2549 Vdd.n797 Vdd.n776 0.00430496
R2550 Vdd.n1026 comparator_no_offsetcal_0.x4.VDD 0.00371429
R2551 SARlogic_0.dffrs_5.vdd Vdd.n950 0.00349428
R2552 SARlogic_0.dffrs_4.vdd Vdd.n912 0.00349428
R2553 SARlogic_0.dffrs_3.vdd Vdd.n873 0.00349428
R2554 SARlogic_0.dffrs_2.vdd Vdd.n835 0.00349428
R2555 SARlogic_0.dffrs_1.vdd Vdd.n797 0.00349428
R2556 SARlogic_0.dffrs_0.vdd Vdd.n758 0.00349428
R2557 Vdd.n770 Vdd.n769 0.00291569
R2558 Vdd.n737 Vdd.n736 0.00285324
R2559 Vdd.n522 Vdd.n260 0.00265596
R2560 Vdd.n776 Vdd.n770 0.00263457
R2561 Vdd.n961 SARlogic_0.dffrs_5.vdd 0.00236325
R2562 Vdd.n923 SARlogic_0.dffrs_4.vdd 0.00236325
R2563 Vdd.n846 SARlogic_0.dffrs_2.vdd 0.00236325
R2564 Vdd.n808 SARlogic_0.dffrs_1.vdd 0.00236325
R2565 Vdd.n769 SARlogic_0.dffrs_0.vdd 0.00236325
R2566 Vdd.n258 Vdd.n257 0.00228481
R2567 Vdd.n885 Vdd.n874 0.0014349
R2568 Vdd.n874 SARlogic_0.dffrs_3.vdd 0.00142836
R2569 Vdd.n974 Vdd.n961 0.0008465
R2570 Vdd.n78 Vdd.n72 0.000518182
R2571 Vdd.n151 Vdd.n145 0.000518182
R2572 Vdd.n583 Vdd.n577 0.000518182
R2573 Vdd.n591 Vdd.n584 0.000518182
R2574 Vdd.n652 Vdd.n646 0.000518182
R2575 Vdd.n1093 Vdd.n1087 0.000518182
R2576 Vdd.n999 Vdd.n993 0.000517689
R2577 Vdd.n736 Vdd.n730 0.000515182
R2578 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t6 41.0041
R2579 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t5 40.6313
R2580 SARlogic_0.dffrs_4.d.n1 SARlogic_0.dffrs_4.d.t4 27.3166
R2581 SARlogic_0.dffrs_4.d.n0 SARlogic_0.dffrs_4.d.t7 26.9438
R2582 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d 17.5382
R2583 SARlogic_0.dffrs_4.d.n3 SARlogic_0.dffrs_4.d.n2 14.0582
R2584 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.t1 10.0473
R2585 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.t0 6.51042
R2586 SARlogic_0.dffrs_4.d.n5 SARlogic_0.dffrs_4.d.n4 6.04952
R2587 SARlogic_0.dffrs_4.nand3_8.A SARlogic_0.dffrs_4.d.n0 5.7755
R2588 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_4.d.n1 5.13907
R2589 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n6 4.72925
R2590 SARlogic_0.dffrs_4.d SARlogic_0.dffrs_4.nand3_8.A 0.784786
R2591 SARlogic_0.dffrs_4.d.n6 SARlogic_0.dffrs_4.d.n5 0.732092
R2592 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t2 0.7285
R2593 SARlogic_0.dffrs_4.d.n4 SARlogic_0.dffrs_4.d.t3 0.7285
R2594 SARlogic_0.dffrs_3.nand3_2.Z SARlogic_0.dffrs_4.d.n3 0.166901
R2595 SARlogic_0.dffrs_4.d.n2 SARlogic_0.dffrs_3.nand3_7.C 0.0455
R2596 Vss.n1495 Vss.n1494 1.11127e+06
R2597 Vss.n1498 Vss.n1496 1.11127e+06
R2598 Vss.n1473 Vss.n1472 1.03768e+06
R2599 Vss.n1491 Vss.n1490 653018
R2600 Vss.n1489 Vss.n1488 533628
R2601 Vss.n1493 Vss.n1492 511643
R2602 Vss.n1700 Vss.n107 149958
R2603 Vss.n1473 Vss.n291 136500
R2604 Vss.n1490 Vss.n1489 106786
R2605 Vss.n1492 Vss.n1491 106786
R2606 Vss.n1552 Vss.n243 106554
R2607 Vss.n892 Vss.n891 50714
R2608 Vss.n1744 Vss.n117 50260.2
R2609 Vss.n1608 Vss.n190 47256
R2610 Vss.n1488 Vss.n1487 42535.5
R2611 Vss.n1617 Vss.n1616 41697.6
R2612 Vss.n1475 Vss.n280 32884
R2613 Vss.n688 Vss.n560 32356.2
R2614 Vss.n1616 Vss.n1615 26779.4
R2615 Vss.n1205 Vss.n1204 24208.9
R2616 Vss.n24 Vss.n16 22665.9
R2617 Vss.n623 Vss.n622 22665.9
R2618 Vss.t105 Vss.n108 18167.5
R2619 Vss.n329 Vss.n280 17319
R2620 Vss.n889 Vss.n877 17088.9
R2621 Vss.n1204 Vss.n371 16547
R2622 Vss.n688 Vss.n687 16547
R2623 Vss.n1496 Vss.n70 16020.5
R2624 Vss.n1502 Vss.n1496 16020.5
R2625 Vss.n624 Vss.n623 15733.7
R2626 Vss.n1870 Vss.n24 15733.7
R2627 Vss.n1182 Vss.n392 15356.8
R2628 Vss.n1487 Vss.n280 14805.6
R2629 Vss.n876 Vss.n875 13656.9
R2630 Vss.n1295 Vss.n1274 13507.5
R2631 Vss.n1259 Vss.n1258 13264.1
R2632 Vss.n393 Vss.n371 12982.5
R2633 Vss.n1323 Vss.n1310 11672.3
R2634 Vss.n1883 Vss.n13 11672.3
R2635 Vss.n1213 Vss.n1212 11670.6
R2636 Vss.n724 Vss.n721 11510.4
R2637 Vss.n1212 Vss.n368 11510.4
R2638 Vss.n1758 Vss.n1755 11510.4
R2639 Vss.n1753 Vss.n1752 11510.4
R2640 Vss.n1310 Vss.n1306 11510.4
R2641 Vss.n751 Vss.n13 11510.4
R2642 Vss.n890 Vss.n889 11510.4
R2643 Vss.n721 Vss.n720 11510.4
R2644 Vss.n1179 Vss.n397 10562.5
R2645 Vss.n1616 Vss.n190 10357.6
R2646 Vss.n1608 Vss.t256 10202.1
R2647 Vss.t222 Vss.n1553 9747.75
R2648 Vss.n1492 Vss.n275 9694.18
R2649 Vss.n272 Vss.n70 9694.18
R2650 Vss.n1492 Vss.n272 9687.98
R2651 Vss.n1502 Vss.n1501 9687.98
R2652 Vss.n876 Vss.n394 9486.49
R2653 Vss.n899 Vss.n533 9213.04
R2654 Vss.n758 Vss.n541 9213.04
R2655 Vss.n1343 Vss.n1342 8696.91
R2656 Vss.n1325 Vss.n1258 7467.21
R2657 Vss.n319 Vss.n290 7154.22
R2658 Vss.n591 Vss.n576 7143.16
R2659 Vss.n839 Vss.n838 7143.16
R2660 Vss.n875 Vss.n840 7143.16
R2661 Vss.n623 Vss.n540 7082.44
R2662 Vss.n532 Vss.n24 7082.44
R2663 Vss.n353 Vss.n352 6961.73
R2664 Vss.n1294 Vss.n1272 6961.73
R2665 Vss.n874 Vss.n391 6961.73
R2666 Vss.n836 Vss.n835 6961.73
R2667 Vss.n602 Vss.n601 6961.73
R2668 Vss.n663 Vss.n643 6925.27
R2669 Vss.n1323 Vss.n1322 6921.73
R2670 Vss.n1883 Vss.n14 6921.73
R2671 Vss.n740 Vss.n739 6921.73
R2672 Vss.n243 Vss.n242 6841.13
R2673 Vss.n1475 Vss.n279 6737.81
R2674 Vss.n1343 Vss.n121 6393.51
R2675 Vss.n1750 Vss.n1744 6375
R2676 Vss.n1488 Vss.n279 6373.63
R2677 Vss.n1609 Vss.n1608 6317.73
R2678 Vss.n797 Vss.n394 6190.48
R2679 Vss.n1213 Vss.n317 6190.48
R2680 Vss.n1412 Vss.n1257 6157.34
R2681 Vss.n1182 Vss.n1181 5894.95
R2682 Vss.n1784 Vss.n1783 5751.62
R2683 Vss.n1177 Vss.n399 5557.62
R2684 Vss.n469 Vss.n451 5557.62
R2685 Vss.n472 Vss.n471 5557.62
R2686 Vss.n1713 Vss.n101 5557.62
R2687 Vss.n1810 Vss.n83 5557.62
R2688 Vss.n1809 Vss.n85 5557.62
R2689 Vss.n1424 Vss.n60 5557.62
R2690 Vss.n1834 Vss.n61 5557.62
R2691 Vss.n1725 Vss.n1724 5557.62
R2692 Vss.n1402 Vss.n144 5557.62
R2693 Vss.n1038 Vss.n502 5557.62
R2694 Vss.n955 Vss.n395 5557.62
R2695 Vss.n665 Vss.n664 5557.62
R2696 Vss.n602 Vss.n589 5551.58
R2697 Vss.n835 Vss.n804 5551.58
R2698 Vss.n981 Vss.n502 5551.58
R2699 Vss.n1724 Vss.n145 5551.58
R2700 Vss.n1132 Vss.n472 5551.58
R2701 Vss.n1122 Vss.n61 5551.58
R2702 Vss.n471 Vss.n469 5551.58
R2703 Vss.n1332 Vss.n1272 5551.58
R2704 Vss.n353 Vss.n340 5551.58
R2705 Vss.n1192 Vss.n391 5551.58
R2706 Vss.n1713 Vss.n1712 5551.58
R2707 Vss.n1535 Vss.n85 5551.58
R2708 Vss.n1810 Vss.n1809 5551.58
R2709 Vss.n1834 Vss.n60 5551.58
R2710 Vss.n1725 Vss.n144 5551.58
R2711 Vss.n1038 Vss.n399 5551.58
R2712 Vss.n956 Vss.n955 5551.58
R2713 Vss.n665 Vss.n566 5551.58
R2714 Vss.n1213 Vss.n367 5418.32
R2715 Vss.n1323 Vss.n291 5416.67
R2716 Vss.n1883 Vss.n11 5416.67
R2717 Vss.n876 Vss.n392 5243.79
R2718 Vss.n1783 Vss.n1782 4925
R2719 Vss.n1581 Vss.n241 4797.83
R2720 Vss.n1783 Vss.n108 4745.41
R2721 Vss.n1179 Vss.n1178 4485.19
R2722 Vss.n974 Vss.n973 4456.62
R2723 Vss.n1401 Vss.n1400 4448.54
R2724 Vss.n720 Vss.n719 4366.67
R2725 Vss.n397 Vss.n372 4316.58
R2726 Vss.n575 Vss.n574 4273.71
R2727 Vss.n1181 Vss.n394 4229.5
R2728 Vss.n1259 Vss.n122 4107.2
R2729 Vss.n1553 Vss.n241 3983.8
R2730 Vss.n397 Vss.n393 3889.63
R2731 Vss.n1181 Vss.n1180 3784.25
R2732 Vss.n907 Vss.n906 3765.76
R2733 Vss.n764 Vss.n763 3765.76
R2734 Vss.n664 Vss.n575 3568.02
R2735 Vss.n1600 Vss.t304 3463.67
R2736 Vss.n1794 Vss.n100 3217.05
R2737 Vss.n1633 Vss.n1632 3214.99
R2738 Vss.n1751 Vss.n122 3201.53
R2739 Vss.n1751 Vss.n1750 3178.74
R2740 Vss.n1150 Vss.n1148 3157.03
R2741 Vss.n1162 Vss.n408 3157.03
R2742 Vss.n438 Vss.n407 3157.03
R2743 Vss.n1821 Vss.n73 3157.03
R2744 Vss.n1414 Vss.n75 3157.03
R2745 Vss.n1447 Vss.n1446 3157.03
R2746 Vss.n1847 Vss.n1846 3157.03
R2747 Vss.n1515 Vss.n252 3157.03
R2748 Vss.n1682 Vss.n226 3157.03
R2749 Vss.n510 Vss.n398 3157.03
R2750 Vss.n477 Vss.n419 3155.01
R2751 Vss.n1100 Vss.n1099 3155.01
R2752 Vss.n1163 Vss.n1162 3155.01
R2753 Vss.n1653 Vss.n1652 3155.01
R2754 Vss.n1821 Vss.n1820 3155.01
R2755 Vss.n1445 Vss.n252 3155.01
R2756 Vss.n1150 Vss.n48 3155.01
R2757 Vss.n1518 Vss.n1516 3155.01
R2758 Vss.n1684 Vss.n1683 3155.01
R2759 Vss.n1359 Vss.n226 3148.94
R2760 Vss.n1411 Vss.n1357 3122.83
R2761 Vss.n692 Vss.n690 2945.66
R2762 Vss.n366 Vss.n365 2944.88
R2763 Vss.n1297 Vss.n1296 2944.88
R2764 Vss.n837 Vss.n15 2944.88
R2765 Vss.n642 Vss.n641 2944.88
R2766 Vss.n1616 Vss.n1553 2850.36
R2767 Vss.n1617 Vss.n242 2846.85
R2768 Vss.n1499 Vss.n243 2814.38
R2769 Vss.n439 Vss.n385 2720.84
R2770 Vss.t222 Vss.n1562 2698.96
R2771 Vss.t304 Vss.n1562 2698.96
R2772 Vss.n366 Vss.n319 2677.48
R2773 Vss.n365 Vss.n318 2677.48
R2774 Vss.n1296 Vss.n1295 2677.48
R2775 Vss.n1324 Vss.n1297 2677.48
R2776 Vss.n838 Vss.n837 2677.48
R2777 Vss.n1882 Vss.n15 2677.48
R2778 Vss.n642 Vss.n576 2677.48
R2779 Vss.n641 Vss.n547 2677.48
R2780 Vss.n1777 Vss.n1776 2575.98
R2781 Vss.n1750 Vss.t254 2437.5
R2782 Vss.n352 Vss.n319 2353.3
R2783 Vss.n1295 Vss.n1294 2353.3
R2784 Vss.n875 Vss.n874 2353.3
R2785 Vss.n838 Vss.n836 2353.3
R2786 Vss.n601 Vss.n576 2353.3
R2787 Vss.n1411 Vss.n1259 2306.19
R2788 Vss.n1274 Vss.n121 2303.4
R2789 Vss.n1476 Vss.n1474 2267.8
R2790 Vss.n862 Vss.n370 2257.8
R2791 Vss.n625 Vss.n611 2257.8
R2792 Vss.n1871 Vss.n23 2257.8
R2793 Vss.n1412 Vss.n1411 2253.62
R2794 Vss.n1752 Vss.n108 2145.4
R2795 Vss.n330 Vss.n318 2028.48
R2796 Vss.n1326 Vss.n1324 2027.23
R2797 Vss.n1882 Vss.n1881 2027.23
R2798 Vss.n617 Vss.n547 2027.23
R2799 Vss.n1651 Vss.n236 1972.34
R2800 Vss.n1651 Vss.n1650 1972.34
R2801 Vss.n1685 Vss.n191 1972.34
R2802 Vss.n1641 Vss.n1640 1953.93
R2803 Vss.n1640 Vss.n1639 1953.93
R2804 Vss.t98 Vss.n1753 1950
R2805 Vss.n1213 Vss.n318 1891.48
R2806 Vss.n1324 Vss.n1323 1890.32
R2807 Vss.n1883 Vss.n1882 1890.32
R2808 Vss.n739 Vss.n547 1890.32
R2809 Vss.n451 Vss.n449 1883.67
R2810 Vss.n1413 Vss.n83 1883.67
R2811 Vss.n1491 Vss.n276 1883.67
R2812 Vss.n1424 Vss.n47 1883.67
R2813 Vss.n1178 Vss.n1177 1883.67
R2814 Vss.n1793 Vss.n101 1861.56
R2815 Vss.n385 Vss.n384 1775.77
R2816 Vss.n877 Vss.n876 1732.36
R2817 Vss.n1685 Vss.n190 1726.87
R2818 Vss.n862 Vss.n367 1659.81
R2819 Vss.n611 Vss.n11 1659.81
R2820 Vss.n877 Vss.n23 1659.81
R2821 Vss.t98 Vss.t105 1657.5
R2822 Vss.n1412 Vss.n1258 1579.08
R2823 Vss.n1260 Vss.n1258 1476.63
R2824 Vss.n1413 Vss.n1412 1450.15
R2825 Vss.n1472 Vss.n279 1392.86
R2826 Vss.n941 Vss.n398 1336.79
R2827 Vss.n438 Vss.n437 1336.79
R2828 Vss.n1848 Vss.n1847 1336.79
R2829 Vss.n1448 Vss.n1447 1336.79
R2830 Vss.n1415 Vss.n1414 1336.79
R2831 Vss.n1100 Vss.n483 1336.25
R2832 Vss.n477 Vss.n476 1336.25
R2833 Vss.n1684 Vss.n192 1336.25
R2834 Vss.n1652 Vss.n234 1336.25
R2835 Vss.n1795 Vss.n1794 1314.68
R2836 Vss.n1633 Vss.n1630 1314.15
R2837 Vss.n1600 Vss.n168 1303.34
R2838 Vss.n1566 Vss.n168 1223
R2839 Vss.n651 Vss.n575 1212.42
R2840 Vss.n1473 Vss.n290 1205.38
R2841 Vss.n313 Vss.n47 1201.62
R2842 Vss.n1203 Vss.n385 1200.6
R2843 Vss.n1752 Vss.n1751 1153.88
R2844 Vss.n449 Vss.n438 1095.12
R2845 Vss.n1794 Vss.n1793 1095.12
R2846 Vss.n1414 Vss.n1413 1095.12
R2847 Vss.n1847 Vss.n47 1095.12
R2848 Vss.n1178 Vss.n398 1095.12
R2849 Vss.n1115 Vss.n477 1094.63
R2850 Vss.n1102 Vss.n1100 1094.63
R2851 Vss.n1640 Vss.n1633 1094.63
R2852 Vss.n1652 Vss.n1651 1094.63
R2853 Vss.n1685 Vss.n1684 1094.63
R2854 Vss.n642 Vss.n546 1086.49
R2855 Vss.n1474 Vss.n1473 1062.42
R2856 Vss.n1413 Vss.n1256 1055.77
R2857 Vss.n739 Vss.n546 1048.57
R2858 Vss.n1181 Vss.n393 996.898
R2859 Vss.n1411 Vss.n1401 933.769
R2860 Vss.n1700 Vss.n169 928.572
R2861 Vss.n1016 Vss.n974 927.706
R2862 Vss.n664 Vss.n663 897.806
R2863 Vss.n1499 Vss.n1498 885.807
R2864 Vss.n1205 Vss.n369 873.918
R2865 Vss.n719 Vss.n713 873.918
R2866 Vss.n1777 Vss.t554 857.144
R2867 Vss.n1781 Vss.t554 857.144
R2868 Vss.t65 Vss.n30 849.126
R2869 Vss.n775 Vss.t130 849.126
R2870 Vss.t254 Vss.n1745 847.827
R2871 Vss.n1755 Vss.t98 847.827
R2872 Vss.n1776 Vss.t105 847.827
R2873 Vss.n1322 Vss.t559 847.827
R2874 Vss.t559 Vss.n1257 847.827
R2875 Vss.t561 Vss.n14 847.827
R2876 Vss.n533 Vss.t561 847.827
R2877 Vss.t149 Vss.n907 847.827
R2878 Vss.n916 Vss.t149 847.827
R2879 Vss.n915 Vss.t111 847.827
R2880 Vss.n912 Vss.t111 847.827
R2881 Vss.n911 Vss.t65 847.827
R2882 Vss.n740 Vss.t446 847.827
R2883 Vss.t446 Vss.n541 847.827
R2884 Vss.n764 Vss.t200 847.827
R2885 Vss.n767 Vss.t200 847.827
R2886 Vss.t238 Vss.n768 847.827
R2887 Vss.n773 Vss.t238 847.827
R2888 Vss.t130 Vss.n774 847.827
R2889 Vss.n994 Vss.n502 832.22
R2890 Vss.n420 Vss.n61 832.22
R2891 Vss.n1090 Vss.n472 832.22
R2892 Vss.n469 Vss.n458 832.22
R2893 Vss.n353 Vss.n341 832.22
R2894 Vss.n1714 Vss.n1713 832.22
R2895 Vss.n1283 Vss.n1272 832.22
R2896 Vss.n1661 Vss.n85 832.22
R2897 Vss.n1811 Vss.n1810 832.22
R2898 Vss.n60 Vss.n59 832.22
R2899 Vss.n1724 Vss.n146 832.22
R2900 Vss.n1360 Vss.n144 832.22
R2901 Vss.n931 Vss.n399 832.22
R2902 Vss.n852 Vss.n391 832.22
R2903 Vss.n955 Vss.n953 832.22
R2904 Vss.n835 Vss.n805 832.22
R2905 Vss.n602 Vss.n590 832.22
R2906 Vss.n665 Vss.n573 832.22
R2907 Vss.n502 Vss.n501 832.101
R2908 Vss.n425 Vss.n61 832.101
R2909 Vss.n491 Vss.n472 832.101
R2910 Vss.n469 Vss.n468 832.101
R2911 Vss.n354 Vss.n353 832.101
R2912 Vss.n1713 Vss.n155 832.101
R2913 Vss.n1272 Vss.n1271 832.101
R2914 Vss.n1668 Vss.n85 832.101
R2915 Vss.n1810 Vss.n84 832.101
R2916 Vss.n1427 Vss.n60 832.101
R2917 Vss.n1724 Vss.n1723 832.101
R2918 Vss.n1389 Vss.n144 832.101
R2919 Vss.n406 Vss.n399 832.101
R2920 Vss.n861 Vss.n391 832.101
R2921 Vss.n955 Vss.n954 832.101
R2922 Vss.n835 Vss.n834 832.101
R2923 Vss.n603 Vss.n602 832.101
R2924 Vss.n666 Vss.n665 832.101
R2925 Vss.n1178 Vss.n385 829.364
R2926 Vss.n1501 Vss.n1500 814.398
R2927 Vss.n272 Vss.n271 814.398
R2928 Vss.n1260 Vss.t544 812.5
R2929 Vss.n1357 Vss.t214 812.5
R2930 Vss.n899 Vss.t422 812.5
R2931 Vss.n758 Vss.t369 812.5
R2932 Vss.n1486 Vss.n281 798.088
R2933 Vss.n689 Vss.n688 767.827
R2934 Vss.n1753 Vss.n120 755.625
R2935 Vss.n282 Vss.n47 750.922
R2936 Vss.n1476 Vss.n1475 748.735
R2937 Vss.t98 Vss.t105 720.653
R2938 Vss.n916 Vss.n915 720.653
R2939 Vss.n912 Vss.n911 720.653
R2940 Vss.n768 Vss.n767 720.653
R2941 Vss.n774 Vss.n773 720.653
R2942 Vss.n1618 Vss.n1617 702.332
R2943 Vss.n1447 Vss.n276 698.639
R2944 Vss.n340 Vss.n339 693.082
R2945 Vss.n627 Vss.n589 692.747
R2946 Vss.n1333 Vss.n1332 692.747
R2947 Vss.n804 Vss.n803 692.747
R2948 Vss.n1615 Vss.t344 676.471
R2949 Vss.n1562 Vss.t344 676.471
R2950 Vss.n1562 Vss.t162 676.471
R2951 Vss.n1609 Vss.t162 676.471
R2952 Vss.n384 Vss.t137 670.104
R2953 Vss.t137 Vss.n383 670.104
R2954 Vss.n380 Vss.t449 670.104
R2955 Vss.n377 Vss.t449 670.104
R2956 Vss.n376 Vss.t646 670.104
R2957 Vss.t646 Vss.n369 670.104
R2958 Vss.n690 Vss.t644 670.104
R2959 Vss.n704 Vss.t644 670.104
R2960 Vss.n705 Vss.t301 670.104
R2961 Vss.n709 Vss.t301 670.104
R2962 Vss.t401 Vss.n712 670.104
R2963 Vss.n713 Vss.t401 670.104
R2964 Vss.n1205 Vss.n370 665.564
R2965 Vss.n625 Vss.n624 665.564
R2966 Vss.n1871 Vss.n1870 665.564
R2967 Vss.n1494 Vss.n272 662.646
R2968 Vss.n340 Vss.n338 662.074
R2969 Vss.n1332 Vss.n1331 661.665
R2970 Vss.n804 Vss.n802 661.665
R2971 Vss.n621 Vss.n589 661.665
R2972 Vss.t544 Vss.t523 650
R2973 Vss.t523 Vss.t214 650
R2974 Vss.t467 Vss.t140 650
R2975 Vss.t497 Vss.t144 650
R2976 Vss.t674 Vss.n1203 642.183
R2977 Vss.t603 Vss.n689 642.183
R2978 Vss.n693 Vss.t38 642.183
R2979 Vss.n1782 Vss.n1781 607.144
R2980 Vss.n840 Vss.n367 597.985
R2981 Vss.n591 Vss.n11 597.985
R2982 Vss.n877 Vss.n839 597.985
R2983 Vss.n1342 Vss.n122 596.029
R2984 Vss.n1749 Vss.t563 590.91
R2985 Vss.t254 Vss.n1749 590.91
R2986 Vss.t607 Vss.n1206 590.909
R2987 Vss.n1210 Vss.t607 590.909
R2988 Vss.t550 Vss.n1210 590.909
R2989 Vss.n1212 Vss.t558 590.909
R2990 Vss.n1212 Vss.t210 590.909
R2991 Vss.n1214 Vss.t212 590.909
R2992 Vss.n1471 Vss.t337 590.909
R2993 Vss.n1309 Vss.t337 590.909
R2994 Vss.t445 Vss.n1309 590.909
R2995 Vss.n1310 Vss.t557 590.909
R2996 Vss.t27 Vss.n1310 590.909
R2997 Vss.n1318 Vss.t25 590.909
R2998 Vss.n616 Vss.t605 590.909
R2999 Vss.t605 Vss.n615 590.909
R3000 Vss.n615 Vss.t551 590.909
R3001 Vss.t564 Vss.n13 590.909
R3002 Vss.n13 Vss.t198 590.909
R3003 Vss.n1884 Vss.t186 590.909
R3004 Vss.n1869 Vss.t20 590.909
R3005 Vss.n880 Vss.t20 590.909
R3006 Vss.t556 Vss.n880 590.909
R3007 Vss.n889 Vss.t444 590.909
R3008 Vss.n889 Vss.t281 590.909
R3009 Vss.t285 Vss.n888 590.909
R3010 Vss.n718 Vss.t580 590.909
R3011 Vss.t580 Vss.n717 590.909
R3012 Vss.n717 Vss.t441 590.909
R3013 Vss.n721 Vss.t549 590.909
R3014 Vss.n721 Vss.t388 590.909
R3015 Vss.n738 Vss.t392 590.909
R3016 Vss.n1147 Vss.t311 582.165
R3017 Vss.n420 Vss.t506 582.165
R3018 Vss.n1091 Vss.t613 582.165
R3019 Vss.t485 Vss.n1090 582.165
R3020 Vss.n452 Vss.t535 582.165
R3021 Vss.n458 Vss.t307 582.165
R3022 Vss.n364 Vss.t22 582.165
R3023 Vss.n341 Vss.t461 582.165
R3024 Vss.n1715 Vss.t672 582.165
R3025 Vss.t317 Vss.n1714 582.165
R3026 Vss.t637 Vss.n1273 582.165
R3027 Vss.n1283 Vss.t473 582.165
R3028 Vss.n1662 Vss.t379 582.165
R3029 Vss.t457 Vss.n1661 582.165
R3030 Vss.n1812 Vss.t414 582.165
R3031 Vss.t151 Vss.n1811 582.165
R3032 Vss.n1426 Vss.t188 582.165
R3033 Vss.t375 Vss.n273 582.165
R3034 Vss.n1845 Vss.t57 582.165
R3035 Vss.n59 Vss.t631 582.165
R3036 Vss.n1514 Vss.t628 582.165
R3037 Vss.n1497 Vss.t487 582.165
R3038 Vss.n1681 Vss.t153 582.165
R3039 Vss.t493 Vss.n146 582.165
R3040 Vss.n1399 Vss.t157 582.165
R3041 Vss.n1360 Vss.t668 582.165
R3042 Vss.n932 Vss.t94 582.165
R3043 Vss.t246 Vss.n931 582.165
R3044 Vss.n1015 Vss.t329 582.165
R3045 Vss.n994 Vss.t489 582.165
R3046 Vss.t394 Vss.n851 582.165
R3047 Vss.n852 Vss.t463 582.165
R3048 Vss.n799 Vss.t385 582.165
R3049 Vss.n953 Vss.t327 582.165
R3050 Vss.n816 Vss.t395 582.165
R3051 Vss.t491 Vss.n805 582.165
R3052 Vss.n640 Vss.t660 582.165
R3053 Vss.n590 Vss.t498 582.165
R3054 Vss.n651 Vss.t374 582.165
R3055 Vss.t514 Vss.n573 582.165
R3056 Vss.n627 Vss.t589 581.712
R3057 Vss.t528 Vss.n626 581.712
R3058 Vss.t662 Vss.n396 581.712
R3059 Vss.n941 Vss.t325 581.712
R3060 Vss.n1176 Vss.t430 581.712
R3061 Vss.n437 Vss.t614 581.712
R3062 Vss.n1153 Vss.t8 581.712
R3063 Vss.t90 Vss.n1152 581.712
R3064 Vss.n1080 Vss.t40 581.712
R3065 Vss.t455 Vss.n417 581.712
R3066 Vss.t134 Vss.n499 581.712
R3067 Vss.n1028 Vss.t427 581.712
R3068 Vss.n983 Vss.t136 581.712
R3069 Vss.t536 Vss.n483 581.712
R3070 Vss.t538 Vss.n500 581.712
R3071 Vss.n1001 Vss.t481 581.712
R3072 Vss.n501 Vss.t49 581.712
R3073 Vss.n1098 Vss.t386 581.712
R3074 Vss.n1123 Vss.t418 581.712
R3075 Vss.t332 Vss.n250 581.712
R3076 Vss.n1131 Vss.t334 581.712
R3077 Vss.n476 Vss.t598 581.712
R3078 Vss.n425 Vss.t51 581.712
R3079 Vss.t147 Vss.n251 581.712
R3080 Vss.n491 Vss.t431 581.712
R3081 Vss.t69 Vss.n490 581.712
R3082 Vss.n468 Vss.t202 581.712
R3083 Vss.n460 Vss.t75 581.712
R3084 Vss.n450 Vss.t88 581.712
R3085 Vss.n1848 Vss.t309 581.712
R3086 Vss.t659 Vss.n1425 581.712
R3087 Vss.n1448 Vss.t95 581.712
R3088 Vss.n1293 Vss.t524 581.712
R3089 Vss.n1275 Vss.t520 581.712
R3090 Vss.n354 Vss.t440 581.712
R3091 Vss.t279 Vss.n289 581.712
R3092 Vss.n351 Vss.t275 581.712
R3093 Vss.n342 Vss.t511 581.712
R3094 Vss.n339 Vss.t117 581.712
R3095 Vss.n1477 Vss.t277 581.712
R3096 Vss.t609 Vss.n1193 581.712
R3097 Vss.n1194 Vss.t586 581.712
R3098 Vss.n139 Vss.t158 581.712
R3099 Vss.t372 Vss.n123 581.712
R3100 Vss.n1796 Vss.t44 581.712
R3101 Vss.t477 Vss.n1795 581.712
R3102 Vss.n1626 Vss.t119 581.712
R3103 Vss.n1630 Vss.t41 581.712
R3104 Vss.n1711 Vss.t548 581.712
R3105 Vss.n170 Vss.t601 581.712
R3106 Vss.n180 Vss.t597 581.712
R3107 Vss.t362 Vss.n171 581.712
R3108 Vss.t438 Vss.n155 581.712
R3109 Vss.n1699 Vss.t227 581.712
R3110 Vss.n1271 Vss.t36 581.712
R3111 Vss.n1344 Vss.t420 581.712
R3112 Vss.n1333 Vss.t649 581.712
R3113 Vss.n1341 Vss.t525 581.712
R3114 Vss.n1370 Vss.t625 581.712
R3115 Vss.t154 Vss.n1358 581.712
R3116 Vss.t29 Vss.n274 581.712
R3117 Vss.n1415 Vss.t377 581.712
R3118 Vss.t160 Vss.n87 581.712
R3119 Vss.n216 Vss.t626 581.712
R3120 Vss.t219 Vss.n88 581.712
R3121 Vss.n222 Vss.t500 581.712
R3122 Vss.n1824 Vss.t252 581.712
R3123 Vss.t31 Vss.n1823 581.712
R3124 Vss.n1503 Vss.t381 581.712
R3125 Vss.t518 Vss.n71 581.712
R3126 Vss.n1536 Vss.t146 581.712
R3127 Vss.t217 Vss.n192 581.712
R3128 Vss.n1500 Vss.t433 581.712
R3129 Vss.n1654 Vss.t339 581.712
R3130 Vss.n1543 Vss.t165 581.712
R3131 Vss.t382 Vss.n234 581.712
R3132 Vss.n1668 Vss.t48 581.712
R3133 Vss.t321 Vss.n193 581.712
R3134 Vss.t640 Vss.n84 581.712
R3135 Vss.n1379 Vss.t323 581.712
R3136 Vss.n271 Vss.t230 581.712
R3137 Vss.n1819 Vss.t260 581.712
R3138 Vss.n1427 Vss.t453 581.712
R3139 Vss.n1444 Vss.t225 581.712
R3140 Vss.n1832 Vss.t127 581.712
R3141 Vss.n1060 Vss.t657 581.712
R3142 Vss.t331 Vss.n63 581.712
R3143 Vss.n1068 Vss.t479 581.712
R3144 Vss.n1723 Vss.t54 581.712
R3145 Vss.n1631 Vss.t451 581.712
R3146 Vss.n1389 Vss.t616 581.712
R3147 Vss.t55 Vss.n125 581.712
R3148 Vss.n1738 Vss.t371 581.712
R3149 Vss.t670 Vss.n126 581.712
R3150 Vss.t380 Vss.n406 581.712
R3151 Vss.n1164 Vss.t346 581.712
R3152 Vss.n522 Vss.t545 581.712
R3153 Vss.t663 Vss.n509 581.712
R3154 Vss.n873 Vss.t417 581.712
R3155 Vss.n841 Vss.t516 581.712
R3156 Vss.t35 Vss.n861 581.712
R3157 Vss.n863 Vss.t266 581.712
R3158 Vss.n954 Vss.t108 581.712
R3159 Vss.n972 Vss.t67 581.712
R3160 Vss.n801 Vss.t622 581.712
R3161 Vss.t483 Vss.n800 581.712
R3162 Vss.n834 Vss.t184 581.712
R3163 Vss.n806 Vss.t576 581.712
R3164 Vss.n603 Vss.t629 581.712
R3165 Vss.n610 Vss.t578 581.712
R3166 Vss.n600 Vss.t530 581.712
R3167 Vss.n592 Vss.t495 581.712
R3168 Vss.n678 Vss.t259 581.712
R3169 Vss.t123 Vss.n677 581.712
R3170 Vss.n803 Vss.t120 581.712
R3171 Vss.n1872 Vss.t620 581.712
R3172 Vss.t37 Vss.n666 581.712
R3173 Vss.n667 Vss.t92 581.712
R3174 Vss.n662 Vss.t604 581.712
R3175 Vss.n644 Vss.t503 581.712
R3176 Vss.n383 Vss.n380 569.588
R3177 Vss.n377 Vss.n376 569.588
R3178 Vss.n705 Vss.n704 569.588
R3179 Vss.n712 Vss.n709 569.588
R3180 Vss.n1751 Vss.n121 565.155
R3181 Vss.t140 Vss.n532 561.686
R3182 Vss.t144 Vss.n540 561.686
R3183 Vss.n1177 Vss.n1176 548.236
R3184 Vss.n451 Vss.n450 548.236
R3185 Vss.n1425 Vss.n1424 548.236
R3186 Vss.n180 Vss.n101 548.236
R3187 Vss.n1370 Vss.n83 548.236
R3188 Vss.n1123 Vss.n1122 548.058
R3189 Vss.n1132 Vss.n1131 548.058
R3190 Vss.n1193 Vss.n1192 548.058
R3191 Vss.n1626 Vss.n145 548.058
R3192 Vss.n1712 Vss.n1711 548.058
R3193 Vss.n1536 Vss.n1535 548.058
R3194 Vss.n678 Vss.n566 548.058
R3195 Vss.t633 Vss.t460 513.746
R3196 Vss.t460 Vss.t674 513.746
R3197 Vss.t505 Vss.t603 513.746
R3198 Vss.t38 Vss.t505 513.746
R3199 Vss.t558 Vss.t550 502.274
R3200 Vss.t210 Vss.t212 502.274
R3201 Vss.t563 Vss.t448 502.274
R3202 Vss.t557 Vss.t445 502.274
R3203 Vss.t25 Vss.t27 502.274
R3204 Vss.t551 Vss.t564 502.274
R3205 Vss.t198 Vss.t186 502.274
R3206 Vss.t444 Vss.t556 502.274
R3207 Vss.t281 Vss.t285 502.274
R3208 Vss.t441 Vss.t549 502.274
R3209 Vss.t388 Vss.t392 502.274
R3210 Vss.n1122 Vss.n1121 484.702
R3211 Vss.n1133 Vss.n1132 484.702
R3212 Vss.n1192 Vss.n1191 484.702
R3213 Vss.n1712 Vss.n156 484.702
R3214 Vss.n1535 Vss.n1534 484.702
R3215 Vss.n1687 Vss.n145 484.702
R3216 Vss.n686 Vss.n566 484.702
R3217 Vss.t330 Vss.t311 465.733
R3218 Vss.t506 Vss.t330 465.733
R3219 Vss.t613 Vss.t600 465.733
R3220 Vss.t600 Vss.t485 465.733
R3221 Vss.t535 Vss.t89 465.733
R3222 Vss.t89 Vss.t307 465.733
R3223 Vss.t276 Vss.t22 465.733
R3224 Vss.t461 Vss.t276 465.733
R3225 Vss.t672 Vss.t596 465.733
R3226 Vss.t596 Vss.t317 465.733
R3227 Vss.t527 Vss.t637 465.733
R3228 Vss.t473 Vss.t527 465.733
R3229 Vss.t379 Vss.t220 465.733
R3230 Vss.t220 Vss.t457 465.733
R3231 Vss.t414 Vss.t624 465.733
R3232 Vss.t624 Vss.t151 465.733
R3233 Vss.t188 Vss.t30 465.733
R3234 Vss.t30 Vss.t375 465.733
R3235 Vss.t656 Vss.t57 465.733
R3236 Vss.t631 Vss.t656 465.733
R3237 Vss.t384 Vss.t628 465.733
R3238 Vss.t487 Vss.t384 465.733
R3239 Vss.t153 Vss.t43 465.733
R3240 Vss.t43 Vss.t493 465.733
R3241 Vss.t370 Vss.t157 465.733
R3242 Vss.t668 Vss.t370 465.733
R3243 Vss.t94 Vss.t429 465.733
R3244 Vss.t429 Vss.t246 465.733
R3245 Vss.t539 Vss.t329 465.733
R3246 Vss.t489 Vss.t539 465.733
R3247 Vss.t588 Vss.t394 465.733
R3248 Vss.t463 Vss.t588 465.733
R3249 Vss.t385 Vss.t661 465.733
R3250 Vss.t661 Vss.t327 465.733
R3251 Vss.t395 Vss.t623 465.733
R3252 Vss.t623 Vss.t491 465.733
R3253 Vss.t531 Vss.t660 465.733
R3254 Vss.t498 Vss.t531 465.733
R3255 Vss.t374 Vss.t122 465.733
R3256 Vss.t122 Vss.t514 465.733
R3257 Vss.t589 Vss.t245 465.37
R3258 Vss.t245 Vss.t528 465.37
R3259 Vss.t546 Vss.t662 465.37
R3260 Vss.t325 Vss.t546 465.37
R3261 Vss.t135 Vss.t430 465.37
R3262 Vss.t614 Vss.t135 465.37
R3263 Vss.t8 Vss.t203 465.37
R3264 Vss.t203 Vss.t90 465.37
R3265 Vss.t40 Vss.t335 465.37
R3266 Vss.t335 Vss.t455 465.37
R3267 Vss.t406 Vss.t134 465.37
R3268 Vss.t427 Vss.t406 465.37
R3269 Vss.t136 Vss.t52 465.37
R3270 Vss.t52 Vss.t536 465.37
R3271 Vss.t118 Vss.t538 465.37
R3272 Vss.t481 Vss.t118 465.37
R3273 Vss.t49 Vss.t365 465.37
R3274 Vss.t365 Vss.t386 465.37
R3275 Vss.t418 Vss.t439 465.37
R3276 Vss.t439 Vss.t332 465.37
R3277 Vss.t437 Vss.t334 465.37
R3278 Vss.t598 Vss.t437 465.37
R3279 Vss.t51 Vss.t357 465.37
R3280 Vss.t357 Vss.t147 465.37
R3281 Vss.t431 Vss.t291 465.37
R3282 Vss.t291 Vss.t69 465.37
R3283 Vss.t358 Vss.t202 465.37
R3284 Vss.t75 Vss.t358 465.37
R3285 Vss.t88 Vss.t9 465.37
R3286 Vss.t9 Vss.t309 465.37
R3287 Vss.t126 Vss.t659 465.37
R3288 Vss.t95 Vss.t126 465.37
R3289 Vss.t648 Vss.t524 465.37
R3290 Vss.t520 Vss.t648 465.37
R3291 Vss.t440 Vss.t469 465.37
R3292 Vss.t469 Vss.t279 465.37
R3293 Vss.t216 Vss.t275 465.37
R3294 Vss.t511 Vss.t216 465.37
R3295 Vss.t117 Vss.t242 465.37
R3296 Vss.t242 Vss.t277 465.37
R3297 Vss.t185 Vss.t609 465.37
R3298 Vss.t586 Vss.t185 465.37
R3299 Vss.t158 Vss.t174 465.37
R3300 Vss.t174 Vss.t372 465.37
R3301 Vss.t44 Vss.t573 465.37
R3302 Vss.t573 Vss.t477 465.37
R3303 Vss.t119 Vss.t434 465.37
R3304 Vss.t434 Vss.t41 465.37
R3305 Vss.t432 Vss.t548 465.37
R3306 Vss.t601 Vss.t432 465.37
R3307 Vss.t597 Vss.t547 465.37
R3308 Vss.t547 Vss.t362 465.37
R3309 Vss.t522 Vss.t438 465.37
R3310 Vss.t227 Vss.t522 465.37
R3311 Vss.t36 Vss.t466 465.37
R3312 Vss.t466 Vss.t420 465.37
R3313 Vss.t649 Vss.t244 465.37
R3314 Vss.t244 Vss.t525 465.37
R3315 Vss.t625 Vss.t161 465.37
R3316 Vss.t161 Vss.t154 465.37
R3317 Vss.t253 Vss.t29 465.37
R3318 Vss.t377 Vss.t253 465.37
R3319 Vss.t639 Vss.t160 465.37
R3320 Vss.t626 Vss.t639 465.37
R3321 Vss.t13 Vss.t219 465.37
R3322 Vss.t500 Vss.t13 465.37
R3323 Vss.t252 Vss.t232 465.37
R3324 Vss.t232 Vss.t31 465.37
R3325 Vss.t381 Vss.t164 465.37
R3326 Vss.t164 Vss.t518 465.37
R3327 Vss.t146 Vss.t50 465.37
R3328 Vss.t50 Vss.t217 465.37
R3329 Vss.t433 Vss.t312 465.37
R3330 Vss.t312 Vss.t339 465.37
R3331 Vss.t165 Vss.t53 465.37
R3332 Vss.t53 Vss.t382 465.37
R3333 Vss.t48 Vss.t316 465.37
R3334 Vss.t316 Vss.t321 465.37
R3335 Vss.t295 Vss.t640 465.37
R3336 Vss.t323 Vss.t295 465.37
R3337 Vss.t230 Vss.t290 465.37
R3338 Vss.t290 Vss.t260 465.37
R3339 Vss.t453 Vss.t313 465.37
R3340 Vss.t313 Vss.t225 465.37
R3341 Vss.t454 Vss.t127 465.37
R3342 Vss.t657 Vss.t454 465.37
R3343 Vss.t419 Vss.t331 465.37
R3344 Vss.t479 Vss.t419 465.37
R3345 Vss.t296 Vss.t54 465.37
R3346 Vss.t451 Vss.t296 465.37
R3347 Vss.t616 Vss.t361 465.37
R3348 Vss.t361 Vss.t55 465.37
R3349 Vss.t371 Vss.t159 465.37
R3350 Vss.t159 Vss.t670 465.37
R3351 Vss.t348 Vss.t380 465.37
R3352 Vss.t346 Vss.t348 465.37
R3353 Vss.t545 Vss.t101 465.37
R3354 Vss.t101 Vss.t663 465.37
R3355 Vss.t610 Vss.t417 465.37
R3356 Vss.t516 Vss.t610 465.37
R3357 Vss.t470 Vss.t35 465.37
R3358 Vss.t266 Vss.t470 465.37
R3359 Vss.t108 Vss.t366 465.37
R3360 Vss.t366 Vss.t67 465.37
R3361 Vss.t622 Vss.t121 465.37
R3362 Vss.t121 Vss.t483 465.37
R3363 Vss.t475 Vss.t184 465.37
R3364 Vss.t576 Vss.t475 465.37
R3365 Vss.t629 Vss.t508 465.37
R3366 Vss.t508 Vss.t578 465.37
R3367 Vss.t590 Vss.t530 465.37
R3368 Vss.t495 Vss.t590 465.37
R3369 Vss.t259 Vss.t243 465.37
R3370 Vss.t243 Vss.t123 465.37
R3371 Vss.t120 Vss.t630 465.37
R3372 Vss.t630 Vss.t620 465.37
R3373 Vss.t513 Vss.t37 465.37
R3374 Vss.t92 Vss.t513 465.37
R3375 Vss.t258 Vss.t604 465.37
R3376 Vss.t503 Vss.t258 465.37
R3377 Vss.n338 Vss.t208 462.849
R3378 Vss.n1331 Vss.t23 462.562
R3379 Vss.n802 Vss.t196 462.562
R3380 Vss.t390 Vss.n621 462.562
R3381 Vss.n1103 Vss.n1102 443.358
R3382 Vss.n1102 Vss.n482 443.358
R3383 Vss.n1115 Vss.n1113 443.358
R3384 Vss.n1115 Vss.n1114 443.358
R3385 Vss.n1162 Vss.n1161 435.214
R3386 Vss.n1821 Vss.n74 435.214
R3387 Vss.n1150 Vss.n1149 435.214
R3388 Vss.n265 Vss.n252 435.214
R3389 Vss.n226 Vss.n225 435.012
R3390 Vss.n1594 Vss.n1565 414.478
R3391 Vss.n1162 Vss.n409 404.991
R3392 Vss.n1822 Vss.n1821 404.991
R3393 Vss.n1151 Vss.n1150 404.991
R3394 Vss.n1069 Vss.n252 404.991
R3395 Vss.n226 Vss.n224 404.803
R3396 Vss.n1204 Vss.n372 402.062
R3397 Vss.t569 Vss.t567 384.214
R3398 Vss.n757 Vss.n749 383.418
R3399 Vss.n757 Vss.n756 383.418
R3400 Vss.n898 Vss.n788 383.418
R3401 Vss.n898 Vss.n897 383.418
R3402 Vss.t465 Vss.t176 370.279
R3403 Vss.t176 Vss.t208 370.279
R3404 Vss.t509 Vss.t673 370.05
R3405 Vss.t673 Vss.t23 370.05
R3406 Vss.t142 Vss.t476 370.05
R3407 Vss.t196 Vss.t142 370.05
R3408 Vss.t510 Vss.t143 370.05
R3409 Vss.t143 Vss.t390 370.05
R3410 Vss.n898 Vss.t467 367.392
R3411 Vss.n757 Vss.t497 367.392
R3412 Vss.n330 Vss.n329 366.255
R3413 Vss.n1047 Vss.t425 366.243
R3414 Vss.t190 Vss.n418 366.243
R3415 Vss.t416 Vss.n1040 366.243
R3416 Vss.n1041 Vss.t166 366.243
R3417 Vss.n1807 Vss.t415 366.243
R3418 Vss.n223 Vss.t58 366.243
R3419 Vss.n264 Vss.t426 366.243
R3420 Vss.t250 Vss.n72 366.243
R3421 Vss.t423 Vss.n62 366.243
R3422 Vss.n1070 Vss.t33 366.243
R3423 Vss.n1326 Vss.n1325 366.027
R3424 Vss.n1881 Vss.n16 366.027
R3425 Vss.n622 Vss.n617 366.027
R3426 Vss.n197 Vss.t424 365.705
R3427 Vss.t533 Vss.n124 365.705
R3428 Vss.t448 Vss.n120 361.933
R3429 Vss.t256 Vss.n1557 350.313
R3430 Vss.n1116 Vss.t349 338.849
R3431 Vss.n1121 Vss.t618 338.849
R3432 Vss.n1101 Vss.t293 338.849
R3433 Vss.n1133 Vss.t114 338.849
R3434 Vss.n1183 Vss.t472 338.849
R3435 Vss.n1638 Vss.t468 338.849
R3436 Vss.t591 Vss.n156 338.849
R3437 Vss.t350 Vss.n235 338.849
R3438 Vss.n1534 Vss.t17 338.849
R3439 Vss.t351 Vss.n1686 338.849
R3440 Vss.n1687 Vss.t2 338.849
R3441 Vss.n574 Vss.t471 338.849
R3442 Vss.t14 Vss.n686 338.849
R3443 Vss.n692 Vss.n691 330.211
R3444 Vss.n1755 Vss.n120 328.534
R3445 Vss.n643 Vss.n642 307.176
R3446 Vss.t425 Vss.t364 292.995
R3447 Vss.t364 Vss.t190 292.995
R3448 Vss.t359 Vss.t416 292.995
R3449 Vss.t166 Vss.t359 292.995
R3450 Vss.t300 Vss.t415 292.995
R3451 Vss.t58 Vss.t300 292.995
R3452 Vss.t426 Vss.t297 292.995
R3453 Vss.t297 Vss.t250 292.995
R3454 Vss.t319 Vss.t423 292.995
R3455 Vss.t33 Vss.t319 292.995
R3456 Vss.t424 Vss.t287 292.565
R3457 Vss.t287 Vss.t533 292.565
R3458 Vss.t422 Vss.n898 282.61
R3459 Vss.t369 Vss.n757 282.61
R3460 Vss.t565 Vss.n1602 282.512
R3461 Vss.n1618 Vss.t16 282.289
R3462 Vss.t665 Vss.n236 282.289
R3463 Vss.n1650 Vss.t676 282.289
R3464 Vss.n237 Vss.t342 282.289
R3465 Vss.t593 Vss.n191 282.289
R3466 Vss.n1641 Vss.t11 282.289
R3467 Vss.n1639 Vss.t110 282.289
R3468 Vss.n1701 Vss.t6 282.289
R3469 Vss.t349 Vss.t77 271.079
R3470 Vss.t77 Vss.t618 271.079
R3471 Vss.t293 Vss.t396 271.079
R3472 Vss.t396 Vss.t114 271.079
R3473 Vss.t472 Vss.t248 271.079
R3474 Vss.t248 Vss.t283 271.079
R3475 Vss.t468 Vss.t634 271.079
R3476 Vss.t634 Vss.t591 271.079
R3477 Vss.t341 Vss.t350 271.079
R3478 Vss.t17 Vss.t341 271.079
R3479 Vss.t10 Vss.t351 271.079
R3480 Vss.t2 Vss.t10 271.079
R3481 Vss.t19 Vss.t14 271.079
R3482 Vss.n1792 Vss.n102 266.082
R3483 Vss.n1603 Vss.t565 259.911
R3484 Vss.n1700 Vss.n102 250.827
R3485 Vss.n906 Vss.n532 250.815
R3486 Vss.n763 Vss.n540 250.815
R3487 Vss.n1017 Vss.n1016 247.475
R3488 Vss.t256 Vss.n1607 246.108
R3489 Vss.n237 Vss.n190 245.469
R3490 Vss.n1204 Vss.t633 240.12
R3491 Vss.n1494 Vss.n1493 232.143
R3492 Vss.n1496 Vss.n1495 232.143
R3493 Vss.n1489 Vss.n278 229.095
R3494 Vss.n1300 Vss.t46 228.071
R3495 Vss.n1300 Vss.t175 228.071
R3496 Vss.n1306 Vss.t173 228.071
R3497 Vss.n1306 Vss.t61 228.071
R3498 Vss.t63 Vss.n1256 228.071
R3499 Vss.t654 Vss.n439 228.004
R3500 Vss.n448 Vss.t638 228.004
R3501 Vss.t641 Vss.n368 228.004
R3502 Vss.t542 Vss.n368 228.004
R3503 Vss.n443 Vss.t540 228.004
R3504 Vss.t571 Vss.n1600 226.008
R3505 Vss.t16 Vss.t354 225.832
R3506 Vss.t354 Vss.t665 225.832
R3507 Vss.t314 Vss.t676 225.832
R3508 Vss.t342 Vss.t314 225.832
R3509 Vss.t292 Vss.t593 225.832
R3510 Vss.t11 Vss.t292 225.832
R3511 Vss.t502 Vss.t6 225.832
R3512 Vss.n1744 Vss.n1743 225.304
R3513 Vss.n687 Vss.t19 220.988
R3514 Vss.n1191 Vss.n371 213.623
R3515 Vss.n1745 Vss.n1744 211.958
R3516 Vss.n1584 Vss.n1570 205.139
R3517 Vss.n1570 Vss.n1564 205.139
R3518 Vss.n1585 Vss.n1564 205.139
R3519 Vss.n1585 Vss.n1584 205.139
R3520 Vss.n1518 Vss.n1517 200.773
R3521 Vss.t175 Vss.t173 193.861
R3522 Vss.t61 Vss.t63 193.861
R3523 Vss.t638 Vss.t641 193.804
R3524 Vss.t540 Vss.t542 193.804
R3525 Vss.n1583 Vss.n1581 193.476
R3526 Vss.n1587 Vss.n1566 193.476
R3527 Vss.n277 Vss.n275 191.959
R3528 Vss.n1519 Vss.n1518 186.831
R3529 Vss.n316 Vss.t552 179.683
R3530 Vss.n313 Vss.t552 179.683
R3531 Vss.t273 Vss.n281 179.683
R3532 Vss.n1233 Vss.t273 179.683
R3533 Vss.n1238 Vss.t236 179.683
R3534 Vss.n1239 Vss.t635 179.683
R3535 Vss.t635 Vss.n278 179.683
R3536 Vss.n1116 Vss.n1115 178.264
R3537 Vss.n1102 Vss.n1101 178.264
R3538 Vss.n1651 Vss.n235 178.264
R3539 Vss.n1686 Vss.n1685 178.264
R3540 Vss.n282 Vss.t125 172.196
R3541 Vss.t128 Vss.n1742 170.268
R3542 Vss.n1743 Vss.t128 170.268
R3543 Vss.n443 Vss.n317 167.056
R3544 Vss.n1579 Vss.n1572 166.989
R3545 Vss.n1592 Vss.n1567 166.989
R3546 Vss.n449 Vss.n448 166.254
R3547 Vss.n471 Vss.n470 165.725
R3548 Vss.n1809 Vss.n86 165.725
R3549 Vss.n1835 Vss.n1834 165.725
R3550 Vss.n1038 Vss.n1037 165.725
R3551 Vss.n1726 Vss.n1725 165.648
R3552 Vss.n1296 Vss.n291 161.839
R3553 Vss.n837 Vss.n11 161.839
R3554 Vss.n367 Vss.n366 160.189
R3555 Vss.n1640 Vss.n1638 156.166
R3556 Vss.n317 Vss.n316 154.976
R3557 Vss.n1234 Vss.n1233 152.731
R3558 Vss.n1239 Vss.n1238 152.731
R3559 Vss.n1148 Vss.n1147 151.869
R3560 Vss.n1091 Vss.n408 151.869
R3561 Vss.n452 Vss.n407 151.869
R3562 Vss.n365 Vss.n364 151.869
R3563 Vss.n1715 Vss.n100 151.869
R3564 Vss.n1297 Vss.n1273 151.869
R3565 Vss.n1662 Vss.n73 151.869
R3566 Vss.n1812 Vss.n75 151.869
R3567 Vss.n1446 Vss.n1426 151.869
R3568 Vss.n1493 Vss.n273 151.869
R3569 Vss.n1846 Vss.n1845 151.869
R3570 Vss.n1515 Vss.n1514 151.869
R3571 Vss.n1498 Vss.n1497 151.869
R3572 Vss.n1682 Vss.n1681 151.869
R3573 Vss.n1400 Vss.n1399 151.869
R3574 Vss.n932 Vss.n510 151.869
R3575 Vss.n1016 Vss.n1015 151.869
R3576 Vss.n851 Vss.n392 151.869
R3577 Vss.n891 Vss.n799 151.869
R3578 Vss.n816 Vss.n15 151.869
R3579 Vss.n641 Vss.n640 151.869
R3580 Vss.n626 Vss.n625 151.751
R3581 Vss.n1179 Vss.n396 151.751
R3582 Vss.n1153 Vss.n416 151.751
R3583 Vss.n1152 Vss.n1151 151.751
R3584 Vss.n1080 Vss.n416 151.751
R3585 Vss.n1151 Vss.n417 151.751
R3586 Vss.n1039 Vss.n499 151.751
R3587 Vss.n1028 Vss.n409 151.751
R3588 Vss.n983 Vss.n982 151.751
R3589 Vss.n1039 Vss.n500 151.751
R3590 Vss.n1001 Vss.n409 151.751
R3591 Vss.n1099 Vss.n1098 151.751
R3592 Vss.n1519 Vss.n250 151.751
R3593 Vss.n1516 Vss.n251 151.751
R3594 Vss.n490 Vss.n419 151.751
R3595 Vss.n460 Vss.n48 151.751
R3596 Vss.n1294 Vss.n1293 151.751
R3597 Vss.n1275 Vss.n1274 151.751
R3598 Vss.n1474 Vss.n289 151.751
R3599 Vss.n352 Vss.n351 151.751
R3600 Vss.n342 Vss.n290 151.751
R3601 Vss.n1477 Vss.n1476 151.751
R3602 Vss.n1194 Vss.n370 151.751
R3603 Vss.n139 Vss.n99 151.751
R3604 Vss.n1744 Vss.n123 151.751
R3605 Vss.n1796 Vss.n99 151.751
R3606 Vss.n1700 Vss.n170 151.751
R3607 Vss.n1700 Vss.n171 151.751
R3608 Vss.n1700 Vss.n1699 151.751
R3609 Vss.n1344 Vss.n1343 151.751
R3610 Vss.n1342 Vss.n1341 151.751
R3611 Vss.n1401 Vss.n1358 151.751
R3612 Vss.n1492 Vss.n274 151.751
R3613 Vss.n1808 Vss.n87 151.751
R3614 Vss.n224 Vss.n216 151.751
R3615 Vss.n1808 Vss.n88 151.751
R3616 Vss.n224 Vss.n222 151.751
R3617 Vss.n1824 Vss.n70 151.751
R3618 Vss.n1823 Vss.n1822 151.751
R3619 Vss.n1503 Vss.n1502 151.751
R3620 Vss.n1822 Vss.n71 151.751
R3621 Vss.n1654 Vss.n1653 151.751
R3622 Vss.n1543 Vss.n242 151.751
R3623 Vss.n1683 Vss.n193 151.751
R3624 Vss.n1379 Vss.n1359 151.751
R3625 Vss.n1820 Vss.n1819 151.751
R3626 Vss.n1445 Vss.n1444 151.751
R3627 Vss.n1833 Vss.n1832 151.751
R3628 Vss.n1069 Vss.n1060 151.751
R3629 Vss.n1833 Vss.n63 151.751
R3630 Vss.n1069 Vss.n1068 151.751
R3631 Vss.n1632 Vss.n1631 151.751
R3632 Vss.n1744 Vss.n125 151.751
R3633 Vss.n1739 Vss.n1738 151.751
R3634 Vss.n1744 Vss.n126 151.751
R3635 Vss.n1164 Vss.n1163 151.751
R3636 Vss.n524 Vss.n522 151.751
R3637 Vss.n974 Vss.n509 151.751
R3638 Vss.n874 Vss.n873 151.751
R3639 Vss.n841 Vss.n840 151.751
R3640 Vss.n863 Vss.n862 151.751
R3641 Vss.n973 Vss.n972 151.751
R3642 Vss.n836 Vss.n801 151.751
R3643 Vss.n839 Vss.n800 151.751
R3644 Vss.n806 Vss.n23 151.751
R3645 Vss.n611 Vss.n610 151.751
R3646 Vss.n601 Vss.n600 151.751
R3647 Vss.n592 Vss.n591 151.751
R3648 Vss.n677 Vss.n545 151.751
R3649 Vss.n1872 Vss.n1871 151.751
R3650 Vss.n667 Vss.n546 151.751
R3651 Vss.n663 Vss.n662 151.751
R3652 Vss.n644 Vss.n643 151.751
R3653 Vss.n1206 Vss.n1205 147.727
R3654 Vss.n1214 Vss.n1213 147.727
R3655 Vss.n1472 Vss.n1471 147.727
R3656 Vss.n1323 Vss.n1318 147.727
R3657 Vss.n624 Vss.n616 147.727
R3658 Vss.n1884 Vss.n1883 147.727
R3659 Vss.n1870 Vss.n1869 147.727
R3660 Vss.n888 Vss.n394 147.727
R3661 Vss.n719 Vss.n718 147.727
R3662 Vss.n739 Vss.n738 147.727
R3663 Vss.n1234 Vss.n276 143.746
R3664 Vss.t125 Vss.t459 137.756
R3665 Vss.t459 Vss.t169 137.756
R3666 Vss.n471 Vss.n416 135.501
R3667 Vss.n1809 Vss.n1808 135.501
R3668 Vss.n1834 Vss.n1833 135.501
R3669 Vss.n1039 Vss.n1038 135.501
R3670 Vss.n1725 Vss.n99 135.439
R3671 Vss.n1749 Vss.n1748 129.76
R3672 Vss.t283 Vss.n371 125.228
R3673 Vss.n1603 Vss.t569 124.305
R3674 Vss.t110 Vss.n169 120.279
R3675 Vss.n796 Vss.t442 119.157
R3676 Vss.n793 Vss.t442 119.157
R3677 Vss.n1589 Vss.n1569 118.222
R3678 Vss.n1161 Vss.t353 115.856
R3679 Vss.n470 Vss.t582 115.856
R3680 Vss.t367 Vss.n74 115.856
R3681 Vss.n86 Vss.t171 115.856
R3682 Vss.n1149 Vss.t360 115.856
R3683 Vss.n1835 Vss.t233 115.856
R3684 Vss.n265 Vss.t356 115.856
R3685 Vss.n270 Vss.t642 115.856
R3686 Vss.n975 Vss.t289 115.856
R3687 Vss.n1037 Vss.t206 115.856
R3688 Vss.n225 Vss.t320 115.802
R3689 Vss.n1726 Vss.t86 115.802
R3690 Vss.n1410 Vss.t132 114.944
R3691 Vss.t132 Vss.n1409 114.944
R3692 Vss.n1406 Vss.t240 114.944
R3693 Vss.n1487 Vss.t169 113.799
R3694 Vss.n793 Vss.n395 113.695
R3695 Vss.n1180 Vss.n1179 108.731
R3696 Vss.t156 Vss.t177 108.138
R3697 Vss.t192 Vss.t272 108.138
R3698 Vss.t181 Vss.t271 108.138
R3699 Vss.t195 Vss.t306 108.138
R3700 Vss.t221 Vss.t182 108.138
R3701 Vss.t229 Vss.t179 108.138
R3702 Vss.t224 Vss.t194 108.138
R3703 Vss.t336 Vss.t368 108.138
R3704 Vss.n169 Vss.t502 105.552
R3705 Vss.n797 Vss.n796 102.773
R3706 Vss.n1602 Vss.t571 101.704
R3707 Vss.t435 Vss.t183 99.0183
R3708 Vss.t178 Vss.t435 99.0183
R3709 Vss.n1409 Vss.n1406 97.7016
R3710 Vss.n329 Vss.t465 96.5949
R3711 Vss.n1325 Vss.t509 96.5352
R3712 Vss.t476 Vss.n16 96.5352
R3713 Vss.n622 Vss.t510 96.5352
R3714 Vss.n1047 Vss.n416 95.5419
R3715 Vss.n1151 Vss.n418 95.5419
R3716 Vss.n1040 Vss.n1039 95.5419
R3717 Vss.n1041 Vss.n409 95.5419
R3718 Vss.n1808 Vss.n1807 95.5419
R3719 Vss.n224 Vss.n223 95.5419
R3720 Vss.n1496 Vss.n264 95.5419
R3721 Vss.n1822 Vss.n72 95.5419
R3722 Vss.n1833 Vss.n62 95.5419
R3723 Vss.n1070 Vss.n1069 95.5419
R3724 Vss.n197 Vss.n99 95.4017
R3725 Vss.n1744 Vss.n124 95.4017
R3726 Vss.t189 Vss.t353 92.6849
R3727 Vss.t582 Vss.t189 92.6849
R3728 Vss.t60 Vss.t367 92.6849
R3729 Vss.t171 Vss.t60 92.6849
R3730 Vss.t360 Vss.t45 92.6849
R3731 Vss.t45 Vss.t233 92.6849
R3732 Vss.t356 Vss.t249 92.6849
R3733 Vss.t249 Vss.t642 92.6849
R3734 Vss.t289 Vss.t168 92.6849
R3735 Vss.t168 Vss.t206 92.6849
R3736 Vss.t320 Vss.t532 92.6419
R3737 Vss.t532 Vss.t86 92.6419
R3738 Vss.t177 Vss.t192 89.8983
R3739 Vss.t272 Vss.t181 89.8983
R3740 Vss.t271 Vss.t195 89.8983
R3741 Vss.t306 Vss.t180 89.8983
R3742 Vss.t193 Vss.t221 89.8983
R3743 Vss.t182 Vss.t229 89.8983
R3744 Vss.t179 Vss.t224 89.8983
R3745 Vss.t194 Vss.t336 89.8983
R3746 Vss.n1183 Vss.n1182 88.3958
R3747 Vss.n737 Vss.n548 87.3061
R3748 Vss.n737 Vss.n549 87.3061
R3749 Vss.n787 Vss.n534 87.3061
R3750 Vss.n787 Vss.n535 87.3061
R3751 Vss.n748 Vss.n542 87.3061
R3752 Vss.n748 Vss.n543 87.3061
R3753 Vss.n887 Vss.n882 87.3061
R3754 Vss.n887 Vss.n883 87.3061
R3755 Vss.n1885 Vss.n9 87.3061
R3756 Vss.n1885 Vss.n10 87.3061
R3757 Vss.n444 Vss.n442 87.3061
R3758 Vss.n445 Vss.n444 87.3061
R3759 Vss.n1303 Vss.n1298 87.3061
R3760 Vss.n1304 Vss.n1303 87.3061
R3761 Vss.n1317 Vss.n1311 87.3061
R3762 Vss.n1317 Vss.n1312 87.3061
R3763 Vss.n1215 Vss.n310 87.3061
R3764 Vss.n1215 Vss.n311 87.3061
R3765 Vss.n892 Vss.n791 87.3061
R3766 Vss.n893 Vss.n892 87.3061
R3767 Vss.n1775 Vss.n109 87.3061
R3768 Vss.n1775 Vss.n110 87.3061
R3769 Vss.n1791 Vss.n103 87.3061
R3770 Vss.n1791 Vss.n104 87.3061
R3771 Vss.n1411 Vss.n1410 86.8248
R3772 Vss.n1583 Vss.t156 80.7782
R3773 Vss.n1582 Vss.t303 80.7782
R3774 Vss.n1588 Vss.t139 80.7782
R3775 Vss.t368 Vss.n1587 80.7782
R3776 Vss.n1572 Vss.n1567 80.5005
R3777 Vss.n981 Vss.n980 76.452
R3778 Vss.n1701 Vss.n1700 73.641
R3779 Vss.n891 Vss.n797 72.984
R3780 Vss.t303 Vss.t116 69.0524
R3781 Vss.t139 Vss.t399 69.0524
R3782 Vss.n714 Vss.n552 67.4727
R3783 Vss.n715 Vss.n552 67.4727
R3784 Vss.n752 Vss.n538 67.4727
R3785 Vss.n753 Vss.n538 67.4727
R3786 Vss.n557 Vss.n556 67.4727
R3787 Vss.n558 Vss.n556 67.4727
R3788 Vss.n1868 Vss.n25 67.4727
R3789 Vss.n1868 Vss.n26 67.4727
R3790 Vss.n612 Vss.n6 67.4727
R3791 Vss.n613 Vss.n6 67.4727
R3792 Vss.n440 Vss.n303 67.4727
R3793 Vss.n446 Vss.n303 67.4727
R3794 Vss.n1299 Vss.n1242 67.4727
R3795 Vss.n1302 Vss.n1242 67.4727
R3796 Vss.n1470 Vss.n292 67.4727
R3797 Vss.n1470 Vss.n293 67.4727
R3798 Vss.n1207 Vss.n307 67.4727
R3799 Vss.n1208 Vss.n307 67.4727
R3800 Vss.n789 Vss.n31 67.4727
R3801 Vss.n894 Vss.n31 67.4727
R3802 Vss.n1746 Vss.n113 67.4727
R3803 Vss.n1747 Vss.n113 67.4727
R3804 Vss.n118 Vss.n117 67.4727
R3805 Vss.n119 Vss.n117 67.4727
R3806 Vss.n1739 Vss.n127 67.0503
R3807 Vss.n714 Vss.n548 66.5005
R3808 Vss.n715 Vss.n549 66.5005
R3809 Vss.n752 Vss.n534 66.5005
R3810 Vss.n753 Vss.n535 66.5005
R3811 Vss.n557 Vss.n542 66.5005
R3812 Vss.n558 Vss.n543 66.5005
R3813 Vss.n882 Vss.n25 66.5005
R3814 Vss.n883 Vss.n26 66.5005
R3815 Vss.n612 Vss.n9 66.5005
R3816 Vss.n613 Vss.n10 66.5005
R3817 Vss.n442 Vss.n440 66.5005
R3818 Vss.n446 Vss.n445 66.5005
R3819 Vss.n1299 Vss.n1298 66.5005
R3820 Vss.n1304 Vss.n1302 66.5005
R3821 Vss.n1311 Vss.n292 66.5005
R3822 Vss.n1312 Vss.n293 66.5005
R3823 Vss.n1207 Vss.n310 66.5005
R3824 Vss.n1208 Vss.n311 66.5005
R3825 Vss.n791 Vss.n789 66.5005
R3826 Vss.n894 Vss.n893 66.5005
R3827 Vss.n1746 Vss.n109 66.5005
R3828 Vss.n1747 Vss.n110 66.5005
R3829 Vss.n118 Vss.n103 66.5005
R3830 Vss.n119 Vss.n104 66.5005
R3831 Vss.n1614 Vss.n1554 65.5283
R3832 Vss.n1610 Vss.n1554 65.5283
R3833 Vss.n1610 Vss.n1555 65.5283
R3834 Vss.n1614 Vss.n1555 65.5283
R3835 Vss.n979 Vss.t113 63.4555
R3836 Vss.n1103 Vss.t403 63.4555
R3837 Vss.n482 Vss.t617 63.4555
R3838 Vss.n1113 Vss.t397 63.4555
R3839 Vss.n1114 Vss.t268 63.4555
R3840 Vss.n1520 Vss.t78 63.4555
R3841 Vss.n982 Vss.n981 62.5094
R3842 Vss.n1402 Vss.n127 61.7821
R3843 Vss.n449 Vss.t654 61.7514
R3844 Vss.n985 Vss.n984 61.0571
R3845 Vss.n1002 Vss.n999 61.0571
R3846 Vss.n1097 Vss.n484 61.0571
R3847 Vss.n1292 Vss.n1276 61.0571
R3848 Vss.n350 Vss.n343 61.0571
R3849 Vss.n1190 Vss.n1184 61.0571
R3850 Vss.n1710 Vss.n157 61.0571
R3851 Vss.n182 Vss.n181 61.0571
R3852 Vss.n1818 Vss.n76 61.0571
R3853 Vss.n1737 Vss.n128 61.0571
R3854 Vss.n872 Vss.n842 61.0571
R3855 Vss.n952 Vss.n525 61.0571
R3856 Vss.n825 Vss.n824 61.0571
R3857 Vss.n599 Vss.n593 61.0571
R3858 Vss.n661 Vss.n645 61.0571
R3859 Vss.n668 Vss.n572 61.0561
R3860 Vss.n620 Vss.n618 61.0561
R3861 Vss.n762 Vss.n759 61.0561
R3862 Vss.n1873 Vss.n21 61.0561
R3863 Vss.n1880 Vss.n17 61.0561
R3864 Vss.n905 Vss.n900 61.0561
R3865 Vss.n609 Vss.n604 61.0561
R3866 Vss.n628 Vss.n588 61.0561
R3867 Vss.n833 Vss.n807 61.0561
R3868 Vss.n817 Vss.n815 61.0561
R3869 Vss.n971 Vss.n511 61.0561
R3870 Vss.n864 Vss.n860 61.0561
R3871 Vss.n853 Vss.n850 61.0561
R3872 Vss.n1202 Vss.n386 61.0561
R3873 Vss.n943 Vss.n942 61.0561
R3874 Vss.n1018 Vss.n508 61.0561
R3875 Vss.n1014 Vss.n995 61.0561
R3876 Vss.n992 Vss.n976 61.0561
R3877 Vss.n1036 Vss.n503 61.0561
R3878 Vss.n1165 Vss.n405 61.0561
R3879 Vss.n933 Vss.n930 61.0561
R3880 Vss.n1390 Vss.n1388 61.0561
R3881 Vss.n1398 Vss.n1361 61.0561
R3882 Vss.n1727 Vss.n143 61.0561
R3883 Vss.n1722 Vss.n147 61.0561
R3884 Vss.n1680 Vss.n227 61.0561
R3885 Vss.n1688 Vss.n189 61.0561
R3886 Vss.n1702 Vss.n167 61.0561
R3887 Vss.n1643 Vss.n1642 61.0561
R3888 Vss.n1649 Vss.n238 61.0561
R3889 Vss.n1620 Vss.n1619 61.0561
R3890 Vss.n1550 Vss.n244 61.0561
R3891 Vss.n1513 Vss.n253 61.0561
R3892 Vss.n269 Vss.n266 61.0561
R3893 Vss.n1072 Vss.n1071 61.0561
R3894 Vss.n1067 Vss.n1061 61.0561
R3895 Vss.n1831 Vss.n64 61.0561
R3896 Vss.n1836 Vss.n58 61.0561
R3897 Vss.n1443 Vss.n1428 61.0561
R3898 Vss.n1844 Vss.n49 61.0561
R3899 Vss.n1849 Vss.n46 61.0561
R3900 Vss.n1175 Vss.n400 61.0561
R3901 Vss.n1160 Vss.n410 61.0561
R3902 Vss.n1049 Vss.n1048 61.0561
R3903 Vss.n1081 Vss.n1079 61.0561
R3904 Vss.n1154 Vss.n415 61.0561
R3905 Vss.n1042 Vss.n498 61.0561
R3906 Vss.n1030 Vss.n1029 61.0561
R3907 Vss.n492 Vss.n489 61.0561
R3908 Vss.n1092 Vss.n1089 61.0561
R3909 Vss.n1134 Vss.n436 61.0561
R3910 Vss.n1521 Vss.n249 61.0561
R3911 Vss.n1112 Vss.n478 61.0561
R3912 Vss.n1104 Vss.n481 61.0561
R3913 Vss.n1120 Vss.n1117 61.0561
R3914 Vss.n1124 Vss.n475 61.0561
R3915 Vss.n1130 Vss.n473 61.0561
R3916 Vss.n427 Vss.n426 61.0561
R3917 Vss.n1146 Vss.n421 61.0561
R3918 Vss.n467 Vss.n461 61.0561
R3919 Vss.n457 Vss.n453 61.0561
R3920 Vss.n1485 Vss.n283 61.0561
R3921 Vss.n1449 Vss.n1423 61.0561
R3922 Vss.n1438 Vss.n1437 61.0561
R3923 Vss.n1356 Vss.n1261 61.0561
R3924 Vss.n1340 Vss.n1334 61.0561
R3925 Vss.n1330 Vss.n1327 61.0561
R3926 Vss.n1345 Vss.n1270 61.0561
R3927 Vss.n1285 Vss.n1284 61.0561
R3928 Vss.n337 Vss.n331 61.0561
R3929 Vss.n1478 Vss.n288 61.0561
R3930 Vss.n355 Vss.n328 61.0561
R3931 Vss.n363 Vss.n320 61.0561
R3932 Vss.n1195 Vss.n390 61.0561
R3933 Vss.n199 Vss.n198 61.0561
R3934 Vss.n140 Vss.n138 61.0561
R3935 Vss.n1797 Vss.n98 61.0561
R3936 Vss.n1637 Vss.n1634 61.0561
R3937 Vss.n1629 Vss.n1627 61.0561
R3938 Vss.n1698 Vss.n172 61.0561
R3939 Vss.n1716 Vss.n154 61.0561
R3940 Vss.n1371 Vss.n1369 61.0561
R3941 Vss.n1417 Vss.n1416 61.0561
R3942 Vss.n204 Vss.n203 61.0561
R3943 Vss.n1806 Vss.n89 61.0561
R3944 Vss.n221 Vss.n217 61.0561
R3945 Vss.n215 Vss.n194 61.0561
R3946 Vss.n1055 Vss.n1054 61.0561
R3947 Vss.n1504 Vss.n263 61.0561
R3948 Vss.n1825 Vss.n69 61.0561
R3949 Vss.n1670 Vss.n1669 61.0561
R3950 Vss.n1663 Vss.n1660 61.0561
R3951 Vss.n1533 Vss.n1530 61.0561
R3952 Vss.n1537 Vss.n1529 61.0561
R3953 Vss.n1544 Vss.n1542 61.0561
R3954 Vss.n1655 Vss.n233 61.0561
R3955 Vss.n1381 Vss.n1380 61.0561
R3956 Vss.n1813 Vss.n82 61.0561
R3957 Vss.n521 Vss.n517 61.0561
R3958 Vss.n958 Vss.n516 61.0561
R3959 Vss.n639 Vss.n577 61.0561
R3960 Vss.n694 Vss.n565 61.0561
R3961 Vss.n685 Vss.n567 61.0561
R3962 Vss.n679 Vss.n676 61.0561
R3963 Vss.n653 Vss.n652 61.0561
R3964 Vss.n1759 Vss.t411 60.019
R3965 Vss.n1759 Vss.t84 60.019
R3966 Vss.t85 Vss.n1758 60.019
R3967 Vss.n1758 Vss.t650 60.019
R3968 Vss.t652 Vss.n1792 60.019
R3969 Vss.n1487 Vss.n1486 58.3972
R3970 Vss.n1490 Vss.n277 57.018
R3971 Vss.n1744 Vss.t411 54.0171
R3972 Vss.n1517 Vss.t315 53.4468
R3973 Vss.n1551 Vss.t269 53.4468
R3974 Vss.n993 Vss.t288 53.4468
R3975 Vss.n980 Vss.t409 53.4468
R3976 Vss.t240 Vss.n1402 53.1614
R3977 Vss.t84 Vss.t85 51.0162
R3978 Vss.t113 Vss.t352 50.7645
R3979 Vss.t352 Vss.t403 50.7645
R3980 Vss.t617 Vss.t298 50.7645
R3981 Vss.t298 Vss.t397 50.7645
R3982 Vss.t268 Vss.t299 50.7645
R3983 Vss.t299 Vss.t78 50.7645
R3984 Vss.n687 Vss.t471 50.0912
R3985 Vss.n1742 Vss.n1739 45.4054
R3986 Vss.n957 Vss.n956 45.3808
R3987 Vss.n1741 Vss.n116 44.1404
R3988 Vss.n708 Vss.n706 44.1404
R3989 Vss.n711 Vss.n555 44.1404
R3990 Vss.n775 Vss.n539 44.1394
R3991 Vss.n772 Vss.n4 44.1394
R3992 Vss.n766 Vss.n765 44.1394
R3993 Vss.n742 Vss.n741 44.1394
R3994 Vss.n910 Vss.n30 44.1394
R3995 Vss.n914 Vss.n913 44.1394
R3996 Vss.n917 Vss.n531 44.1394
R3997 Vss.n782 Vss.n781 44.1394
R3998 Vss.n795 Vss.n794 44.1394
R3999 Vss.n375 Vss.n304 44.1394
R4000 Vss.n379 Vss.n378 44.1394
R4001 Vss.n382 Vss.n36 44.1394
R4002 Vss.n1405 Vss.n1404 44.1394
R4003 Vss.n1408 Vss.n1247 44.1394
R4004 Vss.n1241 Vss.n1240 44.1394
R4005 Vss.n1237 Vss.n1235 44.1394
R4006 Vss.n1232 Vss.n298 44.1394
R4007 Vss.n315 Vss.n314 44.1394
R4008 Vss.n1321 Vss.n1320 44.1394
R4009 Vss.n1780 Vss.n1778 44.1394
R4010 Vss.n1785 Vss.n107 44.1394
R4011 Vss.n703 Vss.n561 44.1394
R4012 Vss.t315 Vss.t667 42.7575
R4013 Vss.t667 Vss.t269 42.7575
R4014 Vss.t405 Vss.t288 42.7575
R4015 Vss.t409 Vss.t405 42.7575
R4016 Vss.n720 Vss.n560 42.4436
R4017 Vss.n964 Vss.t681 41.0041
R4018 Vss.n1021 Vss.t677 41.0041
R4019 Vss.n164 Vss.t680 41.0041
R4020 Vss.n965 Vss.t679 40.8177
R4021 Vss.n1793 Vss.t650 38.0122
R4022 Vss.n956 Vss.n524 37.1047
R4023 Vss.t46 Vss.n275 36.1116
R4024 Vss.t236 Vss.n276 35.9369
R4025 Vss.n523 Vss.t103 35.0024
R4026 Vss.n1017 Vss.t4 35.0024
R4027 Vss.n1771 Vss.t678 34.1066
R4028 Vss.t567 Vss.n1557 33.9022
R4029 Vss.n798 Vss.t355 31.7253
R4030 Vss.n957 Vss.t407 31.7253
R4031 Vss.n693 Vss.n692 30.7136
R4032 Vss.n1586 Vss.n1570 30.5283
R4033 Vss.n1586 Vss.n1585 30.5283
R4034 Vss.n1495 Vss.n270 30.2237
R4035 Vss.n1016 Vss.n975 30.2237
R4036 Vss.n1604 Vss.n1603 29.4859
R4037 Vss.t103 Vss.t294 28.002
R4038 Vss.t294 Vss.t4 28.002
R4039 Vss.n1602 Vss.n1601 27.3737
R4040 Vss.t180 Vss.n1582 27.3607
R4041 Vss.n1588 Vss.t193 27.3607
R4042 Vss.n965 Vss.t100 27.1302
R4043 Vss.n964 Vss.t107 26.9438
R4044 Vss.n1021 Vss.t102 26.9438
R4045 Vss.n164 Vss.t109 26.9438
R4046 Vss.t355 Vss.t413 25.3804
R4047 Vss.t413 Vss.t407 25.3804
R4048 Vss.n1784 Vss.t0 24.9198
R4049 Vss.n1180 Vss.n395 24.8248
R4050 Vss.n691 Vss.t611 24.1401
R4051 Vss.n725 Vss.t611 24.1401
R4052 Vss.n725 Vss.t204 24.1401
R4053 Vss.t205 Vss.n724 24.1401
R4054 Vss.n724 Vss.t80 24.1401
R4055 Vss.n749 Vss.t82 24.1401
R4056 Vss.n756 Vss.t594 24.1401
R4057 Vss.t594 Vss.n755 24.1401
R4058 Vss.n755 Vss.t585 24.1401
R4059 Vss.t584 Vss.n751 24.1401
R4060 Vss.n751 Vss.t264 24.1401
R4061 Vss.n788 Vss.t262 24.1401
R4062 Vss.n897 Vss.t574 24.1401
R4063 Vss.t574 Vss.n896 24.1401
R4064 Vss.n896 Vss.t235 24.1401
R4065 Vss.n890 Vss.t231 24.1401
R4066 Vss.t71 Vss.n890 24.1401
R4067 Vss.t116 Vss.t183 20.8464
R4068 Vss.t399 Vss.t178 20.8464
R4069 Vss.n559 Vss.n548 20.8061
R4070 Vss.n559 Vss.n549 20.8061
R4071 Vss.n716 Vss.n714 20.8061
R4072 Vss.n716 Vss.n715 20.8061
R4073 Vss.n750 Vss.n534 20.8061
R4074 Vss.n750 Vss.n535 20.8061
R4075 Vss.n754 Vss.n752 20.8061
R4076 Vss.n754 Vss.n753 20.8061
R4077 Vss.n723 Vss.n542 20.8061
R4078 Vss.n723 Vss.n543 20.8061
R4079 Vss.n726 Vss.n557 20.8061
R4080 Vss.n726 Vss.n558 20.8061
R4081 Vss.n882 Vss.n881 20.8061
R4082 Vss.n883 Vss.n881 20.8061
R4083 Vss.n879 Vss.n25 20.8061
R4084 Vss.n879 Vss.n26 20.8061
R4085 Vss.n12 Vss.n9 20.8061
R4086 Vss.n12 Vss.n10 20.8061
R4087 Vss.n614 Vss.n612 20.8061
R4088 Vss.n614 Vss.n613 20.8061
R4089 Vss.n442 Vss.n441 20.8061
R4090 Vss.n445 Vss.n441 20.8061
R4091 Vss.n447 Vss.n440 20.8061
R4092 Vss.n447 Vss.n446 20.8061
R4093 Vss.n1305 Vss.n1298 20.8061
R4094 Vss.n1305 Vss.n1304 20.8061
R4095 Vss.n1301 Vss.n1299 20.8061
R4096 Vss.n1302 Vss.n1301 20.8061
R4097 Vss.n1313 Vss.n1311 20.8061
R4098 Vss.n1313 Vss.n1312 20.8061
R4099 Vss.n1308 Vss.n292 20.8061
R4100 Vss.n1308 Vss.n293 20.8061
R4101 Vss.n1209 Vss.n1207 20.8061
R4102 Vss.n1209 Vss.n1208 20.8061
R4103 Vss.n1211 Vss.n310 20.8061
R4104 Vss.n1211 Vss.n311 20.8061
R4105 Vss.n895 Vss.n789 20.8061
R4106 Vss.n895 Vss.n894 20.8061
R4107 Vss.n791 Vss.n790 20.8061
R4108 Vss.n893 Vss.n790 20.8061
R4109 Vss.n1754 Vss.n109 20.8061
R4110 Vss.n1754 Vss.n110 20.8061
R4111 Vss.n1748 Vss.n1746 20.8061
R4112 Vss.n1748 Vss.n1747 20.8061
R4113 Vss.n1561 Vss.n1554 20.8061
R4114 Vss.n1561 Vss.n1555 20.8061
R4115 Vss.n1757 Vss.n103 20.8061
R4116 Vss.n1757 Vss.n104 20.8061
R4117 Vss.n1760 Vss.n118 20.8061
R4118 Vss.n1760 Vss.n119 20.8061
R4119 Vss.t204 Vss.t205 20.5192
R4120 Vss.t80 Vss.t82 20.5192
R4121 Vss.t585 Vss.t584 20.5192
R4122 Vss.t264 Vss.t262 20.5192
R4123 Vss.t231 Vss.t235 20.5192
R4124 Vss.t73 Vss.t71 20.5192
R4125 Vss.n1617 Vss.n241 19.8869
R4126 Vss.n1770 Vss.t97 19.673
R4127 Vss.n1770 Vss.t104 19.4007
R4128 Vss.n1589 Vss.n1567 18.8616
R4129 Vss.n1572 Vss.n1569 18.8616
R4130 Vss.n1700 Vss.t0 18.5862
R4131 Vss.n560 Vss.n545 18.022
R4132 comparator_no_offsetcal_0.x3.avss Vss.n1597 17.8218
R4133 Vss.n1605 Vss.n1557 17.4164
R4134 Vss.n1576 comparator_no_offsetcal_0.x5.avss 16.7565
R4135 Vss.n982 Vss.n979 16.554
R4136 Vss.n1520 Vss.n1519 16.554
R4137 Vss.n1782 Vss.n102 16.1938
R4138 Vss.n1552 Vss.n1551 15.5696
R4139 Vss.n891 Vss.t73 14.6854
R4140 Vss.n1773 Vss.n1772 14.6135
R4141 Vss.n1016 Vss.n993 13.943
R4142 Vss.n165 SARlogic_0.dffrs_13.d 13.7563
R4143 Vss.n967 SARlogic_0.dffrs_12.clk 13.599
R4144 Vss.n1022 SARlogic_0.dffrs_12.d 13.599
R4145 Vss.n1793 Vss.t652 13.0045
R4146 Vss.n1590 Vss.n1568 11.0305
R4147 Vss.n524 Vss.n523 9.13142
R4148 Vss.n1576 Vss.n1573 9.05474
R4149 Vss.n1704 Vss.n165 9.04466
R4150 Vss.n1022 Vss.n1020 9.04027
R4151 Vss.n978 Vss.n480 9.03475
R4152 Vss.n507 Vss.n506 9.03475
R4153 Vss.n586 Vss.n583 9.0005
R4154 Vss.n832 Vss.n831 9.0005
R4155 Vss.n901 Vss.n20 9.0005
R4156 Vss.n1877 Vss.n1876 9.0005
R4157 Vss.n859 Vss.n858 9.0005
R4158 Vss.n945 Vss.n944 9.0005
R4159 Vss.n1167 Vss.n403 9.0005
R4160 Vss.n1063 Vss.n1062 9.0005
R4161 Vss.n989 Vss.n988 9.0005
R4162 Vss.n1006 Vss.n1005 9.0005
R4163 Vss.n1008 Vss.n485 9.0005
R4164 Vss.n1013 Vss.n1012 9.0005
R4165 Vss.n1011 Vss.n997 9.0005
R4166 Vss.n431 Vss.n430 9.0005
R4167 Vss.n1144 Vss.n1142 9.0005
R4168 Vss.n466 Vss.n465 9.0005
R4169 Vss.n45 Vss.n42 9.0005
R4170 Vss.n455 Vss.n402 9.0005
R4171 Vss.n1430 Vss.n1429 9.0005
R4172 Vss.n53 Vss.n51 9.0005
R4173 Vss.n1422 Vss.n1252 9.0005
R4174 Vss.n1269 Vss.n1268 9.0005
R4175 Vss.n1291 Vss.n1290 9.0005
R4176 Vss.n1278 Vss.n1267 9.0005
R4177 Vss.n332 Vss.n284 9.0005
R4178 Vss.n349 Vss.n348 9.0005
R4179 Vss.n347 Vss.n345 9.0005
R4180 Vss.n362 Vss.n321 9.0005
R4181 Vss.n361 Vss.n359 9.0005
R4182 Vss.n357 Vss.n356 9.0005
R4183 Vss.n326 Vss.n325 9.0005
R4184 Vss.n1483 Vss.n1482 9.0005
R4185 Vss.n333 Vss.n287 9.0005
R4186 Vss.n1481 Vss.n1480 9.0005
R4187 Vss.n1185 Vss.n387 9.0005
R4188 Vss.n1186 Vss.n389 9.0005
R4189 Vss.n1198 Vss.n1197 9.0005
R4190 Vss.n1200 Vss.n1199 9.0005
R4191 Vss.n174 Vss.n173 9.0005
R4192 Vss.n163 Vss.n159 9.0005
R4193 Vss.n179 Vss.n178 9.0005
R4194 Vss.n185 Vss.n184 9.0005
R4195 Vss.n1696 Vss.n1695 9.0005
R4196 Vss.n175 Vss.n152 9.0005
R4197 Vss.n1335 Vss.n1262 9.0005
R4198 Vss.n1337 Vss.n1336 9.0005
R4199 Vss.n1338 Vss.n1264 9.0005
R4200 Vss.n1354 Vss.n1353 9.0005
R4201 Vss.n1348 Vss.n1347 9.0005
R4202 Vss.n1287 Vss.n1286 9.0005
R4203 Vss.n1281 Vss.n1280 9.0005
R4204 Vss.n218 Vss.n92 9.0005
R4205 Vss.n1674 Vss.n1673 9.0005
R4206 Vss.n1658 Vss.n230 9.0005
R4207 Vss.n1432 Vss.n77 9.0005
R4208 Vss.n1435 Vss.n1434 9.0005
R4209 Vss.n1736 Vss.n1735 9.0005
R4210 Vss.n1734 Vss.n130 9.0005
R4211 Vss.n1396 Vss.n1394 9.0005
R4212 Vss.n1392 Vss.n1391 9.0005
R4213 Vss.n1386 Vss.n132 9.0005
R4214 Vss.n136 Vss.n133 9.0005
R4215 Vss.n202 Vss.n201 9.0005
R4216 Vss.n1720 Vss.n1718 9.0005
R4217 Vss.n1718 Vss.n1717 9.0005
R4218 Vss.n149 Vss.n96 9.0005
R4219 Vss.n1706 Vss.n166 9.0005
R4220 Vss.n1706 Vss.n1705 9.0005
R4221 Vss.n1708 Vss.n161 9.0005
R4222 Vss.n1709 Vss.n1708 9.0005
R4223 Vss.n1647 Vss.n1645 9.0005
R4224 Vss.n1645 Vss.n1644 9.0005
R4225 Vss.n1527 Vss.n188 9.0005
R4226 Vss.n1625 Vss.n188 9.0005
R4227 Vss.n1672 Vss.n228 9.0005
R4228 Vss.n1679 Vss.n228 9.0005
R4229 Vss.n219 Vss.n93 9.0005
R4230 Vss.n1678 Vss.n1676 9.0005
R4231 Vss.n1721 Vss.n148 9.0005
R4232 Vss.n1799 Vss.n1798 9.0005
R4233 Vss.n1804 Vss.n1802 9.0005
R4234 Vss.n196 Vss.n91 9.0005
R4235 Vss.n213 Vss.n212 9.0005
R4236 Vss.n142 Vss.n141 9.0005
R4237 Vss.n1377 Vss.n1376 9.0005
R4238 Vss.n1397 Vss.n1362 9.0005
R4239 Vss.n1367 Vss.n1363 9.0005
R4240 Vss.n1364 Vss.n80 9.0005
R4241 Vss.n1383 Vss.n1382 9.0005
R4242 Vss.n1373 Vss.n1372 9.0005
R4243 Vss.n1419 Vss.n1418 9.0005
R4244 Vss.n1816 Vss.n1815 9.0005
R4245 Vss.n1815 Vss.n1814 9.0005
R4246 Vss.n1254 Vss.n1253 9.0005
R4247 Vss.n1052 Vss.n90 9.0005
R4248 Vss.n1805 Vss.n90 9.0005
R4249 Vss.n208 Vss.n67 9.0005
R4250 Vss.n208 Vss.n195 9.0005
R4251 Vss.n1665 Vss.n1657 9.0005
R4252 Vss.n1665 Vss.n1664 9.0005
R4253 Vss.n261 Vss.n260 9.0005
R4254 Vss.n1623 Vss.n1622 9.0005
R4255 Vss.n1648 Vss.n1623 9.0005
R4256 Vss.n1540 Vss.n1539 9.0005
R4257 Vss.n1539 Vss.n1538 9.0005
R4258 Vss.n1524 Vss.n1523 9.0005
R4259 Vss.n1524 Vss.n240 9.0005
R4260 Vss.n1546 Vss.n246 9.0005
R4261 Vss.n1546 Vss.n1545 9.0005
R4262 Vss.n429 Vss.n254 9.0005
R4263 Vss.n1512 Vss.n254 9.0005
R4264 Vss.n1065 Vss.n1064 9.0005
R4265 Vss.n1511 Vss.n1509 9.0005
R4266 Vss.n257 Vss.n232 9.0005
R4267 Vss.n1506 Vss.n1505 9.0005
R4268 Vss.n1058 Vss.n1057 9.0005
R4269 Vss.n1057 Vss.n1056 9.0005
R4270 Vss.n1829 Vss.n1827 9.0005
R4271 Vss.n1827 Vss.n1826 9.0005
R4272 Vss.n1441 Vss.n1440 9.0005
R4273 Vss.n1440 Vss.n1439 9.0005
R4274 Vss.n1452 Vss.n1451 9.0005
R4275 Vss.n1842 Vss.n52 9.0005
R4276 Vss.n1843 Vss.n1842 9.0005
R4277 Vss.n1852 Vss.n1851 9.0005
R4278 Vss.n1074 Vss.n1051 9.0005
R4279 Vss.n1074 Vss.n1073 9.0005
R4280 Vss.n413 Vss.n57 9.0005
R4281 Vss.n1830 Vss.n57 9.0005
R4282 Vss.n487 Vss.n422 9.0005
R4283 Vss.n1145 Vss.n422 9.0005
R4284 Vss.n1077 Vss.n1076 9.0005
R4285 Vss.n1110 Vss.n1109 9.0005
R4286 Vss.n1109 Vss.n248 9.0005
R4287 Vss.n1128 Vss.n1126 9.0005
R4288 Vss.n1126 Vss.n1125 9.0005
R4289 Vss.n1107 Vss.n1106 9.0005
R4290 Vss.n1108 Vss.n1107 9.0005
R4291 Vss.n987 Vss.n435 9.0005
R4292 Vss.n1129 Vss.n435 9.0005
R4293 Vss.n1095 Vss.n1094 9.0005
R4294 Vss.n1094 Vss.n1093 9.0005
R4295 Vss.n1004 Vss.n1000 9.0005
R4296 Vss.n1087 Vss.n1086 9.0005
R4297 Vss.n494 Vss.n493 9.0005
R4298 Vss.n1083 Vss.n1082 9.0005
R4299 Vss.n1045 Vss.n1044 9.0005
R4300 Vss.n1046 Vss.n1045 9.0005
R4301 Vss.n1156 Vss.n411 9.0005
R4302 Vss.n1156 Vss.n1155 9.0005
R4303 Vss.n454 Vss.n403 9.0005
R4304 Vss.n1173 Vss.n1171 9.0005
R4305 Vss.n1174 Vss.n401 9.0005
R4306 Vss.n1169 Vss.n1168 9.0005
R4307 Vss.n928 Vss.n926 9.0005
R4308 Vss.n871 Vss.n870 9.0005
R4309 Vss.n869 Vss.n844 9.0005
R4310 Vss.n867 Vss.n866 9.0005
R4311 Vss.n849 Vss.n848 9.0005
R4312 Vss.n856 Vss.n855 9.0005
R4313 Vss.n527 Vss.n526 9.0005
R4314 Vss.n950 Vss.n949 9.0005
R4315 Vss.n947 Vss.n512 9.0005
R4316 Vss.n520 Vss.n515 9.0005
R4317 Vss.n519 Vss.n505 9.0005
R4318 Vss.n969 Vss.n968 9.0005
R4319 Vss.n939 Vss.n938 9.0005
R4320 Vss.n1024 Vss.n497 9.0005
R4321 Vss.n1032 Vss.n1031 9.0005
R4322 Vss.n935 Vss.n934 9.0005
R4323 Vss.n903 Vss.n902 9.0005
R4324 Vss.n1875 Vss.n22 9.0005
R4325 Vss.n823 Vss.n822 9.0005
R4326 Vss.n828 Vss.n827 9.0005
R4327 Vss.n830 Vss.n809 9.0005
R4328 Vss.n819 Vss.n818 9.0005
R4329 Vss.n813 Vss.n812 9.0005
R4330 Vss.n598 Vss.n597 9.0005
R4331 Vss.n596 Vss.n595 9.0005
R4332 Vss.n638 Vss.n578 9.0005
R4333 Vss.n637 Vss.n635 9.0005
R4334 Vss.n605 Vss.n580 9.0005
R4335 Vss.n607 Vss.n606 9.0005
R4336 Vss.n630 Vss.n629 9.0005
R4337 Vss.n681 Vss.n680 9.0005
R4338 Vss.n660 Vss.n659 9.0005
R4339 Vss.n647 Vss.n569 9.0005
R4340 Vss.n650 Vss.n649 9.0005
R4341 Vss.n656 Vss.n655 9.0005
R4342 Vss.n571 Vss.n570 9.0005
R4343 Vss.n671 Vss.n670 9.0005
R4344 Vss.n674 Vss.n563 9.0005
R4345 Vss.n564 Vss.n562 9.0005
R4346 Vss.n697 Vss.n696 9.0005
R4347 Vss.n1601 Vss.t572 8.70131
R4348 Vss.n891 Vss.n798 8.27654
R4349 Vss.n1400 Vss.n1359 8.08508
R4350 Vss.n1365 Vss.n1249 8.05717
R4351 Vss.n1596 Vss.n1595 7.7564
R4352 Vss.n1577 Vss.n1571 7.59387
R4353 Vss.n1501 Vss.n1499 7.29099
R4354 Vss.n618 Vss.n584 6.9012
R4355 Vss.n1880 Vss.n1879 6.9012
R4356 Vss.n1034 Vss.n503 6.9012
R4357 Vss.n1729 Vss.n143 6.9012
R4358 Vss.n1690 Vss.n189 6.9012
R4359 Vss.n1548 Vss.n244 6.9012
R4360 Vss.n267 Vss.n266 6.9012
R4361 Vss.n1838 Vss.n58 6.9012
R4362 Vss.n1160 Vss.n1159 6.9012
R4363 Vss.n1136 Vss.n436 6.9012
R4364 Vss.n992 Vss.n991 6.9012
R4365 Vss.n1118 Vss.n1117 6.9012
R4366 Vss.n335 Vss.n331 6.9012
R4367 Vss.n1188 Vss.n1184 6.9012
R4368 Vss.n1637 Vss.n1636 6.9012
R4369 Vss.n1328 Vss.n1327 6.9012
R4370 Vss.n206 Vss.n203 6.9012
R4371 Vss.n1531 Vss.n1530 6.9012
R4372 Vss.n960 Vss.n516 6.9012
R4373 Vss.n683 Vss.n567 6.9012
R4374 Vss.n760 Vss.n759 6.90005
R4375 Vss.n1579 Vss.n1578 6.64904
R4376 Vss.n1606 Vss.n1558 6.5795
R4377 Vss.n1560 Vss.n1559 6.5795
R4378 Vss.n572 Vss.n571 6.46296
R4379 Vss.n605 Vss.n604 6.46296
R4380 Vss.n629 Vss.n628 6.46296
R4381 Vss.n833 Vss.n832 6.46296
R4382 Vss.n1876 Vss.n21 6.46296
R4383 Vss.n512 Vss.n511 6.46296
R4384 Vss.n860 Vss.n859 6.46296
R4385 Vss.n1168 Vss.n405 6.46296
R4386 Vss.n1391 Vss.n1390 6.46296
R4387 Vss.n1398 Vss.n1397 6.46296
R4388 Vss.n1722 Vss.n1721 6.46296
R4389 Vss.n1680 Vss.n1679 6.46296
R4390 Vss.n1513 Vss.n1512 6.46296
R4391 Vss.n1831 Vss.n1830 6.46296
R4392 Vss.n1155 Vss.n1154 6.46296
R4393 Vss.n1031 Vss.n1030 6.46296
R4394 Vss.n493 Vss.n492 6.46296
R4395 Vss.n1093 Vss.n1092 6.46296
R4396 Vss.n988 Vss.n984 6.46296
R4397 Vss.n485 Vss.n484 6.46296
R4398 Vss.n1014 Vss.n1013 6.46296
R4399 Vss.n1125 Vss.n1124 6.46296
R4400 Vss.n1130 Vss.n1129 6.46296
R4401 Vss.n430 Vss.n426 6.46296
R4402 Vss.n1146 Vss.n1145 6.46296
R4403 Vss.n467 Vss.n466 6.46296
R4404 Vss.n454 Vss.n453 6.46296
R4405 Vss.n1430 Vss.n1428 6.46296
R4406 Vss.n1844 Vss.n1843 6.46296
R4407 Vss.n1270 Vss.n1269 6.46296
R4408 Vss.n356 Vss.n355 6.46296
R4409 Vss.n363 Vss.n362 6.46296
R4410 Vss.n288 Vss.n287 6.46296
R4411 Vss.n390 Vss.n389 6.46296
R4412 Vss.n141 Vss.n140 6.46296
R4413 Vss.n1627 Vss.n1625 6.46296
R4414 Vss.n173 Vss.n172 6.46296
R4415 Vss.n1710 Vss.n1709 6.46296
R4416 Vss.n1717 Vss.n1716 6.46296
R4417 Vss.n1337 Vss.n1334 6.46296
R4418 Vss.n1286 Vss.n1285 6.46296
R4419 Vss.n195 Vss.n194 6.46296
R4420 Vss.n1826 Vss.n1825 6.46296
R4421 Vss.n1673 Vss.n1669 6.46296
R4422 Vss.n1664 Vss.n1663 6.46296
R4423 Vss.n1538 Vss.n1537 6.46296
R4424 Vss.n1545 Vss.n1544 6.46296
R4425 Vss.n233 Vss.n232 6.46296
R4426 Vss.n1382 Vss.n1381 6.46296
R4427 Vss.n1814 Vss.n1813 6.46296
R4428 Vss.n77 Vss.n76 6.46296
R4429 Vss.n1439 Vss.n1438 6.46296
R4430 Vss.n934 Vss.n933 6.46296
R4431 Vss.n521 Vss.n520 6.46296
R4432 Vss.n850 Vss.n849 6.46296
R4433 Vss.n526 Vss.n525 6.46296
R4434 Vss.n818 Vss.n817 6.46296
R4435 Vss.n639 Vss.n638 6.46296
R4436 Vss.n680 Vss.n679 6.46296
R4437 Vss.n652 Vss.n650 6.46296
R4438 Vss.n901 Vss.n900 6.4618
R4439 Vss.n944 Vss.n943 6.4618
R4440 Vss.n508 Vss.n507 6.4618
R4441 Vss.n1644 Vss.n1643 6.4618
R4442 Vss.n1649 Vss.n1648 6.4618
R4443 Vss.n1619 Vss.n240 6.4618
R4444 Vss.n1073 Vss.n1072 6.4618
R4445 Vss.n1063 Vss.n1061 6.4618
R4446 Vss.n1175 Vss.n1174 6.4618
R4447 Vss.n1048 Vss.n1046 6.4618
R4448 Vss.n1082 Vss.n1081 6.4618
R4449 Vss.n498 Vss.n497 6.4618
R4450 Vss.n249 Vss.n248 6.4618
R4451 Vss.n1108 Vss.n478 6.4618
R4452 Vss.n1005 Vss.n999 6.4618
R4453 Vss.n481 Vss.n480 6.4618
R4454 Vss.n46 Vss.n45 6.4618
R4455 Vss.n1423 Vss.n1422 6.4618
R4456 Vss.n1292 Vss.n1291 6.4618
R4457 Vss.n284 Vss.n283 6.4618
R4458 Vss.n350 Vss.n349 6.4618
R4459 Vss.n387 Vss.n386 6.4618
R4460 Vss.n198 Vss.n196 6.4618
R4461 Vss.n1798 Vss.n1797 6.4618
R4462 Vss.n1705 Vss.n167 6.4618
R4463 Vss.n181 Vss.n179 6.4618
R4464 Vss.n1262 Vss.n1261 6.4618
R4465 Vss.n1372 Vss.n1371 6.4618
R4466 Vss.n1418 Vss.n1417 6.4618
R4467 Vss.n1806 Vss.n1805 6.4618
R4468 Vss.n218 Vss.n217 6.4618
R4469 Vss.n1056 Vss.n1055 6.4618
R4470 Vss.n1505 Vss.n1504 6.4618
R4471 Vss.n1737 Vss.n1736 6.4618
R4472 Vss.n872 Vss.n871 6.4618
R4473 Vss.n824 Vss.n823 6.4618
R4474 Vss.n599 Vss.n598 6.4618
R4475 Vss.n565 Vss.n564 6.4618
R4476 Vss.n661 Vss.n660 6.4618
R4477 Vss.n1595 Vss.n1564 6.33584
R4478 Vss.n1584 Vss.n1571 6.32806
R4479 Vss.n1590 Vss.n1589 6.23383
R4480 SARlogic_0.dffrs_12.nand3_1.A Vss.n964 5.7755
R4481 SARlogic_0.dffrs_12.nand3_8.A Vss.n1021 5.7755
R4482 SARlogic_0.dffrs_13.nand3_8.A Vss.n164 5.7755
R4483 SARlogic_0.dffrs_12.nand3_6.B Vss.n965 5.47979
R4484 Vss.n1879 Vss.n18 5.47239
R4485 Vss.n1035 Vss.n1034 5.47239
R4486 Vss.n1729 Vss.n1728 5.47239
R4487 Vss.n1690 Vss.n1689 5.47239
R4488 Vss.n1549 Vss.n1548 5.47239
R4489 Vss.n268 Vss.n267 5.47239
R4490 Vss.n1838 Vss.n1837 5.47239
R4491 Vss.n1159 Vss.n1158 5.47239
R4492 Vss.n1136 Vss.n1135 5.47239
R4493 Vss.n991 Vss.n977 5.47239
R4494 Vss.n1119 Vss.n1118 5.47239
R4495 Vss.n336 Vss.n335 5.47239
R4496 Vss.n1189 Vss.n1188 5.47239
R4497 Vss.n1636 Vss.n1635 5.47239
R4498 Vss.n1329 Vss.n1328 5.47239
R4499 Vss.n206 Vss.n205 5.47239
R4500 Vss.n1532 Vss.n1531 5.47239
R4501 Vss.n960 Vss.n959 5.47239
R4502 Vss.n619 Vss.n584 5.47239
R4503 Vss.n761 Vss.n760 5.47239
R4504 Vss.n684 Vss.n683 5.47239
R4505 Vss.n1772 Vss.n1771 5.18044
R4506 Vss.n670 Vss.n669 5.03414
R4507 Vss.n608 Vss.n607 5.03414
R4508 Vss.n587 Vss.n586 5.03414
R4509 Vss.n814 Vss.n813 5.03414
R4510 Vss.n809 Vss.n808 5.03414
R4511 Vss.n904 Vss.n903 5.03414
R4512 Vss.n1875 Vss.n1874 5.03414
R4513 Vss.n970 Vss.n969 5.03414
R4514 Vss.n855 Vss.n854 5.03414
R4515 Vss.n866 Vss.n865 5.03414
R4516 Vss.n940 Vss.n939 5.03414
R4517 Vss.n1020 Vss.n1019 5.03414
R4518 Vss.n929 Vss.n928 5.03414
R4519 Vss.n1167 Vss.n1166 5.03414
R4520 Vss.n1387 Vss.n1386 5.03414
R4521 Vss.n1396 Vss.n1395 5.03414
R4522 Vss.n1720 Vss.n1719 5.03414
R4523 Vss.n1678 Vss.n1677 5.03414
R4524 Vss.n1624 Vss.n166 5.03414
R4525 Vss.n1647 Vss.n1646 5.03414
R4526 Vss.n1622 Vss.n1621 5.03414
R4527 Vss.n1511 Vss.n1510 5.03414
R4528 Vss.n1059 Vss.n1058 5.03414
R4529 Vss.n1066 Vss.n1065 5.03414
R4530 Vss.n1829 Vss.n1828 5.03414
R4531 Vss.n1173 Vss.n1172 5.03414
R4532 Vss.n1051 Vss.n1050 5.03414
R4533 Vss.n1078 Vss.n1077 5.03414
R4534 Vss.n414 Vss.n413 5.03414
R4535 Vss.n1044 Vss.n1043 5.03414
R4536 Vss.n1027 Vss.n411 5.03414
R4537 Vss.n488 Vss.n487 5.03414
R4538 Vss.n1088 Vss.n1087 5.03414
R4539 Vss.n1523 Vss.n1522 5.03414
R4540 Vss.n1111 Vss.n1110 5.03414
R4541 Vss.n1106 Vss.n1105 5.03414
R4542 Vss.n987 Vss.n986 5.03414
R4543 Vss.n1004 Vss.n1003 5.03414
R4544 Vss.n1096 Vss.n1095 5.03414
R4545 Vss.n997 Vss.n996 5.03414
R4546 Vss.n474 Vss.n246 5.03414
R4547 Vss.n1128 Vss.n1127 5.03414
R4548 Vss.n1144 Vss.n1143 5.03414
R4549 Vss.n429 Vss.n428 5.03414
R4550 Vss.n456 Vss.n455 5.03414
R4551 Vss.n459 Vss.n52 5.03414
R4552 Vss.n1851 Vss.n1850 5.03414
R4553 Vss.n1451 Vss.n1450 5.03414
R4554 Vss.n1442 Vss.n1441 5.03414
R4555 Vss.n51 Vss.n50 5.03414
R4556 Vss.n1436 Vss.n1435 5.03414
R4557 Vss.n1282 Vss.n1281 5.03414
R4558 Vss.n1347 Vss.n1346 5.03414
R4559 Vss.n1278 Vss.n1277 5.03414
R4560 Vss.n1480 Vss.n1479 5.03414
R4561 Vss.n1484 Vss.n1483 5.03414
R4562 Vss.n327 Vss.n326 5.03414
R4563 Vss.n361 Vss.n360 5.03414
R4564 Vss.n345 Vss.n344 5.03414
R4565 Vss.n1201 Vss.n1200 5.03414
R4566 Vss.n1197 Vss.n1196 5.03414
R4567 Vss.n201 Vss.n200 5.03414
R4568 Vss.n137 Vss.n136 5.03414
R4569 Vss.n97 Vss.n96 5.03414
R4570 Vss.n1628 Vss.n161 5.03414
R4571 Vss.n153 Vss.n152 5.03414
R4572 Vss.n1697 Vss.n1696 5.03414
R4573 Vss.n159 Vss.n158 5.03414
R4574 Vss.n1704 Vss.n1703 5.03414
R4575 Vss.n184 Vss.n183 5.03414
R4576 Vss.n1355 Vss.n1354 5.03414
R4577 Vss.n1339 Vss.n1338 5.03414
R4578 Vss.n1368 Vss.n1367 5.03414
R4579 Vss.n1255 Vss.n1254 5.03414
R4580 Vss.n1804 Vss.n1803 5.03414
R4581 Vss.n220 Vss.n219 5.03414
R4582 Vss.n214 Vss.n213 5.03414
R4583 Vss.n1053 Vss.n1052 5.03414
R4584 Vss.n262 Vss.n261 5.03414
R4585 Vss.n68 Vss.n67 5.03414
R4586 Vss.n1659 Vss.n1658 5.03414
R4587 Vss.n1672 Vss.n1671 5.03414
R4588 Vss.n1528 Vss.n1527 5.03414
R4589 Vss.n1541 Vss.n1540 5.03414
R4590 Vss.n1657 Vss.n1656 5.03414
R4591 Vss.n1378 Vss.n1377 5.03414
R4592 Vss.n81 Vss.n80 5.03414
R4593 Vss.n1817 Vss.n1816 5.03414
R4594 Vss.n130 Vss.n129 5.03414
R4595 Vss.n519 Vss.n518 5.03414
R4596 Vss.n844 Vss.n843 5.03414
R4597 Vss.n951 Vss.n950 5.03414
R4598 Vss.n827 Vss.n826 5.03414
R4599 Vss.n637 Vss.n636 5.03414
R4600 Vss.n595 Vss.n594 5.03414
R4601 Vss.n696 Vss.n695 5.03414
R4602 Vss.n675 Vss.n674 5.03414
R4603 Vss.n655 Vss.n654 5.03414
R4604 Vss.n647 Vss.n646 5.03414
R4605 Vss.n909 Vss.t66 4.84702
R4606 Vss.n908 Vss.t112 4.84702
R4607 Vss.n374 Vss.t647 4.84702
R4608 Vss.n373 Vss.t450 4.84702
R4609 Vss.n297 Vss.t636 4.84702
R4610 Vss.n1236 Vss.t237 4.84702
R4611 Vss.n1740 Vss.t129 4.84702
R4612 Vss.n1403 Vss.t241 4.84702
R4613 Vss.n710 Vss.t402 4.84702
R4614 Vss.n707 Vss.t302 4.84702
R4615 Vss.n769 Vss.t131 4.84702
R4616 Vss.n771 Vss.t239 4.84702
R4617 Vss.n1700 Vss.n168 4.79462
R4618 Vss.n669 Vss.t93 4.7885
R4619 Vss.n780 Vss.t562 4.7885
R4620 Vss.n761 Vss.t145 4.7885
R4621 Vss.n619 Vss.t391 4.7885
R4622 Vss.n608 Vss.t579 4.7885
R4623 Vss.n587 Vss.t529 4.7885
R4624 Vss.n7 Vss.t606 4.7885
R4625 Vss.n8 Vss.t199 4.7885
R4626 Vss.n1886 Vss.t187 4.7885
R4627 Vss.n814 Vss.t492 4.7885
R4628 Vss.n808 Vss.t577 4.7885
R4629 Vss.n904 Vss.t141 4.7885
R4630 Vss.n1874 Vss.t621 4.7885
R4631 Vss.n18 Vss.t197 4.7885
R4632 Vss.n970 Vss.t68 4.7885
R4633 Vss.n854 Vss.t464 4.7885
R4634 Vss.n865 Vss.t267 4.7885
R4635 Vss.n940 Vss.t326 4.7885
R4636 Vss.n1019 Vss.t5 4.7885
R4637 Vss.n1035 Vss.t207 4.7885
R4638 Vss.n929 Vss.t247 4.7885
R4639 Vss.n1166 Vss.t347 4.7885
R4640 Vss.n1387 Vss.t56 4.7885
R4641 Vss.n1395 Vss.t669 4.7885
R4642 Vss.n1728 Vss.t87 4.7885
R4643 Vss.n1719 Vss.t452 4.7885
R4644 Vss.n1677 Vss.t494 4.7885
R4645 Vss.n1689 Vss.t3 4.7885
R4646 Vss.n1624 Vss.t12 4.7885
R4647 Vss.n1646 Vss.t343 4.7885
R4648 Vss.n1621 Vss.t666 4.7885
R4649 Vss.n1549 Vss.t270 4.7885
R4650 Vss.n1510 Vss.t488 4.7885
R4651 Vss.n268 Vss.t643 4.7885
R4652 Vss.n1059 Vss.t34 4.7885
R4653 Vss.n1066 Vss.t480 4.7885
R4654 Vss.n1828 Vss.t658 4.7885
R4655 Vss.n1837 Vss.t234 4.7885
R4656 Vss.n1172 Vss.t615 4.7885
R4657 Vss.n1158 Vss.t583 4.7885
R4658 Vss.n1050 Vss.t191 4.7885
R4659 Vss.n1078 Vss.t456 4.7885
R4660 Vss.n414 Vss.t91 4.7885
R4661 Vss.n1043 Vss.t167 4.7885
R4662 Vss.n1027 Vss.t428 4.7885
R4663 Vss.n488 Vss.t70 4.7885
R4664 Vss.n1088 Vss.t486 4.7885
R4665 Vss.n1135 Vss.t115 4.7885
R4666 Vss.n1522 Vss.t79 4.7885
R4667 Vss.n1111 Vss.t398 4.7885
R4668 Vss.n1105 Vss.t404 4.7885
R4669 Vss.n986 Vss.t537 4.7885
R4670 Vss.n977 Vss.t410 4.7885
R4671 Vss.n1003 Vss.t482 4.7885
R4672 Vss.n1096 Vss.t387 4.7885
R4673 Vss.n996 Vss.t490 4.7885
R4674 Vss.n1119 Vss.t619 4.7885
R4675 Vss.n474 Vss.t333 4.7885
R4676 Vss.n1127 Vss.t599 4.7885
R4677 Vss.n1143 Vss.t507 4.7885
R4678 Vss.n428 Vss.t148 4.7885
R4679 Vss.n456 Vss.t308 4.7885
R4680 Vss.n459 Vss.t76 4.7885
R4681 Vss.n1850 Vss.t310 4.7885
R4682 Vss.n1450 Vss.t96 4.7885
R4683 Vss.n1442 Vss.t226 4.7885
R4684 Vss.n50 Vss.t632 4.7885
R4685 Vss.n1436 Vss.t376 4.7885
R4686 Vss.n1282 Vss.t474 4.7885
R4687 Vss.n1346 Vss.t421 4.7885
R4688 Vss.n1277 Vss.t521 4.7885
R4689 Vss.n1307 Vss.t338 4.7885
R4690 Vss.n1314 Vss.t28 4.7885
R4691 Vss.n1316 Vss.t26 4.7885
R4692 Vss.n309 Vss.t211 4.7885
R4693 Vss.n308 Vss.t608 4.7885
R4694 Vss.n1479 Vss.t278 4.7885
R4695 Vss.n336 Vss.t209 4.7885
R4696 Vss.n1484 Vss.t170 4.7885
R4697 Vss.n327 Vss.t280 4.7885
R4698 Vss.n360 Vss.t462 4.7885
R4699 Vss.n344 Vss.t512 4.7885
R4700 Vss.n1216 Vss.t213 4.7885
R4701 Vss.n1201 Vss.t675 4.7885
R4702 Vss.n1196 Vss.t587 4.7885
R4703 Vss.n1189 Vss.t284 4.7885
R4704 Vss.n878 Vss.t21 4.7885
R4705 Vss.n884 Vss.t282 4.7885
R4706 Vss.n886 Vss.t286 4.7885
R4707 Vss.n918 Vss.t150 4.7885
R4708 Vss.n32 Vss.t575 4.7885
R4709 Vss.n33 Vss.t72 4.7885
R4710 Vss.n34 Vss.t74 4.7885
R4711 Vss.n792 Vss.t443 4.7885
R4712 Vss.n381 Vss.t138 4.7885
R4713 Vss.n302 Vss.t655 4.7885
R4714 Vss.n301 Vss.t543 4.7885
R4715 Vss.n300 Vss.t541 4.7885
R4716 Vss.n312 Vss.t553 4.7885
R4717 Vss.n1231 Vss.t274 4.7885
R4718 Vss.n1243 Vss.t47 4.7885
R4719 Vss.n1244 Vss.t62 4.7885
R4720 Vss.n1245 Vss.t64 4.7885
R4721 Vss.n1319 Vss.t560 4.7885
R4722 Vss.n1407 Vss.t133 4.7885
R4723 Vss.n200 Vss.t534 4.7885
R4724 Vss.n137 Vss.t373 4.7885
R4725 Vss.n112 Vss.t255 4.7885
R4726 Vss.n111 Vss.t99 4.7885
R4727 Vss.n1774 Vss.t106 4.7885
R4728 Vss.n1613 Vss.t345 4.7885
R4729 Vss.n1611 Vss.t163 4.7885
R4730 Vss.n97 Vss.t478 4.7885
R4731 Vss.n1635 Vss.t592 4.7885
R4732 Vss.n1628 Vss.t42 4.7885
R4733 Vss.n153 Vss.t318 4.7885
R4734 Vss.n1697 Vss.t228 4.7885
R4735 Vss.n158 Vss.t602 4.7885
R4736 Vss.n1703 Vss.t7 4.7885
R4737 Vss.n1786 Vss.t1 4.7885
R4738 Vss.n1761 Vss.t412 4.7885
R4739 Vss.n1756 Vss.t651 4.7885
R4740 Vss.n1790 Vss.t653 4.7885
R4741 Vss.n1779 Vss.t555 4.7885
R4742 Vss.n183 Vss.t363 4.7885
R4743 Vss.n1355 Vss.t215 4.7885
R4744 Vss.n1339 Vss.t526 4.7885
R4745 Vss.n1329 Vss.t24 4.7885
R4746 Vss.n1368 Vss.t155 4.7885
R4747 Vss.n1255 Vss.t378 4.7885
R4748 Vss.n205 Vss.t172 4.7885
R4749 Vss.n1803 Vss.t59 4.7885
R4750 Vss.n220 Vss.t501 4.7885
R4751 Vss.n214 Vss.t627 4.7885
R4752 Vss.n1053 Vss.t251 4.7885
R4753 Vss.n262 Vss.t519 4.7885
R4754 Vss.n68 Vss.t32 4.7885
R4755 Vss.n1659 Vss.t458 4.7885
R4756 Vss.n1671 Vss.t322 4.7885
R4757 Vss.n1532 Vss.t18 4.7885
R4758 Vss.n1528 Vss.t218 4.7885
R4759 Vss.n1541 Vss.t383 4.7885
R4760 Vss.n1656 Vss.t340 4.7885
R4761 Vss.n1378 Vss.t324 4.7885
R4762 Vss.n81 Vss.t152 4.7885
R4763 Vss.n1817 Vss.t261 4.7885
R4764 Vss.n129 Vss.t671 4.7885
R4765 Vss.n518 Vss.t664 4.7885
R4766 Vss.n959 Vss.t408 4.7885
R4767 Vss.n843 Vss.t517 4.7885
R4768 Vss.n951 Vss.t328 4.7885
R4769 Vss.n826 Vss.t484 4.7885
R4770 Vss.n636 Vss.t499 4.7885
R4771 Vss.n594 Vss.t496 4.7885
R4772 Vss.n551 Vss.t581 4.7885
R4773 Vss.n550 Vss.t389 4.7885
R4774 Vss.n736 Vss.t393 4.7885
R4775 Vss.n702 Vss.t645 4.7885
R4776 Vss.n695 Vss.t39 4.7885
R4777 Vss.n675 Vss.t124 4.7885
R4778 Vss.n684 Vss.t15 4.7885
R4779 Vss.n727 Vss.t612 4.7885
R4780 Vss.n722 Vss.t81 4.7885
R4781 Vss.n747 Vss.t83 4.7885
R4782 Vss.n743 Vss.t447 4.7885
R4783 Vss.n3 Vss.t201 4.7885
R4784 Vss.n537 Vss.t595 4.7885
R4785 Vss.n536 Vss.t265 4.7885
R4786 Vss.n786 Vss.t263 4.7885
R4787 Vss.n654 Vss.t515 4.7885
R4788 Vss.n646 Vss.t504 4.7885
R4789 Vss.n760 Vss.n0 4.28213
R4790 Vss.n631 Vss.n584 4.28213
R4791 Vss.n1879 Vss.n1878 4.28213
R4792 Vss.n991 Vss.n990 4.28213
R4793 Vss.n335 Vss.n334 4.28213
R4794 Vss.n1188 Vss.n1187 4.28213
R4795 Vss.n1328 Vss.n1266 4.28213
R4796 Vss.n1636 Vss.n160 4.28213
R4797 Vss.n1691 Vss.n1690 4.28213
R4798 Vss.n1730 Vss.n1729 4.28213
R4799 Vss.n207 Vss.n206 4.28213
R4800 Vss.n1531 Vss.n1526 4.28213
R4801 Vss.n1548 Vss.n1547 4.28213
R4802 Vss.n267 Vss.n65 4.28213
R4803 Vss.n1839 Vss.n1838 4.28213
R4804 Vss.n1118 Vss.n432 4.28213
R4805 Vss.n1137 Vss.n1136 4.28213
R4806 Vss.n1159 Vss.n1157 4.28213
R4807 Vss.n961 Vss.n960 4.28213
R4808 Vss.n1034 Vss.n1033 4.28213
R4809 Vss.n683 Vss.n682 4.28213
R4810 Vss.n1592 Vss.n1591 3.8722
R4811 Vss.n1571 Vss.n1565 3.52248
R4812 Vss.n1595 Vss.n1594 3.51469
R4813 Vss.n1469 Vss.n1468 3.51467
R4814 Vss.n1220 Vss.n1219 3.51467
R4815 Vss.n1867 Vss.n1866 3.51467
R4816 Vss.n1767 Vss.n1766 3.51467
R4817 Vss.n733 Vss.n732 3.51467
R4818 Vss.n1890 Vss.n1889 3.51467
R4819 Vss.n1574 Vss.t222 3.46717
R4820 Vss.t304 Vss.n1599 3.46717
R4821 Vss.n1575 Vss.t223 2.9111
R4822 Vss.n1598 Vss.t305 2.9111
R4823 Vss.n1351 Vss.n1350 2.45741
R4824 Vss.n1351 Vss.n1250 2.21573
R4825 Vss.n966 SARlogic_0.dffrs_12.nand3_6.B 2.17818
R4826 Vss.n1632 Vss.n100 2.06007
R4827 Vss.n1889 Vss.n6 2.06002
R4828 Vss.n1470 Vss.n1469 2.06002
R4829 Vss.n1219 Vss.n307 2.06002
R4830 Vss.n1868 Vss.n1867 2.06002
R4831 Vss.n1767 Vss.n113 2.06002
R4832 Vss.n733 Vss.n552 2.06002
R4833 Vss.n1568 Vss.t436 2.048
R4834 Vss.n1568 Vss.t400 2.048
R4835 Vss.n1558 Vss.t257 2.03874
R4836 Vss.n1558 Vss.t568 2.03874
R4837 Vss.n1559 Vss.t570 2.03874
R4838 Vss.n1559 Vss.t566 2.03874
R4839 Vss.n1148 Vss.n419 2.02164
R4840 Vss.n1099 Vss.n408 2.02164
R4841 Vss.n1163 Vss.n407 2.02164
R4842 Vss.n1653 Vss.n73 2.02164
R4843 Vss.n1820 Vss.n75 2.02164
R4844 Vss.n1446 Vss.n1445 2.02164
R4845 Vss.n1846 Vss.n48 2.02164
R4846 Vss.n1516 Vss.n1515 2.02164
R4847 Vss.n1683 Vss.n1682 2.02164
R4848 Vss.n973 Vss.n510 2.02164
R4849 Vss.n700 Vss.n561 1.92616
R4850 Vss.n531 Vss.n530 1.90702
R4851 Vss.n914 Vss.n28 1.90702
R4852 Vss.n1864 Vss.n30 1.90702
R4853 Vss.n1863 Vss.n31 1.90702
R4854 Vss.n795 Vss.n35 1.90702
R4855 Vss.n1858 Vss.n36 1.90702
R4856 Vss.n379 Vss.n306 1.90702
R4857 Vss.n1222 Vss.n304 1.90702
R4858 Vss.n1223 Vss.n303 1.90702
R4859 Vss.n315 Vss.n299 1.90702
R4860 Vss.n1228 Vss.n298 1.90702
R4861 Vss.n1235 Vss.n295 1.90702
R4862 Vss.n1466 Vss.n1241 1.90702
R4863 Vss.n1465 Vss.n1242 1.90702
R4864 Vss.n1321 Vss.n1246 1.90702
R4865 Vss.n1460 Vss.n1247 1.90702
R4866 Vss.n1405 Vss.n114 1.90702
R4867 Vss.n1763 Vss.n117 1.90702
R4868 Vss.n1778 Vss.n106 1.90702
R4869 Vss.n1787 Vss.n107 1.90702
R4870 Vss.n1764 Vss.n116 1.90702
R4871 Vss.n706 Vss.n553 1.90702
R4872 Vss.n730 Vss.n555 1.90702
R4873 Vss.n729 Vss.n556 1.90702
R4874 Vss.n744 Vss.n741 1.90702
R4875 Vss.n765 Vss.n2 1.90702
R4876 Vss.n1891 Vss.n4 1.90702
R4877 Vss.n776 Vss.n775 1.90702
R4878 Vss.n777 Vss.n538 1.90702
R4879 Vss.n783 Vss.n782 1.90702
R4880 Vss.n1582 Vss.n1569 1.73383
R4881 Vss.n1589 Vss.n1588 1.73383
R4882 Vss.n1574 Vss.n1556 1.70279
R4883 Vss.n1599 Vss.n1556 1.62925
R4884 Vss.n1617 Vss.n1552 1.62713
R4885 Vss.n1772 adc_PISO_0.2inmux_0.Bit 1.54251
R4886 Vss.n966 SARlogic_0.dffrs_12.nand3_1.A 1.34729
R4887 Vss.n628 Vss.n627 1.3005
R4888 Vss.n588 Vss.n587 1.3005
R4889 Vss.n626 Vss.n588 1.3005
R4890 Vss.n943 Vss.n396 1.3005
R4891 Vss.n942 Vss.n940 1.3005
R4892 Vss.n942 Vss.n941 1.3005
R4893 Vss.n1176 Vss.n1175 1.3005
R4894 Vss.n1172 Vss.n400 1.3005
R4895 Vss.n437 Vss.n400 1.3005
R4896 Vss.n1154 Vss.n1153 1.3005
R4897 Vss.n415 Vss.n414 1.3005
R4898 Vss.n1152 Vss.n415 1.3005
R4899 Vss.n1081 Vss.n1080 1.3005
R4900 Vss.n1079 Vss.n1078 1.3005
R4901 Vss.n1079 Vss.n417 1.3005
R4902 Vss.n1048 Vss.n1047 1.3005
R4903 Vss.n1050 Vss.n1049 1.3005
R4904 Vss.n1049 Vss.n418 1.3005
R4905 Vss.n1030 Vss.n499 1.3005
R4906 Vss.n1029 Vss.n1027 1.3005
R4907 Vss.n1029 Vss.n1028 1.3005
R4908 Vss.n1040 Vss.n498 1.3005
R4909 Vss.n1043 Vss.n1042 1.3005
R4910 Vss.n1042 Vss.n1041 1.3005
R4911 Vss.n986 Vss.n985 1.3005
R4912 Vss.n985 Vss.n483 1.3005
R4913 Vss.n984 Vss.n983 1.3005
R4914 Vss.n1003 Vss.n1002 1.3005
R4915 Vss.n1002 Vss.n1001 1.3005
R4916 Vss.n999 Vss.n500 1.3005
R4917 Vss.n1097 Vss.n1096 1.3005
R4918 Vss.n1098 Vss.n1097 1.3005
R4919 Vss.n501 Vss.n484 1.3005
R4920 Vss.n1124 Vss.n1123 1.3005
R4921 Vss.n475 Vss.n474 1.3005
R4922 Vss.n475 Vss.n250 1.3005
R4923 Vss.n1131 Vss.n1130 1.3005
R4924 Vss.n1127 Vss.n473 1.3005
R4925 Vss.n476 Vss.n473 1.3005
R4926 Vss.n1147 Vss.n1146 1.3005
R4927 Vss.n1143 Vss.n421 1.3005
R4928 Vss.n421 Vss.n420 1.3005
R4929 Vss.n426 Vss.n425 1.3005
R4930 Vss.n428 Vss.n427 1.3005
R4931 Vss.n427 Vss.n251 1.3005
R4932 Vss.n1117 Vss.n1116 1.3005
R4933 Vss.n1120 Vss.n1119 1.3005
R4934 Vss.n1121 Vss.n1120 1.3005
R4935 Vss.n979 Vss.n481 1.3005
R4936 Vss.n1105 Vss.n1104 1.3005
R4937 Vss.n1104 Vss.n1103 1.3005
R4938 Vss.n482 Vss.n478 1.3005
R4939 Vss.n1112 Vss.n1111 1.3005
R4940 Vss.n1113 Vss.n1112 1.3005
R4941 Vss.n1114 Vss.n249 1.3005
R4942 Vss.n1522 Vss.n1521 1.3005
R4943 Vss.n1521 Vss.n1520 1.3005
R4944 Vss.n1101 Vss.n436 1.3005
R4945 Vss.n1135 Vss.n1134 1.3005
R4946 Vss.n1134 Vss.n1133 1.3005
R4947 Vss.n1092 Vss.n1091 1.3005
R4948 Vss.n1089 Vss.n1088 1.3005
R4949 Vss.n1090 Vss.n1089 1.3005
R4950 Vss.n492 Vss.n491 1.3005
R4951 Vss.n489 Vss.n488 1.3005
R4952 Vss.n490 Vss.n489 1.3005
R4953 Vss.n453 Vss.n452 1.3005
R4954 Vss.n457 Vss.n456 1.3005
R4955 Vss.n458 Vss.n457 1.3005
R4956 Vss.n468 Vss.n467 1.3005
R4957 Vss.n461 Vss.n459 1.3005
R4958 Vss.n461 Vss.n460 1.3005
R4959 Vss.n1161 Vss.n1160 1.3005
R4960 Vss.n1158 Vss.n410 1.3005
R4961 Vss.n470 Vss.n410 1.3005
R4962 Vss.n450 Vss.n46 1.3005
R4963 Vss.n1850 Vss.n1849 1.3005
R4964 Vss.n1849 Vss.n1848 1.3005
R4965 Vss.n1425 Vss.n1423 1.3005
R4966 Vss.n1450 Vss.n1449 1.3005
R4967 Vss.n1449 Vss.n1448 1.3005
R4968 Vss.n1277 Vss.n1276 1.3005
R4969 Vss.n1276 Vss.n1275 1.3005
R4970 Vss.n1293 Vss.n1292 1.3005
R4971 Vss.n364 Vss.n363 1.3005
R4972 Vss.n360 Vss.n320 1.3005
R4973 Vss.n341 Vss.n320 1.3005
R4974 Vss.n355 Vss.n354 1.3005
R4975 Vss.n328 Vss.n327 1.3005
R4976 Vss.n328 Vss.n289 1.3005
R4977 Vss.n344 Vss.n343 1.3005
R4978 Vss.n343 Vss.n342 1.3005
R4979 Vss.n351 Vss.n350 1.3005
R4980 Vss.n339 Vss.n288 1.3005
R4981 Vss.n1479 Vss.n1478 1.3005
R4982 Vss.n1478 Vss.n1477 1.3005
R4983 Vss.n331 Vss.n330 1.3005
R4984 Vss.n337 Vss.n336 1.3005
R4985 Vss.n338 Vss.n337 1.3005
R4986 Vss.n1209 Vss.n308 1.3005
R4987 Vss.n1210 Vss.n1209 1.3005
R4988 Vss.n1206 Vss.n307 1.3005
R4989 Vss.n1211 Vss.n309 1.3005
R4990 Vss.n1212 Vss.n1211 1.3005
R4991 Vss.n1216 Vss.n1215 1.3005
R4992 Vss.n1215 Vss.n1214 1.3005
R4993 Vss.n1193 Vss.n390 1.3005
R4994 Vss.n1196 Vss.n1195 1.3005
R4995 Vss.n1195 Vss.n1194 1.3005
R4996 Vss.n1190 Vss.n1189 1.3005
R4997 Vss.n1191 Vss.n1190 1.3005
R4998 Vss.n1184 Vss.n1183 1.3005
R4999 Vss.n892 Vss.n34 1.3005
R5000 Vss.n140 Vss.n139 1.3005
R5001 Vss.n138 Vss.n137 1.3005
R5002 Vss.n138 Vss.n123 1.3005
R5003 Vss.n198 Vss.n197 1.3005
R5004 Vss.n200 Vss.n199 1.3005
R5005 Vss.n199 Vss.n124 1.3005
R5006 Vss.n1614 Vss.n1613 1.3005
R5007 Vss.n1615 Vss.n1614 1.3005
R5008 Vss.n1562 Vss.n1561 1.3005
R5009 Vss.n1611 Vss.n1610 1.3005
R5010 Vss.n1610 Vss.n1609 1.3005
R5011 Vss.n1797 Vss.n1796 1.3005
R5012 Vss.n98 Vss.n97 1.3005
R5013 Vss.n1795 Vss.n98 1.3005
R5014 Vss.n1627 Vss.n1626 1.3005
R5015 Vss.n1629 Vss.n1628 1.3005
R5016 Vss.n1630 Vss.n1629 1.3005
R5017 Vss.n158 Vss.n157 1.3005
R5018 Vss.n170 Vss.n157 1.3005
R5019 Vss.n1711 Vss.n1710 1.3005
R5020 Vss.n1786 Vss.n1785 1.3005
R5021 Vss.n1785 Vss.n1784 1.3005
R5022 Vss.n183 Vss.n182 1.3005
R5023 Vss.n182 Vss.n171 1.3005
R5024 Vss.n181 Vss.n180 1.3005
R5025 Vss.n1716 Vss.n1715 1.3005
R5026 Vss.n154 Vss.n153 1.3005
R5027 Vss.n1714 Vss.n154 1.3005
R5028 Vss.n172 Vss.n155 1.3005
R5029 Vss.n1698 Vss.n1697 1.3005
R5030 Vss.n1699 Vss.n1698 1.3005
R5031 Vss.n1638 Vss.n1637 1.3005
R5032 Vss.n1635 Vss.n1634 1.3005
R5033 Vss.n1634 Vss.n156 1.3005
R5034 Vss.n1761 Vss.n1760 1.3005
R5035 Vss.n1760 Vss.n1759 1.3005
R5036 Vss.n1757 Vss.n1756 1.3005
R5037 Vss.n1758 Vss.n1757 1.3005
R5038 Vss.n1791 Vss.n1790 1.3005
R5039 Vss.n1792 Vss.n1791 1.3005
R5040 Vss.n1778 Vss.n1777 1.3005
R5041 Vss.n1780 Vss.n1779 1.3005
R5042 Vss.n1781 Vss.n1780 1.3005
R5043 Vss.n1745 Vss.n113 1.3005
R5044 Vss.n1748 Vss.n112 1.3005
R5045 Vss.n1754 Vss.n111 1.3005
R5046 Vss.n1755 Vss.n1754 1.3005
R5047 Vss.n1775 Vss.n1774 1.3005
R5048 Vss.n1776 Vss.n1775 1.3005
R5049 Vss.n1741 Vss.n1740 1.3005
R5050 Vss.n1742 Vss.n1741 1.3005
R5051 Vss.n1743 Vss.n116 1.3005
R5052 Vss.n1285 Vss.n1273 1.3005
R5053 Vss.n1284 Vss.n1282 1.3005
R5054 Vss.n1284 Vss.n1283 1.3005
R5055 Vss.n1271 Vss.n1270 1.3005
R5056 Vss.n1346 Vss.n1345 1.3005
R5057 Vss.n1345 Vss.n1344 1.3005
R5058 Vss.n1471 Vss.n1470 1.3005
R5059 Vss.n1308 Vss.n1307 1.3005
R5060 Vss.n1309 Vss.n1308 1.3005
R5061 Vss.n1314 Vss.n1313 1.3005
R5062 Vss.n1313 Vss.n1310 1.3005
R5063 Vss.n1317 Vss.n1316 1.3005
R5064 Vss.n1318 Vss.n1317 1.3005
R5065 Vss.n1327 Vss.n1326 1.3005
R5066 Vss.n1330 Vss.n1329 1.3005
R5067 Vss.n1331 Vss.n1330 1.3005
R5068 Vss.n1334 Vss.n1333 1.3005
R5069 Vss.n1340 Vss.n1339 1.3005
R5070 Vss.n1341 Vss.n1340 1.3005
R5071 Vss.n1322 Vss.n1321 1.3005
R5072 Vss.n1320 Vss.n1319 1.3005
R5073 Vss.n1320 Vss.n1257 1.3005
R5074 Vss.n1261 Vss.n1260 1.3005
R5075 Vss.n1356 Vss.n1355 1.3005
R5076 Vss.n1357 Vss.n1356 1.3005
R5077 Vss.n1371 Vss.n1370 1.3005
R5078 Vss.n1369 Vss.n1368 1.3005
R5079 Vss.n1369 Vss.n1358 1.3005
R5080 Vss.n1417 Vss.n274 1.3005
R5081 Vss.n1416 Vss.n1255 1.3005
R5082 Vss.n1416 Vss.n1415 1.3005
R5083 Vss.n194 Vss.n87 1.3005
R5084 Vss.n215 Vss.n214 1.3005
R5085 Vss.n216 Vss.n215 1.3005
R5086 Vss.n217 Vss.n88 1.3005
R5087 Vss.n221 Vss.n220 1.3005
R5088 Vss.n222 Vss.n221 1.3005
R5089 Vss.n1807 Vss.n1806 1.3005
R5090 Vss.n1803 Vss.n89 1.3005
R5091 Vss.n223 Vss.n89 1.3005
R5092 Vss.n1825 Vss.n1824 1.3005
R5093 Vss.n69 Vss.n68 1.3005
R5094 Vss.n1823 Vss.n69 1.3005
R5095 Vss.n1504 Vss.n1503 1.3005
R5096 Vss.n263 Vss.n262 1.3005
R5097 Vss.n263 Vss.n71 1.3005
R5098 Vss.n1055 Vss.n264 1.3005
R5099 Vss.n1054 Vss.n1053 1.3005
R5100 Vss.n1054 Vss.n72 1.3005
R5101 Vss.n1537 Vss.n1536 1.3005
R5102 Vss.n1529 Vss.n1528 1.3005
R5103 Vss.n1529 Vss.n192 1.3005
R5104 Vss.n1500 Vss.n233 1.3005
R5105 Vss.n1656 Vss.n1655 1.3005
R5106 Vss.n1655 Vss.n1654 1.3005
R5107 Vss.n1544 Vss.n1543 1.3005
R5108 Vss.n1542 Vss.n1541 1.3005
R5109 Vss.n1542 Vss.n234 1.3005
R5110 Vss.n1530 Vss.n235 1.3005
R5111 Vss.n1533 Vss.n1532 1.3005
R5112 Vss.n1534 Vss.n1533 1.3005
R5113 Vss.n1663 Vss.n1662 1.3005
R5114 Vss.n1660 Vss.n1659 1.3005
R5115 Vss.n1661 Vss.n1660 1.3005
R5116 Vss.n1669 Vss.n1668 1.3005
R5117 Vss.n1671 Vss.n1670 1.3005
R5118 Vss.n1670 Vss.n193 1.3005
R5119 Vss.n1813 Vss.n1812 1.3005
R5120 Vss.n82 Vss.n81 1.3005
R5121 Vss.n1811 Vss.n82 1.3005
R5122 Vss.n1381 Vss.n84 1.3005
R5123 Vss.n1380 Vss.n1378 1.3005
R5124 Vss.n1380 Vss.n1379 1.3005
R5125 Vss.n203 Vss.n74 1.3005
R5126 Vss.n205 Vss.n204 1.3005
R5127 Vss.n204 Vss.n86 1.3005
R5128 Vss.n1242 Vss.n277 1.3005
R5129 Vss.n1301 Vss.n1243 1.3005
R5130 Vss.n1301 Vss.n1300 1.3005
R5131 Vss.n1305 Vss.n1244 1.3005
R5132 Vss.n1306 Vss.n1305 1.3005
R5133 Vss.n1303 Vss.n1245 1.3005
R5134 Vss.n1303 Vss.n1256 1.3005
R5135 Vss.n1818 Vss.n1817 1.3005
R5136 Vss.n1819 Vss.n1818 1.3005
R5137 Vss.n271 Vss.n76 1.3005
R5138 Vss.n1438 Vss.n1426 1.3005
R5139 Vss.n1437 Vss.n1436 1.3005
R5140 Vss.n1437 Vss.n273 1.3005
R5141 Vss.n316 Vss.n315 1.3005
R5142 Vss.n314 Vss.n312 1.3005
R5143 Vss.n314 Vss.n313 1.3005
R5144 Vss.n283 Vss.n282 1.3005
R5145 Vss.n1485 Vss.n1484 1.3005
R5146 Vss.n1486 Vss.n1485 1.3005
R5147 Vss.n298 Vss.n281 1.3005
R5148 Vss.n1232 Vss.n1231 1.3005
R5149 Vss.n1233 Vss.n1232 1.3005
R5150 Vss.n1235 Vss.n1234 1.3005
R5151 Vss.n1237 Vss.n1236 1.3005
R5152 Vss.n1238 Vss.n1237 1.3005
R5153 Vss.n1240 Vss.n297 1.3005
R5154 Vss.n1240 Vss.n1239 1.3005
R5155 Vss.n1241 Vss.n278 1.3005
R5156 Vss.n1845 Vss.n1844 1.3005
R5157 Vss.n50 Vss.n49 1.3005
R5158 Vss.n59 Vss.n49 1.3005
R5159 Vss.n1428 Vss.n1427 1.3005
R5160 Vss.n1443 Vss.n1442 1.3005
R5161 Vss.n1444 Vss.n1443 1.3005
R5162 Vss.n1149 Vss.n58 1.3005
R5163 Vss.n1837 Vss.n1836 1.3005
R5164 Vss.n1836 Vss.n1835 1.3005
R5165 Vss.n1832 Vss.n1831 1.3005
R5166 Vss.n1828 Vss.n64 1.3005
R5167 Vss.n1060 Vss.n64 1.3005
R5168 Vss.n1061 Vss.n63 1.3005
R5169 Vss.n1067 Vss.n1066 1.3005
R5170 Vss.n1068 Vss.n1067 1.3005
R5171 Vss.n1072 Vss.n62 1.3005
R5172 Vss.n1071 Vss.n1059 1.3005
R5173 Vss.n1071 Vss.n1070 1.3005
R5174 Vss.n266 Vss.n265 1.3005
R5175 Vss.n269 Vss.n268 1.3005
R5176 Vss.n270 Vss.n269 1.3005
R5177 Vss.n1514 Vss.n1513 1.3005
R5178 Vss.n1510 Vss.n253 1.3005
R5179 Vss.n1497 Vss.n253 1.3005
R5180 Vss.n1517 Vss.n244 1.3005
R5181 Vss.n1550 Vss.n1549 1.3005
R5182 Vss.n1551 Vss.n1550 1.3005
R5183 Vss.n1619 Vss.n1618 1.3005
R5184 Vss.n1621 Vss.n1620 1.3005
R5185 Vss.n1620 Vss.n236 1.3005
R5186 Vss.n1650 Vss.n1649 1.3005
R5187 Vss.n1646 Vss.n238 1.3005
R5188 Vss.n238 Vss.n237 1.3005
R5189 Vss.n1643 Vss.n191 1.3005
R5190 Vss.n1642 Vss.n1624 1.3005
R5191 Vss.n1642 Vss.n1641 1.3005
R5192 Vss.n1639 Vss.n167 1.3005
R5193 Vss.n1703 Vss.n1702 1.3005
R5194 Vss.n1702 Vss.n1701 1.3005
R5195 Vss.n1686 Vss.n189 1.3005
R5196 Vss.n1689 Vss.n1688 1.3005
R5197 Vss.n1688 Vss.n1687 1.3005
R5198 Vss.n1681 Vss.n1680 1.3005
R5199 Vss.n1677 Vss.n227 1.3005
R5200 Vss.n227 Vss.n146 1.3005
R5201 Vss.n1723 Vss.n1722 1.3005
R5202 Vss.n1719 Vss.n147 1.3005
R5203 Vss.n1631 Vss.n147 1.3005
R5204 Vss.n225 Vss.n143 1.3005
R5205 Vss.n1728 Vss.n1727 1.3005
R5206 Vss.n1727 Vss.n1726 1.3005
R5207 Vss.n1399 Vss.n1398 1.3005
R5208 Vss.n1395 Vss.n1361 1.3005
R5209 Vss.n1361 Vss.n1360 1.3005
R5210 Vss.n1390 Vss.n1389 1.3005
R5211 Vss.n1388 Vss.n1387 1.3005
R5212 Vss.n1388 Vss.n125 1.3005
R5213 Vss.n1410 Vss.n1247 1.3005
R5214 Vss.n1408 Vss.n1407 1.3005
R5215 Vss.n1409 Vss.n1408 1.3005
R5216 Vss.n1406 Vss.n1405 1.3005
R5217 Vss.n1404 Vss.n1403 1.3005
R5218 Vss.n1404 Vss.n127 1.3005
R5219 Vss.n129 Vss.n128 1.3005
R5220 Vss.n128 Vss.n126 1.3005
R5221 Vss.n1738 Vss.n1737 1.3005
R5222 Vss.n933 Vss.n932 1.3005
R5223 Vss.n930 Vss.n929 1.3005
R5224 Vss.n931 Vss.n930 1.3005
R5225 Vss.n406 Vss.n405 1.3005
R5226 Vss.n1166 Vss.n1165 1.3005
R5227 Vss.n1165 Vss.n1164 1.3005
R5228 Vss.n975 Vss.n503 1.3005
R5229 Vss.n1036 Vss.n1035 1.3005
R5230 Vss.n1037 Vss.n1036 1.3005
R5231 Vss.n993 Vss.n992 1.3005
R5232 Vss.n977 Vss.n976 1.3005
R5233 Vss.n980 Vss.n976 1.3005
R5234 Vss.n1015 Vss.n1014 1.3005
R5235 Vss.n996 Vss.n995 1.3005
R5236 Vss.n995 Vss.n994 1.3005
R5237 Vss.n522 Vss.n521 1.3005
R5238 Vss.n518 Vss.n517 1.3005
R5239 Vss.n517 Vss.n509 1.3005
R5240 Vss.n798 Vss.n516 1.3005
R5241 Vss.n959 Vss.n958 1.3005
R5242 Vss.n958 Vss.n957 1.3005
R5243 Vss.n523 Vss.n508 1.3005
R5244 Vss.n1019 Vss.n1018 1.3005
R5245 Vss.n1018 Vss.n1017 1.3005
R5246 Vss.n439 Vss.n303 1.3005
R5247 Vss.n447 Vss.n302 1.3005
R5248 Vss.n448 Vss.n447 1.3005
R5249 Vss.n441 Vss.n301 1.3005
R5250 Vss.n441 Vss.n368 1.3005
R5251 Vss.n444 Vss.n300 1.3005
R5252 Vss.n444 Vss.n443 1.3005
R5253 Vss.n386 Vss.n372 1.3005
R5254 Vss.n1202 Vss.n1201 1.3005
R5255 Vss.n1203 Vss.n1202 1.3005
R5256 Vss.n384 Vss.n36 1.3005
R5257 Vss.n382 Vss.n381 1.3005
R5258 Vss.n383 Vss.n382 1.3005
R5259 Vss.n380 Vss.n379 1.3005
R5260 Vss.n378 Vss.n373 1.3005
R5261 Vss.n378 Vss.n377 1.3005
R5262 Vss.n375 Vss.n374 1.3005
R5263 Vss.n376 Vss.n375 1.3005
R5264 Vss.n369 Vss.n304 1.3005
R5265 Vss.n843 Vss.n842 1.3005
R5266 Vss.n842 Vss.n841 1.3005
R5267 Vss.n873 Vss.n872 1.3005
R5268 Vss.n851 Vss.n850 1.3005
R5269 Vss.n854 Vss.n853 1.3005
R5270 Vss.n853 Vss.n852 1.3005
R5271 Vss.n861 Vss.n860 1.3005
R5272 Vss.n865 Vss.n864 1.3005
R5273 Vss.n864 Vss.n863 1.3005
R5274 Vss.n796 Vss.n795 1.3005
R5275 Vss.n794 Vss.n792 1.3005
R5276 Vss.n794 Vss.n793 1.3005
R5277 Vss.n954 Vss.n511 1.3005
R5278 Vss.n971 Vss.n970 1.3005
R5279 Vss.n972 Vss.n971 1.3005
R5280 Vss.n952 Vss.n951 1.3005
R5281 Vss.n953 Vss.n952 1.3005
R5282 Vss.n799 Vss.n525 1.3005
R5283 Vss.n826 Vss.n825 1.3005
R5284 Vss.n825 Vss.n800 1.3005
R5285 Vss.n824 Vss.n801 1.3005
R5286 Vss.n817 Vss.n816 1.3005
R5287 Vss.n815 Vss.n814 1.3005
R5288 Vss.n815 Vss.n805 1.3005
R5289 Vss.n834 Vss.n833 1.3005
R5290 Vss.n808 Vss.n807 1.3005
R5291 Vss.n807 Vss.n806 1.3005
R5292 Vss.n616 Vss.n6 1.3005
R5293 Vss.n614 Vss.n7 1.3005
R5294 Vss.n615 Vss.n614 1.3005
R5295 Vss.n12 Vss.n8 1.3005
R5296 Vss.n13 Vss.n12 1.3005
R5297 Vss.n1886 Vss.n1885 1.3005
R5298 Vss.n1885 Vss.n1884 1.3005
R5299 Vss.n640 Vss.n639 1.3005
R5300 Vss.n636 Vss.n577 1.3005
R5301 Vss.n590 Vss.n577 1.3005
R5302 Vss.n604 Vss.n603 1.3005
R5303 Vss.n609 Vss.n608 1.3005
R5304 Vss.n610 Vss.n609 1.3005
R5305 Vss.n594 Vss.n593 1.3005
R5306 Vss.n593 Vss.n592 1.3005
R5307 Vss.n600 Vss.n599 1.3005
R5308 Vss.n679 Vss.n678 1.3005
R5309 Vss.n676 Vss.n675 1.3005
R5310 Vss.n677 Vss.n676 1.3005
R5311 Vss.n574 Vss.n567 1.3005
R5312 Vss.n685 Vss.n684 1.3005
R5313 Vss.n686 Vss.n685 1.3005
R5314 Vss.n689 Vss.n565 1.3005
R5315 Vss.n695 Vss.n694 1.3005
R5316 Vss.n694 Vss.n693 1.3005
R5317 Vss.n690 Vss.n561 1.3005
R5318 Vss.n703 Vss.n702 1.3005
R5319 Vss.n704 Vss.n703 1.3005
R5320 Vss.n706 Vss.n705 1.3005
R5321 Vss.n708 Vss.n707 1.3005
R5322 Vss.n709 Vss.n708 1.3005
R5323 Vss.n711 Vss.n710 1.3005
R5324 Vss.n712 Vss.n711 1.3005
R5325 Vss.n713 Vss.n555 1.3005
R5326 Vss.n782 Vss.n14 1.3005
R5327 Vss.n781 Vss.n780 1.3005
R5328 Vss.n781 Vss.n533 1.3005
R5329 Vss.n900 Vss.n899 1.3005
R5330 Vss.n905 Vss.n904 1.3005
R5331 Vss.n906 Vss.n905 1.3005
R5332 Vss.n907 Vss.n531 1.3005
R5333 Vss.n918 Vss.n917 1.3005
R5334 Vss.n917 Vss.n916 1.3005
R5335 Vss.n915 Vss.n914 1.3005
R5336 Vss.n913 Vss.n908 1.3005
R5337 Vss.n913 Vss.n912 1.3005
R5338 Vss.n910 Vss.n909 1.3005
R5339 Vss.n911 Vss.n910 1.3005
R5340 Vss.n1881 Vss.n1880 1.3005
R5341 Vss.n18 Vss.n17 1.3005
R5342 Vss.n802 Vss.n17 1.3005
R5343 Vss.n803 Vss.n21 1.3005
R5344 Vss.n1874 Vss.n1873 1.3005
R5345 Vss.n1873 Vss.n1872 1.3005
R5346 Vss.n1869 Vss.n1868 1.3005
R5347 Vss.n879 Vss.n878 1.3005
R5348 Vss.n880 Vss.n879 1.3005
R5349 Vss.n884 Vss.n881 1.3005
R5350 Vss.n889 Vss.n881 1.3005
R5351 Vss.n887 Vss.n886 1.3005
R5352 Vss.n888 Vss.n887 1.3005
R5353 Vss.n691 Vss.n556 1.3005
R5354 Vss.n727 Vss.n726 1.3005
R5355 Vss.n726 Vss.n725 1.3005
R5356 Vss.n723 Vss.n722 1.3005
R5357 Vss.n724 Vss.n723 1.3005
R5358 Vss.n748 Vss.n747 1.3005
R5359 Vss.n749 Vss.n748 1.3005
R5360 Vss.n756 Vss.n538 1.3005
R5361 Vss.n754 Vss.n537 1.3005
R5362 Vss.n755 Vss.n754 1.3005
R5363 Vss.n750 Vss.n536 1.3005
R5364 Vss.n751 Vss.n750 1.3005
R5365 Vss.n787 Vss.n786 1.3005
R5366 Vss.n788 Vss.n787 1.3005
R5367 Vss.n897 Vss.n31 1.3005
R5368 Vss.n895 Vss.n32 1.3005
R5369 Vss.n896 Vss.n895 1.3005
R5370 Vss.n790 Vss.n33 1.3005
R5371 Vss.n890 Vss.n790 1.3005
R5372 Vss.n741 Vss.n740 1.3005
R5373 Vss.n743 Vss.n742 1.3005
R5374 Vss.n742 Vss.n541 1.3005
R5375 Vss.n759 Vss.n758 1.3005
R5376 Vss.n762 Vss.n761 1.3005
R5377 Vss.n763 Vss.n762 1.3005
R5378 Vss.n765 Vss.n764 1.3005
R5379 Vss.n766 Vss.n3 1.3005
R5380 Vss.n767 Vss.n766 1.3005
R5381 Vss.n768 Vss.n4 1.3005
R5382 Vss.n772 Vss.n771 1.3005
R5383 Vss.n773 Vss.n772 1.3005
R5384 Vss.n769 Vss.n539 1.3005
R5385 Vss.n774 Vss.n539 1.3005
R5386 Vss.n618 Vss.n617 1.3005
R5387 Vss.n620 Vss.n619 1.3005
R5388 Vss.n621 Vss.n620 1.3005
R5389 Vss.n718 Vss.n552 1.3005
R5390 Vss.n716 Vss.n551 1.3005
R5391 Vss.n717 Vss.n716 1.3005
R5392 Vss.n559 Vss.n550 1.3005
R5393 Vss.n721 Vss.n559 1.3005
R5394 Vss.n737 Vss.n736 1.3005
R5395 Vss.n738 Vss.n737 1.3005
R5396 Vss.n652 Vss.n651 1.3005
R5397 Vss.n654 Vss.n653 1.3005
R5398 Vss.n653 Vss.n573 1.3005
R5399 Vss.n666 Vss.n572 1.3005
R5400 Vss.n669 Vss.n668 1.3005
R5401 Vss.n668 Vss.n667 1.3005
R5402 Vss.n646 Vss.n645 1.3005
R5403 Vss.n645 Vss.n644 1.3005
R5404 Vss.n662 Vss.n661 1.3005
R5405 Vss.n1612 Vss.n1556 1.29323
R5406 Vss.n1613 Vss.n1612 1.00923
R5407 Vss.n1593 Vss.n1592 0.999917
R5408 Vss.n1580 Vss.n1565 0.999917
R5409 Vss.n1580 Vss.n1579 0.999917
R5410 Vss.n1594 Vss.n1593 0.999917
R5411 Vss.n784 Vss.n530 0.990409
R5412 Vss.n1859 Vss.n1858 0.990409
R5413 Vss.n1228 Vss.n1227 0.990409
R5414 Vss.n1461 Vss.n1460 0.990409
R5415 Vss.n745 Vss.n2 0.990409
R5416 Vss.n1612 Vss.n1611 0.984484
R5417 Vss.n1591 Vss.n1563 0.949529
R5418 Vss.n670 Vss.n571 0.92075
R5419 Vss.n607 Vss.n605 0.92075
R5420 Vss.n629 Vss.n586 0.92075
R5421 Vss.n832 Vss.n809 0.92075
R5422 Vss.n903 Vss.n901 0.92075
R5423 Vss.n1876 Vss.n1875 0.92075
R5424 Vss.n969 Vss.n512 0.92075
R5425 Vss.n866 Vss.n859 0.92075
R5426 Vss.n944 Vss.n939 0.92075
R5427 Vss.n1020 Vss.n507 0.92075
R5428 Vss.n1168 Vss.n1167 0.92075
R5429 Vss.n1391 Vss.n1386 0.92075
R5430 Vss.n1397 Vss.n1396 0.92075
R5431 Vss.n1721 Vss.n1720 0.92075
R5432 Vss.n1679 Vss.n1678 0.92075
R5433 Vss.n1644 Vss.n166 0.92075
R5434 Vss.n1648 Vss.n1647 0.92075
R5435 Vss.n1622 Vss.n240 0.92075
R5436 Vss.n1512 Vss.n1511 0.92075
R5437 Vss.n1073 Vss.n1058 0.92075
R5438 Vss.n1065 Vss.n1063 0.92075
R5439 Vss.n1830 Vss.n1829 0.92075
R5440 Vss.n1174 Vss.n1173 0.92075
R5441 Vss.n1051 Vss.n1046 0.92075
R5442 Vss.n1082 Vss.n1077 0.92075
R5443 Vss.n1155 Vss.n413 0.92075
R5444 Vss.n1044 Vss.n497 0.92075
R5445 Vss.n1031 Vss.n411 0.92075
R5446 Vss.n493 Vss.n487 0.92075
R5447 Vss.n1093 Vss.n1087 0.92075
R5448 Vss.n1523 Vss.n248 0.92075
R5449 Vss.n1110 Vss.n1108 0.92075
R5450 Vss.n988 Vss.n987 0.92075
R5451 Vss.n1005 Vss.n1004 0.92075
R5452 Vss.n1095 Vss.n485 0.92075
R5453 Vss.n1013 Vss.n997 0.92075
R5454 Vss.n1106 Vss.n480 0.92075
R5455 Vss.n1125 Vss.n246 0.92075
R5456 Vss.n1129 Vss.n1128 0.92075
R5457 Vss.n430 Vss.n429 0.92075
R5458 Vss.n1145 Vss.n1144 0.92075
R5459 Vss.n466 Vss.n52 0.92075
R5460 Vss.n1851 Vss.n45 0.92075
R5461 Vss.n455 Vss.n454 0.92075
R5462 Vss.n1441 Vss.n1430 0.92075
R5463 Vss.n1843 Vss.n51 0.92075
R5464 Vss.n1451 Vss.n1422 0.92075
R5465 Vss.n1347 Vss.n1269 0.92075
R5466 Vss.n1291 Vss.n1278 0.92075
R5467 Vss.n1483 Vss.n284 0.92075
R5468 Vss.n356 Vss.n326 0.92075
R5469 Vss.n362 Vss.n361 0.92075
R5470 Vss.n349 Vss.n345 0.92075
R5471 Vss.n1480 Vss.n287 0.92075
R5472 Vss.n1200 Vss.n387 0.92075
R5473 Vss.n1197 Vss.n389 0.92075
R5474 Vss.n201 Vss.n196 0.92075
R5475 Vss.n141 Vss.n136 0.92075
R5476 Vss.n1798 Vss.n96 0.92075
R5477 Vss.n1625 Vss.n161 0.92075
R5478 Vss.n1696 Vss.n173 0.92075
R5479 Vss.n1709 Vss.n159 0.92075
R5480 Vss.n1705 Vss.n1704 0.92075
R5481 Vss.n184 Vss.n179 0.92075
R5482 Vss.n1717 Vss.n152 0.92075
R5483 Vss.n1354 Vss.n1262 0.92075
R5484 Vss.n1338 Vss.n1337 0.92075
R5485 Vss.n1286 Vss.n1281 0.92075
R5486 Vss.n1372 Vss.n1367 0.92075
R5487 Vss.n1418 Vss.n1254 0.92075
R5488 Vss.n1805 Vss.n1804 0.92075
R5489 Vss.n219 Vss.n218 0.92075
R5490 Vss.n213 Vss.n195 0.92075
R5491 Vss.n1056 Vss.n1052 0.92075
R5492 Vss.n1505 Vss.n261 0.92075
R5493 Vss.n1826 Vss.n67 0.92075
R5494 Vss.n1673 Vss.n1672 0.92075
R5495 Vss.n1664 Vss.n1658 0.92075
R5496 Vss.n1538 Vss.n1527 0.92075
R5497 Vss.n1545 Vss.n1540 0.92075
R5498 Vss.n1657 Vss.n232 0.92075
R5499 Vss.n1382 Vss.n1377 0.92075
R5500 Vss.n1814 Vss.n80 0.92075
R5501 Vss.n1816 Vss.n77 0.92075
R5502 Vss.n1439 Vss.n1435 0.92075
R5503 Vss.n1736 Vss.n130 0.92075
R5504 Vss.n934 Vss.n928 0.92075
R5505 Vss.n520 Vss.n519 0.92075
R5506 Vss.n871 Vss.n844 0.92075
R5507 Vss.n855 Vss.n849 0.92075
R5508 Vss.n950 Vss.n526 0.92075
R5509 Vss.n827 Vss.n823 0.92075
R5510 Vss.n818 Vss.n813 0.92075
R5511 Vss.n638 Vss.n637 0.92075
R5512 Vss.n598 Vss.n595 0.92075
R5513 Vss.n696 Vss.n564 0.92075
R5514 Vss.n680 Vss.n674 0.92075
R5515 Vss.n655 Vss.n650 0.92075
R5516 Vss.n660 Vss.n647 0.92075
R5517 Vss.n1578 Vss.n1563 0.907842
R5518 Vss.n1584 Vss.n1583 0.867167
R5519 Vss.t435 Vss.n1586 0.867167
R5520 Vss.n1587 Vss.n1564 0.867167
R5521 SARlogic_0.dffrs_12.d SARlogic_0.dffrs_12.nand3_8.A 0.784786
R5522 SARlogic_0.dffrs_13.d SARlogic_0.dffrs_13.nand3_8.A 0.784786
R5523 Vss.n202 Vss.n95 0.780467
R5524 Vss.n1887 Vss.n1886 0.771017
R5525 Vss.n1316 Vss.n1315 0.771017
R5526 Vss.n1217 Vss.n1216 0.771017
R5527 Vss.n886 Vss.n885 0.771017
R5528 Vss.n736 Vss.n735 0.771017
R5529 adc_PISO_0.avss Vss.n1787 0.762138
R5530 Vss.n1573 Vss.n1 0.714636
R5531 Vss.n1787 Vss.n1786 0.679217
R5532 Vss.n1229 Vss.n41 0.669813
R5533 Vss.n1857 Vss.n1856 0.669683
R5534 Vss.n921 Vss.n920 0.669683
R5535 Vss.n1591 comparator_no_offsetcal_0.no_offsetLatch_0.VSS 0.664071
R5536 Vss.n1894 Vss.n1893 0.651683
R5537 Vss.n739 Vss.n545 0.63255
R5538 SARlogic_0.dffrs_12.clk Vss.n966 0.611214
R5539 Vss.n700 Vss.n699 0.601415
R5540 Vss.n1459 Vss.n1458 0.600912
R5541 Vss.n1774 Vss.n1773 0.471317
R5542 Vss.n783 Vss.n780 0.463217
R5543 Vss.n1888 Vss.n7 0.463217
R5544 Vss.n1887 Vss.n8 0.463217
R5545 Vss.n1307 Vss.n294 0.463217
R5546 Vss.n1315 Vss.n1314 0.463217
R5547 Vss.n1217 Vss.n309 0.463217
R5548 Vss.n1218 Vss.n308 0.463217
R5549 Vss.n878 Vss.n27 0.463217
R5550 Vss.n885 Vss.n884 0.463217
R5551 Vss.n919 Vss.n918 0.463217
R5552 Vss.n1862 Vss.n32 0.463217
R5553 Vss.n1861 Vss.n33 0.463217
R5554 Vss.n1860 Vss.n34 0.463217
R5555 Vss.n792 Vss.n35 0.463217
R5556 Vss.n381 Vss.n37 0.463217
R5557 Vss.n1224 Vss.n302 0.463217
R5558 Vss.n1225 Vss.n301 0.463217
R5559 Vss.n1226 Vss.n300 0.463217
R5560 Vss.n312 Vss.n299 0.463217
R5561 Vss.n1231 Vss.n1230 0.463217
R5562 Vss.n1464 Vss.n1243 0.463217
R5563 Vss.n1463 Vss.n1244 0.463217
R5564 Vss.n1462 Vss.n1245 0.463217
R5565 Vss.n1319 Vss.n1246 0.463217
R5566 Vss.n1407 Vss.n1248 0.463217
R5567 Vss.n1768 Vss.n112 0.463217
R5568 Vss.n1769 Vss.n111 0.463217
R5569 Vss.n1762 Vss.n1761 0.463217
R5570 Vss.n1756 Vss.n105 0.463217
R5571 Vss.n1790 Vss.n1789 0.463217
R5572 Vss.n1779 Vss.n106 0.463217
R5573 Vss.n734 Vss.n551 0.463217
R5574 Vss.n735 Vss.n550 0.463217
R5575 Vss.n702 Vss.n701 0.463217
R5576 Vss.n728 Vss.n727 0.463217
R5577 Vss.n722 Vss.n544 0.463217
R5578 Vss.n747 Vss.n746 0.463217
R5579 Vss.n744 Vss.n743 0.463217
R5580 Vss.n1892 Vss.n3 0.463217
R5581 Vss.n778 Vss.n537 0.463217
R5582 Vss.n779 Vss.n536 0.463217
R5583 Vss.n786 Vss.n785 0.463217
R5584 Vss.n925 Vss.n39 0.441453
R5585 Vss.n1597 comparator_no_offsetcal_0.VSS 0.404079
R5586 Vss.n699 Vss.n1 0.328611
R5587 Vss.n1888 Vss.n1887 0.3083
R5588 Vss.n1315 Vss.n294 0.3083
R5589 Vss.n1218 Vss.n1217 0.3083
R5590 Vss.n885 Vss.n27 0.3083
R5591 Vss.n1862 Vss.n1861 0.3083
R5592 Vss.n1861 Vss.n1860 0.3083
R5593 Vss.n1225 Vss.n1224 0.3083
R5594 Vss.n1226 Vss.n1225 0.3083
R5595 Vss.n1464 Vss.n1463 0.3083
R5596 Vss.n1463 Vss.n1462 0.3083
R5597 Vss.n1769 Vss.n1768 0.3083
R5598 Vss.n1762 Vss.n105 0.3083
R5599 Vss.n1789 Vss.n105 0.3083
R5600 Vss.n735 Vss.n734 0.3083
R5601 Vss.n728 Vss.n544 0.3083
R5602 Vss.n746 Vss.n544 0.3083
R5603 Vss.n779 Vss.n778 0.3083
R5604 Vss.n785 Vss.n779 0.3083
R5605 Vss.n1773 Vss.n1769 0.3002
R5606 Vss.n922 Vss.n921 0.284919
R5607 Vss.n1771 Vss.n1770 0.252687
R5608 Vss.n1597 Vss.n1596 0.238053
R5609 Vss.n1863 Vss.n1862 0.2165
R5610 Vss.n1224 Vss.n1223 0.2165
R5611 Vss.n1465 Vss.n1464 0.2165
R5612 Vss.n1763 Vss.n1762 0.2165
R5613 Vss.n729 Vss.n728 0.2165
R5614 Vss.n778 Vss.n777 0.2165
R5615 Vss.n1577 Vss.n1576 0.211763
R5616 Vss.n937 Vss.n925 0.195855
R5617 comparator_no_offsetcal_0.x5.avss Vss.n1575 0.188808
R5618 Vss.n1598 comparator_no_offsetcal_0.x3.avss 0.188808
R5619 Vss.n1860 Vss.n1859 0.1748
R5620 Vss.n1462 Vss.n1461 0.1748
R5621 Vss.n746 Vss.n745 0.1748
R5622 Vss.n785 Vss.n784 0.1748
R5623 Vss.n1227 Vss.n1226 0.17465
R5624 Vss.n1596 Vss.n1563 0.163684
R5625 comparator_no_offsetcal_0.no_offsetLatch_0.VSS Vss.n1590 0.1605
R5626 Vss.n1789 Vss.n1788 0.1598
R5627 Vss.n1605 Vss.n1604 0.154786
R5628 Vss.n1788 Vss.n106 0.152487
R5629 Vss.n1864 Vss.n1863 0.148459
R5630 Vss.n1223 Vss.n1222 0.148459
R5631 Vss.n1466 Vss.n1465 0.148459
R5632 Vss.n1764 Vss.n1763 0.148459
R5633 Vss.n730 Vss.n729 0.148459
R5634 Vss.n777 Vss.n776 0.148459
R5635 Vss.n1855 Vss.n1854 0.145432
R5636 Vss.n1455 Vss.n1454 0.145432
R5637 Vss.n211 Vss.n133 0.143322
R5638 Vss.n937 Vss.n936 0.140365
R5639 Vss.n1227 Vss.n299 0.13865
R5640 Vss.n1859 Vss.n35 0.1385
R5641 Vss.n1461 Vss.n1246 0.1385
R5642 Vss.n745 Vss.n744 0.1385
R5643 Vss.n784 Vss.n783 0.1385
R5644 Vss.n1456 Vss.n1455 0.136253
R5645 Vss.n1601 Vss.n1560 0.1355
R5646 Vss.n1575 Vss.n1574 0.128901
R5647 Vss.n1599 Vss.n1598 0.127885
R5648 Vss.n946 Vss.n528 0.122607
R5649 Vss.n1007 Vss.n998 0.122607
R5650 Vss.n1289 Vss.n1288 0.122607
R5651 Vss.n323 Vss.n322 0.122607
R5652 Vss.n847 Vss.n845 0.122607
R5653 Vss.n821 Vss.n820 0.122607
R5654 Vss.n581 Vss.n579 0.122607
R5655 Vss.n658 Vss.n648 0.122607
R5656 Vss.n936 Vss.n935 0.118169
R5657 Vss.n1707 Vss.n163 0.115241
R5658 Vss.n1578 Vss.n1577 0.112526
R5659 Vss.n1607 Vss.n1606 0.109786
R5660 Vss.n1854 Vss.n41 0.104592
R5661 Vss.n632 Vss.n582 0.10457
R5662 Vss.n346 Vss.n286 0.10457
R5663 Vss.n868 Vss.n388 0.10457
R5664 Vss.n1694 Vss.n1693 0.10457
R5665 Vss.n1733 Vss.n1732 0.10457
R5666 Vss.n829 Vss.n19 0.10457
R5667 Vss.n673 Vss.n672 0.10457
R5668 SARlogic_0.dffrs_14.vss Vss.n1801 0.102612
R5669 SARlogic_0.dffrs_8.vss Vss.n258 0.102537
R5670 SARlogic_0.dffrs_10.vss Vss.n495 0.102537
R5671 Vss.n259 SARlogic_0.dffrs_7.vss 0.101537
R5672 Vss.n1075 SARlogic_0.dffrs_9.vss 0.101537
R5673 Vss.n1856 Vss.n1855 0.0911096
R5674 Vss.n967 Vss.n963 0.078611
R5675 Vss.n935 Vss.n927 0.0781858
R5676 Vss.n1455 Vss.n1251 0.0776599
R5677 Vss.n1454 Vss.n1453 0.0776599
R5678 Vss.n1855 Vss.n40 0.0776599
R5679 Vss.n1854 Vss.n1853 0.0776599
R5680 Vss.n1865 Vss.n29 0.073981
R5681 Vss.n1221 Vss.n305 0.073981
R5682 Vss.n1467 Vss.n296 0.073981
R5683 Vss.n1765 Vss.n115 0.073981
R5684 Vss.n731 Vss.n554 0.073981
R5685 Vss.n770 Vss.n5 0.073981
R5686 Vss.n1877 Vss.n20 0.0679983
R5687 Vss.n333 Vss.n332 0.0679983
R5688 Vss.n1186 Vss.n1185 0.0679983
R5689 Vss.n1336 Vss.n1335 0.0679983
R5690 Vss.n681 Vss.n562 0.0679983
R5691 Vss.n285 Vss.n41 0.0673674
R5692 Vss.n1856 Vss.n38 0.0673025
R5693 Vss.n921 Vss.n529 0.0673025
R5694 Vss.n1350 Vss.n1349 0.0665049
R5695 Vss.n1026 Vss.n1023 0.0660086
R5696 Vss.n1026 Vss.n1025 0.0655096
R5697 Vss.n989 Vss.n978 0.0645882
R5698 Vss.n515 Vss.n506 0.0645882
R5699 Vss.n1889 Vss.n1888 0.0635
R5700 Vss.n1469 Vss.n294 0.0635
R5701 Vss.n1219 Vss.n1218 0.0635
R5702 Vss.n1867 Vss.n27 0.0635
R5703 Vss.n1768 Vss.n1767 0.0635
R5704 Vss.n734 Vss.n733 0.0635
R5705 Vss.n150 Vss.n149 0.0625376
R5706 Vss.n648 Vss.n568 0.0622481
R5707 Vss.n820 Vss.n811 0.0622481
R5708 Vss.n1009 Vss.n998 0.0622481
R5709 Vss.n324 Vss.n323 0.0622481
R5710 Vss.n847 Vss.n846 0.0622481
R5711 Vss.n1288 Vss.n1265 0.0622481
R5712 Vss.n528 Vss.n514 0.0622481
R5713 Vss.n633 Vss.n581 0.0622481
R5714 Vss.n1675 Vss.n93 0.0616538
R5715 Vss.n1253 Vss.n78 0.0616538
R5716 Vss.n260 Vss.n231 0.0616538
R5717 Vss.n1064 Vss.n255 0.0616538
R5718 Vss.n1452 Vss.n1421 0.0616538
R5719 Vss.n1852 Vss.n44 0.0616538
R5720 Vss.n1076 Vss.n423 0.0616538
R5721 Vss.n1000 Vss.n486 0.0616538
R5722 Vss.n1171 Vss.n1170 0.0616538
R5723 Vss.n1385 Vss.n1363 0.0615256
R5724 Vss.n1894 Vss.n1 0.0600636
R5725 Vss.n1482 Vss.n1481 0.0568904
R5726 Vss.n1199 Vss.n1198 0.0568904
R5727 Vss.n902 Vss.n22 0.0568904
R5728 Vss.n697 Vss.n563 0.0568904
R5729 Vss.n1350 Vss.n1264 0.0566774
R5730 Vss.n1458 Vss.n1457 0.0561349
R5731 Vss.n923 Vss.n922 0.0551896
R5732 Vss.n937 Vss.n513 0.0551896
R5733 Vss.n632 Vss.n583 0.054837
R5734 Vss.n1481 Vss.n286 0.054837
R5735 Vss.n1198 Vss.n388 0.054837
R5736 Vss.n1693 Vss.n163 0.054837
R5737 Vss.n1732 Vss.n133 0.054837
R5738 Vss.n22 Vss.n19 0.054837
R5739 Vss.n673 Vss.n563 0.054837
R5740 Vss.n1856 Vss.n39 0.0521009
R5741 Vss.n585 Vss.n583 0.0502328
R5742 Vss.n1458 Vss.n1249 0.0480028
R5743 Vss.n1075 Vss.n424 0.0478478
R5744 Vss.n462 Vss.n40 0.0478478
R5745 Vss.n1853 Vss.n43 0.0478478
R5746 Vss.n177 Vss.n95 0.0478478
R5747 Vss.n259 Vss.n229 0.0478478
R5748 Vss.n1365 Vss.n131 0.0478478
R5749 Vss.n1801 Vss.n1800 0.0478478
R5750 Vss.n1374 Vss.n1251 0.0478478
R5751 Vss.n1453 Vss.n1420 0.0478478
R5752 Vss.n1507 Vss.n258 0.0478478
R5753 Vss.n1084 Vss.n495 0.0478478
R5754 Vss.n925 Vss.n924 0.0478478
R5755 Vss.n585 Vss.n0 0.0467
R5756 Vss.n347 Vss.n346 0.0466843
R5757 Vss.n1694 Vss.n185 0.0466843
R5758 Vss.n1734 Vss.n1733 0.0466843
R5759 Vss.n869 Vss.n868 0.0466843
R5760 Vss.n829 Vss.n828 0.0466843
R5761 Vss.n596 Vss.n582 0.0466843
R5762 Vss.n672 Vss.n569 0.0466843
R5763 Vss.n938 Vss.n923 0.0465106
R5764 Vss.n968 Vss.n513 0.0465106
R5765 Vss.n963 Vss.n505 0.0465106
R5766 Vss.n209 Vss.n208 0.0465022
R5767 Vss.n1827 Vss.n66 0.0465022
R5768 Vss.n496 Vss.n57 0.0465022
R5769 Vss.n1156 Vss.n412 0.0465022
R5770 Vss.n212 Vss.n211 0.0464521
R5771 Vss.n1606 Vss.n1605 0.0455
R5772 Vss.n811 Vss.n19 0.0415307
R5773 Vss.n1009 Vss.n433 0.0415307
R5774 Vss.n324 Vss.n286 0.0415307
R5775 Vss.n846 Vss.n388 0.0415307
R5776 Vss.n1350 Vss.n1265 0.0415307
R5777 Vss.n962 Vss.n514 0.0415307
R5778 Vss.n633 Vss.n632 0.0415307
R5779 Vss.n673 Vss.n568 0.0415307
R5780 Vss.n1454 Vss.n41 0.0413406
R5781 Vss.n1012 Vss.n1011 0.0405109
R5782 Vss.n1290 Vss.n1267 0.0405109
R5783 Vss.n348 Vss.n347 0.0405109
R5784 Vss.n359 Vss.n321 0.0405109
R5785 Vss.n357 Vss.n325 0.0405109
R5786 Vss.n185 Vss.n178 0.0405109
R5787 Vss.n1695 Vss.n174 0.0405109
R5788 Vss.n1287 Vss.n1280 0.0405109
R5789 Vss.n1348 Vss.n1268 0.0405109
R5790 Vss.n1735 Vss.n1734 0.0405109
R5791 Vss.n1392 Vss.n132 0.0405109
R5792 Vss.n870 Vss.n869 0.0405109
R5793 Vss.n856 Vss.n848 0.0405109
R5794 Vss.n867 Vss.n858 0.0405109
R5795 Vss.n949 Vss.n527 0.0405109
R5796 Vss.n828 Vss.n822 0.0405109
R5797 Vss.n819 Vss.n812 0.0405109
R5798 Vss.n831 Vss.n830 0.0405109
R5799 Vss.n597 Vss.n596 0.0405109
R5800 Vss.n635 Vss.n578 0.0405109
R5801 Vss.n606 Vss.n580 0.0405109
R5802 Vss.n659 Vss.n569 0.0405109
R5803 Vss.n656 Vss.n649 0.0405109
R5804 Vss.n671 Vss.n570 0.0405109
R5805 Vss.n927 Vss.n504 0.040346
R5806 Vss.n1865 Vss.n1864 0.0389018
R5807 Vss.n1222 Vss.n1221 0.0389018
R5808 Vss.n1467 Vss.n1466 0.0389018
R5809 Vss.n1765 Vss.n1764 0.0389018
R5810 Vss.n731 Vss.n730 0.0389018
R5811 Vss.n776 Vss.n5 0.0389018
R5812 Vss.n1708 Vss.n1707 0.0368083
R5813 Vss.n188 Vss.n162 0.036505
R5814 Vss.n1539 Vss.n239 0.036505
R5815 Vss.n1546 Vss.n1525 0.036505
R5816 Vss.n1126 Vss.n247 0.036505
R5817 Vss.n479 Vss.n435 0.036505
R5818 Vss.n1142 Vss.n423 0.0361576
R5819 Vss.n1170 Vss.n402 0.0361576
R5820 Vss.n53 Vss.n44 0.0361576
R5821 Vss.n175 Vss.n150 0.0361576
R5822 Vss.n231 Vss.n230 0.0361576
R5823 Vss.n1434 Vss.n1421 0.0361576
R5824 Vss.n1394 Vss.n1385 0.0361576
R5825 Vss.n1676 Vss.n1675 0.0361576
R5826 Vss.n1364 Vss.n78 0.0361576
R5827 Vss.n1509 Vss.n255 0.0361576
R5828 Vss.n1086 Vss.n486 0.0361576
R5829 Vss.n936 Vss.n926 0.0361576
R5830 Vss.n332 Vss.n285 0.035635
R5831 Vss.n1185 Vss.n38 0.035635
R5832 Vss.n529 Vss.n20 0.035635
R5833 Vss.n698 Vss.n562 0.035635
R5834 Vss.n699 Vss.n698 0.0352182
R5835 Vss.n1878 Vss.n19 0.0349747
R5836 Vss.n990 Vss.n433 0.0349747
R5837 Vss.n334 Vss.n286 0.0349747
R5838 Vss.n1187 Vss.n388 0.0349747
R5839 Vss.n1350 Vss.n1266 0.0349747
R5840 Vss.n962 Vss.n961 0.0349747
R5841 Vss.n632 Vss.n631 0.0349747
R5842 Vss.n682 Vss.n673 0.0349747
R5843 Vss.n1335 Vss.n1263 0.0346145
R5844 Vss.n1718 Vss.n150 0.0340549
R5845 Vss.n1033 Vss.n504 0.0339793
R5846 Vss.n1675 Vss.n228 0.0335769
R5847 Vss.n1366 Vss.n1363 0.0335769
R5848 Vss.n1253 Vss.n1251 0.0335769
R5849 Vss.n1815 Vss.n78 0.0335769
R5850 Vss.n1665 Vss.n231 0.0335769
R5851 Vss.n255 Vss.n254 0.0335769
R5852 Vss.n1453 Vss.n1452 0.0335769
R5853 Vss.n1440 Vss.n1421 0.0335769
R5854 Vss.n1853 Vss.n1852 0.0335769
R5855 Vss.n1842 Vss.n44 0.0335769
R5856 Vss.n423 Vss.n422 0.0335769
R5857 Vss.n1094 Vss.n486 0.0335769
R5858 Vss.n1171 Vss.n40 0.0335769
R5859 Vss.n1170 Vss.n403 0.0335769
R5860 Vss.n1384 Vss.n1362 0.0334487
R5861 Vss.n811 Vss.n810 0.0322085
R5862 Vss.n948 Vss.n946 0.0322085
R5863 Vss.n1085 Vss.n434 0.0322085
R5864 Vss.n1508 Vss.n256 0.0322085
R5865 Vss.n187 Vss.n94 0.0322085
R5866 Vss.n1141 Vss.n424 0.0322085
R5867 Vss.n1010 Vss.n1007 0.0322085
R5868 Vss.n1010 Vss.n1009 0.0322085
R5869 Vss.n464 Vss.n462 0.0322085
R5870 Vss.n464 Vss.n463 0.0322085
R5871 Vss.n54 Vss.n43 0.0322085
R5872 Vss.n1289 Vss.n1279 0.0322085
R5873 Vss.n358 Vss.n322 0.0322085
R5874 Vss.n358 Vss.n324 0.0322085
R5875 Vss.n857 Vss.n846 0.0322085
R5876 Vss.n177 Vss.n176 0.0322085
R5877 Vss.n1279 Vss.n1265 0.0322085
R5878 Vss.n1667 Vss.n229 0.0322085
R5879 Vss.n1433 Vss.n1420 0.0322085
R5880 Vss.n1433 Vss.n1431 0.0322085
R5881 Vss.n1393 Vss.n131 0.0322085
R5882 Vss.n1393 Vss.n134 0.0322085
R5883 Vss.n176 Vss.n151 0.0322085
R5884 Vss.n1800 Vss.n94 0.0322085
R5885 Vss.n1375 Vss.n1374 0.0322085
R5886 Vss.n1375 Vss.n79 0.0322085
R5887 Vss.n1667 Vss.n1666 0.0322085
R5888 Vss.n1508 Vss.n1507 0.0322085
R5889 Vss.n1841 Vss.n54 0.0322085
R5890 Vss.n1141 Vss.n1140 0.0322085
R5891 Vss.n1085 Vss.n1084 0.0322085
R5892 Vss.n924 Vss.n404 0.0322085
R5893 Vss.n927 Vss.n404 0.0322085
R5894 Vss.n857 Vss.n845 0.0322085
R5895 Vss.n948 Vss.n514 0.0322085
R5896 Vss.n821 Vss.n810 0.0322085
R5897 Vss.n634 Vss.n579 0.0322085
R5898 Vss.n634 Vss.n633 0.0322085
R5899 Vss.n658 Vss.n657 0.0322085
R5900 Vss.n657 Vss.n568 0.0322085
R5901 Vss.n1457 Vss.n1250 0.0317776
R5902 Vss.n938 Vss.n937 0.0308765
R5903 Vss.n1457 Vss.n1456 0.0306923
R5904 Vss.n945 Vss.n923 0.0268641
R5905 Vss.n1062 Vss.n258 0.0268641
R5906 Vss.n1006 Vss.n495 0.0268641
R5907 Vss.n1008 Vss.n486 0.0268641
R5908 Vss.n431 Vss.n255 0.0268641
R5909 Vss.n1853 Vss.n42 0.0268641
R5910 Vss.n465 Vss.n44 0.0268641
R5911 Vss.n1429 Vss.n1421 0.0268641
R5912 Vss.n1453 Vss.n1252 0.0268641
R5913 Vss.n1801 Vss.n92 0.0268641
R5914 Vss.n1675 Vss.n1674 0.0268641
R5915 Vss.n1432 Vss.n78 0.0268641
R5916 Vss.n150 Vss.n148 0.0268641
R5917 Vss.n1799 Vss.n95 0.0268641
R5918 Vss.n1384 Vss.n1383 0.0268641
R5919 Vss.n1373 Vss.n1366 0.0268641
R5920 Vss.n1419 Vss.n1251 0.0268641
R5921 Vss.n257 Vss.n231 0.0268641
R5922 Vss.n1506 Vss.n259 0.0268641
R5923 Vss.n494 Vss.n423 0.0268641
R5924 Vss.n1083 Vss.n1075 0.0268641
R5925 Vss.n401 Vss.n40 0.0268641
R5926 Vss.n1170 Vss.n1169 0.0268641
R5927 Vss.n947 Vss.n513 0.0268641
R5928 Vss.n211 Vss.n202 0.0263346
R5929 Vss.n908 Vss.n29 0.0258591
R5930 Vss.n909 Vss.n29 0.0258591
R5931 Vss.n373 Vss.n305 0.0258591
R5932 Vss.n374 Vss.n305 0.0258591
R5933 Vss.n1236 Vss.n296 0.0258591
R5934 Vss.n297 Vss.n296 0.0258591
R5935 Vss.n1403 Vss.n115 0.0258591
R5936 Vss.n1740 Vss.n115 0.0258591
R5937 Vss.n707 Vss.n554 0.0258591
R5938 Vss.n710 Vss.n554 0.0258591
R5939 Vss.n771 Vss.n770 0.0258591
R5940 Vss.n770 Vss.n769 0.0258591
R5941 Vss.n1693 Vss.n151 0.0237454
R5942 Vss.n1692 Vss.n187 0.0235512
R5943 Vss.n1732 Vss.n134 0.0235512
R5944 Vss.n135 Vss.n79 0.0235512
R5945 Vss.n1666 Vss.n186 0.0235512
R5946 Vss.n256 Vss.n245 0.0235512
R5947 Vss.n1431 Vss.n56 0.0235512
R5948 Vss.n1841 Vss.n1840 0.0235512
R5949 Vss.n1140 Vss.n1139 0.0235512
R5950 Vss.n1138 Vss.n434 0.0235512
R5951 Vss.n463 Vss.n55 0.0235512
R5952 Vss.n630 Vss.n585 0.0232899
R5953 Vss.n1866 Vss.n1865 0.023066
R5954 Vss.n1221 Vss.n1220 0.023066
R5955 Vss.n1468 Vss.n1467 0.023066
R5956 Vss.n1766 Vss.n1765 0.023066
R5957 Vss.n732 Vss.n731 0.023066
R5958 Vss.n1890 Vss.n5 0.023066
R5959 Vss.n1718 Vss.n151 0.0226532
R5960 Vss.n963 Vss.n962 0.0225109
R5961 Vss.n504 Vss.n55 0.0225109
R5962 Vss.n1840 Vss.n55 0.0225109
R5963 Vss.n1840 Vss.n56 0.0225109
R5964 Vss.n135 Vss.n56 0.0225109
R5965 Vss.n1731 Vss.n135 0.0225109
R5966 Vss.n1693 Vss.n1692 0.0225109
R5967 Vss.n1692 Vss.n186 0.0225109
R5968 Vss.n245 Vss.n186 0.0225109
R5969 Vss.n1139 Vss.n245 0.0225109
R5970 Vss.n1139 Vss.n1138 0.0225109
R5971 Vss.n1138 Vss.n433 0.0225109
R5972 Vss.n479 Vss.n247 0.0223682
R5973 Vss.n1525 Vss.n247 0.0223682
R5974 Vss.n1525 Vss.n239 0.0223682
R5975 Vss.n239 Vss.n162 0.0223682
R5976 Vss.n1707 Vss.n162 0.0223682
R5977 Vss.n978 Vss.n479 0.0223682
R5978 Vss.n1023 Vss.n506 0.0223682
R5979 Vss.n228 Vss.n187 0.0223376
R5980 Vss.n1815 Vss.n79 0.0223376
R5981 Vss.n1666 Vss.n1665 0.0223376
R5982 Vss.n256 Vss.n254 0.0223376
R5983 Vss.n1440 Vss.n1431 0.0223376
R5984 Vss.n1842 Vss.n1841 0.0223376
R5985 Vss.n1140 Vss.n422 0.0223376
R5986 Vss.n1094 Vss.n434 0.0223376
R5987 Vss.n463 Vss.n403 0.0223376
R5988 Vss.n1376 Vss.n134 0.0222094
R5989 Vss.n1581 Vss.n1580 0.0215413
R5990 Vss.n1593 Vss.n1566 0.0215413
R5991 Vss.n946 Vss.n945 0.0214837
R5992 Vss.n1062 Vss.n424 0.0214837
R5993 Vss.n1007 Vss.n1006 0.0214837
R5994 Vss.n1010 Vss.n1008 0.0214837
R5995 Vss.n1141 Vss.n431 0.0214837
R5996 Vss.n462 Vss.n42 0.0214837
R5997 Vss.n465 Vss.n464 0.0214837
R5998 Vss.n1429 Vss.n54 0.0214837
R5999 Vss.n1252 Vss.n43 0.0214837
R6000 Vss.n1290 Vss.n1289 0.0214837
R6001 Vss.n348 Vss.n322 0.0214837
R6002 Vss.n358 Vss.n357 0.0214837
R6003 Vss.n178 Vss.n177 0.0214837
R6004 Vss.n176 Vss.n174 0.0214837
R6005 Vss.n1279 Vss.n1268 0.0214837
R6006 Vss.n229 Vss.n92 0.0214837
R6007 Vss.n1674 Vss.n1667 0.0214837
R6008 Vss.n1433 Vss.n1432 0.0214837
R6009 Vss.n1735 Vss.n131 0.0214837
R6010 Vss.n1393 Vss.n1392 0.0214837
R6011 Vss.n148 Vss.n94 0.0214837
R6012 Vss.n1800 Vss.n1799 0.0214837
R6013 Vss.n1383 Vss.n1375 0.0214837
R6014 Vss.n1374 Vss.n1373 0.0214837
R6015 Vss.n1420 Vss.n1419 0.0214837
R6016 Vss.n1508 Vss.n257 0.0214837
R6017 Vss.n1507 Vss.n1506 0.0214837
R6018 Vss.n1085 Vss.n494 0.0214837
R6019 Vss.n1084 Vss.n1083 0.0214837
R6020 Vss.n924 Vss.n401 0.0214837
R6021 Vss.n1169 Vss.n404 0.0214837
R6022 Vss.n870 Vss.n845 0.0214837
R6023 Vss.n858 Vss.n857 0.0214837
R6024 Vss.n948 Vss.n947 0.0214837
R6025 Vss.n822 Vss.n821 0.0214837
R6026 Vss.n831 Vss.n810 0.0214837
R6027 Vss.n597 Vss.n579 0.0214837
R6028 Vss.n634 Vss.n580 0.0214837
R6029 Vss.n659 Vss.n658 0.0214837
R6030 Vss.n657 Vss.n570 0.0214837
R6031 Vss.n1026 Vss.n505 0.0204141
R6032 Vss.n1693 Vss.n160 0.0200312
R6033 Vss.n1707 Vss.n1706 0.0199048
R6034 Vss.n1692 Vss.n1691 0.019868
R6035 Vss.n207 Vss.n135 0.019868
R6036 Vss.n1526 Vss.n186 0.019868
R6037 Vss.n1547 Vss.n245 0.019868
R6038 Vss.n65 Vss.n56 0.019868
R6039 Vss.n1840 Vss.n1839 0.019868
R6040 Vss.n1139 Vss.n432 0.019868
R6041 Vss.n1138 Vss.n1137 0.019868
R6042 Vss.n1157 Vss.n55 0.019868
R6043 Vss.n1731 Vss.n1730 0.0197929
R6044 Vss.n1604 Vss.n1560 0.0197857
R6045 Vss.n1645 Vss.n162 0.0197428
R6046 Vss.n1623 Vss.n239 0.0197428
R6047 Vss.n1525 Vss.n1524 0.0197428
R6048 Vss.n1109 Vss.n247 0.0197428
R6049 Vss.n1107 Vss.n479 0.0197428
R6050 Vss.n920 Vss.n530 0.0196349
R6051 Vss.n1858 Vss.n1857 0.0196349
R6052 Vss.n1229 Vss.n1228 0.0196349
R6053 Vss.n1460 Vss.n1459 0.0196349
R6054 Vss.n1893 Vss.n2 0.0196349
R6055 adc_PISO_0.dffrs_4.vss Vss.n1894 0.0170545
R6056 Vss.n1025 Vss.n1024 0.0164817
R6057 Vss.n1866 Vss.n28 0.0163358
R6058 Vss.n1220 Vss.n306 0.0163358
R6059 Vss.n1468 Vss.n295 0.0163358
R6060 Vss.n1766 Vss.n114 0.0163358
R6061 Vss.n732 Vss.n553 0.0163358
R6062 Vss.n1891 Vss.n1890 0.0163358
R6063 Vss.n1025 Vss.n412 0.0157888
R6064 Vss.n496 Vss.n412 0.0157888
R6065 Vss.n496 Vss.n66 0.0157888
R6066 Vss.n209 Vss.n66 0.0157888
R6067 Vss.n210 Vss.n209 0.0157888
R6068 Vss.n1032 Vss.n1026 0.0150091
R6069 Vss.n149 Vss.n95 0.0142428
R6070 Vss.n1801 Vss.n93 0.014047
R6071 Vss.n260 Vss.n259 0.014047
R6072 Vss.n1064 Vss.n258 0.014047
R6073 Vss.n1076 Vss.n1075 0.014047
R6074 Vss.n1000 Vss.n495 0.014047
R6075 Vss.n919 Vss.n28 0.0139604
R6076 Vss.n306 Vss.n37 0.0139604
R6077 Vss.n1230 Vss.n295 0.0139604
R6078 Vss.n1248 Vss.n114 0.0139604
R6079 Vss.n701 Vss.n553 0.0139604
R6080 Vss.n1892 Vss.n1891 0.0139604
R6081 Vss.n920 Vss.n919 0.0130367
R6082 Vss.n1857 Vss.n37 0.0130367
R6083 Vss.n1230 Vss.n1229 0.0130367
R6084 Vss.n1459 Vss.n1248 0.0130367
R6085 Vss.n701 Vss.n700 0.0130367
R6086 Vss.n1893 Vss.n1892 0.0130367
R6087 Vss.n1011 Vss.n1010 0.0121902
R6088 Vss.n1142 Vss.n1141 0.0121902
R6089 Vss.n464 Vss.n402 0.0121902
R6090 Vss.n54 Vss.n53 0.0121902
R6091 Vss.n359 Vss.n358 0.0121902
R6092 Vss.n176 Vss.n175 0.0121902
R6093 Vss.n1280 Vss.n1279 0.0121902
R6094 Vss.n1667 Vss.n230 0.0121902
R6095 Vss.n1434 Vss.n1433 0.0121902
R6096 Vss.n1394 Vss.n1393 0.0121902
R6097 Vss.n1676 Vss.n94 0.0121902
R6098 Vss.n1375 Vss.n1364 0.0121902
R6099 Vss.n1509 Vss.n1508 0.0121902
R6100 Vss.n1086 Vss.n1085 0.0121902
R6101 Vss.n926 Vss.n404 0.0121902
R6102 Vss.n857 Vss.n856 0.0121902
R6103 Vss.n949 Vss.n948 0.0121902
R6104 Vss.n812 Vss.n810 0.0121902
R6105 Vss.n635 Vss.n634 0.0121902
R6106 Vss.n657 Vss.n656 0.0121902
R6107 Vss.n1788 adc_PISO_0.avss 0.0118245
R6108 Vss.n1352 Vss.n1264 0.0110968
R6109 Vss.n1707 Vss.n165 0.0102582
R6110 Vss.n209 Vss.n90 0.00974555
R6111 Vss.n1057 Vss.n66 0.00974555
R6112 Vss.n1074 Vss.n496 0.00974555
R6113 Vss.n1045 Vss.n412 0.00974555
R6114 Vss.n1456 Vss.n1249 0.00967928
R6115 Vss.n210 Vss.n91 0.00967038
R6116 Vss.n1012 Vss.n998 0.00915761
R6117 Vss.n323 Vss.n321 0.00915761
R6118 Vss.n1288 Vss.n1287 0.00915761
R6119 Vss.n848 Vss.n847 0.00915761
R6120 Vss.n528 Vss.n527 0.00915761
R6121 Vss.n820 Vss.n819 0.00915761
R6122 Vss.n581 Vss.n578 0.00915761
R6123 Vss.n649 Vss.n648 0.00915761
R6124 Vss.n1263 Vss.n1250 0.00760526
R6125 Vss.n968 Vss.n967 0.00745509
R6126 Vss.n1024 SARlogic_0.dffrs_11.vss 0.00734312
R6127 Vss.n346 Vss.n325 0.00720109
R6128 Vss.n1695 Vss.n1694 0.00720109
R6129 Vss.n1733 Vss.n132 0.00720109
R6130 Vss.n868 Vss.n867 0.00720109
R6131 Vss.n830 Vss.n829 0.00720109
R6132 Vss.n606 Vss.n582 0.00720109
R6133 Vss.n672 Vss.n671 0.00720109
R6134 Vss.n1023 Vss.n1022 0.00638507
R6135 Vss.n1349 Vss.n1267 0.00617391
R6136 Vss.n1349 Vss.n1348 0.00617391
R6137 Vss.n1353 Vss.n1263 0.00613715
R6138 Vss.n1353 Vss.n1352 0.00613715
R6139 Vss.n1573 Vss 0.00568182
R6140 Vss.n1482 Vss.n285 0.00511663
R6141 Vss.n1199 Vss.n38 0.00511663
R6142 Vss.n902 Vss.n529 0.00511663
R6143 Vss.n698 Vss.n697 0.00511663
R6144 adc_PISO_0.dffrs_4.vss Vss.n0 0.00480909
R6145 Vss.n922 Vss.n39 0.00478552
R6146 SARlogic_0.dffrs_7.vss Vss.n90 0.0044588
R6147 Vss.n1057 SARlogic_0.dffrs_8.vss 0.0044588
R6148 SARlogic_0.dffrs_9.vss Vss.n1074 0.0044588
R6149 Vss.n1045 SARlogic_0.dffrs_10.vss 0.0044588
R6150 Vss.n1802 SARlogic_0.dffrs_14.vss 0.00438363
R6151 Vss.n1607 comparator_no_offsetcal_0.x4.VSS 0.00371429
R6152 Vss.n1352 Vss.n1351 0.00175057
R6153 Vss.n1385 Vss.n1384 0.000628205
R6154 Vss.n1376 Vss.n1362 0.000628205
R6155 Vss.n1732 Vss.n1731 0.000575167
R6156 Vss.n212 Vss.n142 0.000575167
R6157 Vss.n1802 Vss.n91 0.000575167
R6158 Vss.n211 Vss.n210 0.000550111
R6159 Vss.n1878 Vss.n1877 0.000544599
R6160 Vss.n990 Vss.n989 0.000544599
R6161 Vss.n334 Vss.n333 0.000544599
R6162 Vss.n1187 Vss.n1186 0.000544599
R6163 Vss.n1336 Vss.n1266 0.000544599
R6164 Vss.n961 Vss.n515 0.000544599
R6165 Vss.n631 Vss.n630 0.000544599
R6166 Vss.n682 Vss.n681 0.000544599
R6167 Vss.n1033 Vss.n1032 0.000543311
R6168 Vss.n1366 Vss.n1365 0.000542735
R6169 Vss.n1708 Vss.n160 0.000525267
R6170 Vss.n1691 Vss.n188 0.000525056
R6171 Vss.n1730 Vss.n142 0.000525056
R6172 Vss.n208 Vss.n207 0.000525056
R6173 Vss.n1539 Vss.n1526 0.000525056
R6174 Vss.n1547 Vss.n1546 0.000525056
R6175 Vss.n1827 Vss.n65 0.000525056
R6176 Vss.n1839 Vss.n57 0.000525056
R6177 Vss.n1126 Vss.n432 0.000525056
R6178 Vss.n1137 Vss.n435 0.000525056
R6179 Vss.n1157 Vss.n1156 0.000525056
R6180 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t4 41.0041
R6181 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t9 40.8177
R6182 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t8 40.6313
R6183 SARlogic_0.dffrs_12.nand3_6.C.n3 SARlogic_0.dffrs_12.nand3_6.C.t7 27.3166
R6184 SARlogic_0.dffrs_12.nand3_6.C.n0 SARlogic_0.dffrs_12.nand3_6.C.t5 27.1302
R6185 SARlogic_0.dffrs_12.nand3_6.C.n1 SARlogic_0.dffrs_12.nand3_6.C.t6 26.9438
R6186 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.t1 10.0473
R6187 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n4 9.90747
R6188 SARlogic_0.dffrs_12.nand3_6.C.n5 SARlogic_0.dffrs_12.nand3_6.C.n2 9.90116
R6189 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.t2 6.51042
R6190 SARlogic_0.dffrs_12.nand3_6.C.n8 SARlogic_0.dffrs_12.nand3_6.C.n7 6.04952
R6191 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_6.C.n1 5.7305
R6192 SARlogic_0.dffrs_12.nand3_2.B SARlogic_0.dffrs_12.nand3_6.C.n0 5.47979
R6193 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C.n3 5.13907
R6194 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n9 4.72925
R6195 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_6.C.n5 4.5005
R6196 SARlogic_0.dffrs_12.nand3_6.C.n9 SARlogic_0.dffrs_12.nand3_6.C.n8 0.732092
R6197 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t3 0.7285
R6198 SARlogic_0.dffrs_12.nand3_6.C.n7 SARlogic_0.dffrs_12.nand3_6.C.t0 0.7285
R6199 SARlogic_0.dffrs_12.nand3_1.Z SARlogic_0.dffrs_12.nand3_6.C.n6 0.449758
R6200 SARlogic_0.dffrs_12.nand3_6.C.n6 SARlogic_0.dffrs_12.nand3_2.B 0.166901
R6201 SARlogic_0.dffrs_12.nand3_6.C.n2 SARlogic_0.dffrs_12.nand3_0.A 0.0455
R6202 SARlogic_0.dffrs_12.nand3_6.C.n4 SARlogic_0.dffrs_12.nand3_6.C 0.0455
R6203 inv2_0.out.n30 inv2_0.out.t25 34.2529
R6204 inv2_0.out.n24 inv2_0.out.t8 34.2529
R6205 inv2_0.out.n18 inv2_0.out.t13 34.2529
R6206 inv2_0.out.n12 inv2_0.out.t21 34.2529
R6207 inv2_0.out.n6 inv2_0.out.t15 34.2529
R6208 inv2_0.out.n1 inv2_0.out.t28 34.2529
R6209 inv2_0.out.n32 inv2_0.out.t20 34.1797
R6210 inv2_0.out.n26 inv2_0.out.t22 34.1797
R6211 inv2_0.out.n20 inv2_0.out.t17 34.1797
R6212 inv2_0.out.n14 inv2_0.out.t5 34.1797
R6213 inv2_0.out.n8 inv2_0.out.t24 34.1797
R6214 inv2_0.out.n3 inv2_0.out.t7 34.1797
R6215 inv2_0.out.n29 inv2_0.out.t31 19.673
R6216 inv2_0.out.n23 inv2_0.out.t11 19.673
R6217 inv2_0.out.n17 inv2_0.out.t12 19.673
R6218 inv2_0.out.n11 inv2_0.out.t27 19.673
R6219 inv2_0.out.n5 inv2_0.out.t19 19.673
R6220 inv2_0.out.n0 inv2_0.out.t2 19.673
R6221 inv2_0.out.n32 inv2_0.out.t9 19.5798
R6222 inv2_0.out.n26 inv2_0.out.t14 19.5798
R6223 inv2_0.out.n20 inv2_0.out.t6 19.5798
R6224 inv2_0.out.n14 inv2_0.out.t26 19.5798
R6225 inv2_0.out.n8 inv2_0.out.t16 19.5798
R6226 inv2_0.out.n3 inv2_0.out.t30 19.5798
R6227 inv2_0.out.n29 inv2_0.out.t18 19.4007
R6228 inv2_0.out.n23 inv2_0.out.t29 19.4007
R6229 inv2_0.out.n17 inv2_0.out.t3 19.4007
R6230 inv2_0.out.n11 inv2_0.out.t10 19.4007
R6231 inv2_0.out.n5 inv2_0.out.t4 19.4007
R6232 inv2_0.out.n0 inv2_0.out.t23 19.4007
R6233 inv2_0.out.n10 inv2_0.out.n4 15.5531
R6234 inv2_0.out.n36 inv2_0.out.t0 9.6935
R6235 inv2_0.out.n34 inv2_0.out.n33 8.46371
R6236 inv2_0.out.n22 inv2_0.out.n21 8.37371
R6237 inv2_0.out.n28 inv2_0.out.n27 8.32871
R6238 inv2_0.out.n16 inv2_0.out.n15 8.32871
R6239 inv2_0.out.n10 inv2_0.out.n9 8.32871
R6240 inv2_0.out.n31 inv2_0.out.n30 7.87164
R6241 inv2_0.out.n25 inv2_0.out.n24 7.87164
R6242 inv2_0.out.n19 inv2_0.out.n18 7.87164
R6243 inv2_0.out.n13 inv2_0.out.n12 7.87164
R6244 inv2_0.out.n7 inv2_0.out.n6 7.87164
R6245 inv2_0.out.n2 inv2_0.out.n1 7.87164
R6246 inv2_0.out.n34 inv2_0.out.n28 7.26762
R6247 inv2_0.out.n16 inv2_0.out.n10 7.22491
R6248 inv2_0.out.n22 inv2_0.out.n16 7.22491
R6249 inv2_0.out.n28 inv2_0.out.n22 7.22491
R6250 inv2_0.out.n33 inv2_0.out.n32 5.00771
R6251 inv2_0.out.n21 inv2_0.out.n20 5.00771
R6252 inv2_0.out.n27 inv2_0.out.n26 4.96432
R6253 inv2_0.out.n15 inv2_0.out.n14 4.96432
R6254 inv2_0.out.n9 inv2_0.out.n8 4.96432
R6255 inv2_0.out.n4 inv2_0.out.n3 4.96432
R6256 inv2_0.out inv2_0.out.n35 4.85086
R6257 inv2_0.out.n36 inv2_0.out.t1 4.35383
R6258 inv2_0.out.n27 inv2_0.out.n25 2.11068
R6259 inv2_0.out.n15 inv2_0.out.n13 2.11068
R6260 inv2_0.out.n9 inv2_0.out.n7 2.11068
R6261 inv2_0.out.n4 inv2_0.out.n2 2.11068
R6262 inv2_0.out.n33 inv2_0.out.n31 2.06729
R6263 inv2_0.out.n21 inv2_0.out.n19 2.06729
R6264 inv2_0.out inv2_0.out.n36 0.254429
R6265 inv2_0.out.n31 adc_PISO_0.2inmux_0.Load 0.2255
R6266 inv2_0.out.n25 adc_PISO_0.2inmux_2.Load 0.2255
R6267 inv2_0.out.n19 adc_PISO_0.2inmux_3.Load 0.2255
R6268 inv2_0.out.n13 adc_PISO_0.2inmux_4.Load 0.2255
R6269 inv2_0.out.n7 adc_PISO_0.2inmux_5.Load 0.2255
R6270 inv2_0.out.n2 adc_PISO_0.2inmux_1.Load 0.2255
R6271 inv2_0.out.n35 inv2_0.out.n34 0.182025
R6272 inv2_0.out.n30 inv2_0.out.n29 0.106438
R6273 inv2_0.out.n24 inv2_0.out.n23 0.106438
R6274 inv2_0.out.n18 inv2_0.out.n17 0.106438
R6275 inv2_0.out.n12 inv2_0.out.n11 0.106438
R6276 inv2_0.out.n6 inv2_0.out.n5 0.106438
R6277 inv2_0.out.n1 inv2_0.out.n0 0.106438
R6278 inv2_0.out.n35 adc_PISO_0.load 0.0294831
R6279 a_37499_31160.n0 a_37499_31160.t5 34.1797
R6280 a_37499_31160.n0 a_37499_31160.t4 19.5798
R6281 a_37499_31160.n1 a_37499_31160.t2 18.7717
R6282 a_37499_31160.n1 a_37499_31160.t1 9.2885
R6283 a_37499_31160.n2 a_37499_31160.n0 4.93379
R6284 a_37499_31160.t0 a_37499_31160.n3 4.23346
R6285 a_37499_31160.n3 a_37499_31160.t3 3.85546
R6286 a_37499_31160.n2 a_37499_31160.n1 0.4055
R6287 a_37499_31160.n3 a_37499_31160.n2 0.352625
R6288 a_n9429_n2007.n18 a_n9429_n2007.n17 11.2899
R6289 a_n9429_n2007.n17 a_n9429_n2007.n16 8.49339
R6290 a_n9429_n2007.n10 a_n9429_n2007.n9 4.89725
R6291 a_n9429_n2007.n14 a_n9429_n2007.n2 4.89725
R6292 a_n9429_n2007.n13 a_n9429_n2007.n3 4.89725
R6293 a_n9429_n2007.n12 a_n9429_n2007.n5 4.89725
R6294 a_n9429_n2007.n11 a_n9429_n2007.n7 4.89725
R6295 a_n9429_n2007.n13 a_n9429_n2007.n4 4.88712
R6296 a_n9429_n2007.n12 a_n9429_n2007.n6 4.88712
R6297 a_n9429_n2007.n11 a_n9429_n2007.n8 4.88712
R6298 a_n9429_n2007.n1 a_n9429_n2007.n0 4.4
R6299 a_n9429_n2007.n16 a_n9429_n2007.n15 4.35275
R6300 a_n9429_n2007.t0 a_n9429_n2007.n18 2.048
R6301 a_n9429_n2007.n18 a_n9429_n2007.t21 2.048
R6302 a_n9429_n2007.n17 a_n9429_n2007.n1 1.95895
R6303 a_n9429_n2007.n9 a_n9429_n2007.t2 1.0925
R6304 a_n9429_n2007.n9 a_n9429_n2007.t20 1.0925
R6305 a_n9429_n2007.n0 a_n9429_n2007.t17 1.0925
R6306 a_n9429_n2007.n0 a_n9429_n2007.t9 1.0925
R6307 a_n9429_n2007.n2 a_n9429_n2007.t7 1.0925
R6308 a_n9429_n2007.n2 a_n9429_n2007.t16 1.0925
R6309 a_n9429_n2007.n15 a_n9429_n2007.t14 1.0925
R6310 a_n9429_n2007.n15 a_n9429_n2007.t4 1.0925
R6311 a_n9429_n2007.n3 a_n9429_n2007.t11 1.0925
R6312 a_n9429_n2007.n3 a_n9429_n2007.t3 1.0925
R6313 a_n9429_n2007.n4 a_n9429_n2007.t10 1.0925
R6314 a_n9429_n2007.n4 a_n9429_n2007.t18 1.0925
R6315 a_n9429_n2007.n5 a_n9429_n2007.t6 1.0925
R6316 a_n9429_n2007.n5 a_n9429_n2007.t15 1.0925
R6317 a_n9429_n2007.n6 a_n9429_n2007.t13 1.0925
R6318 a_n9429_n2007.n6 a_n9429_n2007.t1 1.0925
R6319 a_n9429_n2007.n7 a_n9429_n2007.t19 1.0925
R6320 a_n9429_n2007.n7 a_n9429_n2007.t5 1.0925
R6321 a_n9429_n2007.n8 a_n9429_n2007.t8 1.0925
R6322 a_n9429_n2007.n8 a_n9429_n2007.t12 1.0925
R6323 a_n9429_n2007.n14 a_n9429_n2007.n13 0.849071
R6324 a_n9429_n2007.n13 a_n9429_n2007.n12 0.849071
R6325 a_n9429_n2007.n12 a_n9429_n2007.n11 0.849071
R6326 a_n9429_n2007.n11 a_n9429_n2007.n10 0.849071
R6327 a_n9429_n2007.n16 a_n9429_n2007.n14 0.534875
R6328 a_n9429_n2007.n10 a_n9429_n2007.n1 0.487625
R6329 SARlogic_0.d1.n3 SARlogic_0.d1.t9 41.0041
R6330 SARlogic_0.d1.n4 SARlogic_0.d1.t7 40.8177
R6331 SARlogic_0.d1.n7 SARlogic_0.d1.t8 40.6313
R6332 SARlogic_0.d1.n1 SARlogic_0.d1.t4 34.2529
R6333 SARlogic_0.d1.n6 SARlogic_0.dffrs_9.clk 33.8765
R6334 SARlogic_0.d1.n7 SARlogic_0.d1.t5 27.3166
R6335 SARlogic_0.d1.n4 SARlogic_0.d1.t12 27.1302
R6336 SARlogic_0.d1.n3 SARlogic_0.d1.t11 26.9438
R6337 SARlogic_0.d1 adc_PISO_0.B2 26.2596
R6338 SARlogic_0.d1.n0 SARlogic_0.d1.t6 19.673
R6339 SARlogic_0.d1.n0 SARlogic_0.d1.t10 19.4007
R6340 SARlogic_0.d1.n9 SARlogic_0.d1.n8 14.0582
R6341 SARlogic_0.d1.n9 SARlogic_0.d1.n6 11.729
R6342 SARlogic_0.d1.n12 SARlogic_0.d1.t2 10.0473
R6343 SARlogic_0.d1.n2 SARlogic_0.d1.n1 8.05164
R6344 SARlogic_0.d1.n11 SARlogic_0.d1.t3 6.51042
R6345 SARlogic_0.d1.n11 SARlogic_0.d1.n10 6.04952
R6346 SARlogic_0.dffrs_9.nand3_1.A SARlogic_0.d1.n3 5.7755
R6347 SARlogic_0.dffrs_9.nand3_6.B SARlogic_0.d1.n4 5.47979
R6348 SARlogic_0.d1.n8 SARlogic_0.d1.n7 5.13907
R6349 SARlogic_0.dffrs_10.nand3_2.Z SARlogic_0.d1.n12 4.72925
R6350 SARlogic_0.d1.n5 SARlogic_0.dffrs_9.nand3_6.B 2.17818
R6351 adc_PISO_0.B2 SARlogic_0.d1.n2 1.87121
R6352 SARlogic_0.d1.n5 SARlogic_0.dffrs_9.nand3_1.A 1.34729
R6353 SARlogic_0.d1.n6 SARlogic_0.d1 0.985679
R6354 SARlogic_0.d1.n12 SARlogic_0.d1.n11 0.732092
R6355 SARlogic_0.d1.n10 SARlogic_0.d1.t0 0.7285
R6356 SARlogic_0.d1.n10 SARlogic_0.d1.t1 0.7285
R6357 SARlogic_0.dffrs_9.clk SARlogic_0.d1.n5 0.610571
R6358 SARlogic_0.dffrs_10.nand3_2.Z SARlogic_0.d1.n9 0.166901
R6359 SARlogic_0.d1.n1 SARlogic_0.d1.n0 0.106438
R6360 SARlogic_0.d1.n8 SARlogic_0.dffrs_10.nand3_7.C 0.0455
R6361 SARlogic_0.d1.n2 adc_PISO_0.2inmux_5.In 0.0455
R6362 a_28027_28820.n0 a_28027_28820.t5 34.1797
R6363 a_28027_28820.n0 a_28027_28820.t4 19.5798
R6364 a_28027_28820.t1 a_28027_28820.n3 18.7717
R6365 a_28027_28820.n3 a_28027_28820.t0 9.2885
R6366 a_28027_28820.n2 a_28027_28820.n0 4.93379
R6367 a_28027_28820.n1 a_28027_28820.t3 4.23346
R6368 a_28027_28820.n1 a_28027_28820.t2 3.85546
R6369 a_28027_28820.n3 a_28027_28820.n2 0.4055
R6370 a_28027_28820.n2 a_28027_28820.n1 0.352625
R6371 Reset.n80 Reset.t25 41.0041
R6372 Reset.n86 Reset.t52 41.0041
R6373 Reset.n66 Reset.t59 41.0041
R6374 Reset.n72 Reset.t1 41.0041
R6375 Reset.n52 Reset.t39 41.0041
R6376 Reset.n58 Reset.t66 41.0041
R6377 Reset.n38 Reset.t48 41.0041
R6378 Reset.n44 Reset.t72 41.0041
R6379 Reset.n24 Reset.t36 41.0041
R6380 Reset.n30 Reset.t64 41.0041
R6381 Reset.n10 Reset.t65 41.0041
R6382 Reset.n16 Reset.t7 41.0041
R6383 Reset.n4 Reset.t38 41.0041
R6384 Reset.n83 Reset.t10 40.8177
R6385 Reset.n82 Reset.t0 40.8177
R6386 Reset.n89 Reset.t26 40.8177
R6387 Reset.n88 Reset.t29 40.8177
R6388 Reset.n69 Reset.t37 40.8177
R6389 Reset.n68 Reset.t28 40.8177
R6390 Reset.n75 Reset.t54 40.8177
R6391 Reset.n74 Reset.t57 40.8177
R6392 Reset.n55 Reset.t30 40.8177
R6393 Reset.n54 Reset.t20 40.8177
R6394 Reset.n61 Reset.t75 40.8177
R6395 Reset.n60 Reset.t51 40.8177
R6396 Reset.n41 Reset.t58 40.8177
R6397 Reset.n40 Reset.t53 40.8177
R6398 Reset.n47 Reset.t42 40.8177
R6399 Reset.n46 Reset.t77 40.8177
R6400 Reset.n27 Reset.t2 40.8177
R6401 Reset.n26 Reset.t78 40.8177
R6402 Reset.n33 Reset.t34 40.8177
R6403 Reset.n32 Reset.t24 40.8177
R6404 Reset.n13 Reset.t76 40.8177
R6405 Reset.n12 Reset.t68 40.8177
R6406 Reset.n19 Reset.t73 40.8177
R6407 Reset.n18 Reset.t13 40.8177
R6408 Reset.n7 Reset.t21 40.8177
R6409 Reset.n6 Reset.t14 40.8177
R6410 Reset.n2 Reset.t63 40.6313
R6411 Reset.n0 Reset.t62 40.6313
R6412 Reset.n2 Reset.t23 27.3166
R6413 Reset.n0 Reset.t79 27.3166
R6414 Reset.n83 Reset.t35 27.1302
R6415 Reset.n82 Reset.t22 27.1302
R6416 Reset.n89 Reset.t45 27.1302
R6417 Reset.n88 Reset.t50 27.1302
R6418 Reset.n69 Reset.t61 27.1302
R6419 Reset.n68 Reset.t49 27.1302
R6420 Reset.n75 Reset.t70 27.1302
R6421 Reset.n74 Reset.t74 27.1302
R6422 Reset.n55 Reset.t55 27.1302
R6423 Reset.n54 Reset.t43 27.1302
R6424 Reset.n61 Reset.t11 27.1302
R6425 Reset.n60 Reset.t67 27.1302
R6426 Reset.n41 Reset.t80 27.1302
R6427 Reset.n40 Reset.t69 27.1302
R6428 Reset.n47 Reset.t60 27.1302
R6429 Reset.n46 Reset.t16 27.1302
R6430 Reset.n27 Reset.t27 27.1302
R6431 Reset.n26 Reset.t17 27.1302
R6432 Reset.n33 Reset.t56 27.1302
R6433 Reset.n32 Reset.t44 27.1302
R6434 Reset.n13 Reset.t18 27.1302
R6435 Reset.n12 Reset.t3 27.1302
R6436 Reset.n19 Reset.t8 27.1302
R6437 Reset.n18 Reset.t31 27.1302
R6438 Reset.n7 Reset.t47 27.1302
R6439 Reset.n6 Reset.t32 27.1302
R6440 Reset.n80 Reset.t81 26.9438
R6441 Reset.n86 Reset.t6 26.9438
R6442 Reset.n66 Reset.t33 26.9438
R6443 Reset.n72 Reset.t5 26.9438
R6444 Reset.n52 Reset.t15 26.9438
R6445 Reset.n58 Reset.t71 26.9438
R6446 Reset.n38 Reset.t19 26.9438
R6447 Reset.n44 Reset.t4 26.9438
R6448 Reset.n24 Reset.t9 26.9438
R6449 Reset.n30 Reset.t46 26.9438
R6450 Reset.n10 Reset.t41 26.9438
R6451 Reset.n16 Reset.t40 26.9438
R6452 Reset.n4 Reset.t12 26.9438
R6453 Reset.n78 SARlogic_0.dffrs_1.resetb 19.0901
R6454 Reset.n64 SARlogic_0.dffrs_2.resetb 19.0901
R6455 Reset.n50 SARlogic_0.dffrs_3.resetb 19.0901
R6456 Reset.n36 SARlogic_0.dffrs_4.resetb 19.0901
R6457 Reset.n22 SARlogic_0.dffrs_5.resetb 19.0901
R6458 Reset.n92 SARlogic_0.dffrs_0.resetb 19.0467
R6459 Reset.n23 SARlogic_0.dffrs_12.resetb 14.0622
R6460 Reset.n84 SARlogic_0.dffrs_14.nand3_1.B 12.1571
R6461 Reset.n90 SARlogic_0.dffrs_0.nand3_1.B 12.1571
R6462 Reset.n70 SARlogic_0.dffrs_7.nand3_1.B 12.1571
R6463 Reset.n76 SARlogic_0.dffrs_1.nand3_1.B 12.1571
R6464 Reset.n56 SARlogic_0.dffrs_8.nand3_1.B 12.1571
R6465 Reset.n62 SARlogic_0.dffrs_2.nand3_1.B 12.1571
R6466 Reset.n42 SARlogic_0.dffrs_9.nand3_1.B 12.1571
R6467 Reset.n48 SARlogic_0.dffrs_3.nand3_1.B 12.1571
R6468 Reset.n28 SARlogic_0.dffrs_10.nand3_1.B 12.1571
R6469 Reset.n34 SARlogic_0.dffrs_4.nand3_1.B 12.1571
R6470 Reset.n14 SARlogic_0.dffrs_11.nand3_1.B 12.1571
R6471 Reset.n20 SARlogic_0.dffrs_5.nand3_1.B 12.1571
R6472 Reset.n8 SARlogic_0.dffrs_12.nand3_1.B 12.1571
R6473 Reset.n3 Reset.n1 9.22229
R6474 Reset.n94 Reset.n93 7.9889
R6475 Reset.n85 Reset.n81 7.75389
R6476 Reset.n91 Reset.n87 7.75389
R6477 Reset.n71 Reset.n67 7.75389
R6478 Reset.n77 Reset.n73 7.75389
R6479 Reset.n57 Reset.n53 7.75389
R6480 Reset.n63 Reset.n59 7.75389
R6481 Reset.n43 Reset.n39 7.75389
R6482 Reset.n49 Reset.n45 7.75389
R6483 Reset.n29 Reset.n25 7.75389
R6484 Reset.n35 Reset.n31 7.75389
R6485 Reset.n15 Reset.n11 7.75389
R6486 Reset.n21 Reset.n17 7.75389
R6487 Reset.n9 Reset.n5 7.75389
R6488 Reset.n94 SARlogic_0.dffrs_13.setb 6.43164
R6489 Reset.n85 Reset.n84 5.93546
R6490 Reset.n91 Reset.n90 5.93546
R6491 Reset.n71 Reset.n70 5.93546
R6492 Reset.n77 Reset.n76 5.93546
R6493 Reset.n57 Reset.n56 5.93546
R6494 Reset.n63 Reset.n62 5.93546
R6495 Reset.n43 Reset.n42 5.93546
R6496 Reset.n49 Reset.n48 5.93546
R6497 Reset.n29 Reset.n28 5.93546
R6498 Reset.n35 Reset.n34 5.93546
R6499 Reset.n15 Reset.n14 5.93546
R6500 Reset.n21 Reset.n20 5.93546
R6501 Reset.n9 Reset.n8 5.93546
R6502 Reset.n78 SARlogic_0.dffrs_7.resetb 5.93246
R6503 Reset.n64 SARlogic_0.dffrs_8.resetb 5.93246
R6504 Reset.n50 SARlogic_0.dffrs_9.resetb 5.93246
R6505 Reset.n36 SARlogic_0.dffrs_10.resetb 5.93246
R6506 Reset.n22 SARlogic_0.dffrs_11.resetb 5.93246
R6507 Reset.n92 SARlogic_0.dffrs_14.resetb 5.88425
R6508 Reset.n81 Reset.n80 5.7305
R6509 Reset.n87 Reset.n86 5.7305
R6510 Reset.n67 Reset.n66 5.7305
R6511 Reset.n73 Reset.n72 5.7305
R6512 Reset.n53 Reset.n52 5.7305
R6513 Reset.n59 Reset.n58 5.7305
R6514 Reset.n39 Reset.n38 5.7305
R6515 Reset.n45 Reset.n44 5.7305
R6516 Reset.n25 Reset.n24 5.7305
R6517 Reset.n31 Reset.n30 5.7305
R6518 Reset.n11 Reset.n10 5.7305
R6519 Reset.n17 Reset.n16 5.7305
R6520 Reset.n5 Reset.n4 5.7305
R6521 SARlogic_0.dffrs_14.nand3_8.B Reset.n83 5.47979
R6522 SARlogic_0.dffrs_14.nand3_1.B Reset.n82 5.47979
R6523 SARlogic_0.dffrs_0.nand3_8.B Reset.n89 5.47979
R6524 SARlogic_0.dffrs_0.nand3_1.B Reset.n88 5.47979
R6525 SARlogic_0.dffrs_7.nand3_8.B Reset.n69 5.47979
R6526 SARlogic_0.dffrs_7.nand3_1.B Reset.n68 5.47979
R6527 SARlogic_0.dffrs_1.nand3_8.B Reset.n75 5.47979
R6528 SARlogic_0.dffrs_1.nand3_1.B Reset.n74 5.47979
R6529 SARlogic_0.dffrs_8.nand3_8.B Reset.n55 5.47979
R6530 SARlogic_0.dffrs_8.nand3_1.B Reset.n54 5.47979
R6531 SARlogic_0.dffrs_2.nand3_8.B Reset.n61 5.47979
R6532 SARlogic_0.dffrs_2.nand3_1.B Reset.n60 5.47979
R6533 SARlogic_0.dffrs_9.nand3_8.B Reset.n41 5.47979
R6534 SARlogic_0.dffrs_9.nand3_1.B Reset.n40 5.47979
R6535 SARlogic_0.dffrs_3.nand3_8.B Reset.n47 5.47979
R6536 SARlogic_0.dffrs_3.nand3_1.B Reset.n46 5.47979
R6537 SARlogic_0.dffrs_10.nand3_8.B Reset.n27 5.47979
R6538 SARlogic_0.dffrs_10.nand3_1.B Reset.n26 5.47979
R6539 SARlogic_0.dffrs_4.nand3_8.B Reset.n33 5.47979
R6540 SARlogic_0.dffrs_4.nand3_1.B Reset.n32 5.47979
R6541 SARlogic_0.dffrs_11.nand3_8.B Reset.n13 5.47979
R6542 SARlogic_0.dffrs_11.nand3_1.B Reset.n12 5.47979
R6543 SARlogic_0.dffrs_5.nand3_8.B Reset.n19 5.47979
R6544 SARlogic_0.dffrs_5.nand3_1.B Reset.n18 5.47979
R6545 SARlogic_0.dffrs_12.nand3_8.B Reset.n7 5.47979
R6546 SARlogic_0.dffrs_12.nand3_1.B Reset.n6 5.47979
R6547 Reset.n3 Reset.n2 5.14711
R6548 Reset.n1 Reset.n0 5.13907
R6549 Reset.n84 SARlogic_0.dffrs_14.nand3_8.B 5.09593
R6550 Reset.n90 SARlogic_0.dffrs_0.nand3_8.B 5.09593
R6551 Reset.n70 SARlogic_0.dffrs_7.nand3_8.B 5.09593
R6552 Reset.n76 SARlogic_0.dffrs_1.nand3_8.B 5.09593
R6553 Reset.n56 SARlogic_0.dffrs_8.nand3_8.B 5.09593
R6554 Reset.n62 SARlogic_0.dffrs_2.nand3_8.B 5.09593
R6555 Reset.n42 SARlogic_0.dffrs_9.nand3_8.B 5.09593
R6556 Reset.n48 SARlogic_0.dffrs_3.nand3_8.B 5.09593
R6557 Reset.n28 SARlogic_0.dffrs_10.nand3_8.B 5.09593
R6558 Reset.n34 SARlogic_0.dffrs_4.nand3_8.B 5.09593
R6559 Reset.n14 SARlogic_0.dffrs_11.nand3_8.B 5.09593
R6560 Reset.n20 SARlogic_0.dffrs_5.nand3_8.B 5.09593
R6561 Reset.n8 SARlogic_0.dffrs_12.nand3_8.B 5.09593
R6562 Reset.n23 Reset.n22 4.5005
R6563 Reset.n37 Reset.n36 4.5005
R6564 Reset.n51 Reset.n50 4.5005
R6565 Reset.n65 Reset.n64 4.5005
R6566 Reset.n79 Reset.n78 4.5005
R6567 Reset.n93 Reset.n92 4.5005
R6568 Reset.n37 Reset.n23 3.6383
R6569 Reset.n51 Reset.n37 3.6383
R6570 Reset.n65 Reset.n51 3.6383
R6571 Reset.n79 Reset.n65 3.6383
R6572 Reset.n93 Reset.n79 3.6113
R6573 SARlogic_0.dffrs_13.setb SARlogic_0.dffrs_13.nand3_0.C 0.783821
R6574 SARlogic_0.reset Reset 0.18425
R6575 SARlogic_0.reset Reset.n94 0.13775
R6576 SARlogic_0.dffrs_14.resetb Reset.n85 0.136036
R6577 SARlogic_0.dffrs_0.resetb Reset.n91 0.136036
R6578 SARlogic_0.dffrs_7.resetb Reset.n71 0.136036
R6579 SARlogic_0.dffrs_1.resetb Reset.n77 0.136036
R6580 SARlogic_0.dffrs_8.resetb Reset.n57 0.136036
R6581 SARlogic_0.dffrs_2.resetb Reset.n63 0.136036
R6582 SARlogic_0.dffrs_9.resetb Reset.n43 0.136036
R6583 SARlogic_0.dffrs_3.resetb Reset.n49 0.136036
R6584 SARlogic_0.dffrs_10.resetb Reset.n29 0.136036
R6585 SARlogic_0.dffrs_4.resetb Reset.n35 0.136036
R6586 SARlogic_0.dffrs_11.resetb Reset.n15 0.136036
R6587 SARlogic_0.dffrs_5.resetb Reset.n21 0.136036
R6588 SARlogic_0.dffrs_12.resetb Reset.n9 0.136036
R6589 Reset.n1 SARlogic_0.dffrs_13.nand3_2.C 0.0455
R6590 Reset.n81 SARlogic_0.dffrs_14.nand3_7.A 0.0455
R6591 Reset.n87 SARlogic_0.dffrs_0.nand3_7.A 0.0455
R6592 Reset.n67 SARlogic_0.dffrs_7.nand3_7.A 0.0455
R6593 Reset.n73 SARlogic_0.dffrs_1.nand3_7.A 0.0455
R6594 Reset.n53 SARlogic_0.dffrs_8.nand3_7.A 0.0455
R6595 Reset.n59 SARlogic_0.dffrs_2.nand3_7.A 0.0455
R6596 Reset.n39 SARlogic_0.dffrs_9.nand3_7.A 0.0455
R6597 Reset.n45 SARlogic_0.dffrs_3.nand3_7.A 0.0455
R6598 Reset.n25 SARlogic_0.dffrs_10.nand3_7.A 0.0455
R6599 Reset.n31 SARlogic_0.dffrs_4.nand3_7.A 0.0455
R6600 Reset.n11 SARlogic_0.dffrs_11.nand3_7.A 0.0455
R6601 Reset.n17 SARlogic_0.dffrs_5.nand3_7.A 0.0455
R6602 Reset.n5 SARlogic_0.dffrs_12.nand3_7.A 0.0455
R6603 SARlogic_0.dffrs_13.nand3_0.C Reset.n3 0.0374643
R6604 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t5 41.0041
R6605 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t4 40.8177
R6606 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t9 40.6313
R6607 SARlogic_0.dffrs_14.nand3_6.C.n3 SARlogic_0.dffrs_14.nand3_6.C.t8 27.3166
R6608 SARlogic_0.dffrs_14.nand3_6.C.n0 SARlogic_0.dffrs_14.nand3_6.C.t6 27.1302
R6609 SARlogic_0.dffrs_14.nand3_6.C.n1 SARlogic_0.dffrs_14.nand3_6.C.t7 26.9438
R6610 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.t3 10.0473
R6611 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n4 9.90747
R6612 SARlogic_0.dffrs_14.nand3_6.C.n5 SARlogic_0.dffrs_14.nand3_6.C.n2 9.90116
R6613 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.t2 6.51042
R6614 SARlogic_0.dffrs_14.nand3_6.C.n8 SARlogic_0.dffrs_14.nand3_6.C.n7 6.04952
R6615 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_6.C.n1 5.7305
R6616 SARlogic_0.dffrs_14.nand3_2.B SARlogic_0.dffrs_14.nand3_6.C.n0 5.47979
R6617 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C.n3 5.13907
R6618 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n9 4.72925
R6619 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_6.C.n5 4.5005
R6620 SARlogic_0.dffrs_14.nand3_6.C.n9 SARlogic_0.dffrs_14.nand3_6.C.n8 0.732092
R6621 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t1 0.7285
R6622 SARlogic_0.dffrs_14.nand3_6.C.n7 SARlogic_0.dffrs_14.nand3_6.C.t0 0.7285
R6623 SARlogic_0.dffrs_14.nand3_1.Z SARlogic_0.dffrs_14.nand3_6.C.n6 0.449758
R6624 SARlogic_0.dffrs_14.nand3_6.C.n6 SARlogic_0.dffrs_14.nand3_2.B 0.166901
R6625 SARlogic_0.dffrs_14.nand3_6.C.n2 SARlogic_0.dffrs_14.nand3_0.A 0.0455
R6626 SARlogic_0.dffrs_14.nand3_6.C.n4 SARlogic_0.dffrs_14.nand3_6.C 0.0455
R6627 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t8 41.0041
R6628 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t7 40.8177
R6629 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t6 40.6313
R6630 SARlogic_0.dffrs_2.nand3_6.C.n3 SARlogic_0.dffrs_2.nand3_6.C.t5 27.3166
R6631 SARlogic_0.dffrs_2.nand3_6.C.n0 SARlogic_0.dffrs_2.nand3_6.C.t9 27.1302
R6632 SARlogic_0.dffrs_2.nand3_6.C.n1 SARlogic_0.dffrs_2.nand3_6.C.t4 26.9438
R6633 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.t3 10.0473
R6634 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n4 9.90747
R6635 SARlogic_0.dffrs_2.nand3_6.C.n5 SARlogic_0.dffrs_2.nand3_6.C.n2 9.90116
R6636 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.t0 6.51042
R6637 SARlogic_0.dffrs_2.nand3_6.C.n8 SARlogic_0.dffrs_2.nand3_6.C.n7 6.04952
R6638 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_6.C.n1 5.7305
R6639 SARlogic_0.dffrs_2.nand3_2.B SARlogic_0.dffrs_2.nand3_6.C.n0 5.47979
R6640 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C.n3 5.13907
R6641 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n9 4.72925
R6642 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_6.C.n5 4.5005
R6643 SARlogic_0.dffrs_2.nand3_6.C.n9 SARlogic_0.dffrs_2.nand3_6.C.n8 0.732092
R6644 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t1 0.7285
R6645 SARlogic_0.dffrs_2.nand3_6.C.n7 SARlogic_0.dffrs_2.nand3_6.C.t2 0.7285
R6646 SARlogic_0.dffrs_2.nand3_1.Z SARlogic_0.dffrs_2.nand3_6.C.n6 0.449758
R6647 SARlogic_0.dffrs_2.nand3_6.C.n6 SARlogic_0.dffrs_2.nand3_2.B 0.166901
R6648 SARlogic_0.dffrs_2.nand3_6.C.n2 SARlogic_0.dffrs_2.nand3_0.A 0.0455
R6649 SARlogic_0.dffrs_2.nand3_6.C.n4 SARlogic_0.dffrs_2.nand3_6.C 0.0455
R6650 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t4 40.6313
R6651 SARlogic_0.dffrs_2.nand3_1.C.n0 SARlogic_0.dffrs_2.nand3_1.C.t5 27.3166
R6652 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n1 14.2854
R6653 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.t3 10.0473
R6654 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.t2 6.51042
R6655 SARlogic_0.dffrs_2.nand3_1.C.n3 SARlogic_0.dffrs_2.nand3_1.C.n2 6.04952
R6656 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C.n0 5.13907
R6657 SARlogic_0.dffrs_2.nand3_0.Z SARlogic_0.dffrs_2.nand3_1.C.n4 4.72925
R6658 SARlogic_0.dffrs_2.nand3_1.C.n4 SARlogic_0.dffrs_2.nand3_1.C.n3 0.732092
R6659 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t0 0.7285
R6660 SARlogic_0.dffrs_2.nand3_1.C.n2 SARlogic_0.dffrs_2.nand3_1.C.t1 0.7285
R6661 SARlogic_0.dffrs_2.nand3_1.C.n1 SARlogic_0.dffrs_2.nand3_1.C 0.0455
R6662 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t8 41.0041
R6663 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t5 40.6313
R6664 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t4 40.6313
R6665 SARlogic_0.dffrs_1.Qb SARlogic_0.dffrs_8.setb 28.021
R6666 SARlogic_0.dffrs_1.Qb.n4 SARlogic_0.dffrs_1.Qb.t7 27.3166
R6667 SARlogic_0.dffrs_1.Qb.n2 SARlogic_0.dffrs_1.Qb.t6 27.3166
R6668 SARlogic_0.dffrs_1.Qb.n0 SARlogic_0.dffrs_1.Qb.t9 26.9438
R6669 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.t1 10.0473
R6670 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb.n1 9.84255
R6671 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n3 9.22229
R6672 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.t2 6.51042
R6673 SARlogic_0.dffrs_1.Qb.n8 SARlogic_0.dffrs_1.Qb.n7 6.04952
R6674 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.Qb.n0 5.7305
R6675 SARlogic_0.dffrs_1.Qb.n5 SARlogic_0.dffrs_1.Qb.n4 5.14711
R6676 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_1.Qb.n2 5.13907
R6677 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n6 4.94976
R6678 SARlogic_0.dffrs_1.nand3_7.Z SARlogic_0.dffrs_1.Qb.n9 4.72925
R6679 SARlogic_0.dffrs_8.setb SARlogic_0.dffrs_8.nand3_0.C 0.784786
R6680 SARlogic_0.dffrs_1.Qb.n9 SARlogic_0.dffrs_1.Qb.n8 0.732092
R6681 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t3 0.7285
R6682 SARlogic_0.dffrs_1.Qb.n7 SARlogic_0.dffrs_1.Qb.t0 0.7285
R6683 SARlogic_0.dffrs_1.Qb.n6 SARlogic_0.dffrs_1.Qb 0.175225
R6684 SARlogic_0.dffrs_1.Qb.n1 SARlogic_0.dffrs_1.nand3_2.A 0.0455
R6685 SARlogic_0.dffrs_1.Qb.n3 SARlogic_0.dffrs_8.nand3_2.C 0.0455
R6686 SARlogic_0.dffrs_8.nand3_0.C SARlogic_0.dffrs_1.Qb.n5 0.0374643
R6687 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t6 41.0041
R6688 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t5 40.8177
R6689 SARlogic_0.dffrs_4.nand3_8.Z.n1 SARlogic_0.dffrs_4.nand3_8.Z.t7 27.1302
R6690 SARlogic_0.dffrs_4.nand3_8.Z.n0 SARlogic_0.dffrs_4.nand3_8.Z.t4 26.9438
R6691 SARlogic_0.dffrs_4.nand3_6.A SARlogic_0.dffrs_4.nand3_0.B 17.0041
R6692 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n2 14.8493
R6693 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.t2 10.0473
R6694 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.t3 6.51042
R6695 SARlogic_0.dffrs_4.nand3_8.Z.n4 SARlogic_0.dffrs_4.nand3_8.Z.n3 6.04952
R6696 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_8.Z.n0 5.7305
R6697 SARlogic_0.dffrs_4.nand3_0.B SARlogic_0.dffrs_4.nand3_8.Z.n1 5.47979
R6698 SARlogic_0.dffrs_4.nand3_8.Z SARlogic_0.dffrs_4.nand3_8.Z.n5 4.72925
R6699 SARlogic_0.dffrs_4.nand3_8.Z.n5 SARlogic_0.dffrs_4.nand3_8.Z.n4 0.732092
R6700 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t0 0.7285
R6701 SARlogic_0.dffrs_4.nand3_8.Z.n3 SARlogic_0.dffrs_4.nand3_8.Z.t1 0.7285
R6702 SARlogic_0.dffrs_4.nand3_8.Z.n2 SARlogic_0.dffrs_4.nand3_6.A 0.0455
R6703 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t7 40.8177
R6704 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t5 40.6313
R6705 SARlogic_0.dffrs_4.nand3_8.C.n1 SARlogic_0.dffrs_4.nand3_8.C.t6 27.3166
R6706 SARlogic_0.dffrs_4.nand3_8.C.n0 SARlogic_0.dffrs_4.nand3_8.C.t4 27.1302
R6707 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_8.C.n2 14.119
R6708 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.t0 10.0473
R6709 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.t1 6.51042
R6710 SARlogic_0.dffrs_4.nand3_8.C.n5 SARlogic_0.dffrs_4.nand3_8.C.n4 6.04952
R6711 SARlogic_0.dffrs_4.nand3_7.B SARlogic_0.dffrs_4.nand3_8.C.n0 5.47979
R6712 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C.n1 5.13907
R6713 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n6 4.72925
R6714 SARlogic_0.dffrs_4.nand3_8.C.n6 SARlogic_0.dffrs_4.nand3_8.C.n5 0.732092
R6715 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t2 0.7285
R6716 SARlogic_0.dffrs_4.nand3_8.C.n4 SARlogic_0.dffrs_4.nand3_8.C.t3 0.7285
R6717 SARlogic_0.dffrs_4.nand3_8.C.n3 SARlogic_0.dffrs_4.nand3_7.B 0.438233
R6718 SARlogic_0.dffrs_4.nand3_6.Z SARlogic_0.dffrs_4.nand3_8.C.n3 0.166901
R6719 SARlogic_0.dffrs_4.nand3_8.C.n2 SARlogic_0.dffrs_4.nand3_8.C 0.0455
R6720 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t4 40.8177
R6721 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t6 40.6313
R6722 SARlogic_0.dffrs_1.nand3_8.C.n1 SARlogic_0.dffrs_1.nand3_8.C.t7 27.3166
R6723 SARlogic_0.dffrs_1.nand3_8.C.n0 SARlogic_0.dffrs_1.nand3_8.C.t5 27.1302
R6724 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_8.C.n2 14.119
R6725 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.t1 10.0473
R6726 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.t0 6.51042
R6727 SARlogic_0.dffrs_1.nand3_8.C.n5 SARlogic_0.dffrs_1.nand3_8.C.n4 6.04952
R6728 SARlogic_0.dffrs_1.nand3_7.B SARlogic_0.dffrs_1.nand3_8.C.n0 5.47979
R6729 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C.n1 5.13907
R6730 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n6 4.72925
R6731 SARlogic_0.dffrs_1.nand3_8.C.n6 SARlogic_0.dffrs_1.nand3_8.C.n5 0.732092
R6732 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t3 0.7285
R6733 SARlogic_0.dffrs_1.nand3_8.C.n4 SARlogic_0.dffrs_1.nand3_8.C.t2 0.7285
R6734 SARlogic_0.dffrs_1.nand3_8.C.n3 SARlogic_0.dffrs_1.nand3_7.B 0.438233
R6735 SARlogic_0.dffrs_1.nand3_6.Z SARlogic_0.dffrs_1.nand3_8.C.n3 0.166901
R6736 SARlogic_0.dffrs_1.nand3_8.C.n2 SARlogic_0.dffrs_1.nand3_8.C 0.0455
R6737 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t6 40.8177
R6738 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t7 40.6313
R6739 SARlogic_0.dffrs_5.nand3_8.C.n1 SARlogic_0.dffrs_5.nand3_8.C.t4 27.3166
R6740 SARlogic_0.dffrs_5.nand3_8.C.n0 SARlogic_0.dffrs_5.nand3_8.C.t5 27.1302
R6741 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_8.C.n2 14.119
R6742 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.t1 10.0473
R6743 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.t2 6.51042
R6744 SARlogic_0.dffrs_5.nand3_8.C.n5 SARlogic_0.dffrs_5.nand3_8.C.n4 6.04952
R6745 SARlogic_0.dffrs_5.nand3_7.B SARlogic_0.dffrs_5.nand3_8.C.n0 5.47979
R6746 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C.n1 5.13907
R6747 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n6 4.72925
R6748 SARlogic_0.dffrs_5.nand3_8.C.n6 SARlogic_0.dffrs_5.nand3_8.C.n5 0.732092
R6749 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t0 0.7285
R6750 SARlogic_0.dffrs_5.nand3_8.C.n4 SARlogic_0.dffrs_5.nand3_8.C.t3 0.7285
R6751 SARlogic_0.dffrs_5.nand3_8.C.n3 SARlogic_0.dffrs_5.nand3_7.B 0.438233
R6752 SARlogic_0.dffrs_5.nand3_6.Z SARlogic_0.dffrs_5.nand3_8.C.n3 0.166901
R6753 SARlogic_0.dffrs_5.nand3_8.C.n2 SARlogic_0.dffrs_5.nand3_8.C 0.0455
R6754 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t4 41.0041
R6755 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t7 40.8177
R6756 SARlogic_0.dffrs_3.nand3_8.Z.n1 SARlogic_0.dffrs_3.nand3_8.Z.t6 27.1302
R6757 SARlogic_0.dffrs_3.nand3_8.Z.n0 SARlogic_0.dffrs_3.nand3_8.Z.t5 26.9438
R6758 SARlogic_0.dffrs_3.nand3_6.A SARlogic_0.dffrs_3.nand3_0.B 17.0041
R6759 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n2 14.8493
R6760 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.t2 10.0473
R6761 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.t3 6.51042
R6762 SARlogic_0.dffrs_3.nand3_8.Z.n4 SARlogic_0.dffrs_3.nand3_8.Z.n3 6.04952
R6763 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_8.Z.n0 5.7305
R6764 SARlogic_0.dffrs_3.nand3_0.B SARlogic_0.dffrs_3.nand3_8.Z.n1 5.47979
R6765 SARlogic_0.dffrs_3.nand3_8.Z SARlogic_0.dffrs_3.nand3_8.Z.n5 4.72925
R6766 SARlogic_0.dffrs_3.nand3_8.Z.n5 SARlogic_0.dffrs_3.nand3_8.Z.n4 0.732092
R6767 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t0 0.7285
R6768 SARlogic_0.dffrs_3.nand3_8.Z.n3 SARlogic_0.dffrs_3.nand3_8.Z.t1 0.7285
R6769 SARlogic_0.dffrs_3.nand3_8.Z.n2 SARlogic_0.dffrs_3.nand3_6.A 0.0455
R6770 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t7 40.8177
R6771 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t5 40.6313
R6772 SARlogic_0.dffrs_3.nand3_8.C.n1 SARlogic_0.dffrs_3.nand3_8.C.t6 27.3166
R6773 SARlogic_0.dffrs_3.nand3_8.C.n0 SARlogic_0.dffrs_3.nand3_8.C.t4 27.1302
R6774 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_8.C.n2 14.119
R6775 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.t0 10.0473
R6776 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.t1 6.51042
R6777 SARlogic_0.dffrs_3.nand3_8.C.n5 SARlogic_0.dffrs_3.nand3_8.C.n4 6.04952
R6778 SARlogic_0.dffrs_3.nand3_7.B SARlogic_0.dffrs_3.nand3_8.C.n0 5.47979
R6779 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C.n1 5.13907
R6780 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n6 4.72925
R6781 SARlogic_0.dffrs_3.nand3_8.C.n6 SARlogic_0.dffrs_3.nand3_8.C.n5 0.732092
R6782 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t3 0.7285
R6783 SARlogic_0.dffrs_3.nand3_8.C.n4 SARlogic_0.dffrs_3.nand3_8.C.t2 0.7285
R6784 SARlogic_0.dffrs_3.nand3_8.C.n3 SARlogic_0.dffrs_3.nand3_7.B 0.438233
R6785 SARlogic_0.dffrs_3.nand3_6.Z SARlogic_0.dffrs_3.nand3_8.C.n3 0.166901
R6786 SARlogic_0.dffrs_3.nand3_8.C.n2 SARlogic_0.dffrs_3.nand3_8.C 0.0455
R6787 a_33257_31423.n1 a_33257_31423.t5 41.0041
R6788 a_33257_31423.n0 a_33257_31423.t6 40.8177
R6789 a_33257_31423.n2 a_33257_31423.t9 40.6313
R6790 a_33257_31423.n2 a_33257_31423.t4 27.3166
R6791 a_33257_31423.n0 a_33257_31423.t8 27.1302
R6792 a_33257_31423.n1 a_33257_31423.t7 26.9438
R6793 a_33257_31423.n3 a_33257_31423.n1 15.6312
R6794 a_33257_31423.n3 a_33257_31423.n2 15.046
R6795 a_33257_31423.n5 a_33257_31423.t3 10.0473
R6796 a_33257_31423.n6 a_33257_31423.t2 6.51042
R6797 a_33257_31423.n7 a_33257_31423.n6 6.04952
R6798 a_33257_31423.n4 a_33257_31423.n0 5.64619
R6799 a_33257_31423.n5 a_33257_31423.n4 5.17851
R6800 a_33257_31423.n4 a_33257_31423.n3 4.5005
R6801 a_33257_31423.n6 a_33257_31423.n5 0.732092
R6802 a_33257_31423.t0 a_33257_31423.n7 0.7285
R6803 a_33257_31423.n7 a_33257_31423.t1 0.7285
R6804 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t8 41.0041
R6805 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t7 40.8177
R6806 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t4 40.6313
R6807 SARlogic_0.dffrs_5.nand3_6.C.n3 SARlogic_0.dffrs_5.nand3_6.C.t5 27.3166
R6808 SARlogic_0.dffrs_5.nand3_6.C.n0 SARlogic_0.dffrs_5.nand3_6.C.t9 27.1302
R6809 SARlogic_0.dffrs_5.nand3_6.C.n1 SARlogic_0.dffrs_5.nand3_6.C.t6 26.9438
R6810 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.t0 10.0473
R6811 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n4 9.90747
R6812 SARlogic_0.dffrs_5.nand3_6.C.n5 SARlogic_0.dffrs_5.nand3_6.C.n2 9.90116
R6813 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.t3 6.51042
R6814 SARlogic_0.dffrs_5.nand3_6.C.n8 SARlogic_0.dffrs_5.nand3_6.C.n7 6.04952
R6815 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_6.C.n1 5.7305
R6816 SARlogic_0.dffrs_5.nand3_2.B SARlogic_0.dffrs_5.nand3_6.C.n0 5.47979
R6817 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C.n3 5.13907
R6818 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n9 4.72925
R6819 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_6.C.n5 4.5005
R6820 SARlogic_0.dffrs_5.nand3_6.C.n9 SARlogic_0.dffrs_5.nand3_6.C.n8 0.732092
R6821 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t1 0.7285
R6822 SARlogic_0.dffrs_5.nand3_6.C.n7 SARlogic_0.dffrs_5.nand3_6.C.t2 0.7285
R6823 SARlogic_0.dffrs_5.nand3_1.Z SARlogic_0.dffrs_5.nand3_6.C.n6 0.449758
R6824 SARlogic_0.dffrs_5.nand3_6.C.n6 SARlogic_0.dffrs_5.nand3_2.B 0.166901
R6825 SARlogic_0.dffrs_5.nand3_6.C.n2 SARlogic_0.dffrs_5.nand3_0.A 0.0455
R6826 SARlogic_0.dffrs_5.nand3_6.C.n4 SARlogic_0.dffrs_5.nand3_6.C 0.0455
R6827 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t6 40.8177
R6828 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t5 40.6313
R6829 SARlogic_0.dffrs_12.nand3_8.C.n1 SARlogic_0.dffrs_12.nand3_8.C.t7 27.3166
R6830 SARlogic_0.dffrs_12.nand3_8.C.n0 SARlogic_0.dffrs_12.nand3_8.C.t4 27.1302
R6831 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_8.C.n2 14.119
R6832 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.t2 10.0473
R6833 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.t3 6.51042
R6834 SARlogic_0.dffrs_12.nand3_8.C.n5 SARlogic_0.dffrs_12.nand3_8.C.n4 6.04952
R6835 SARlogic_0.dffrs_12.nand3_7.B SARlogic_0.dffrs_12.nand3_8.C.n0 5.47979
R6836 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C.n1 5.13907
R6837 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n6 4.72925
R6838 SARlogic_0.dffrs_12.nand3_8.C.n6 SARlogic_0.dffrs_12.nand3_8.C.n5 0.732092
R6839 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t1 0.7285
R6840 SARlogic_0.dffrs_12.nand3_8.C.n4 SARlogic_0.dffrs_12.nand3_8.C.t0 0.7285
R6841 SARlogic_0.dffrs_12.nand3_8.C.n3 SARlogic_0.dffrs_12.nand3_7.B 0.438233
R6842 SARlogic_0.dffrs_12.nand3_6.Z SARlogic_0.dffrs_12.nand3_8.C.n3 0.166901
R6843 SARlogic_0.dffrs_12.nand3_8.C.n2 SARlogic_0.dffrs_12.nand3_8.C 0.0455
R6844 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t16 49.7997
R6845 comparator_no_offsetcal_0.x3.in comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t11 31.5367
R6846 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t9 19.735
R6847 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 18.0852
R6848 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t0 16.9998
R6849 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t15 14.5537
R6850 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 14.2885
R6851 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t17 13.6729
R6852 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t12 13.3844
R6853 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t14 13.3445
R6854 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 11.24
R6855 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 7.16477
R6856 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 6.95627
R6857 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 6.75194
R6858 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 6.32624
R6859 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t10 5.04666
R6860 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t13 4.84137
R6861 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 2.836
R6862 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n10 2.75432
R6863 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t2 1.8205
R6864 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t3 1.8205
R6865 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t5 1.8205
R6866 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t7 1.8205
R6867 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t1 0.8195
R6868 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t4 0.8195
R6869 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t8 0.8195
R6870 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.t6 0.8195
R6871 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n12 0.733357
R6872 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n6 0.440894
R6873 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n3 0.426875
R6874 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n4 0.289009
R6875 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n7 0.0607115
R6876 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1.n0 comparator_no_offsetcal_0.x3.in 0.014
R6877 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t16 49.7997
R6878 comparator_no_offsetcal_0.x5.in comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t12 31.5367
R6879 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t10 19.735
R6880 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t9 18.9075
R6881 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t1 16.9998
R6882 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t14 13.6729
R6883 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t11 13.3844
R6884 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t17 13.3445
R6885 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 12.247
R6886 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 11.2403
R6887 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 9.4181
R6888 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 7.4449
R6889 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 6.95074
R6890 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 6.75194
R6891 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 6.32761
R6892 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t15 5.04666
R6893 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 4.94262
R6894 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t13 4.84137
R6895 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 2.836
R6896 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n1 2.75432
R6897 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t7 1.8205
R6898 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t6 1.8205
R6899 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t8 1.8205
R6900 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t5 1.8205
R6901 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t2 0.8195
R6902 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t3 0.8195
R6903 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t4 0.8195
R6904 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.t0 0.8195
R6905 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n12 0.733357
R6906 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n7 0.5315
R6907 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n5 0.289009
R6908 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n9 0.184462
R6909 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2.n0 comparator_no_offsetcal_0.x5.in 0.014
R6910 Clk.n0 Clk.t23 41.0041
R6911 Clk.n22 Clk.t5 41.0041
R6912 Clk.n18 Clk.t24 41.0041
R6913 Clk.n14 Clk.t14 41.0041
R6914 Clk.n10 Clk.t1 41.0041
R6915 Clk.n6 Clk.t10 41.0041
R6916 Clk.n3 Clk.t28 41.0041
R6917 Clk.n1 Clk.t25 40.8177
R6918 Clk.n23 Clk.t8 40.8177
R6919 Clk.n19 Clk.t20 40.8177
R6920 Clk.n15 Clk.t17 40.8177
R6921 Clk.n11 Clk.t29 40.8177
R6922 Clk.n7 Clk.t6 40.8177
R6923 Clk.n4 Clk.t2 40.8177
R6924 Clk.n1 Clk.t19 27.1302
R6925 Clk.n23 Clk.t26 27.1302
R6926 Clk.n19 Clk.t4 27.1302
R6927 Clk.n15 Clk.t15 27.1302
R6928 Clk.n11 Clk.t32 27.1302
R6929 Clk.n7 Clk.t30 27.1302
R6930 Clk.n4 Clk.t13 27.1302
R6931 Clk.n0 Clk.t31 26.9438
R6932 Clk.n22 Clk.t16 26.9438
R6933 Clk.n18 Clk.t0 26.9438
R6934 Clk.n14 Clk.t21 26.9438
R6935 Clk.n10 Clk.t7 26.9438
R6936 Clk.n6 Clk.t18 26.9438
R6937 Clk.n3 Clk.t3 26.9438
R6938 Clk.n31 Clk.t12 21.1483
R6939 Clk.n30 Clk.t11 21.1483
R6940 Clk.n29 Clk.t22 21.1483
R6941 Clk.n28 Clk.t9 21.1483
R6942 Clk.n27 Clk.t27 20.5929
R6943 Clk.n9 SARlogic_0.dffrs_5.clk 20.5278
R6944 Clk.n28 Clk.n27 19.1491
R6945 Clk.n21 SARlogic_0.dffrs_1.clk 16.89
R6946 Clk.n17 SARlogic_0.dffrs_2.clk 16.89
R6947 Clk.n13 SARlogic_0.dffrs_3.clk 16.89
R6948 Clk.n9 SARlogic_0.dffrs_4.clk 16.89
R6949 Clk.n25 SARlogic_0.dffrs_0.clk 16.8417
R6950 Clk.n32 Clk.n31 15.5861
R6951 Clk.n26 SARlogic_0.dffrs_13.clk 12.2453
R6952 SARlogic_0.clk Clk.n33 11.0885
R6953 Clk.n26 Clk.n25 8.1113
R6954 SARlogic_0.dffrs_13.nand3_1.A Clk.n0 5.7755
R6955 SARlogic_0.dffrs_0.nand3_1.A Clk.n22 5.7755
R6956 SARlogic_0.dffrs_1.nand3_1.A Clk.n18 5.7755
R6957 SARlogic_0.dffrs_2.nand3_1.A Clk.n14 5.7755
R6958 SARlogic_0.dffrs_3.nand3_1.A Clk.n10 5.7755
R6959 SARlogic_0.dffrs_4.nand3_1.A Clk.n6 5.7755
R6960 SARlogic_0.dffrs_5.nand3_1.A Clk.n3 5.7755
R6961 SARlogic_0.dffrs_13.nand3_6.B Clk.n1 5.47979
R6962 SARlogic_0.dffrs_0.nand3_6.B Clk.n23 5.47979
R6963 SARlogic_0.dffrs_1.nand3_6.B Clk.n19 5.47979
R6964 SARlogic_0.dffrs_2.nand3_6.B Clk.n15 5.47979
R6965 SARlogic_0.dffrs_3.nand3_6.B Clk.n11 5.47979
R6966 SARlogic_0.dffrs_4.nand3_6.B Clk.n7 5.47979
R6967 SARlogic_0.dffrs_5.nand3_6.B Clk.n4 5.47979
R6968 Clk.n33 comparator_no_offsetcal_0.CLK 5.11456
R6969 Clk.n30 Clk.n29 4.47208
R6970 Clk.n13 Clk.n9 3.6383
R6971 Clk.n17 Clk.n13 3.6383
R6972 Clk.n21 Clk.n17 3.6383
R6973 Clk.n25 Clk.n21 3.6113
R6974 Clk.n32 Clk.n27 3.56405
R6975 Clk.n2 SARlogic_0.dffrs_13.nand3_6.B 2.17818
R6976 Clk.n24 SARlogic_0.dffrs_0.nand3_6.B 2.17818
R6977 Clk.n20 SARlogic_0.dffrs_1.nand3_6.B 2.17818
R6978 Clk.n16 SARlogic_0.dffrs_2.nand3_6.B 2.17818
R6979 Clk.n12 SARlogic_0.dffrs_3.nand3_6.B 2.17818
R6980 Clk.n8 SARlogic_0.dffrs_4.nand3_6.B 2.17818
R6981 Clk.n5 SARlogic_0.dffrs_5.nand3_6.B 2.17818
R6982 comparator_no_offsetcal_0.CLK Clk.n32 1.60543
R6983 Clk.n2 SARlogic_0.dffrs_13.nand3_1.A 1.34729
R6984 Clk.n24 SARlogic_0.dffrs_0.nand3_1.A 1.34729
R6985 Clk.n20 SARlogic_0.dffrs_1.nand3_1.A 1.34729
R6986 Clk.n16 SARlogic_0.dffrs_2.nand3_1.A 1.34729
R6987 Clk.n12 SARlogic_0.dffrs_3.nand3_1.A 1.34729
R6988 Clk.n8 SARlogic_0.dffrs_4.nand3_1.A 1.34729
R6989 Clk.n5 SARlogic_0.dffrs_5.nand3_1.A 1.34729
R6990 Clk.n29 Clk.n28 1.01892
R6991 Clk.n31 Clk.n30 1.01892
R6992 SARlogic_0.dffrs_13.clk Clk.n2 0.611214
R6993 SARlogic_0.dffrs_0.clk Clk.n24 0.611214
R6994 SARlogic_0.dffrs_1.clk Clk.n20 0.611214
R6995 SARlogic_0.dffrs_2.clk Clk.n16 0.611214
R6996 SARlogic_0.dffrs_3.clk Clk.n12 0.611214
R6997 SARlogic_0.dffrs_4.clk Clk.n8 0.611214
R6998 SARlogic_0.dffrs_5.clk Clk.n5 0.611214
R6999 Clk.n33 Clk 0.514034
R7000 SARlogic_0.clk Clk.n26 0.13775
R7001 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t8 41.0041
R7002 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t6 40.8177
R7003 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t7 40.6313
R7004 SARlogic_0.dffrs_1.nand3_6.C.n3 SARlogic_0.dffrs_1.nand3_6.C.t4 27.3166
R7005 SARlogic_0.dffrs_1.nand3_6.C.n0 SARlogic_0.dffrs_1.nand3_6.C.t9 27.1302
R7006 SARlogic_0.dffrs_1.nand3_6.C.n1 SARlogic_0.dffrs_1.nand3_6.C.t5 26.9438
R7007 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.t1 10.0473
R7008 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n4 9.90747
R7009 SARlogic_0.dffrs_1.nand3_6.C.n5 SARlogic_0.dffrs_1.nand3_6.C.n2 9.90116
R7010 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.t2 6.51042
R7011 SARlogic_0.dffrs_1.nand3_6.C.n8 SARlogic_0.dffrs_1.nand3_6.C.n7 6.04952
R7012 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_6.C.n1 5.7305
R7013 SARlogic_0.dffrs_1.nand3_2.B SARlogic_0.dffrs_1.nand3_6.C.n0 5.47979
R7014 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C.n3 5.13907
R7015 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n9 4.72925
R7016 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_6.C.n5 4.5005
R7017 SARlogic_0.dffrs_1.nand3_6.C.n9 SARlogic_0.dffrs_1.nand3_6.C.n8 0.732092
R7018 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t0 0.7285
R7019 SARlogic_0.dffrs_1.nand3_6.C.n7 SARlogic_0.dffrs_1.nand3_6.C.t3 0.7285
R7020 SARlogic_0.dffrs_1.nand3_1.Z SARlogic_0.dffrs_1.nand3_6.C.n6 0.449758
R7021 SARlogic_0.dffrs_1.nand3_6.C.n6 SARlogic_0.dffrs_1.nand3_2.B 0.166901
R7022 SARlogic_0.dffrs_1.nand3_6.C.n2 SARlogic_0.dffrs_1.nand3_0.A 0.0455
R7023 SARlogic_0.dffrs_1.nand3_6.C.n4 SARlogic_0.dffrs_1.nand3_6.C 0.0455
R7024 SARlogic_0.d2.n3 SARlogic_0.d2.t5 41.0041
R7025 SARlogic_0.d2.n4 SARlogic_0.d2.t11 40.8177
R7026 SARlogic_0.d2.n7 SARlogic_0.d2.t4 40.6313
R7027 SARlogic_0.d2.n1 SARlogic_0.d2.t6 34.2529
R7028 SARlogic_0.d2.n6 SARlogic_0.dffrs_8.clk 34.1594
R7029 SARlogic_0.d2.n7 SARlogic_0.d2.t10 27.3166
R7030 SARlogic_0.d2.n4 SARlogic_0.d2.t9 27.1302
R7031 SARlogic_0.d2.n3 SARlogic_0.d2.t7 26.9438
R7032 SARlogic_0.d2.n0 SARlogic_0.d2.t8 19.673
R7033 SARlogic_0.d2.n0 SARlogic_0.d2.t12 19.4007
R7034 SARlogic_0.d2 adc_PISO_0.B3 17.5376
R7035 SARlogic_0.d2.n9 SARlogic_0.d2.n8 14.0582
R7036 SARlogic_0.d2.n9 SARlogic_0.d2.n6 12.0118
R7037 SARlogic_0.d2.n12 SARlogic_0.d2.t0 10.0473
R7038 SARlogic_0.d2.n2 SARlogic_0.d2.n1 8.05164
R7039 SARlogic_0.d2.n11 SARlogic_0.d2.t1 6.51042
R7040 SARlogic_0.d2.n11 SARlogic_0.d2.n10 6.04952
R7041 SARlogic_0.dffrs_8.nand3_1.A SARlogic_0.d2.n3 5.7755
R7042 SARlogic_0.dffrs_8.nand3_6.B SARlogic_0.d2.n4 5.47979
R7043 SARlogic_0.d2.n8 SARlogic_0.d2.n7 5.13907
R7044 SARlogic_0.dffrs_9.nand3_2.Z SARlogic_0.d2.n12 4.72925
R7045 SARlogic_0.d2.n5 SARlogic_0.dffrs_8.nand3_6.B 2.17818
R7046 adc_PISO_0.B3 SARlogic_0.d2.n2 1.87121
R7047 SARlogic_0.d2.n5 SARlogic_0.dffrs_8.nand3_1.A 1.34729
R7048 SARlogic_0.d2.n12 SARlogic_0.d2.n11 0.732092
R7049 SARlogic_0.d2.n10 SARlogic_0.d2.t3 0.7285
R7050 SARlogic_0.d2.n10 SARlogic_0.d2.t2 0.7285
R7051 SARlogic_0.d2.n6 SARlogic_0.d2 0.698
R7052 SARlogic_0.dffrs_8.clk SARlogic_0.d2.n5 0.610571
R7053 SARlogic_0.dffrs_9.nand3_2.Z SARlogic_0.d2.n9 0.166901
R7054 SARlogic_0.d2.n1 SARlogic_0.d2.n0 0.106438
R7055 SARlogic_0.d2.n8 SARlogic_0.dffrs_9.nand3_7.C 0.0455
R7056 SARlogic_0.d2.n2 adc_PISO_0.2inmux_4.In 0.0455
R7057 a_4841_31422.n1 a_4841_31422.t4 41.0041
R7058 a_4841_31422.n0 a_4841_31422.t6 40.8177
R7059 a_4841_31422.n2 a_4841_31422.t7 40.6313
R7060 a_4841_31422.n2 a_4841_31422.t9 27.3166
R7061 a_4841_31422.n0 a_4841_31422.t8 27.1302
R7062 a_4841_31422.n1 a_4841_31422.t5 26.9438
R7063 a_4841_31422.n3 a_4841_31422.n1 15.6312
R7064 a_4841_31422.n3 a_4841_31422.n2 15.046
R7065 a_4841_31422.n5 a_4841_31422.t2 10.0473
R7066 a_4841_31422.t0 a_4841_31422.n7 6.51042
R7067 a_4841_31422.n7 a_4841_31422.n6 6.04952
R7068 a_4841_31422.n4 a_4841_31422.n0 5.64619
R7069 a_4841_31422.n5 a_4841_31422.n4 5.17851
R7070 a_4841_31422.n4 a_4841_31422.n3 4.5005
R7071 a_4841_31422.n7 a_4841_31422.n5 0.732092
R7072 a_4841_31422.n6 a_4841_31422.t3 0.7285
R7073 a_4841_31422.n6 a_4841_31422.t1 0.7285
R7074 a_4841_33627.n0 a_4841_33627.t4 40.6313
R7075 a_4841_33627.n0 a_4841_33627.t5 27.3166
R7076 a_4841_33627.n1 a_4841_33627.n0 24.1527
R7077 a_4841_33627.n1 a_4841_33627.t2 10.0473
R7078 a_4841_33627.n2 a_4841_33627.t3 6.51042
R7079 a_4841_33627.n3 a_4841_33627.n2 6.04952
R7080 a_4841_33627.n2 a_4841_33627.n1 0.732092
R7081 a_4841_33627.t0 a_4841_33627.n3 0.7285
R7082 a_4841_33627.n3 a_4841_33627.t1 0.7285
R7083 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t6 40.6313
R7084 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.t4 34.1066
R7085 adc_PISO_0.2inmux_1.Bit.n3 adc_PISO_0.2inmux_1.Bit.t7 27.3166
R7086 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t5 19.673
R7087 adc_PISO_0.2inmux_1.Bit.n0 adc_PISO_0.2inmux_1.Bit.t8 19.4007
R7088 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n3 14.6967
R7089 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.t2 10.0473
R7090 adc_PISO_0.2inmux_1.Bit.n7 adc_PISO_0.2inmux_1.Bit.n6 9.39565
R7091 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit.n1 6.70486
R7092 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.t3 6.51042
R7093 adc_PISO_0.2inmux_1.Bit.n5 adc_PISO_0.2inmux_1.Bit.n4 6.04952
R7094 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n2 5.81514
R7095 adc_PISO_0.2inmux_1.Bit.n6 adc_PISO_0.2inmux_1.Bit.n5 0.732092
R7096 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t0 0.7285
R7097 adc_PISO_0.2inmux_1.Bit.n4 adc_PISO_0.2inmux_1.Bit.t1 0.7285
R7098 adc_PISO_0.dffrs_4.Q adc_PISO_0.2inmux_1.Bit.n7 0.458082
R7099 adc_PISO_0.2inmux_1.Bit.n1 adc_PISO_0.2inmux_1.Bit.n0 0.252687
R7100 adc_PISO_0.2inmux_1.Bit.n2 adc_PISO_0.2inmux_1.Bit 0.0519286
R7101 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t4 40.6313
R7102 SARlogic_0.dffrs_5.nand3_1.C.n0 SARlogic_0.dffrs_5.nand3_1.C.t5 27.3166
R7103 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n1 14.2854
R7104 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.t0 10.0473
R7105 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.t1 6.51042
R7106 SARlogic_0.dffrs_5.nand3_1.C.n3 SARlogic_0.dffrs_5.nand3_1.C.n2 6.04952
R7107 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C.n0 5.13907
R7108 SARlogic_0.dffrs_5.nand3_0.Z SARlogic_0.dffrs_5.nand3_1.C.n4 4.72925
R7109 SARlogic_0.dffrs_5.nand3_1.C.n4 SARlogic_0.dffrs_5.nand3_1.C.n3 0.732092
R7110 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t2 0.7285
R7111 SARlogic_0.dffrs_5.nand3_1.C.n2 SARlogic_0.dffrs_5.nand3_1.C.t3 0.7285
R7112 SARlogic_0.dffrs_5.nand3_1.C.n1 SARlogic_0.dffrs_5.nand3_1.C 0.0455
R7113 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t5 41.0041
R7114 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t6 40.8177
R7115 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t4 40.6313
R7116 SARlogic_0.dffrs_3.nand3_6.C.n3 SARlogic_0.dffrs_3.nand3_6.C.t9 27.3166
R7117 SARlogic_0.dffrs_3.nand3_6.C.n0 SARlogic_0.dffrs_3.nand3_6.C.t7 27.1302
R7118 SARlogic_0.dffrs_3.nand3_6.C.n1 SARlogic_0.dffrs_3.nand3_6.C.t8 26.9438
R7119 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.t1 10.0473
R7120 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n4 9.90747
R7121 SARlogic_0.dffrs_3.nand3_6.C.n5 SARlogic_0.dffrs_3.nand3_6.C.n2 9.90116
R7122 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.t2 6.51042
R7123 SARlogic_0.dffrs_3.nand3_6.C.n8 SARlogic_0.dffrs_3.nand3_6.C.n7 6.04952
R7124 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_6.C.n1 5.7305
R7125 SARlogic_0.dffrs_3.nand3_2.B SARlogic_0.dffrs_3.nand3_6.C.n0 5.47979
R7126 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C.n3 5.13907
R7127 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n9 4.72925
R7128 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_6.C.n5 4.5005
R7129 SARlogic_0.dffrs_3.nand3_6.C.n9 SARlogic_0.dffrs_3.nand3_6.C.n8 0.732092
R7130 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t0 0.7285
R7131 SARlogic_0.dffrs_3.nand3_6.C.n7 SARlogic_0.dffrs_3.nand3_6.C.t3 0.7285
R7132 SARlogic_0.dffrs_3.nand3_1.Z SARlogic_0.dffrs_3.nand3_6.C.n6 0.449758
R7133 SARlogic_0.dffrs_3.nand3_6.C.n6 SARlogic_0.dffrs_3.nand3_2.B 0.166901
R7134 SARlogic_0.dffrs_3.nand3_6.C.n2 SARlogic_0.dffrs_3.nand3_0.A 0.0455
R7135 SARlogic_0.dffrs_3.nand3_6.C.n4 SARlogic_0.dffrs_3.nand3_6.C 0.0455
R7136 a_33337_30170.n0 a_33337_30170.t7 41.0041
R7137 a_33337_30170.n1 a_33337_30170.t4 40.8177
R7138 a_33337_30170.n1 a_33337_30170.t6 27.1302
R7139 a_33337_30170.n0 a_33337_30170.t5 26.9438
R7140 a_33337_30170.n2 a_33337_30170.n1 22.5284
R7141 a_33337_30170.n3 a_33337_30170.n2 19.5781
R7142 a_33337_30170.n3 a_33337_30170.t2 10.0473
R7143 a_33337_30170.t0 a_33337_30170.n5 6.51042
R7144 a_33337_30170.n5 a_33337_30170.n4 6.04952
R7145 a_33337_30170.n2 a_33337_30170.n0 5.7305
R7146 a_33337_30170.n5 a_33337_30170.n3 0.732092
R7147 a_33337_30170.n4 a_33337_30170.t3 0.7285
R7148 a_33337_30170.n4 a_33337_30170.t1 0.7285
R7149 a_33257_33628.n2 a_33257_33628.t4 40.6313
R7150 a_33257_33628.n2 a_33257_33628.t5 27.3166
R7151 a_33257_33628.n3 a_33257_33628.n2 24.1527
R7152 a_33257_33628.t0 a_33257_33628.n3 10.0473
R7153 a_33257_33628.n1 a_33257_33628.t1 6.51042
R7154 a_33257_33628.n1 a_33257_33628.n0 6.04952
R7155 a_33257_33628.n3 a_33257_33628.n1 0.732092
R7156 a_33257_33628.n0 a_33257_33628.t2 0.7285
R7157 a_33257_33628.n0 a_33257_33628.t3 0.7285
R7158 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t5 41.0041
R7159 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t4 40.6313
R7160 SARlogic_0.dffrs_0.d.n1 SARlogic_0.dffrs_0.d.t6 27.3166
R7161 SARlogic_0.dffrs_0.d.n0 SARlogic_0.dffrs_0.d.t7 26.9438
R7162 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d 17.5022
R7163 SARlogic_0.dffrs_0.d.n3 SARlogic_0.dffrs_0.d.n2 14.0582
R7164 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.t3 10.0473
R7165 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.t2 6.51042
R7166 SARlogic_0.dffrs_0.d.n5 SARlogic_0.dffrs_0.d.n4 6.04952
R7167 SARlogic_0.dffrs_0.nand3_8.A SARlogic_0.dffrs_0.d.n0 5.7755
R7168 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_0.d.n1 5.13907
R7169 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n6 4.72925
R7170 SARlogic_0.dffrs_0.d SARlogic_0.dffrs_0.nand3_8.A 0.783821
R7171 SARlogic_0.dffrs_0.d.n6 SARlogic_0.dffrs_0.d.n5 0.732092
R7172 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t1 0.7285
R7173 SARlogic_0.dffrs_0.d.n4 SARlogic_0.dffrs_0.d.t0 0.7285
R7174 SARlogic_0.dffrs_13.nand3_2.Z SARlogic_0.dffrs_0.d.n3 0.166901
R7175 SARlogic_0.dffrs_0.d.n2 SARlogic_0.dffrs_13.nand3_7.C 0.0455
R7176 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t7 41.0041
R7177 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t4 40.6313
R7178 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t8 40.6313
R7179 SARlogic_0.dffrs_13.Qb SARlogic_0.dffrs_14.setb 27.9776
R7180 SARlogic_0.dffrs_13.Qb.n4 SARlogic_0.dffrs_13.Qb.t6 27.3166
R7181 SARlogic_0.dffrs_13.Qb.n2 SARlogic_0.dffrs_13.Qb.t5 27.3166
R7182 SARlogic_0.dffrs_13.Qb.n0 SARlogic_0.dffrs_13.Qb.t9 26.9438
R7183 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.t2 10.0473
R7184 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb.n1 9.84255
R7185 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n3 9.22229
R7186 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.t3 6.51042
R7187 SARlogic_0.dffrs_13.Qb.n8 SARlogic_0.dffrs_13.Qb.n7 6.04952
R7188 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.Qb.n0 5.7305
R7189 SARlogic_0.dffrs_13.Qb.n5 SARlogic_0.dffrs_13.Qb.n4 5.14711
R7190 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_13.Qb.n2 5.13907
R7191 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n6 4.94976
R7192 SARlogic_0.dffrs_13.nand3_7.Z SARlogic_0.dffrs_13.Qb.n9 4.72925
R7193 SARlogic_0.dffrs_14.setb SARlogic_0.dffrs_14.nand3_0.C 0.784786
R7194 SARlogic_0.dffrs_13.Qb.n9 SARlogic_0.dffrs_13.Qb.n8 0.732092
R7195 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t0 0.7285
R7196 SARlogic_0.dffrs_13.Qb.n7 SARlogic_0.dffrs_13.Qb.t1 0.7285
R7197 SARlogic_0.dffrs_13.Qb.n6 SARlogic_0.dffrs_13.Qb 0.175225
R7198 SARlogic_0.dffrs_13.Qb.n1 SARlogic_0.dffrs_13.nand3_2.A 0.0455
R7199 SARlogic_0.dffrs_13.Qb.n3 SARlogic_0.dffrs_14.nand3_2.C 0.0455
R7200 SARlogic_0.dffrs_14.nand3_0.C SARlogic_0.dffrs_13.Qb.n5 0.0374643
R7201 Comp_out.n0 Comp_out 11.2807
R7202 Comp_out.n6 Comp_out.n5 6.5435
R7203 Comp_out.n3 Comp_out.n2 6.5435
R7204 comparator_no_offsetcal_0.x4.Y Comp_out.n9 4.5005
R7205 comparator_no_offsetcal_0.x4.Y Comp_out.n0 2.3842
R7206 Comp_out.n7 Comp_out.n4 2.17483
R7207 Comp_out.n5 Comp_out.t1 2.03874
R7208 Comp_out.n5 Comp_out.t2 2.03874
R7209 Comp_out.n2 Comp_out.t0 2.03874
R7210 Comp_out.n2 Comp_out.t3 2.03874
R7211 Comp_out.n9 Comp_out.n1 2.00383
R7212 Comp_out.n1 Comp_out.t7 1.13285
R7213 Comp_out.n1 Comp_out.t6 1.13285
R7214 Comp_out.n4 Comp_out.t4 1.13285
R7215 Comp_out.n4 Comp_out.t5 1.13285
R7216 Comp_out.n6 Comp_out.n3 0.5105
R7217 Comp_out.n8 Comp_out.n7 0.5105
R7218 Comp_out.n0 comparator_no_offsetcal_0.Vout 0.3995
R7219 Comp_out.n8 Comp_out.n3 0.2165
R7220 Comp_out.n7 Comp_out.n6 0.2165
R7221 Comp_out.n9 Comp_out.n8 0.1175
R7222 a_9083_28820.n0 a_9083_28820.t4 34.1797
R7223 a_9083_28820.n0 a_9083_28820.t5 19.5798
R7224 a_9083_28820.n1 a_9083_28820.t2 18.7717
R7225 a_9083_28820.n1 a_9083_28820.t1 9.2885
R7226 a_9083_28820.n2 a_9083_28820.n0 4.93379
R7227 a_9083_28820.t0 a_9083_28820.n3 4.23346
R7228 a_9083_28820.n3 a_9083_28820.t3 3.85546
R7229 a_9083_28820.n2 a_9083_28820.n1 0.4055
R7230 a_9083_28820.n3 a_9083_28820.n2 0.352625
R7231 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t7 41.0041
R7232 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t8 40.8177
R7233 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t6 40.6313
R7234 SARlogic_0.dffrs_9.nand3_6.C.n3 SARlogic_0.dffrs_9.nand3_6.C.t5 27.3166
R7235 SARlogic_0.dffrs_9.nand3_6.C.n0 SARlogic_0.dffrs_9.nand3_6.C.t4 27.1302
R7236 SARlogic_0.dffrs_9.nand3_6.C.n1 SARlogic_0.dffrs_9.nand3_6.C.t9 26.9438
R7237 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.t0 10.0473
R7238 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n4 9.90747
R7239 SARlogic_0.dffrs_9.nand3_6.C.n5 SARlogic_0.dffrs_9.nand3_6.C.n2 9.90116
R7240 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.t1 6.51042
R7241 SARlogic_0.dffrs_9.nand3_6.C.n8 SARlogic_0.dffrs_9.nand3_6.C.n7 6.04952
R7242 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_6.C.n1 5.7305
R7243 SARlogic_0.dffrs_9.nand3_2.B SARlogic_0.dffrs_9.nand3_6.C.n0 5.47979
R7244 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C.n3 5.13907
R7245 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n9 4.72925
R7246 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_6.C.n5 4.5005
R7247 SARlogic_0.dffrs_9.nand3_6.C.n9 SARlogic_0.dffrs_9.nand3_6.C.n8 0.732092
R7248 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t2 0.7285
R7249 SARlogic_0.dffrs_9.nand3_6.C.n7 SARlogic_0.dffrs_9.nand3_6.C.t3 0.7285
R7250 SARlogic_0.dffrs_9.nand3_1.Z SARlogic_0.dffrs_9.nand3_6.C.n6 0.449758
R7251 SARlogic_0.dffrs_9.nand3_6.C.n6 SARlogic_0.dffrs_9.nand3_2.B 0.166901
R7252 SARlogic_0.dffrs_9.nand3_6.C.n2 SARlogic_0.dffrs_9.nand3_0.A 0.0455
R7253 SARlogic_0.dffrs_9.nand3_6.C.n4 SARlogic_0.dffrs_9.nand3_6.C 0.0455
R7254 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t6 40.8177
R7255 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t7 40.6313
R7256 SARlogic_0.dffrs_2.nand3_8.C.n1 SARlogic_0.dffrs_2.nand3_8.C.t4 27.3166
R7257 SARlogic_0.dffrs_2.nand3_8.C.n0 SARlogic_0.dffrs_2.nand3_8.C.t5 27.1302
R7258 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_8.C.n2 14.119
R7259 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.t2 10.0473
R7260 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.t1 6.51042
R7261 SARlogic_0.dffrs_2.nand3_8.C.n5 SARlogic_0.dffrs_2.nand3_8.C.n4 6.04952
R7262 SARlogic_0.dffrs_2.nand3_7.B SARlogic_0.dffrs_2.nand3_8.C.n0 5.47979
R7263 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C.n1 5.13907
R7264 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n6 4.72925
R7265 SARlogic_0.dffrs_2.nand3_8.C.n6 SARlogic_0.dffrs_2.nand3_8.C.n5 0.732092
R7266 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t0 0.7285
R7267 SARlogic_0.dffrs_2.nand3_8.C.n4 SARlogic_0.dffrs_2.nand3_8.C.t3 0.7285
R7268 SARlogic_0.dffrs_2.nand3_8.C.n3 SARlogic_0.dffrs_2.nand3_7.B 0.438233
R7269 SARlogic_0.dffrs_2.nand3_6.Z SARlogic_0.dffrs_2.nand3_8.C.n3 0.166901
R7270 SARlogic_0.dffrs_2.nand3_8.C.n2 SARlogic_0.dffrs_2.nand3_8.C 0.0455
R7271 a_30255_29264.n0 a_30255_29264.t5 34.1797
R7272 a_30255_29264.n0 a_30255_29264.t4 19.5798
R7273 a_30255_29264.t0 a_30255_29264.n3 10.3401
R7274 a_30255_29264.n3 a_30255_29264.t1 9.2885
R7275 a_30255_29264.n2 a_30255_29264.n0 4.93379
R7276 a_30255_29264.n1 a_30255_29264.t2 4.09202
R7277 a_30255_29264.n1 a_30255_29264.t3 3.95079
R7278 a_30255_29264.n3 a_30255_29264.n2 0.599711
R7279 a_30255_29264.n2 a_30255_29264.n1 0.296375
R7280 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t3 41.0041
R7281 adc_PISO_0.2inmux_5.OUT.n0 adc_PISO_0.2inmux_5.OUT.t2 26.9438
R7282 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t0 9.6935
R7283 adc_PISO_0.dffrs_4.d adc_PISO_0.2inmux_5.OUT.n0 6.55979
R7284 adc_PISO_0.2inmux_5.OUT adc_PISO_0.dffrs_4.d 4.883
R7285 adc_PISO_0.2inmux_5.OUT.n1 adc_PISO_0.2inmux_5.OUT.t1 4.35383
R7286 adc_PISO_0.2inmux_5.OUT adc_PISO_0.2inmux_5.OUT.n1 0.350857
R7287 SARlogic_0.d0.n3 SARlogic_0.d0.t4 41.0041
R7288 SARlogic_0.d0.n4 SARlogic_0.d0.t10 40.8177
R7289 SARlogic_0.d0.n7 SARlogic_0.d0.t5 40.6313
R7290 SARlogic_0.d0.n6 adc_PISO_0.B1 36.2544
R7291 SARlogic_0.d0.n1 SARlogic_0.d0.t9 34.2529
R7292 SARlogic_0.d0.n6 SARlogic_0.dffrs_10.clk 33.5936
R7293 SARlogic_0.d0.n7 SARlogic_0.d0.t12 27.3166
R7294 SARlogic_0.d0.n4 SARlogic_0.d0.t7 27.1302
R7295 SARlogic_0.d0.n3 SARlogic_0.d0.t6 26.9438
R7296 SARlogic_0.d0.n0 SARlogic_0.d0.t11 19.673
R7297 SARlogic_0.d0.n0 SARlogic_0.d0.t8 19.4007
R7298 SARlogic_0.d0.n9 SARlogic_0.d0.n8 14.0582
R7299 SARlogic_0.d0.n9 SARlogic_0.d0.n6 11.4461
R7300 SARlogic_0.d0.n12 SARlogic_0.d0.t0 10.0473
R7301 SARlogic_0.d0.n2 SARlogic_0.d0.n1 8.05164
R7302 SARlogic_0.d0.n11 SARlogic_0.d0.t1 6.51042
R7303 SARlogic_0.d0.n11 SARlogic_0.d0.n10 6.04952
R7304 SARlogic_0.dffrs_10.nand3_1.A SARlogic_0.d0.n3 5.7755
R7305 SARlogic_0.dffrs_10.nand3_6.B SARlogic_0.d0.n4 5.47979
R7306 SARlogic_0.d0.n8 SARlogic_0.d0.n7 5.13907
R7307 SARlogic_0.dffrs_11.nand3_2.Z SARlogic_0.d0.n12 4.72925
R7308 SARlogic_0.d0.n5 SARlogic_0.dffrs_10.nand3_6.B 2.17818
R7309 adc_PISO_0.B1 SARlogic_0.d0.n2 1.87121
R7310 SARlogic_0.d0.n5 SARlogic_0.dffrs_10.nand3_1.A 1.34729
R7311 SARlogic_0.d0.n12 SARlogic_0.d0.n11 0.732092
R7312 SARlogic_0.d0.n10 SARlogic_0.d0.t2 0.7285
R7313 SARlogic_0.d0.n10 SARlogic_0.d0.t3 0.7285
R7314 SARlogic_0.dffrs_10.clk SARlogic_0.d0.n5 0.610571
R7315 SARlogic_0.dffrs_11.nand3_2.Z SARlogic_0.d0.n9 0.166901
R7316 SARlogic_0.d0.n1 SARlogic_0.d0.n0 0.106438
R7317 SARlogic_0.d0.n8 SARlogic_0.dffrs_11.nand3_7.C 0.0455
R7318 SARlogic_0.d0.n2 adc_PISO_0.2inmux_1.In 0.0455
R7319 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t4 41.0041
R7320 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t5 40.8177
R7321 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t9 40.6313
R7322 SARlogic_0.dffrs_10.nand3_6.C.n3 SARlogic_0.dffrs_10.nand3_6.C.t8 27.3166
R7323 SARlogic_0.dffrs_10.nand3_6.C.n0 SARlogic_0.dffrs_10.nand3_6.C.t7 27.1302
R7324 SARlogic_0.dffrs_10.nand3_6.C.n1 SARlogic_0.dffrs_10.nand3_6.C.t6 26.9438
R7325 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.t2 10.0473
R7326 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n4 9.90747
R7327 SARlogic_0.dffrs_10.nand3_6.C.n5 SARlogic_0.dffrs_10.nand3_6.C.n2 9.90116
R7328 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.t3 6.51042
R7329 SARlogic_0.dffrs_10.nand3_6.C.n8 SARlogic_0.dffrs_10.nand3_6.C.n7 6.04952
R7330 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_6.C.n1 5.7305
R7331 SARlogic_0.dffrs_10.nand3_2.B SARlogic_0.dffrs_10.nand3_6.C.n0 5.47979
R7332 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C.n3 5.13907
R7333 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n9 4.72925
R7334 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_6.C.n5 4.5005
R7335 SARlogic_0.dffrs_10.nand3_6.C.n9 SARlogic_0.dffrs_10.nand3_6.C.n8 0.732092
R7336 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t0 0.7285
R7337 SARlogic_0.dffrs_10.nand3_6.C.n7 SARlogic_0.dffrs_10.nand3_6.C.t1 0.7285
R7338 SARlogic_0.dffrs_10.nand3_1.Z SARlogic_0.dffrs_10.nand3_6.C.n6 0.449758
R7339 SARlogic_0.dffrs_10.nand3_6.C.n6 SARlogic_0.dffrs_10.nand3_2.B 0.166901
R7340 SARlogic_0.dffrs_10.nand3_6.C.n2 SARlogic_0.dffrs_10.nand3_0.A 0.0455
R7341 SARlogic_0.dffrs_10.nand3_6.C.n4 SARlogic_0.dffrs_10.nand3_6.C 0.0455
R7342 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t8 41.0041
R7343 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t5 40.6313
R7344 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t4 40.6313
R7345 SARlogic_0.dffrs_3.Qb SARlogic_0.dffrs_10.setb 28.021
R7346 SARlogic_0.dffrs_3.Qb.n4 SARlogic_0.dffrs_3.Qb.t7 27.3166
R7347 SARlogic_0.dffrs_3.Qb.n2 SARlogic_0.dffrs_3.Qb.t6 27.3166
R7348 SARlogic_0.dffrs_3.Qb.n0 SARlogic_0.dffrs_3.Qb.t9 26.9438
R7349 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.t0 10.0473
R7350 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb.n1 9.84255
R7351 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n3 9.22229
R7352 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.t1 6.51042
R7353 SARlogic_0.dffrs_3.Qb.n8 SARlogic_0.dffrs_3.Qb.n7 6.04952
R7354 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.Qb.n0 5.7305
R7355 SARlogic_0.dffrs_3.Qb.n5 SARlogic_0.dffrs_3.Qb.n4 5.14711
R7356 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_3.Qb.n2 5.13907
R7357 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n6 4.94976
R7358 SARlogic_0.dffrs_3.nand3_7.Z SARlogic_0.dffrs_3.Qb.n9 4.72925
R7359 SARlogic_0.dffrs_10.setb SARlogic_0.dffrs_10.nand3_0.C 0.784786
R7360 SARlogic_0.dffrs_3.Qb.n9 SARlogic_0.dffrs_3.Qb.n8 0.732092
R7361 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t3 0.7285
R7362 SARlogic_0.dffrs_3.Qb.n7 SARlogic_0.dffrs_3.Qb.t2 0.7285
R7363 SARlogic_0.dffrs_3.Qb.n6 SARlogic_0.dffrs_3.Qb 0.175225
R7364 SARlogic_0.dffrs_3.Qb.n1 SARlogic_0.dffrs_3.nand3_2.A 0.0455
R7365 SARlogic_0.dffrs_3.Qb.n3 SARlogic_0.dffrs_10.nand3_2.C 0.0455
R7366 SARlogic_0.dffrs_10.nand3_0.C SARlogic_0.dffrs_3.Qb.n5 0.0374643
R7367 a_14313_33628.n2 a_14313_33628.t5 40.6313
R7368 a_14313_33628.n2 a_14313_33628.t4 27.3166
R7369 a_14313_33628.n3 a_14313_33628.n2 24.1527
R7370 a_14313_33628.t0 a_14313_33628.n3 10.0473
R7371 a_14313_33628.n1 a_14313_33628.t2 6.51042
R7372 a_14313_33628.n1 a_14313_33628.n0 6.04952
R7373 a_14313_33628.n3 a_14313_33628.n1 0.732092
R7374 a_14313_33628.n0 a_14313_33628.t3 0.7285
R7375 a_14313_33628.n0 a_14313_33628.t1 0.7285
R7376 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t8 41.0041
R7377 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t4 40.6313
R7378 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t5 40.6313
R7379 SARlogic_0.dffrs_5.Qb SARlogic_0.dffrs_12.setb 28.013
R7380 SARlogic_0.dffrs_5.Qb.n4 SARlogic_0.dffrs_5.Qb.t6 27.3166
R7381 SARlogic_0.dffrs_5.Qb.n2 SARlogic_0.dffrs_5.Qb.t7 27.3166
R7382 SARlogic_0.dffrs_5.Qb.n0 SARlogic_0.dffrs_5.Qb.t9 26.9438
R7383 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.t0 10.0473
R7384 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb.n1 9.84255
R7385 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n3 9.22229
R7386 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.t1 6.51042
R7387 SARlogic_0.dffrs_5.Qb.n8 SARlogic_0.dffrs_5.Qb.n7 6.04952
R7388 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.Qb.n0 5.7305
R7389 SARlogic_0.dffrs_5.Qb.n5 SARlogic_0.dffrs_5.Qb.n4 5.14711
R7390 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_5.Qb.n2 5.13907
R7391 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n6 4.94976
R7392 SARlogic_0.dffrs_5.nand3_7.Z SARlogic_0.dffrs_5.Qb.n9 4.72925
R7393 SARlogic_0.dffrs_12.setb SARlogic_0.dffrs_12.nand3_0.C 0.784786
R7394 SARlogic_0.dffrs_5.Qb.n9 SARlogic_0.dffrs_5.Qb.n8 0.732092
R7395 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t3 0.7285
R7396 SARlogic_0.dffrs_5.Qb.n7 SARlogic_0.dffrs_5.Qb.t2 0.7285
R7397 SARlogic_0.dffrs_5.Qb.n6 SARlogic_0.dffrs_5.Qb 0.175225
R7398 SARlogic_0.dffrs_5.Qb.n1 SARlogic_0.dffrs_5.nand3_2.A 0.0455
R7399 SARlogic_0.dffrs_5.Qb.n3 SARlogic_0.dffrs_12.nand3_2.C 0.0455
R7400 SARlogic_0.dffrs_12.nand3_0.C SARlogic_0.dffrs_5.Qb.n5 0.0374643
R7401 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t4 40.6313
R7402 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.t8 34.1066
R7403 adc_PISO_0.dffrs_1.Q.n3 adc_PISO_0.dffrs_1.Q.t5 27.3166
R7404 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t6 19.673
R7405 adc_PISO_0.dffrs_1.Q.n0 adc_PISO_0.dffrs_1.Q.t7 19.4007
R7406 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n3 14.6967
R7407 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.t0 10.0473
R7408 adc_PISO_0.dffrs_1.Q.n7 adc_PISO_0.dffrs_1.Q.n6 9.39565
R7409 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.dffrs_1.Q.n1 6.70486
R7410 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.t1 6.51042
R7411 adc_PISO_0.dffrs_1.Q.n5 adc_PISO_0.dffrs_1.Q.n4 6.04952
R7412 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n2 5.81354
R7413 adc_PISO_0.dffrs_1.Q.n6 adc_PISO_0.dffrs_1.Q.n5 0.732092
R7414 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t3 0.7285
R7415 adc_PISO_0.dffrs_1.Q.n4 adc_PISO_0.dffrs_1.Q.t2 0.7285
R7416 adc_PISO_0.dffrs_1.Q adc_PISO_0.dffrs_1.Q.n7 0.458082
R7417 adc_PISO_0.dffrs_1.Q.n1 adc_PISO_0.dffrs_1.Q.n0 0.252687
R7418 adc_PISO_0.dffrs_1.Q.n2 adc_PISO_0.2inmux_3.Bit 0.0519286
R7419 SARlogic_0.d5.n3 SARlogic_0.d5.t4 40.6313
R7420 SARlogic_0.d5.n1 SARlogic_0.d5.t6 34.2529
R7421 SARlogic_0.d5.n3 SARlogic_0.d5.t8 27.3166
R7422 SARlogic_0.d5.n5 adc_PISO_0.B6 23.5656
R7423 SARlogic_0.d5.n0 SARlogic_0.d5.t7 19.673
R7424 SARlogic_0.d5.n0 SARlogic_0.d5.t5 19.4007
R7425 SARlogic_0.d5.n5 SARlogic_0.d5.n4 14.0582
R7426 SARlogic_0.d5.n8 SARlogic_0.d5.t1 10.0473
R7427 SARlogic_0.d5.n2 SARlogic_0.d5.n1 8.05164
R7428 SARlogic_0.d5.n7 SARlogic_0.d5.t2 6.51042
R7429 SARlogic_0.d5.n7 SARlogic_0.d5.n6 6.04952
R7430 SARlogic_0.d5.n4 SARlogic_0.d5.n3 5.13907
R7431 SARlogic_0.dffrs_14.nand3_2.Z SARlogic_0.d5.n8 4.72925
R7432 adc_PISO_0.B6 SARlogic_0.d5.n2 1.87121
R7433 SARlogic_0.d5.n8 SARlogic_0.d5.n7 0.732092
R7434 SARlogic_0.d5.n6 SARlogic_0.d5.t0 0.7285
R7435 SARlogic_0.d5.n6 SARlogic_0.d5.t3 0.7285
R7436 SARlogic_0.dffrs_14.nand3_2.Z SARlogic_0.d5.n5 0.166901
R7437 SARlogic_0.d5.n1 SARlogic_0.d5.n0 0.106438
R7438 SARlogic_0.d5.n4 SARlogic_0.dffrs_14.nand3_7.C 0.0455
R7439 SARlogic_0.d5.n2 adc_PISO_0.2inmux_0.In 0.0455
R7440 a_33257_29218.n0 a_33257_29218.t4 40.8177
R7441 a_33257_29218.n1 a_33257_29218.t7 40.6313
R7442 a_33257_29218.n1 a_33257_29218.t6 27.3166
R7443 a_33257_29218.n0 a_33257_29218.t5 27.1302
R7444 a_33257_29218.n2 a_33257_29218.n1 19.2576
R7445 a_33257_29218.n3 a_33257_29218.t2 10.0473
R7446 a_33257_29218.n4 a_33257_29218.t3 6.51042
R7447 a_33257_29218.n5 a_33257_29218.n4 6.04952
R7448 a_33257_29218.n2 a_33257_29218.n0 5.91752
R7449 a_33257_29218.n3 a_33257_29218.n2 4.89565
R7450 a_33257_29218.n4 a_33257_29218.n3 0.732092
R7451 a_33257_29218.t0 a_33257_29218.n5 0.7285
R7452 a_33257_29218.n5 a_33257_29218.t1 0.7285
R7453 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t5 41.0041
R7454 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t6 40.6313
R7455 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t4 40.6313
R7456 SARlogic_0.dffrs_0.Qb SARlogic_0.dffrs_7.setb 28.021
R7457 SARlogic_0.dffrs_0.Qb.n4 SARlogic_0.dffrs_0.Qb.t9 27.3166
R7458 SARlogic_0.dffrs_0.Qb.n2 SARlogic_0.dffrs_0.Qb.t7 27.3166
R7459 SARlogic_0.dffrs_0.Qb.n0 SARlogic_0.dffrs_0.Qb.t8 26.9438
R7460 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.t3 10.0473
R7461 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb.n1 9.84255
R7462 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n3 9.22229
R7463 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.t2 6.51042
R7464 SARlogic_0.dffrs_0.Qb.n8 SARlogic_0.dffrs_0.Qb.n7 6.04952
R7465 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.Qb.n0 5.7305
R7466 SARlogic_0.dffrs_0.Qb.n5 SARlogic_0.dffrs_0.Qb.n4 5.14711
R7467 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_0.Qb.n2 5.13907
R7468 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n6 4.94976
R7469 SARlogic_0.dffrs_0.nand3_7.Z SARlogic_0.dffrs_0.Qb.n9 4.72925
R7470 SARlogic_0.dffrs_7.setb SARlogic_0.dffrs_7.nand3_0.C 0.784786
R7471 SARlogic_0.dffrs_0.Qb.n9 SARlogic_0.dffrs_0.Qb.n8 0.732092
R7472 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t1 0.7285
R7473 SARlogic_0.dffrs_0.Qb.n7 SARlogic_0.dffrs_0.Qb.t0 0.7285
R7474 SARlogic_0.dffrs_0.Qb.n6 SARlogic_0.dffrs_0.Qb 0.175225
R7475 SARlogic_0.dffrs_0.Qb.n1 SARlogic_0.dffrs_0.nand3_2.A 0.0455
R7476 SARlogic_0.dffrs_0.Qb.n3 SARlogic_0.dffrs_7.nand3_2.C 0.0455
R7477 SARlogic_0.dffrs_7.nand3_0.C SARlogic_0.dffrs_0.Qb.n5 0.0374643
R7478 a_9083_31160.n0 a_9083_31160.t5 34.1797
R7479 a_9083_31160.n0 a_9083_31160.t4 19.5798
R7480 a_9083_31160.n1 a_9083_31160.t2 18.7717
R7481 a_9083_31160.n1 a_9083_31160.t3 9.2885
R7482 a_9083_31160.n2 a_9083_31160.n0 4.93379
R7483 a_9083_31160.t0 a_9083_31160.n3 4.23346
R7484 a_9083_31160.n3 a_9083_31160.t1 3.85546
R7485 a_9083_31160.n2 a_9083_31160.n1 0.4055
R7486 a_9083_31160.n3 a_9083_31160.n2 0.352625
R7487 a_23785_29218.n2 a_23785_29218.t5 40.8177
R7488 a_23785_29218.n3 a_23785_29218.t4 40.6313
R7489 a_23785_29218.n3 a_23785_29218.t7 27.3166
R7490 a_23785_29218.n2 a_23785_29218.t6 27.1302
R7491 a_23785_29218.n4 a_23785_29218.n3 19.2576
R7492 a_23785_29218.t0 a_23785_29218.n5 10.0473
R7493 a_23785_29218.n1 a_23785_29218.t1 6.51042
R7494 a_23785_29218.n1 a_23785_29218.n0 6.04952
R7495 a_23785_29218.n4 a_23785_29218.n2 5.91752
R7496 a_23785_29218.n5 a_23785_29218.n4 4.89565
R7497 a_23785_29218.n5 a_23785_29218.n1 0.732092
R7498 a_23785_29218.n0 a_23785_29218.t3 0.7285
R7499 a_23785_29218.n0 a_23785_29218.t2 0.7285
R7500 a_23865_30170.n0 a_23865_30170.t7 41.0041
R7501 a_23865_30170.n1 a_23865_30170.t5 40.8177
R7502 a_23865_30170.n1 a_23865_30170.t6 27.1302
R7503 a_23865_30170.n0 a_23865_30170.t4 26.9438
R7504 a_23865_30170.n2 a_23865_30170.n1 22.5284
R7505 a_23865_30170.n3 a_23865_30170.n2 19.5781
R7506 a_23865_30170.n3 a_23865_30170.t1 10.0473
R7507 a_23865_30170.n4 a_23865_30170.t3 6.51042
R7508 a_23865_30170.n5 a_23865_30170.n4 6.04952
R7509 a_23865_30170.n2 a_23865_30170.n0 5.7305
R7510 a_23865_30170.n4 a_23865_30170.n3 0.732092
R7511 a_23865_30170.n5 a_23865_30170.t2 0.7285
R7512 a_23865_30170.t0 a_23865_30170.n5 0.7285
R7513 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t4 40.6313
R7514 SARlogic_0.dffrs_3.nand3_1.C.n0 SARlogic_0.dffrs_3.nand3_1.C.t5 27.3166
R7515 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n1 14.2854
R7516 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.t1 10.0473
R7517 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.t2 6.51042
R7518 SARlogic_0.dffrs_3.nand3_1.C.n3 SARlogic_0.dffrs_3.nand3_1.C.n2 6.04952
R7519 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C.n0 5.13907
R7520 SARlogic_0.dffrs_3.nand3_0.Z SARlogic_0.dffrs_3.nand3_1.C.n4 4.72925
R7521 SARlogic_0.dffrs_3.nand3_1.C.n4 SARlogic_0.dffrs_3.nand3_1.C.n3 0.732092
R7522 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t0 0.7285
R7523 SARlogic_0.dffrs_3.nand3_1.C.n2 SARlogic_0.dffrs_3.nand3_1.C.t3 0.7285
R7524 SARlogic_0.dffrs_3.nand3_1.C.n1 SARlogic_0.dffrs_3.nand3_1.C 0.0455
R7525 a_42729_33628.n0 a_42729_33628.t4 40.6313
R7526 a_42729_33628.n0 a_42729_33628.t5 27.3166
R7527 a_42729_33628.n1 a_42729_33628.n0 24.1527
R7528 a_42729_33628.n1 a_42729_33628.t3 10.0473
R7529 a_42729_33628.n2 a_42729_33628.t2 6.51042
R7530 a_42729_33628.n3 a_42729_33628.n2 6.04952
R7531 a_42729_33628.n2 a_42729_33628.n1 0.732092
R7532 a_42729_33628.t0 a_42729_33628.n3 0.7285
R7533 a_42729_33628.n3 a_42729_33628.t1 0.7285
R7534 a_42729_31423.n3 a_42729_31423.t4 41.0041
R7535 a_42729_31423.n2 a_42729_31423.t5 40.8177
R7536 a_42729_31423.n4 a_42729_31423.t6 40.6313
R7537 a_42729_31423.n4 a_42729_31423.t9 27.3166
R7538 a_42729_31423.n2 a_42729_31423.t8 27.1302
R7539 a_42729_31423.n3 a_42729_31423.t7 26.9438
R7540 a_42729_31423.n5 a_42729_31423.n3 15.6312
R7541 a_42729_31423.n5 a_42729_31423.n4 15.046
R7542 a_42729_31423.t0 a_42729_31423.n7 10.0473
R7543 a_42729_31423.n1 a_42729_31423.t2 6.51042
R7544 a_42729_31423.n1 a_42729_31423.n0 6.04952
R7545 a_42729_31423.n6 a_42729_31423.n2 5.64619
R7546 a_42729_31423.n7 a_42729_31423.n6 5.17851
R7547 a_42729_31423.n6 a_42729_31423.n5 4.5005
R7548 a_42729_31423.n7 a_42729_31423.n1 0.732092
R7549 a_42729_31423.n0 a_42729_31423.t3 0.7285
R7550 a_42729_31423.n0 a_42729_31423.t1 0.7285
R7551 a_28027_31160.n0 a_28027_31160.t4 34.1797
R7552 a_28027_31160.n0 a_28027_31160.t5 19.5798
R7553 a_28027_31160.n1 a_28027_31160.t1 18.7717
R7554 a_28027_31160.n1 a_28027_31160.t2 9.2885
R7555 a_28027_31160.n2 a_28027_31160.n0 4.93379
R7556 a_28027_31160.t0 a_28027_31160.n3 4.23346
R7557 a_28027_31160.n3 a_28027_31160.t3 3.85546
R7558 a_28027_31160.n2 a_28027_31160.n1 0.4055
R7559 a_28027_31160.n3 a_28027_31160.n2 0.352625
R7560 a_23785_31423.n1 a_23785_31423.t5 41.0041
R7561 a_23785_31423.n0 a_23785_31423.t7 40.8177
R7562 a_23785_31423.n2 a_23785_31423.t4 40.6313
R7563 a_23785_31423.n2 a_23785_31423.t6 27.3166
R7564 a_23785_31423.n0 a_23785_31423.t9 27.1302
R7565 a_23785_31423.n1 a_23785_31423.t8 26.9438
R7566 a_23785_31423.n3 a_23785_31423.n1 15.6312
R7567 a_23785_31423.n3 a_23785_31423.n2 15.046
R7568 a_23785_31423.n5 a_23785_31423.t1 10.0473
R7569 a_23785_31423.n6 a_23785_31423.t3 6.51042
R7570 a_23785_31423.n7 a_23785_31423.n6 6.04952
R7571 a_23785_31423.n4 a_23785_31423.n0 5.64619
R7572 a_23785_31423.n5 a_23785_31423.n4 5.17851
R7573 a_23785_31423.n4 a_23785_31423.n3 4.5005
R7574 a_23785_31423.n6 a_23785_31423.n5 0.732092
R7575 a_23785_31423.n7 a_23785_31423.t2 0.7285
R7576 a_23785_31423.t0 a_23785_31423.n7 0.7285
R7577 Vin1.n7 Vin1.n6 23.1032
R7578 Vin1.n3 Vin1.n2 23.1032
R7579 Vin1.n0 Vin1.t8 22.5295
R7580 Vin1.n2 Vin1.t2 16.3641
R7581 Vin1.n6 Vin1.t6 16.3626
R7582 Vin1.n2 Vin1.t7 16.0225
R7583 Vin1.n6 Vin1.t1 16.021
R7584 Vin1.n8 Vin1.t4 11.5195
R7585 Vin1.n5 Vin1.t3 11.5195
R7586 Vin1.n4 Vin1.t9 11.5195
R7587 Vin1.n1 Vin1.t5 11.5195
R7588 Vin1.n0 Vin1.t0 11.5195
R7589 comparator_no_offsetcal_0.Vin1 Vin1 5.6843
R7590 Vin1.n1 Vin1.n0 4.00673
R7591 comparator_no_offsetcal_0.Vin1 Vin1.n8 3.9441
R7592 Vin1.n7 Vin1.n5 3.16619
R7593 Vin1.n3 Vin1.n1 0.650658
R7594 Vin1.n8 Vin1.n7 0.280193
R7595 Vin1.n4 Vin1.n3 0.279681
R7596 Vin1.n5 Vin1.n4 0.231705
R7597 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 19.5626
R7598 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 11.9065
R7599 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 11.2495
R7600 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 11.243
R7601 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 8.80104
R7602 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 6.60725
R7603 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 6.52262
R7604 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 6.386
R7605 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 5.44213
R7606 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 4.36738
R7607 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 4.36738
R7608 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 4.3505
R7609 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n15 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 2.2505
R7610 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n12 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 2.14009
R7611 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n7 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 1.50001
R7612 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n13 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n4 1.49326
R7613 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t12 1.0925
R7614 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n14 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t5 1.0925
R7615 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t10 1.0925
R7616 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n11 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t15 1.0925
R7617 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t6 1.0925
R7618 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n5 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t8 1.0925
R7619 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t14 1.0925
R7620 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n8 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t9 1.0925
R7621 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t16 1.0925
R7622 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n6 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t11 1.0925
R7623 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t7 1.0925
R7624 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n3 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t13 1.0925
R7625 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t2 0.8195
R7626 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n1 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t4 0.8195
R7627 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t3 0.8195
R7628 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n0 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.t1 0.8195
R7629 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n10 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n9 0.314375
R7630 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n16 comparator_no_offsetcal_0.no_offsetLatch_0.Vp.n2 0.16025
R7631 a_n4631_31422.n3 a_n4631_31422.t9 41.0041
R7632 a_n4631_31422.n2 a_n4631_31422.t6 40.8177
R7633 a_n4631_31422.n4 a_n4631_31422.t5 40.6313
R7634 a_n4631_31422.n4 a_n4631_31422.t7 27.3166
R7635 a_n4631_31422.n2 a_n4631_31422.t8 27.1302
R7636 a_n4631_31422.n3 a_n4631_31422.t4 26.9438
R7637 a_n4631_31422.n5 a_n4631_31422.n3 15.6312
R7638 a_n4631_31422.n5 a_n4631_31422.n4 15.046
R7639 a_n4631_31422.t0 a_n4631_31422.n7 10.0473
R7640 a_n4631_31422.n1 a_n4631_31422.t1 6.51042
R7641 a_n4631_31422.n1 a_n4631_31422.n0 6.04952
R7642 a_n4631_31422.n6 a_n4631_31422.n2 5.64619
R7643 a_n4631_31422.n7 a_n4631_31422.n6 5.17851
R7644 a_n4631_31422.n6 a_n4631_31422.n5 4.5005
R7645 a_n4631_31422.n7 a_n4631_31422.n1 0.732092
R7646 a_n4631_31422.n0 a_n4631_31422.t3 0.7285
R7647 a_n4631_31422.n0 a_n4631_31422.t2 0.7285
R7648 a_n4631_33627.n2 a_n4631_33627.t4 40.6313
R7649 a_n4631_33627.n2 a_n4631_33627.t5 27.3166
R7650 a_n4631_33627.n3 a_n4631_33627.n2 24.1527
R7651 a_n4631_33627.t0 a_n4631_33627.n3 10.0473
R7652 a_n4631_33627.n1 a_n4631_33627.t1 6.51042
R7653 a_n4631_33627.n1 a_n4631_33627.n0 6.04952
R7654 a_n4631_33627.n3 a_n4631_33627.n1 0.732092
R7655 a_n4631_33627.n0 a_n4631_33627.t3 0.7285
R7656 a_n4631_33627.n0 a_n4631_33627.t2 0.7285
R7657 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t6 40.8177
R7658 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t7 40.6313
R7659 SARlogic_0.dffrs_11.nand3_8.C.n1 SARlogic_0.dffrs_11.nand3_8.C.t4 27.3166
R7660 SARlogic_0.dffrs_11.nand3_8.C.n0 SARlogic_0.dffrs_11.nand3_8.C.t5 27.1302
R7661 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_8.C.n2 14.119
R7662 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.t0 10.0473
R7663 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.t1 6.51042
R7664 SARlogic_0.dffrs_11.nand3_8.C.n5 SARlogic_0.dffrs_11.nand3_8.C.n4 6.04952
R7665 SARlogic_0.dffrs_11.nand3_7.B SARlogic_0.dffrs_11.nand3_8.C.n0 5.47979
R7666 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C.n1 5.13907
R7667 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n6 4.72925
R7668 SARlogic_0.dffrs_11.nand3_8.C.n6 SARlogic_0.dffrs_11.nand3_8.C.n5 0.732092
R7669 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t2 0.7285
R7670 SARlogic_0.dffrs_11.nand3_8.C.n4 SARlogic_0.dffrs_11.nand3_8.C.t3 0.7285
R7671 SARlogic_0.dffrs_11.nand3_8.C.n3 SARlogic_0.dffrs_11.nand3_7.B 0.438233
R7672 SARlogic_0.dffrs_11.nand3_6.Z SARlogic_0.dffrs_11.nand3_8.C.n3 0.166901
R7673 SARlogic_0.dffrs_11.nand3_8.C.n2 SARlogic_0.dffrs_11.nand3_8.C 0.0455
R7674 SAR_in.n9 SAR_in.t11 41.0041
R7675 SAR_in.n7 SAR_in.t6 41.0041
R7676 SAR_in.n5 SAR_in.t2 41.0041
R7677 SAR_in.n3 SAR_in.t8 41.0041
R7678 SAR_in.n1 SAR_in.t1 41.0041
R7679 SAR_in.n0 SAR_in.t7 41.0041
R7680 SAR_in.n9 SAR_in.t3 26.9438
R7681 SAR_in.n7 SAR_in.t9 26.9438
R7682 SAR_in.n5 SAR_in.t5 26.9438
R7683 SAR_in.n3 SAR_in.t0 26.9438
R7684 SAR_in.n1 SAR_in.t4 26.9438
R7685 SAR_in.n0 SAR_in.t10 26.9438
R7686 SAR_in.n2 SARlogic_0.dffrs_11.d 15.3544
R7687 SAR_in.n8 SARlogic_0.dffrs_7.d 11.7166
R7688 SAR_in.n6 SARlogic_0.dffrs_8.d 11.7166
R7689 SAR_in.n4 SARlogic_0.dffrs_9.d 11.7166
R7690 SAR_in.n2 SARlogic_0.dffrs_10.d 11.7166
R7691 SAR_in.n10 SARlogic_0.dffrs_14.d 11.6732
R7692 SARlogic_0.comp_in SAR_in.n10 7.63655
R7693 SARlogic_0.dffrs_14.nand3_8.A SAR_in.n9 5.7755
R7694 SARlogic_0.dffrs_7.nand3_8.A SAR_in.n7 5.7755
R7695 SARlogic_0.dffrs_8.nand3_8.A SAR_in.n5 5.7755
R7696 SARlogic_0.dffrs_9.nand3_8.A SAR_in.n3 5.7755
R7697 SARlogic_0.dffrs_10.nand3_8.A SAR_in.n1 5.7755
R7698 SARlogic_0.dffrs_11.nand3_8.A SAR_in.n0 5.7755
R7699 SAR_in.n4 SAR_in.n2 3.6383
R7700 SAR_in.n6 SAR_in.n4 3.6383
R7701 SAR_in.n8 SAR_in.n6 3.6383
R7702 SAR_in.n10 SAR_in.n8 3.6113
R7703 SARlogic_0.dffrs_14.d SARlogic_0.dffrs_14.nand3_8.A 0.784786
R7704 SARlogic_0.dffrs_7.d SARlogic_0.dffrs_7.nand3_8.A 0.784786
R7705 SARlogic_0.dffrs_8.d SARlogic_0.dffrs_8.nand3_8.A 0.784786
R7706 SARlogic_0.dffrs_9.d SARlogic_0.dffrs_9.nand3_8.A 0.784786
R7707 SARlogic_0.dffrs_10.d SARlogic_0.dffrs_10.nand3_8.A 0.784786
R7708 SARlogic_0.dffrs_11.d SARlogic_0.dffrs_11.nand3_8.A 0.784786
R7709 SARlogic_0.comp_in SAR_in 0.1775
R7710 a_n9861_31159.n0 a_n9861_31159.t4 34.1797
R7711 a_n9861_31159.n0 a_n9861_31159.t5 19.5798
R7712 a_n9861_31159.n1 a_n9861_31159.t2 18.7717
R7713 a_n9861_31159.n1 a_n9861_31159.t3 9.2885
R7714 a_n9861_31159.n2 a_n9861_31159.n0 4.93379
R7715 a_n9861_31159.t0 a_n9861_31159.n3 4.23346
R7716 a_n9861_31159.n3 a_n9861_31159.t1 3.85546
R7717 a_n9861_31159.n2 a_n9861_31159.n1 0.4055
R7718 a_n9861_31159.n3 a_n9861_31159.n2 0.352625
R7719 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t6 40.8177
R7720 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t7 40.6313
R7721 SARlogic_0.dffrs_14.nand3_8.C.n1 SARlogic_0.dffrs_14.nand3_8.C.t5 27.3166
R7722 SARlogic_0.dffrs_14.nand3_8.C.n0 SARlogic_0.dffrs_14.nand3_8.C.t4 27.1302
R7723 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_8.C.n2 14.119
R7724 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.t1 10.0473
R7725 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.t2 6.51042
R7726 SARlogic_0.dffrs_14.nand3_8.C.n5 SARlogic_0.dffrs_14.nand3_8.C.n4 6.04952
R7727 SARlogic_0.dffrs_14.nand3_7.B SARlogic_0.dffrs_14.nand3_8.C.n0 5.47979
R7728 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C.n1 5.13907
R7729 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n6 4.72925
R7730 SARlogic_0.dffrs_14.nand3_8.C.n6 SARlogic_0.dffrs_14.nand3_8.C.n5 0.732092
R7731 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t3 0.7285
R7732 SARlogic_0.dffrs_14.nand3_8.C.n4 SARlogic_0.dffrs_14.nand3_8.C.t0 0.7285
R7733 SARlogic_0.dffrs_14.nand3_8.C.n3 SARlogic_0.dffrs_14.nand3_7.B 0.438233
R7734 SARlogic_0.dffrs_14.nand3_6.Z SARlogic_0.dffrs_14.nand3_8.C.n3 0.166901
R7735 SARlogic_0.dffrs_14.nand3_8.C.n2 SARlogic_0.dffrs_14.nand3_8.C 0.0455
R7736 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t6 41.0041
R7737 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t7 40.8177
R7738 SARlogic_0.dffrs_13.nand3_8.Z.n1 SARlogic_0.dffrs_13.nand3_8.Z.t4 27.1302
R7739 SARlogic_0.dffrs_13.nand3_8.Z.n0 SARlogic_0.dffrs_13.nand3_8.Z.t5 26.9438
R7740 SARlogic_0.dffrs_13.nand3_6.A SARlogic_0.dffrs_13.nand3_0.B 17.0041
R7741 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n2 14.8493
R7742 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.t1 10.0473
R7743 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.t0 6.51042
R7744 SARlogic_0.dffrs_13.nand3_8.Z.n4 SARlogic_0.dffrs_13.nand3_8.Z.n3 6.04952
R7745 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_8.Z.n0 5.7305
R7746 SARlogic_0.dffrs_13.nand3_0.B SARlogic_0.dffrs_13.nand3_8.Z.n1 5.47979
R7747 SARlogic_0.dffrs_13.nand3_8.Z SARlogic_0.dffrs_13.nand3_8.Z.n5 4.72925
R7748 SARlogic_0.dffrs_13.nand3_8.Z.n5 SARlogic_0.dffrs_13.nand3_8.Z.n4 0.732092
R7749 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t2 0.7285
R7750 SARlogic_0.dffrs_13.nand3_8.Z.n3 SARlogic_0.dffrs_13.nand3_8.Z.t3 0.7285
R7751 SARlogic_0.dffrs_13.nand3_8.Z.n2 SARlogic_0.dffrs_13.nand3_6.A 0.0455
R7752 a_n389_31159.n0 a_n389_31159.t4 34.1797
R7753 a_n389_31159.n0 a_n389_31159.t5 19.5798
R7754 a_n389_31159.n1 a_n389_31159.t2 18.7717
R7755 a_n389_31159.n1 a_n389_31159.t1 9.2885
R7756 a_n389_31159.n2 a_n389_31159.n0 4.93379
R7757 a_n389_31159.t0 a_n389_31159.n3 4.23346
R7758 a_n389_31159.n3 a_n389_31159.t3 3.85546
R7759 a_n389_31159.n2 a_n389_31159.n1 0.4055
R7760 a_n389_31159.n3 a_n389_31159.n2 0.352625
R7761 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t5 40.8177
R7762 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t7 40.6313
R7763 SARlogic_0.dffrs_9.nand3_8.C.n1 SARlogic_0.dffrs_9.nand3_8.C.t4 27.3166
R7764 SARlogic_0.dffrs_9.nand3_8.C.n0 SARlogic_0.dffrs_9.nand3_8.C.t6 27.1302
R7765 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_8.C.n2 14.119
R7766 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.t1 10.0473
R7767 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.t2 6.51042
R7768 SARlogic_0.dffrs_9.nand3_8.C.n5 SARlogic_0.dffrs_9.nand3_8.C.n4 6.04952
R7769 SARlogic_0.dffrs_9.nand3_7.B SARlogic_0.dffrs_9.nand3_8.C.n0 5.47979
R7770 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C.n1 5.13907
R7771 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n6 4.72925
R7772 SARlogic_0.dffrs_9.nand3_8.C.n6 SARlogic_0.dffrs_9.nand3_8.C.n5 0.732092
R7773 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t0 0.7285
R7774 SARlogic_0.dffrs_9.nand3_8.C.n4 SARlogic_0.dffrs_9.nand3_8.C.t3 0.7285
R7775 SARlogic_0.dffrs_9.nand3_8.C.n3 SARlogic_0.dffrs_9.nand3_7.B 0.438233
R7776 SARlogic_0.dffrs_9.nand3_6.Z SARlogic_0.dffrs_9.nand3_8.C.n3 0.166901
R7777 SARlogic_0.dffrs_9.nand3_8.C.n2 SARlogic_0.dffrs_9.nand3_8.C 0.0455
R7778 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t6 41.0041
R7779 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t7 40.8177
R7780 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t4 40.6313
R7781 SARlogic_0.dffrs_0.nand3_6.C.n3 SARlogic_0.dffrs_0.nand3_6.C.t5 27.3166
R7782 SARlogic_0.dffrs_0.nand3_6.C.n0 SARlogic_0.dffrs_0.nand3_6.C.t8 27.1302
R7783 SARlogic_0.dffrs_0.nand3_6.C.n1 SARlogic_0.dffrs_0.nand3_6.C.t9 26.9438
R7784 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.t1 10.0473
R7785 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n4 9.90747
R7786 SARlogic_0.dffrs_0.nand3_6.C.n5 SARlogic_0.dffrs_0.nand3_6.C.n2 9.90116
R7787 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.t2 6.51042
R7788 SARlogic_0.dffrs_0.nand3_6.C.n8 SARlogic_0.dffrs_0.nand3_6.C.n7 6.04952
R7789 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_6.C.n1 5.7305
R7790 SARlogic_0.dffrs_0.nand3_2.B SARlogic_0.dffrs_0.nand3_6.C.n0 5.47979
R7791 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C.n3 5.13907
R7792 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n9 4.72925
R7793 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_6.C.n5 4.5005
R7794 SARlogic_0.dffrs_0.nand3_6.C.n9 SARlogic_0.dffrs_0.nand3_6.C.n8 0.732092
R7795 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t0 0.7285
R7796 SARlogic_0.dffrs_0.nand3_6.C.n7 SARlogic_0.dffrs_0.nand3_6.C.t3 0.7285
R7797 SARlogic_0.dffrs_0.nand3_1.Z SARlogic_0.dffrs_0.nand3_6.C.n6 0.449758
R7798 SARlogic_0.dffrs_0.nand3_6.C.n6 SARlogic_0.dffrs_0.nand3_2.B 0.166901
R7799 SARlogic_0.dffrs_0.nand3_6.C.n2 SARlogic_0.dffrs_0.nand3_0.A 0.0455
R7800 SARlogic_0.dffrs_0.nand3_6.C.n4 SARlogic_0.dffrs_0.nand3_6.C 0.0455
R7801 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t6 40.8177
R7802 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t5 40.6313
R7803 SARlogic_0.dffrs_0.nand3_8.C.n1 SARlogic_0.dffrs_0.nand3_8.C.t7 27.3166
R7804 SARlogic_0.dffrs_0.nand3_8.C.n0 SARlogic_0.dffrs_0.nand3_8.C.t4 27.1302
R7805 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_8.C.n2 14.119
R7806 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.t2 10.0473
R7807 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.t1 6.51042
R7808 SARlogic_0.dffrs_0.nand3_8.C.n5 SARlogic_0.dffrs_0.nand3_8.C.n4 6.04952
R7809 SARlogic_0.dffrs_0.nand3_7.B SARlogic_0.dffrs_0.nand3_8.C.n0 5.47979
R7810 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C.n1 5.13907
R7811 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n6 4.72925
R7812 SARlogic_0.dffrs_0.nand3_8.C.n6 SARlogic_0.dffrs_0.nand3_8.C.n5 0.732092
R7813 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t0 0.7285
R7814 SARlogic_0.dffrs_0.nand3_8.C.n4 SARlogic_0.dffrs_0.nand3_8.C.t3 0.7285
R7815 SARlogic_0.dffrs_0.nand3_8.C.n3 SARlogic_0.dffrs_0.nand3_7.B 0.438233
R7816 SARlogic_0.dffrs_0.nand3_6.Z SARlogic_0.dffrs_0.nand3_8.C.n3 0.166901
R7817 SARlogic_0.dffrs_0.nand3_8.C.n2 SARlogic_0.dffrs_0.nand3_8.C 0.0455
R7818 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t7 41.0041
R7819 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t6 40.8177
R7820 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t5 40.6313
R7821 SARlogic_0.dffrs_11.nand3_6.C.n3 SARlogic_0.dffrs_11.nand3_6.C.t4 27.3166
R7822 SARlogic_0.dffrs_11.nand3_6.C.n0 SARlogic_0.dffrs_11.nand3_6.C.t8 27.1302
R7823 SARlogic_0.dffrs_11.nand3_6.C.n1 SARlogic_0.dffrs_11.nand3_6.C.t9 26.9438
R7824 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.t2 10.0473
R7825 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n4 9.90747
R7826 SARlogic_0.dffrs_11.nand3_6.C.n5 SARlogic_0.dffrs_11.nand3_6.C.n2 9.90116
R7827 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.t3 6.51042
R7828 SARlogic_0.dffrs_11.nand3_6.C.n8 SARlogic_0.dffrs_11.nand3_6.C.n7 6.04952
R7829 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_6.C.n1 5.7305
R7830 SARlogic_0.dffrs_11.nand3_2.B SARlogic_0.dffrs_11.nand3_6.C.n0 5.47979
R7831 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C.n3 5.13907
R7832 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n9 4.72925
R7833 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_6.C.n5 4.5005
R7834 SARlogic_0.dffrs_11.nand3_6.C.n9 SARlogic_0.dffrs_11.nand3_6.C.n8 0.732092
R7835 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t0 0.7285
R7836 SARlogic_0.dffrs_11.nand3_6.C.n7 SARlogic_0.dffrs_11.nand3_6.C.t1 0.7285
R7837 SARlogic_0.dffrs_11.nand3_1.Z SARlogic_0.dffrs_11.nand3_6.C.n6 0.449758
R7838 SARlogic_0.dffrs_11.nand3_6.C.n6 SARlogic_0.dffrs_11.nand3_2.B 0.166901
R7839 SARlogic_0.dffrs_11.nand3_6.C.n2 SARlogic_0.dffrs_11.nand3_0.A 0.0455
R7840 SARlogic_0.dffrs_11.nand3_6.C.n4 SARlogic_0.dffrs_11.nand3_6.C 0.0455
R7841 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t4 41.0041
R7842 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t5 40.8177
R7843 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t9 40.6313
R7844 SARlogic_0.dffrs_8.nand3_6.C.n3 SARlogic_0.dffrs_8.nand3_6.C.t8 27.3166
R7845 SARlogic_0.dffrs_8.nand3_6.C.n0 SARlogic_0.dffrs_8.nand3_6.C.t7 27.1302
R7846 SARlogic_0.dffrs_8.nand3_6.C.n1 SARlogic_0.dffrs_8.nand3_6.C.t6 26.9438
R7847 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.t1 10.0473
R7848 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n4 9.90747
R7849 SARlogic_0.dffrs_8.nand3_6.C.n5 SARlogic_0.dffrs_8.nand3_6.C.n2 9.90116
R7850 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.t2 6.51042
R7851 SARlogic_0.dffrs_8.nand3_6.C.n8 SARlogic_0.dffrs_8.nand3_6.C.n7 6.04952
R7852 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_6.C.n1 5.7305
R7853 SARlogic_0.dffrs_8.nand3_2.B SARlogic_0.dffrs_8.nand3_6.C.n0 5.47979
R7854 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C.n3 5.13907
R7855 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n9 4.72925
R7856 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_6.C.n5 4.5005
R7857 SARlogic_0.dffrs_8.nand3_6.C.n9 SARlogic_0.dffrs_8.nand3_6.C.n8 0.732092
R7858 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t0 0.7285
R7859 SARlogic_0.dffrs_8.nand3_6.C.n7 SARlogic_0.dffrs_8.nand3_6.C.t3 0.7285
R7860 SARlogic_0.dffrs_8.nand3_1.Z SARlogic_0.dffrs_8.nand3_6.C.n6 0.449758
R7861 SARlogic_0.dffrs_8.nand3_6.C.n6 SARlogic_0.dffrs_8.nand3_2.B 0.166901
R7862 SARlogic_0.dffrs_8.nand3_6.C.n2 SARlogic_0.dffrs_8.nand3_0.A 0.0455
R7863 SARlogic_0.dffrs_8.nand3_6.C.n4 SARlogic_0.dffrs_8.nand3_6.C 0.0455
R7864 a_n389_28819.n0 a_n389_28819.t5 34.1797
R7865 a_n389_28819.n0 a_n389_28819.t4 19.5798
R7866 a_n389_28819.n1 a_n389_28819.t1 18.7717
R7867 a_n389_28819.n1 a_n389_28819.t2 9.2885
R7868 a_n389_28819.n2 a_n389_28819.n0 4.93379
R7869 a_n389_28819.t0 a_n389_28819.n3 4.23346
R7870 a_n389_28819.n3 a_n389_28819.t3 3.85546
R7871 a_n389_28819.n2 a_n389_28819.n1 0.4055
R7872 a_n389_28819.n3 a_n389_28819.n2 0.352625
R7873 a_1839_29263.n0 a_1839_29263.t5 34.1797
R7874 a_1839_29263.n0 a_1839_29263.t4 19.5798
R7875 a_1839_29263.n3 a_1839_29263.t3 10.3401
R7876 a_1839_29263.t0 a_1839_29263.n3 9.2885
R7877 a_1839_29263.n2 a_1839_29263.n0 4.93379
R7878 a_1839_29263.n1 a_1839_29263.t1 4.09202
R7879 a_1839_29263.n1 a_1839_29263.t2 3.95079
R7880 a_1839_29263.n3 a_1839_29263.n2 0.599711
R7881 a_1839_29263.n2 a_1839_29263.n1 0.296375
R7882 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t4 40.6313
R7883 SARlogic_0.dffrs_0.nand3_1.C.n0 SARlogic_0.dffrs_0.nand3_1.C.t5 27.3166
R7884 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n1 14.2854
R7885 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.t2 10.0473
R7886 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.t3 6.51042
R7887 SARlogic_0.dffrs_0.nand3_1.C.n3 SARlogic_0.dffrs_0.nand3_1.C.n2 6.04952
R7888 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C.n0 5.13907
R7889 SARlogic_0.dffrs_0.nand3_0.Z SARlogic_0.dffrs_0.nand3_1.C.n4 4.72925
R7890 SARlogic_0.dffrs_0.nand3_1.C.n4 SARlogic_0.dffrs_0.nand3_1.C.n3 0.732092
R7891 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t0 0.7285
R7892 SARlogic_0.dffrs_0.nand3_1.C.n2 SARlogic_0.dffrs_0.nand3_1.C.t1 0.7285
R7893 SARlogic_0.dffrs_0.nand3_1.C.n1 SARlogic_0.dffrs_0.nand3_1.C 0.0455
R7894 a_20783_29264.n0 a_20783_29264.t5 34.1797
R7895 a_20783_29264.n0 a_20783_29264.t4 19.5798
R7896 a_20783_29264.t0 a_20783_29264.n3 10.3401
R7897 a_20783_29264.n3 a_20783_29264.t3 9.2885
R7898 a_20783_29264.n2 a_20783_29264.n0 4.93379
R7899 a_20783_29264.n1 a_20783_29264.t2 4.09202
R7900 a_20783_29264.n1 a_20783_29264.t1 3.95079
R7901 a_20783_29264.n3 a_20783_29264.n2 0.599711
R7902 a_20783_29264.n2 a_20783_29264.n1 0.296375
R7903 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t8 40.6313
R7904 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.t6 34.1066
R7905 adc_PISO_0.2inmux_2.Bit.n3 adc_PISO_0.2inmux_2.Bit.t4 27.3166
R7906 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t7 19.673
R7907 adc_PISO_0.2inmux_2.Bit.n0 adc_PISO_0.2inmux_2.Bit.t5 19.4007
R7908 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n3 14.6967
R7909 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.t2 10.0473
R7910 adc_PISO_0.2inmux_2.Bit.n7 adc_PISO_0.2inmux_2.Bit.n6 9.39565
R7911 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit.n1 6.70486
R7912 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.t3 6.51042
R7913 adc_PISO_0.2inmux_2.Bit.n5 adc_PISO_0.2inmux_2.Bit.n4 6.04952
R7914 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n2 5.81514
R7915 adc_PISO_0.2inmux_2.Bit.n6 adc_PISO_0.2inmux_2.Bit.n5 0.732092
R7916 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t0 0.7285
R7917 adc_PISO_0.2inmux_2.Bit.n4 adc_PISO_0.2inmux_2.Bit.t1 0.7285
R7918 adc_PISO_0.dffrs_0.Q adc_PISO_0.2inmux_2.Bit.n7 0.458082
R7919 adc_PISO_0.2inmux_2.Bit.n1 adc_PISO_0.2inmux_2.Bit.n0 0.252687
R7920 adc_PISO_0.2inmux_2.Bit.n2 adc_PISO_0.2inmux_2.Bit 0.0519286
R7921 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_11.clk 44.4671
R7922 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t7 41.0041
R7923 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t6 40.8177
R7924 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t8 40.6313
R7925 SARlogic_0.dffrs_12.Q.n3 SARlogic_0.dffrs_12.Q.t5 27.3166
R7926 SARlogic_0.dffrs_12.Q.n1 SARlogic_0.dffrs_12.Q.t4 27.1302
R7927 SARlogic_0.dffrs_12.Q.n0 SARlogic_0.dffrs_12.Q.t9 26.9438
R7928 SARlogic_0.dffrs_12.Q.n5 SARlogic_0.dffrs_12.Q.n4 14.0582
R7929 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.t2 10.0473
R7930 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.t3 6.51042
R7931 SARlogic_0.dffrs_12.Q.n7 SARlogic_0.dffrs_12.Q.n6 6.04952
R7932 SARlogic_0.dffrs_11.nand3_1.A SARlogic_0.dffrs_12.Q.n0 5.7755
R7933 SARlogic_0.dffrs_11.nand3_6.B SARlogic_0.dffrs_12.Q.n1 5.47979
R7934 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.Q.n3 5.13907
R7935 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n8 4.72925
R7936 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_6.B 2.17818
R7937 SARlogic_0.dffrs_12.Q.n2 SARlogic_0.dffrs_11.nand3_1.A 1.34729
R7938 SARlogic_0.dffrs_12.Q.n8 SARlogic_0.dffrs_12.Q.n7 0.732092
R7939 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t0 0.7285
R7940 SARlogic_0.dffrs_12.Q.n6 SARlogic_0.dffrs_12.Q.t1 0.7285
R7941 SARlogic_0.dffrs_11.clk SARlogic_0.dffrs_12.Q.n2 0.610571
R7942 SARlogic_0.dffrs_12.nand3_2.Z SARlogic_0.dffrs_12.Q.n5 0.166901
R7943 SARlogic_0.dffrs_12.Q.n4 SARlogic_0.dffrs_12.nand3_7.C 0.0455
R7944 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t3 41.0041
R7945 adc_PISO_0.2inmux_2.OUT.n0 adc_PISO_0.2inmux_2.OUT.t2 26.9438
R7946 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t0 9.6935
R7947 adc_PISO_0.dffrs_1.d adc_PISO_0.2inmux_2.OUT.n0 6.55979
R7948 adc_PISO_0.2inmux_2.OUT adc_PISO_0.dffrs_1.d 4.883
R7949 adc_PISO_0.2inmux_2.OUT.n1 adc_PISO_0.2inmux_2.OUT.t1 4.35383
R7950 adc_PISO_0.2inmux_2.OUT adc_PISO_0.2inmux_2.OUT.n1 0.350857
R7951 a_4921_30169.n2 a_4921_30169.t5 41.0041
R7952 a_4921_30169.n3 a_4921_30169.t6 40.8177
R7953 a_4921_30169.n3 a_4921_30169.t4 27.1302
R7954 a_4921_30169.n2 a_4921_30169.t7 26.9438
R7955 a_4921_30169.n4 a_4921_30169.n3 22.5284
R7956 a_4921_30169.n5 a_4921_30169.n4 19.5781
R7957 a_4921_30169.t0 a_4921_30169.n5 10.0473
R7958 a_4921_30169.n1 a_4921_30169.t1 6.51042
R7959 a_4921_30169.n1 a_4921_30169.n0 6.04952
R7960 a_4921_30169.n4 a_4921_30169.n2 5.7305
R7961 a_4921_30169.n5 a_4921_30169.n1 0.732092
R7962 a_4921_30169.n0 a_4921_30169.t3 0.7285
R7963 a_4921_30169.n0 a_4921_30169.t2 0.7285
R7964 a_n4631_29217.n0 a_n4631_29217.t6 40.8177
R7965 a_n4631_29217.n1 a_n4631_29217.t5 40.6313
R7966 a_n4631_29217.n1 a_n4631_29217.t7 27.3166
R7967 a_n4631_29217.n0 a_n4631_29217.t4 27.1302
R7968 a_n4631_29217.n2 a_n4631_29217.n1 19.2576
R7969 a_n4631_29217.n3 a_n4631_29217.t3 10.0473
R7970 a_n4631_29217.n4 a_n4631_29217.t2 6.51042
R7971 a_n4631_29217.n5 a_n4631_29217.n4 6.04952
R7972 a_n4631_29217.n2 a_n4631_29217.n0 5.91752
R7973 a_n4631_29217.n3 a_n4631_29217.n2 4.89565
R7974 a_n4631_29217.n4 a_n4631_29217.n3 0.732092
R7975 a_n4631_29217.n5 a_n4631_29217.t1 0.7285
R7976 a_n4631_29217.t0 a_n4631_29217.n5 0.7285
R7977 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t6 41.0041
R7978 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t5 40.8177
R7979 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t4 40.6313
R7980 SARlogic_0.dffrs_7.nand3_6.C.n3 SARlogic_0.dffrs_7.nand3_6.C.t9 27.3166
R7981 SARlogic_0.dffrs_7.nand3_6.C.n0 SARlogic_0.dffrs_7.nand3_6.C.t7 27.1302
R7982 SARlogic_0.dffrs_7.nand3_6.C.n1 SARlogic_0.dffrs_7.nand3_6.C.t8 26.9438
R7983 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.t3 10.0473
R7984 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n4 9.90747
R7985 SARlogic_0.dffrs_7.nand3_6.C.n5 SARlogic_0.dffrs_7.nand3_6.C.n2 9.90116
R7986 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.t2 6.51042
R7987 SARlogic_0.dffrs_7.nand3_6.C.n8 SARlogic_0.dffrs_7.nand3_6.C.n7 6.04952
R7988 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_6.C.n1 5.7305
R7989 SARlogic_0.dffrs_7.nand3_2.B SARlogic_0.dffrs_7.nand3_6.C.n0 5.47979
R7990 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C.n3 5.13907
R7991 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n9 4.72925
R7992 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_6.C.n5 4.5005
R7993 SARlogic_0.dffrs_7.nand3_6.C.n9 SARlogic_0.dffrs_7.nand3_6.C.n8 0.732092
R7994 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t0 0.7285
R7995 SARlogic_0.dffrs_7.nand3_6.C.n7 SARlogic_0.dffrs_7.nand3_6.C.t1 0.7285
R7996 SARlogic_0.dffrs_7.nand3_1.Z SARlogic_0.dffrs_7.nand3_6.C.n6 0.449758
R7997 SARlogic_0.dffrs_7.nand3_6.C.n6 SARlogic_0.dffrs_7.nand3_2.B 0.166901
R7998 SARlogic_0.dffrs_7.nand3_6.C.n2 SARlogic_0.dffrs_7.nand3_0.A 0.0455
R7999 SARlogic_0.dffrs_7.nand3_6.C.n4 SARlogic_0.dffrs_7.nand3_6.C 0.0455
R8000 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t2 41.0041
R8001 adc_PISO_0.2inmux_3.OUT.n0 adc_PISO_0.2inmux_3.OUT.t3 26.9438
R8002 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t0 9.6935
R8003 adc_PISO_0.dffrs_2.d adc_PISO_0.2inmux_3.OUT.n0 6.55979
R8004 adc_PISO_0.2inmux_3.OUT adc_PISO_0.dffrs_2.d 4.883
R8005 adc_PISO_0.2inmux_3.OUT.n1 adc_PISO_0.2inmux_3.OUT.t1 4.35383
R8006 adc_PISO_0.2inmux_3.OUT adc_PISO_0.2inmux_3.OUT.n1 0.350857
R8007 a_14393_30170.n2 a_14393_30170.t4 41.0041
R8008 a_14393_30170.n3 a_14393_30170.t6 40.8177
R8009 a_14393_30170.n3 a_14393_30170.t7 27.1302
R8010 a_14393_30170.n2 a_14393_30170.t5 26.9438
R8011 a_14393_30170.n4 a_14393_30170.n3 22.5284
R8012 a_14393_30170.n5 a_14393_30170.n4 19.5781
R8013 a_14393_30170.t0 a_14393_30170.n5 10.0473
R8014 a_14393_30170.n1 a_14393_30170.t1 6.51042
R8015 a_14393_30170.n1 a_14393_30170.n0 6.04952
R8016 a_14393_30170.n4 a_14393_30170.n2 5.7305
R8017 a_14393_30170.n5 a_14393_30170.n1 0.732092
R8018 a_14393_30170.n0 a_14393_30170.t3 0.7285
R8019 a_14393_30170.n0 a_14393_30170.t2 0.7285
R8020 Vin2.n7 Vin2.n6 23.1032
R8021 Vin2.n3 Vin2.n2 23.1032
R8022 Vin2.n0 Vin2.t6 22.8502
R8023 Vin2.n2 Vin2.t5 16.3656
R8024 Vin2.n6 Vin2.t1 16.3641
R8025 Vin2.n2 Vin2.t2 16.021
R8026 Vin2.n6 Vin2.t4 16.0195
R8027 Vin2.n8 Vin2.t8 11.5195
R8028 Vin2.n5 Vin2.t7 11.5195
R8029 Vin2.n4 Vin2.t0 11.5195
R8030 Vin2.n1 Vin2.t9 11.5195
R8031 Vin2.n0 Vin2.t3 11.5195
R8032 comparator_no_offsetcal_0.Vin2 Vin2 5.6819
R8033 comparator_no_offsetcal_0.Vin2 Vin2.n8 3.94555
R8034 Vin2.n7 Vin2.n5 2.53166
R8035 Vin2.n1 Vin2.n0 2.48408
R8036 Vin2.n3 Vin2.n1 1.40666
R8037 Vin2.n8 Vin2.n7 0.647658
R8038 Vin2.n4 Vin2.n3 0.647132
R8039 Vin2.n5 Vin2.n4 0.234605
R8040 Clk_piso.n19 Clk_piso.t9 41.0041
R8041 Clk_piso.n15 Clk_piso.t16 41.0041
R8042 Clk_piso.n11 Clk_piso.t6 41.0041
R8043 Clk_piso.n7 Clk_piso.t2 41.0041
R8044 Clk_piso.n3 Clk_piso.t0 41.0041
R8045 Clk_piso.n0 Clk_piso.t10 41.0041
R8046 Clk_piso.n20 Clk_piso.t13 40.8177
R8047 Clk_piso.n16 Clk_piso.t11 40.8177
R8048 Clk_piso.n12 Clk_piso.t3 40.8177
R8049 Clk_piso.n8 Clk_piso.t1 40.8177
R8050 Clk_piso.n4 Clk_piso.t15 40.8177
R8051 Clk_piso.n1 Clk_piso.t12 40.8177
R8052 Clk_piso.n20 Clk_piso.t21 27.1302
R8053 Clk_piso.n16 Clk_piso.t19 27.1302
R8054 Clk_piso.n12 Clk_piso.t8 27.1302
R8055 Clk_piso.n8 Clk_piso.t5 27.1302
R8056 Clk_piso.n4 Clk_piso.t22 27.1302
R8057 Clk_piso.n1 Clk_piso.t20 27.1302
R8058 Clk_piso.n19 Clk_piso.t17 26.9438
R8059 Clk_piso.n15 Clk_piso.t23 26.9438
R8060 Clk_piso.n11 Clk_piso.t14 26.9438
R8061 Clk_piso.n7 Clk_piso.t7 26.9438
R8062 Clk_piso.n3 Clk_piso.t4 26.9438
R8063 Clk_piso.n0 Clk_piso.t18 26.9438
R8064 Clk_piso.n6 adc_PISO_0.dffrs_5.clk 23.2034
R8065 Clk_piso.n22 Clk_piso.n18 13.9468
R8066 Clk_piso.n18 Clk_piso.n14 13.9463
R8067 Clk_piso.n10 Clk_piso.n6 13.9457
R8068 Clk_piso.n14 Clk_piso.n10 13.9457
R8069 Clk_piso.n23 Clk_piso 13.1341
R8070 Clk_piso.n22 adc_PISO_0.dffrs_0.clk 9.25764
R8071 Clk_piso.n18 adc_PISO_0.dffrs_1.clk 9.25764
R8072 Clk_piso.n14 adc_PISO_0.dffrs_2.clk 9.25764
R8073 Clk_piso.n10 adc_PISO_0.dffrs_3.clk 9.25764
R8074 Clk_piso.n6 adc_PISO_0.dffrs_4.clk 9.25764
R8075 Clk_piso.n21 Clk_piso.n20 7.65746
R8076 Clk_piso.n17 Clk_piso.n16 7.65746
R8077 Clk_piso.n13 Clk_piso.n12 7.65746
R8078 Clk_piso.n9 Clk_piso.n8 7.65746
R8079 Clk_piso.n5 Clk_piso.n4 7.65746
R8080 Clk_piso.n2 Clk_piso.n1 7.65746
R8081 Clk_piso.n21 Clk_piso.n19 7.12229
R8082 Clk_piso.n17 Clk_piso.n15 7.12229
R8083 Clk_piso.n13 Clk_piso.n11 7.12229
R8084 Clk_piso.n9 Clk_piso.n7 7.12229
R8085 Clk_piso.n5 Clk_piso.n3 7.12229
R8086 Clk_piso.n2 Clk_piso.n0 7.12229
R8087 Clk_piso.n23 Clk_piso.n22 3.49505
R8088 adc_PISO_0.dffrs_0.clk Clk_piso.n21 0.611214
R8089 adc_PISO_0.dffrs_1.clk Clk_piso.n17 0.611214
R8090 adc_PISO_0.dffrs_2.clk Clk_piso.n13 0.611214
R8091 adc_PISO_0.dffrs_3.clk Clk_piso.n9 0.611214
R8092 adc_PISO_0.dffrs_4.clk Clk_piso.n5 0.611214
R8093 adc_PISO_0.dffrs_5.clk Clk_piso.n2 0.611214
R8094 adc_PISO_0.clk Clk_piso.n23 0.0336579
R8095 a_14313_29218.n2 a_14313_29218.t6 40.8177
R8096 a_14313_29218.n3 a_14313_29218.t5 40.6313
R8097 a_14313_29218.n3 a_14313_29218.t4 27.3166
R8098 a_14313_29218.n2 a_14313_29218.t7 27.1302
R8099 a_14313_29218.n4 a_14313_29218.n3 19.2576
R8100 a_14313_29218.t0 a_14313_29218.n5 10.0473
R8101 a_14313_29218.n1 a_14313_29218.t1 6.51042
R8102 a_14313_29218.n1 a_14313_29218.n0 6.04952
R8103 a_14313_29218.n4 a_14313_29218.n2 5.91752
R8104 a_14313_29218.n5 a_14313_29218.n4 4.89565
R8105 a_14313_29218.n5 a_14313_29218.n1 0.732092
R8106 a_14313_29218.n0 a_14313_29218.t3 0.7285
R8107 a_14313_29218.n0 a_14313_29218.t2 0.7285
R8108 a_4841_29217.n0 a_4841_29217.t6 40.8177
R8109 a_4841_29217.n1 a_4841_29217.t5 40.6313
R8110 a_4841_29217.n1 a_4841_29217.t7 27.3166
R8111 a_4841_29217.n0 a_4841_29217.t4 27.1302
R8112 a_4841_29217.n2 a_4841_29217.n1 19.2576
R8113 a_4841_29217.n3 a_4841_29217.t1 10.0473
R8114 a_4841_29217.t0 a_4841_29217.n5 6.51042
R8115 a_4841_29217.n5 a_4841_29217.n4 6.04952
R8116 a_4841_29217.n2 a_4841_29217.n0 5.91752
R8117 a_4841_29217.n3 a_4841_29217.n2 4.89565
R8118 a_4841_29217.n5 a_4841_29217.n3 0.732092
R8119 a_4841_29217.n4 a_4841_29217.t3 0.7285
R8120 a_4841_29217.n4 a_4841_29217.t2 0.7285
R8121 SARlogic_0.d4.n3 SARlogic_0.d4.t11 41.0041
R8122 SARlogic_0.d4.n4 SARlogic_0.d4.t12 40.8177
R8123 SARlogic_0.d4.n7 SARlogic_0.d4.t7 40.6313
R8124 SARlogic_0.d4.n1 SARlogic_0.d4.t10 34.2529
R8125 SARlogic_0.d4.n6 SARlogic_0.dffrs_14.clk 33.675
R8126 SARlogic_0.d4.n7 SARlogic_0.d4.t5 27.3166
R8127 SARlogic_0.d4.n4 SARlogic_0.d4.t8 27.1302
R8128 SARlogic_0.d4.n3 SARlogic_0.d4.t4 26.9438
R8129 SARlogic_0.d4.n0 SARlogic_0.d4.t6 19.673
R8130 SARlogic_0.d4.n0 SARlogic_0.d4.t9 19.4007
R8131 SARlogic_0.d4.n9 SARlogic_0.d4.n8 14.0582
R8132 SARlogic_0.d4.n9 SARlogic_0.d4.n6 11.3593
R8133 SARlogic_0.d4.n12 SARlogic_0.d4.t1 10.0473
R8134 SARlogic_0.d4.n2 SARlogic_0.d4.n1 8.05164
R8135 SARlogic_0.d4.n11 SARlogic_0.d4.t2 6.51042
R8136 SARlogic_0.d4.n11 SARlogic_0.d4.n10 6.04952
R8137 SARlogic_0.dffrs_14.nand3_1.A SARlogic_0.d4.n3 5.7755
R8138 SARlogic_0.dffrs_14.nand3_6.B SARlogic_0.d4.n4 5.47979
R8139 SARlogic_0.d4.n8 SARlogic_0.d4.n7 5.13907
R8140 SARlogic_0.dffrs_7.nand3_2.Z SARlogic_0.d4.n12 4.72925
R8141 SARlogic_0.d4.n6 adc_PISO_0.B5 3.49604
R8142 SARlogic_0.d4.n5 SARlogic_0.dffrs_14.nand3_6.B 2.17818
R8143 adc_PISO_0.B5 SARlogic_0.d4.n2 1.87121
R8144 SARlogic_0.d4.n5 SARlogic_0.dffrs_14.nand3_1.A 1.34729
R8145 SARlogic_0.d4.n12 SARlogic_0.d4.n11 0.732092
R8146 SARlogic_0.d4.n10 SARlogic_0.d4.t0 0.7285
R8147 SARlogic_0.d4.n10 SARlogic_0.d4.t3 0.7285
R8148 SARlogic_0.dffrs_14.clk SARlogic_0.d4.n5 0.611214
R8149 SARlogic_0.dffrs_7.nand3_2.Z SARlogic_0.d4.n9 0.166901
R8150 SARlogic_0.d4.n1 SARlogic_0.d4.n0 0.106438
R8151 SARlogic_0.d4.n8 SARlogic_0.dffrs_7.nand3_7.C 0.0455
R8152 SARlogic_0.d4.n2 adc_PISO_0.2inmux_2.In 0.0455
R8153 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t5 41.0041
R8154 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t7 40.6313
R8155 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t8 40.6313
R8156 SARlogic_0.dffrs_4.Qb SARlogic_0.dffrs_11.setb 28.021
R8157 SARlogic_0.dffrs_4.Qb.n4 SARlogic_0.dffrs_4.Qb.t9 27.3166
R8158 SARlogic_0.dffrs_4.Qb.n2 SARlogic_0.dffrs_4.Qb.t4 27.3166
R8159 SARlogic_0.dffrs_4.Qb.n0 SARlogic_0.dffrs_4.Qb.t6 26.9438
R8160 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.t0 10.0473
R8161 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb.n1 9.84255
R8162 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n3 9.22229
R8163 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.t1 6.51042
R8164 SARlogic_0.dffrs_4.Qb.n8 SARlogic_0.dffrs_4.Qb.n7 6.04952
R8165 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.Qb.n0 5.7305
R8166 SARlogic_0.dffrs_4.Qb.n5 SARlogic_0.dffrs_4.Qb.n4 5.14711
R8167 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_4.Qb.n2 5.13907
R8168 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n6 4.94976
R8169 SARlogic_0.dffrs_4.nand3_7.Z SARlogic_0.dffrs_4.Qb.n9 4.72925
R8170 SARlogic_0.dffrs_11.setb SARlogic_0.dffrs_11.nand3_0.C 0.784786
R8171 SARlogic_0.dffrs_4.Qb.n9 SARlogic_0.dffrs_4.Qb.n8 0.732092
R8172 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t3 0.7285
R8173 SARlogic_0.dffrs_4.Qb.n7 SARlogic_0.dffrs_4.Qb.t2 0.7285
R8174 SARlogic_0.dffrs_4.Qb.n6 SARlogic_0.dffrs_4.Qb 0.175225
R8175 SARlogic_0.dffrs_4.Qb.n1 SARlogic_0.dffrs_4.nand3_2.A 0.0455
R8176 SARlogic_0.dffrs_4.Qb.n3 SARlogic_0.dffrs_11.nand3_2.C 0.0455
R8177 SARlogic_0.dffrs_11.nand3_0.C SARlogic_0.dffrs_4.Qb.n5 0.0374643
R8178 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t6 40.8177
R8179 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t5 40.6313
R8180 SARlogic_0.dffrs_8.nand3_8.C.n1 SARlogic_0.dffrs_8.nand3_8.C.t7 27.3166
R8181 SARlogic_0.dffrs_8.nand3_8.C.n0 SARlogic_0.dffrs_8.nand3_8.C.t4 27.1302
R8182 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_8.C.n2 14.119
R8183 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.t1 10.0473
R8184 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.t2 6.51042
R8185 SARlogic_0.dffrs_8.nand3_8.C.n5 SARlogic_0.dffrs_8.nand3_8.C.n4 6.04952
R8186 SARlogic_0.dffrs_8.nand3_7.B SARlogic_0.dffrs_8.nand3_8.C.n0 5.47979
R8187 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C.n1 5.13907
R8188 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n6 4.72925
R8189 SARlogic_0.dffrs_8.nand3_8.C.n6 SARlogic_0.dffrs_8.nand3_8.C.n5 0.732092
R8190 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t0 0.7285
R8191 SARlogic_0.dffrs_8.nand3_8.C.n4 SARlogic_0.dffrs_8.nand3_8.C.t3 0.7285
R8192 SARlogic_0.dffrs_8.nand3_8.C.n3 SARlogic_0.dffrs_8.nand3_7.B 0.438233
R8193 SARlogic_0.dffrs_8.nand3_6.Z SARlogic_0.dffrs_8.nand3_8.C.n3 0.166901
R8194 SARlogic_0.dffrs_8.nand3_8.C.n2 SARlogic_0.dffrs_8.nand3_8.C 0.0455
R8195 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t5 41.0041
R8196 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t6 40.8177
R8197 SARlogic_0.dffrs_2.nand3_8.Z.n1 SARlogic_0.dffrs_2.nand3_8.Z.t4 27.1302
R8198 SARlogic_0.dffrs_2.nand3_8.Z.n0 SARlogic_0.dffrs_2.nand3_8.Z.t7 26.9438
R8199 SARlogic_0.dffrs_2.nand3_6.A SARlogic_0.dffrs_2.nand3_0.B 17.0041
R8200 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n2 14.8493
R8201 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.t1 10.0473
R8202 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.t0 6.51042
R8203 SARlogic_0.dffrs_2.nand3_8.Z.n4 SARlogic_0.dffrs_2.nand3_8.Z.n3 6.04952
R8204 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_8.Z.n0 5.7305
R8205 SARlogic_0.dffrs_2.nand3_0.B SARlogic_0.dffrs_2.nand3_8.Z.n1 5.47979
R8206 SARlogic_0.dffrs_2.nand3_8.Z SARlogic_0.dffrs_2.nand3_8.Z.n5 4.72925
R8207 SARlogic_0.dffrs_2.nand3_8.Z.n5 SARlogic_0.dffrs_2.nand3_8.Z.n4 0.732092
R8208 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t2 0.7285
R8209 SARlogic_0.dffrs_2.nand3_8.Z.n3 SARlogic_0.dffrs_2.nand3_8.Z.t3 0.7285
R8210 SARlogic_0.dffrs_2.nand3_8.Z.n2 SARlogic_0.dffrs_2.nand3_6.A 0.0455
R8211 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t5 40.6313
R8212 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.t6 34.1066
R8213 adc_PISO_0.dffrs_3.Q.n3 adc_PISO_0.dffrs_3.Q.t7 27.3166
R8214 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t8 19.673
R8215 adc_PISO_0.dffrs_3.Q.n0 adc_PISO_0.dffrs_3.Q.t4 19.4007
R8216 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n3 14.6967
R8217 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.t0 10.0473
R8218 adc_PISO_0.dffrs_3.Q.n7 adc_PISO_0.dffrs_3.Q.n6 9.39565
R8219 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.dffrs_3.Q.n1 6.70486
R8220 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.t1 6.51042
R8221 adc_PISO_0.dffrs_3.Q.n5 adc_PISO_0.dffrs_3.Q.n4 6.04952
R8222 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n2 5.81514
R8223 adc_PISO_0.dffrs_3.Q.n6 adc_PISO_0.dffrs_3.Q.n5 0.732092
R8224 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t3 0.7285
R8225 adc_PISO_0.dffrs_3.Q.n4 adc_PISO_0.dffrs_3.Q.t2 0.7285
R8226 adc_PISO_0.dffrs_3.Q adc_PISO_0.dffrs_3.Q.n7 0.458082
R8227 adc_PISO_0.dffrs_3.Q.n1 adc_PISO_0.dffrs_3.Q.n0 0.252687
R8228 adc_PISO_0.dffrs_3.Q.n2 adc_PISO_0.2inmux_5.Bit 0.0519286
R8229 a_39727_29264.n0 a_39727_29264.t5 34.1797
R8230 a_39727_29264.n0 a_39727_29264.t4 19.5798
R8231 a_39727_29264.n3 a_39727_29264.t3 10.3401
R8232 a_39727_29264.t0 a_39727_29264.n3 9.2885
R8233 a_39727_29264.n2 a_39727_29264.n0 4.93379
R8234 a_39727_29264.n1 a_39727_29264.t1 4.09202
R8235 a_39727_29264.n1 a_39727_29264.t2 3.95079
R8236 a_39727_29264.n3 a_39727_29264.n2 0.599711
R8237 a_39727_29264.n2 a_39727_29264.n1 0.296375
R8238 a_42809_30170.n0 a_42809_30170.t5 41.0041
R8239 a_42809_30170.n1 a_42809_30170.t7 40.8177
R8240 a_42809_30170.n1 a_42809_30170.t4 27.1302
R8241 a_42809_30170.n0 a_42809_30170.t6 26.9438
R8242 a_42809_30170.n2 a_42809_30170.n1 22.5284
R8243 a_42809_30170.n3 a_42809_30170.n2 19.5781
R8244 a_42809_30170.n3 a_42809_30170.t3 10.0473
R8245 a_42809_30170.n4 a_42809_30170.t2 6.51042
R8246 a_42809_30170.n5 a_42809_30170.n4 6.04952
R8247 a_42809_30170.n2 a_42809_30170.n0 5.7305
R8248 a_42809_30170.n4 a_42809_30170.n3 0.732092
R8249 a_42809_30170.n5 a_42809_30170.t1 0.7285
R8250 a_42809_30170.t0 a_42809_30170.n5 0.7285
R8251 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t7 40.8177
R8252 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t5 40.6313
R8253 SARlogic_0.dffrs_10.nand3_8.C.n1 SARlogic_0.dffrs_10.nand3_8.C.t6 27.3166
R8254 SARlogic_0.dffrs_10.nand3_8.C.n0 SARlogic_0.dffrs_10.nand3_8.C.t4 27.1302
R8255 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_8.C.n2 14.119
R8256 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.t1 10.0473
R8257 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.t0 6.51042
R8258 SARlogic_0.dffrs_10.nand3_8.C.n5 SARlogic_0.dffrs_10.nand3_8.C.n4 6.04952
R8259 SARlogic_0.dffrs_10.nand3_7.B SARlogic_0.dffrs_10.nand3_8.C.n0 5.47979
R8260 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C.n1 5.13907
R8261 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n6 4.72925
R8262 SARlogic_0.dffrs_10.nand3_8.C.n6 SARlogic_0.dffrs_10.nand3_8.C.n5 0.732092
R8263 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t2 0.7285
R8264 SARlogic_0.dffrs_10.nand3_8.C.n4 SARlogic_0.dffrs_10.nand3_8.C.t3 0.7285
R8265 SARlogic_0.dffrs_10.nand3_8.C.n3 SARlogic_0.dffrs_10.nand3_7.B 0.438233
R8266 SARlogic_0.dffrs_10.nand3_6.Z SARlogic_0.dffrs_10.nand3_8.C.n3 0.166901
R8267 SARlogic_0.dffrs_10.nand3_8.C.n2 SARlogic_0.dffrs_10.nand3_8.C 0.0455
R8268 adc_PISO_0.serial_out Piso_out 68.5339
R8269 Piso_out.n0 Piso_out.t5 40.6313
R8270 Piso_out.n0 Piso_out.t4 27.3166
R8271 Piso_out.n4 Piso_out.n0 14.6967
R8272 Piso_out.n3 Piso_out.t1 10.0473
R8273 Piso_out.n4 Piso_out.n3 9.39565
R8274 Piso_out.n2 Piso_out.t2 6.51042
R8275 Piso_out.n2 Piso_out.n1 6.04952
R8276 adc_PISO_0.serial_out adc_PISO_0.dffrs_5.Q 5.90514
R8277 Piso_out.n3 Piso_out.n2 0.732092
R8278 Piso_out.n1 Piso_out.t0 0.7285
R8279 Piso_out.n1 Piso_out.t3 0.7285
R8280 adc_PISO_0.dffrs_5.Q Piso_out.n4 0.458082
R8281 a_n4551_30169.n0 a_n4551_30169.t5 41.0041
R8282 a_n4551_30169.n1 a_n4551_30169.t7 40.8177
R8283 a_n4551_30169.n1 a_n4551_30169.t4 27.1302
R8284 a_n4551_30169.n0 a_n4551_30169.t6 26.9438
R8285 a_n4551_30169.n2 a_n4551_30169.n1 22.5284
R8286 a_n4551_30169.n3 a_n4551_30169.n2 19.5781
R8287 a_n4551_30169.n3 a_n4551_30169.t3 10.0473
R8288 a_n4551_30169.n4 a_n4551_30169.t1 6.51042
R8289 a_n4551_30169.n5 a_n4551_30169.n4 6.04952
R8290 a_n4551_30169.n2 a_n4551_30169.n0 5.7305
R8291 a_n4551_30169.n4 a_n4551_30169.n3 0.732092
R8292 a_n4551_30169.n5 a_n4551_30169.t2 0.7285
R8293 a_n4551_30169.t0 a_n4551_30169.n5 0.7285
R8294 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t4 41.0041
R8295 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t5 40.8177
R8296 SARlogic_0.dffrs_0.nand3_8.Z.n1 SARlogic_0.dffrs_0.nand3_8.Z.t7 27.1302
R8297 SARlogic_0.dffrs_0.nand3_8.Z.n0 SARlogic_0.dffrs_0.nand3_8.Z.t6 26.9438
R8298 SARlogic_0.dffrs_0.nand3_6.A SARlogic_0.dffrs_0.nand3_0.B 17.0041
R8299 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n2 14.8493
R8300 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.t2 10.0473
R8301 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.t3 6.51042
R8302 SARlogic_0.dffrs_0.nand3_8.Z.n4 SARlogic_0.dffrs_0.nand3_8.Z.n3 6.04952
R8303 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_8.Z.n0 5.7305
R8304 SARlogic_0.dffrs_0.nand3_0.B SARlogic_0.dffrs_0.nand3_8.Z.n1 5.47979
R8305 SARlogic_0.dffrs_0.nand3_8.Z SARlogic_0.dffrs_0.nand3_8.Z.n5 4.72925
R8306 SARlogic_0.dffrs_0.nand3_8.Z.n5 SARlogic_0.dffrs_0.nand3_8.Z.n4 0.732092
R8307 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t0 0.7285
R8308 SARlogic_0.dffrs_0.nand3_8.Z.n3 SARlogic_0.dffrs_0.nand3_8.Z.t1 0.7285
R8309 SARlogic_0.dffrs_0.nand3_8.Z.n2 SARlogic_0.dffrs_0.nand3_6.A 0.0455
R8310 a_11311_29264.n0 a_11311_29264.t5 34.1797
R8311 a_11311_29264.n0 a_11311_29264.t4 19.5798
R8312 a_11311_29264.n3 a_11311_29264.t3 10.3401
R8313 a_11311_29264.t0 a_11311_29264.n3 9.2885
R8314 a_11311_29264.n2 a_11311_29264.n0 4.93379
R8315 a_11311_29264.n1 a_11311_29264.t2 4.09202
R8316 a_11311_29264.n1 a_11311_29264.t1 3.95079
R8317 a_11311_29264.n3 a_11311_29264.n2 0.599711
R8318 a_11311_29264.n2 a_11311_29264.n1 0.296375
R8319 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t7 41.0041
R8320 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t4 40.8177
R8321 SARlogic_0.dffrs_5.nand3_8.Z.n1 SARlogic_0.dffrs_5.nand3_8.Z.t5 27.1302
R8322 SARlogic_0.dffrs_5.nand3_8.Z.n0 SARlogic_0.dffrs_5.nand3_8.Z.t6 26.9438
R8323 SARlogic_0.dffrs_5.nand3_6.A SARlogic_0.dffrs_5.nand3_0.B 17.0041
R8324 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n2 14.8493
R8325 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.t2 10.0473
R8326 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.t1 6.51042
R8327 SARlogic_0.dffrs_5.nand3_8.Z.n4 SARlogic_0.dffrs_5.nand3_8.Z.n3 6.04952
R8328 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_8.Z.n0 5.7305
R8329 SARlogic_0.dffrs_5.nand3_0.B SARlogic_0.dffrs_5.nand3_8.Z.n1 5.47979
R8330 SARlogic_0.dffrs_5.nand3_8.Z SARlogic_0.dffrs_5.nand3_8.Z.n5 4.72925
R8331 SARlogic_0.dffrs_5.nand3_8.Z.n5 SARlogic_0.dffrs_5.nand3_8.Z.n4 0.732092
R8332 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t0 0.7285
R8333 SARlogic_0.dffrs_5.nand3_8.Z.n3 SARlogic_0.dffrs_5.nand3_8.Z.t3 0.7285
R8334 SARlogic_0.dffrs_5.nand3_8.Z.n2 SARlogic_0.dffrs_5.nand3_6.A 0.0455
R8335 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t7 40.8177
R8336 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t5 40.6313
R8337 SARlogic_0.dffrs_13.nand3_8.C.n1 SARlogic_0.dffrs_13.nand3_8.C.t6 27.3166
R8338 SARlogic_0.dffrs_13.nand3_8.C.n0 SARlogic_0.dffrs_13.nand3_8.C.t4 27.1302
R8339 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_8.C.n2 14.119
R8340 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.t1 10.0473
R8341 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.t2 6.51042
R8342 SARlogic_0.dffrs_13.nand3_8.C.n5 SARlogic_0.dffrs_13.nand3_8.C.n4 6.04952
R8343 SARlogic_0.dffrs_13.nand3_7.B SARlogic_0.dffrs_13.nand3_8.C.n0 5.47979
R8344 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C.n1 5.13907
R8345 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n6 4.72925
R8346 SARlogic_0.dffrs_13.nand3_8.C.n6 SARlogic_0.dffrs_13.nand3_8.C.n5 0.732092
R8347 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t0 0.7285
R8348 SARlogic_0.dffrs_13.nand3_8.C.n4 SARlogic_0.dffrs_13.nand3_8.C.t3 0.7285
R8349 SARlogic_0.dffrs_13.nand3_8.C.n3 SARlogic_0.dffrs_13.nand3_7.B 0.438233
R8350 SARlogic_0.dffrs_13.nand3_6.Z SARlogic_0.dffrs_13.nand3_8.C.n3 0.166901
R8351 SARlogic_0.dffrs_13.nand3_8.C.n2 SARlogic_0.dffrs_13.nand3_8.C 0.0455
R8352 a_n7633_29263.n0 a_n7633_29263.t4 34.1797
R8353 a_n7633_29263.n0 a_n7633_29263.t5 19.5798
R8354 a_n7633_29263.t0 a_n7633_29263.n3 10.3401
R8355 a_n7633_29263.n3 a_n7633_29263.t1 9.2885
R8356 a_n7633_29263.n2 a_n7633_29263.n0 4.93379
R8357 a_n7633_29263.n1 a_n7633_29263.t2 4.09202
R8358 a_n7633_29263.n1 a_n7633_29263.t3 3.95079
R8359 a_n7633_29263.n3 a_n7633_29263.n2 0.599711
R8360 a_n7633_29263.n2 a_n7633_29263.n1 0.296375
R8361 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t2 41.0041
R8362 adc_PISO_0.2inmux_0.OUT.n0 adc_PISO_0.2inmux_0.OUT.t3 26.9438
R8363 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t0 9.6935
R8364 adc_PISO_0.dffrs_0.d adc_PISO_0.2inmux_0.OUT.n0 6.55979
R8365 adc_PISO_0.2inmux_0.OUT adc_PISO_0.dffrs_0.d 4.883
R8366 adc_PISO_0.2inmux_0.OUT.n1 adc_PISO_0.2inmux_0.OUT.t1 4.35383
R8367 adc_PISO_0.2inmux_0.OUT adc_PISO_0.2inmux_0.OUT.n1 0.350857
R8368 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t4 41.0041
R8369 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t6 40.6313
R8370 SARlogic_0.dffrs_4.Q.n1 SARlogic_0.dffrs_4.Q.t7 27.3166
R8371 SARlogic_0.dffrs_4.Q.n0 SARlogic_0.dffrs_4.Q.t5 26.9438
R8372 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_5.d 17.5382
R8373 SARlogic_0.dffrs_4.Q.n3 SARlogic_0.dffrs_4.Q.n2 14.0582
R8374 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.t0 10.0473
R8375 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.t1 6.51042
R8376 SARlogic_0.dffrs_4.Q.n5 SARlogic_0.dffrs_4.Q.n4 6.04952
R8377 SARlogic_0.dffrs_5.nand3_8.A SARlogic_0.dffrs_4.Q.n0 5.7755
R8378 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.Q.n1 5.13907
R8379 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n6 4.72925
R8380 SARlogic_0.dffrs_5.d SARlogic_0.dffrs_5.nand3_8.A 0.784786
R8381 SARlogic_0.dffrs_4.Q.n6 SARlogic_0.dffrs_4.Q.n5 0.732092
R8382 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t3 0.7285
R8383 SARlogic_0.dffrs_4.Q.n4 SARlogic_0.dffrs_4.Q.t2 0.7285
R8384 SARlogic_0.dffrs_4.nand3_2.Z SARlogic_0.dffrs_4.Q.n3 0.166901
R8385 SARlogic_0.dffrs_4.Q.n2 SARlogic_0.dffrs_4.nand3_7.C 0.0455
R8386 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t4 41.0041
R8387 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t7 40.6313
R8388 SARlogic_0.dffrs_0.Q.n1 SARlogic_0.dffrs_0.Q.t6 27.3166
R8389 SARlogic_0.dffrs_0.Q.n0 SARlogic_0.dffrs_0.Q.t5 26.9438
R8390 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_1.d 17.5382
R8391 SARlogic_0.dffrs_0.Q.n3 SARlogic_0.dffrs_0.Q.n2 14.0582
R8392 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.t1 10.0473
R8393 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.t2 6.51042
R8394 SARlogic_0.dffrs_0.Q.n5 SARlogic_0.dffrs_0.Q.n4 6.04952
R8395 SARlogic_0.dffrs_1.nand3_8.A SARlogic_0.dffrs_0.Q.n0 5.7755
R8396 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.Q.n1 5.13907
R8397 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n6 4.72925
R8398 SARlogic_0.dffrs_1.d SARlogic_0.dffrs_1.nand3_8.A 0.784786
R8399 SARlogic_0.dffrs_0.Q.n6 SARlogic_0.dffrs_0.Q.n5 0.732092
R8400 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t3 0.7285
R8401 SARlogic_0.dffrs_0.Q.n4 SARlogic_0.dffrs_0.Q.t0 0.7285
R8402 SARlogic_0.dffrs_0.nand3_2.Z SARlogic_0.dffrs_0.Q.n3 0.166901
R8403 SARlogic_0.dffrs_0.Q.n2 SARlogic_0.dffrs_0.nand3_7.C 0.0455
R8404 a_18555_28820.n0 a_18555_28820.t5 34.1797
R8405 a_18555_28820.n0 a_18555_28820.t4 19.5798
R8406 a_18555_28820.n1 a_18555_28820.t3 18.7717
R8407 a_18555_28820.n1 a_18555_28820.t2 9.2885
R8408 a_18555_28820.n2 a_18555_28820.n0 4.93379
R8409 a_18555_28820.t0 a_18555_28820.n3 4.23346
R8410 a_18555_28820.n3 a_18555_28820.t1 3.85546
R8411 a_18555_28820.n2 a_18555_28820.n1 0.4055
R8412 a_18555_28820.n3 a_18555_28820.n2 0.352625
R8413 a_23785_33628.n0 a_23785_33628.t4 40.6313
R8414 a_23785_33628.n0 a_23785_33628.t5 27.3166
R8415 a_23785_33628.n1 a_23785_33628.n0 24.1527
R8416 a_23785_33628.n1 a_23785_33628.t2 10.0473
R8417 a_23785_33628.n2 a_23785_33628.t3 6.51042
R8418 a_23785_33628.n3 a_23785_33628.n2 6.04952
R8419 a_23785_33628.n2 a_23785_33628.n1 0.732092
R8420 a_23785_33628.n3 a_23785_33628.t1 0.7285
R8421 a_23785_33628.t0 a_23785_33628.n3 0.7285
R8422 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t6 41.0041
R8423 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t5 40.8177
R8424 SARlogic_0.dffrs_1.nand3_8.Z.n1 SARlogic_0.dffrs_1.nand3_8.Z.t4 27.1302
R8425 SARlogic_0.dffrs_1.nand3_8.Z.n0 SARlogic_0.dffrs_1.nand3_8.Z.t7 26.9438
R8426 SARlogic_0.dffrs_1.nand3_6.A SARlogic_0.dffrs_1.nand3_0.B 17.0041
R8427 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n2 14.8493
R8428 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.t1 10.0473
R8429 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.t2 6.51042
R8430 SARlogic_0.dffrs_1.nand3_8.Z.n4 SARlogic_0.dffrs_1.nand3_8.Z.n3 6.04952
R8431 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_8.Z.n0 5.7305
R8432 SARlogic_0.dffrs_1.nand3_0.B SARlogic_0.dffrs_1.nand3_8.Z.n1 5.47979
R8433 SARlogic_0.dffrs_1.nand3_8.Z SARlogic_0.dffrs_1.nand3_8.Z.n5 4.72925
R8434 SARlogic_0.dffrs_1.nand3_8.Z.n5 SARlogic_0.dffrs_1.nand3_8.Z.n4 0.732092
R8435 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t0 0.7285
R8436 SARlogic_0.dffrs_1.nand3_8.Z.n3 SARlogic_0.dffrs_1.nand3_8.Z.t3 0.7285
R8437 SARlogic_0.dffrs_1.nand3_8.Z.n2 SARlogic_0.dffrs_1.nand3_6.A 0.0455
R8438 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t4 41.0041
R8439 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t7 40.6313
R8440 SARlogic_0.dffrs_2.d.n1 SARlogic_0.dffrs_2.d.t6 27.3166
R8441 SARlogic_0.dffrs_2.d.n0 SARlogic_0.dffrs_2.d.t5 26.9438
R8442 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d 17.5382
R8443 SARlogic_0.dffrs_2.d.n3 SARlogic_0.dffrs_2.d.n2 14.0582
R8444 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.t1 10.0473
R8445 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.t2 6.51042
R8446 SARlogic_0.dffrs_2.d.n5 SARlogic_0.dffrs_2.d.n4 6.04952
R8447 SARlogic_0.dffrs_2.nand3_8.A SARlogic_0.dffrs_2.d.n0 5.7755
R8448 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_2.d.n1 5.13907
R8449 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n6 4.72925
R8450 SARlogic_0.dffrs_2.d SARlogic_0.dffrs_2.nand3_8.A 0.784786
R8451 SARlogic_0.dffrs_2.d.n6 SARlogic_0.dffrs_2.d.n5 0.732092
R8452 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t0 0.7285
R8453 SARlogic_0.dffrs_2.d.n4 SARlogic_0.dffrs_2.d.t3 0.7285
R8454 SARlogic_0.dffrs_1.nand3_2.Z SARlogic_0.dffrs_2.d.n3 0.166901
R8455 SARlogic_0.dffrs_2.d.n2 SARlogic_0.dffrs_1.nand3_7.C 0.0455
R8456 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t5 40.6313
R8457 SARlogic_0.dffrs_5.Q.n0 SARlogic_0.dffrs_5.Q.t4 27.3166
R8458 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n1 14.2246
R8459 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.t1 10.0473
R8460 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.t2 6.51042
R8461 SARlogic_0.dffrs_5.Q.n3 SARlogic_0.dffrs_5.Q.n2 6.04952
R8462 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.Q.n0 5.13907
R8463 SARlogic_0.dffrs_5.nand3_2.Z SARlogic_0.dffrs_5.Q.n4 4.72925
R8464 SARlogic_0.dffrs_5.Q.n4 SARlogic_0.dffrs_5.Q.n3 0.732092
R8465 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t0 0.7285
R8466 SARlogic_0.dffrs_5.Q.n2 SARlogic_0.dffrs_5.Q.t3 0.7285
R8467 SARlogic_0.dffrs_5.Q.n1 SARlogic_0.dffrs_5.nand3_7.C 0.0455
R8468 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t5 41.0041
R8469 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t6 40.8177
R8470 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t4 40.6313
R8471 SARlogic_0.dffrs_4.nand3_6.C.n3 SARlogic_0.dffrs_4.nand3_6.C.t7 27.3166
R8472 SARlogic_0.dffrs_4.nand3_6.C.n0 SARlogic_0.dffrs_4.nand3_6.C.t8 27.1302
R8473 SARlogic_0.dffrs_4.nand3_6.C.n1 SARlogic_0.dffrs_4.nand3_6.C.t9 26.9438
R8474 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.t2 10.0473
R8475 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n4 9.90747
R8476 SARlogic_0.dffrs_4.nand3_6.C.n5 SARlogic_0.dffrs_4.nand3_6.C.n2 9.90116
R8477 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.t3 6.51042
R8478 SARlogic_0.dffrs_4.nand3_6.C.n8 SARlogic_0.dffrs_4.nand3_6.C.n7 6.04952
R8479 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_6.C.n1 5.7305
R8480 SARlogic_0.dffrs_4.nand3_2.B SARlogic_0.dffrs_4.nand3_6.C.n0 5.47979
R8481 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C.n3 5.13907
R8482 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n9 4.72925
R8483 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_6.C.n5 4.5005
R8484 SARlogic_0.dffrs_4.nand3_6.C.n9 SARlogic_0.dffrs_4.nand3_6.C.n8 0.732092
R8485 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t0 0.7285
R8486 SARlogic_0.dffrs_4.nand3_6.C.n7 SARlogic_0.dffrs_4.nand3_6.C.t1 0.7285
R8487 SARlogic_0.dffrs_4.nand3_1.Z SARlogic_0.dffrs_4.nand3_6.C.n6 0.449758
R8488 SARlogic_0.dffrs_4.nand3_6.C.n6 SARlogic_0.dffrs_4.nand3_2.B 0.166901
R8489 SARlogic_0.dffrs_4.nand3_6.C.n2 SARlogic_0.dffrs_4.nand3_0.A 0.0455
R8490 SARlogic_0.dffrs_4.nand3_6.C.n4 SARlogic_0.dffrs_4.nand3_6.C 0.0455
R8491 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t2 41.0041
R8492 adc_PISO_0.2inmux_1.OUT.n0 adc_PISO_0.2inmux_1.OUT.t3 26.9438
R8493 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t0 9.6935
R8494 adc_PISO_0.dffrs_5.d adc_PISO_0.2inmux_1.OUT.n0 6.55979
R8495 adc_PISO_0.2inmux_1.OUT adc_PISO_0.dffrs_5.d 4.883
R8496 adc_PISO_0.2inmux_1.OUT.n1 adc_PISO_0.2inmux_1.OUT.t1 4.35383
R8497 adc_PISO_0.2inmux_1.OUT adc_PISO_0.2inmux_1.OUT.n1 0.350857
R8498 Load.n0 Load.t1 34.1797
R8499 Load.n0 Load.t0 19.5798
R8500 inv2_0.in Load.n0 4.87271
R8501 inv2_0.in Load 0.868357
R8502 a_42729_29218.n0 a_42729_29218.t5 40.8177
R8503 a_42729_29218.n1 a_42729_29218.t6 40.6313
R8504 a_42729_29218.n1 a_42729_29218.t4 27.3166
R8505 a_42729_29218.n0 a_42729_29218.t7 27.1302
R8506 a_42729_29218.n2 a_42729_29218.n1 19.2576
R8507 a_42729_29218.n3 a_42729_29218.t1 10.0473
R8508 a_42729_29218.n4 a_42729_29218.t2 6.51042
R8509 a_42729_29218.n5 a_42729_29218.n4 6.04952
R8510 a_42729_29218.n2 a_42729_29218.n0 5.91752
R8511 a_42729_29218.n3 a_42729_29218.n2 4.89565
R8512 a_42729_29218.n4 a_42729_29218.n3 0.732092
R8513 a_42729_29218.n5 a_42729_29218.t3 0.7285
R8514 a_42729_29218.t0 a_42729_29218.n5 0.7285
R8515 a_18555_31160.n0 a_18555_31160.t5 34.1797
R8516 a_18555_31160.n0 a_18555_31160.t4 19.5798
R8517 a_18555_31160.n1 a_18555_31160.t1 18.7717
R8518 a_18555_31160.n1 a_18555_31160.t2 9.2885
R8519 a_18555_31160.n2 a_18555_31160.n0 4.93379
R8520 a_18555_31160.t0 a_18555_31160.n3 4.23346
R8521 a_18555_31160.n3 a_18555_31160.t3 3.85546
R8522 a_18555_31160.n2 a_18555_31160.n1 0.4055
R8523 a_18555_31160.n3 a_18555_31160.n2 0.352625
R8524 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t7 41.0041
R8525 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t5 40.8177
R8526 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t6 40.6313
R8527 SARlogic_0.dffrs_13.nand3_6.C.n3 SARlogic_0.dffrs_13.nand3_6.C.t9 27.3166
R8528 SARlogic_0.dffrs_13.nand3_6.C.n0 SARlogic_0.dffrs_13.nand3_6.C.t8 27.1302
R8529 SARlogic_0.dffrs_13.nand3_6.C.n1 SARlogic_0.dffrs_13.nand3_6.C.t4 26.9438
R8530 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.t0 10.0473
R8531 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n4 9.90747
R8532 SARlogic_0.dffrs_13.nand3_6.C.n5 SARlogic_0.dffrs_13.nand3_6.C.n2 9.90116
R8533 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.t1 6.51042
R8534 SARlogic_0.dffrs_13.nand3_6.C.n8 SARlogic_0.dffrs_13.nand3_6.C.n7 6.04952
R8535 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_6.C.n1 5.7305
R8536 SARlogic_0.dffrs_13.nand3_2.B SARlogic_0.dffrs_13.nand3_6.C.n0 5.47979
R8537 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C.n3 5.13907
R8538 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n9 4.72925
R8539 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_6.C.n5 4.5005
R8540 SARlogic_0.dffrs_13.nand3_6.C.n9 SARlogic_0.dffrs_13.nand3_6.C.n8 0.732092
R8541 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t2 0.7285
R8542 SARlogic_0.dffrs_13.nand3_6.C.n7 SARlogic_0.dffrs_13.nand3_6.C.t3 0.7285
R8543 SARlogic_0.dffrs_13.nand3_1.Z SARlogic_0.dffrs_13.nand3_6.C.n6 0.449758
R8544 SARlogic_0.dffrs_13.nand3_6.C.n6 SARlogic_0.dffrs_13.nand3_2.B 0.166901
R8545 SARlogic_0.dffrs_13.nand3_6.C.n2 SARlogic_0.dffrs_13.nand3_0.A 0.0455
R8546 SARlogic_0.dffrs_13.nand3_6.C.n4 SARlogic_0.dffrs_13.nand3_6.C 0.0455
R8547 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t4 40.6313
R8548 SARlogic_0.dffrs_13.nand3_1.C.n0 SARlogic_0.dffrs_13.nand3_1.C.t5 27.3166
R8549 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n1 14.2854
R8550 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.t2 10.0473
R8551 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.t3 6.51042
R8552 SARlogic_0.dffrs_13.nand3_1.C.n3 SARlogic_0.dffrs_13.nand3_1.C.n2 6.04952
R8553 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C.n0 5.13907
R8554 SARlogic_0.dffrs_13.nand3_0.Z SARlogic_0.dffrs_13.nand3_1.C.n4 4.72925
R8555 SARlogic_0.dffrs_13.nand3_1.C.n4 SARlogic_0.dffrs_13.nand3_1.C.n3 0.732092
R8556 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t1 0.7285
R8557 SARlogic_0.dffrs_13.nand3_1.C.n2 SARlogic_0.dffrs_13.nand3_1.C.t0 0.7285
R8558 SARlogic_0.dffrs_13.nand3_1.C.n1 SARlogic_0.dffrs_13.nand3_1.C 0.0455
R8559 a_n9861_28819.n0 a_n9861_28819.t5 34.1797
R8560 a_n9861_28819.n0 a_n9861_28819.t4 19.5798
R8561 a_n9861_28819.n1 a_n9861_28819.t1 18.7717
R8562 a_n9861_28819.n1 a_n9861_28819.t2 9.2885
R8563 a_n9861_28819.n2 a_n9861_28819.n0 4.93379
R8564 a_n9861_28819.n3 a_n9861_28819.t3 4.23346
R8565 a_n9861_28819.t0 a_n9861_28819.n3 3.85546
R8566 a_n9861_28819.n2 a_n9861_28819.n1 0.4055
R8567 a_n9861_28819.n3 a_n9861_28819.n2 0.352625
R8568 a_37499_28820.n0 a_37499_28820.t5 34.1797
R8569 a_37499_28820.n0 a_37499_28820.t4 19.5798
R8570 a_37499_28820.n1 a_37499_28820.t1 18.7717
R8571 a_37499_28820.n1 a_37499_28820.t2 9.2885
R8572 a_37499_28820.n2 a_37499_28820.n0 4.93379
R8573 a_37499_28820.t0 a_37499_28820.n3 4.23346
R8574 a_37499_28820.n3 a_37499_28820.t3 3.85546
R8575 a_37499_28820.n2 a_37499_28820.n1 0.4055
R8576 a_37499_28820.n3 a_37499_28820.n2 0.352625
R8577 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t4 40.6313
R8578 SARlogic_0.dffrs_4.nand3_1.C.n0 SARlogic_0.dffrs_4.nand3_1.C.t5 27.3166
R8579 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n1 14.2854
R8580 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.t2 10.0473
R8581 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.t1 6.51042
R8582 SARlogic_0.dffrs_4.nand3_1.C.n3 SARlogic_0.dffrs_4.nand3_1.C.n2 6.04952
R8583 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C.n0 5.13907
R8584 SARlogic_0.dffrs_4.nand3_0.Z SARlogic_0.dffrs_4.nand3_1.C.n4 4.72925
R8585 SARlogic_0.dffrs_4.nand3_1.C.n4 SARlogic_0.dffrs_4.nand3_1.C.n3 0.732092
R8586 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t0 0.7285
R8587 SARlogic_0.dffrs_4.nand3_1.C.n2 SARlogic_0.dffrs_4.nand3_1.C.t3 0.7285
R8588 SARlogic_0.dffrs_4.nand3_1.C.n1 SARlogic_0.dffrs_4.nand3_1.C 0.0455
R8589 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t5 41.0041
R8590 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t6 40.6313
R8591 SARlogic_0.dffrs_2.Q.n1 SARlogic_0.dffrs_2.Q.t4 27.3166
R8592 SARlogic_0.dffrs_2.Q.n0 SARlogic_0.dffrs_2.Q.t7 26.9438
R8593 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_3.d 17.5382
R8594 SARlogic_0.dffrs_2.Q.n3 SARlogic_0.dffrs_2.Q.n2 14.0582
R8595 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.t2 10.0473
R8596 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.t1 6.51042
R8597 SARlogic_0.dffrs_2.Q.n5 SARlogic_0.dffrs_2.Q.n4 6.04952
R8598 SARlogic_0.dffrs_3.nand3_8.A SARlogic_0.dffrs_2.Q.n0 5.7755
R8599 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.Q.n1 5.13907
R8600 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n6 4.72925
R8601 SARlogic_0.dffrs_3.d SARlogic_0.dffrs_3.nand3_8.A 0.784786
R8602 SARlogic_0.dffrs_2.Q.n6 SARlogic_0.dffrs_2.Q.n5 0.732092
R8603 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t3 0.7285
R8604 SARlogic_0.dffrs_2.Q.n4 SARlogic_0.dffrs_2.Q.t0 0.7285
R8605 SARlogic_0.dffrs_2.nand3_2.Z SARlogic_0.dffrs_2.Q.n3 0.166901
R8606 SARlogic_0.dffrs_2.Q.n2 SARlogic_0.dffrs_2.nand3_7.C 0.0455
R8607 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t6 40.6313
R8608 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.t5 34.1066
R8609 adc_PISO_0.dffrs_2.Q.n3 adc_PISO_0.dffrs_2.Q.t7 27.3166
R8610 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t8 19.673
R8611 adc_PISO_0.dffrs_2.Q.n0 adc_PISO_0.dffrs_2.Q.t4 19.4007
R8612 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n3 14.6967
R8613 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.t0 10.0473
R8614 adc_PISO_0.dffrs_2.Q.n7 adc_PISO_0.dffrs_2.Q.n6 9.39565
R8615 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.dffrs_2.Q.n1 6.70486
R8616 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.t1 6.51042
R8617 adc_PISO_0.dffrs_2.Q.n5 adc_PISO_0.dffrs_2.Q.n4 6.04952
R8618 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n2 5.81514
R8619 adc_PISO_0.dffrs_2.Q.n6 adc_PISO_0.dffrs_2.Q.n5 0.732092
R8620 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t2 0.7285
R8621 adc_PISO_0.dffrs_2.Q.n4 adc_PISO_0.dffrs_2.Q.t3 0.7285
R8622 adc_PISO_0.dffrs_2.Q adc_PISO_0.dffrs_2.Q.n7 0.458082
R8623 adc_PISO_0.dffrs_2.Q.n1 adc_PISO_0.dffrs_2.Q.n0 0.252687
R8624 adc_PISO_0.dffrs_2.Q.n2 adc_PISO_0.2inmux_4.Bit 0.0519286
R8625 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t4 40.6313
R8626 SARlogic_0.dffrs_1.nand3_1.C.n0 SARlogic_0.dffrs_1.nand3_1.C.t5 27.3166
R8627 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n1 14.2854
R8628 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.t0 10.0473
R8629 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.t1 6.51042
R8630 SARlogic_0.dffrs_1.nand3_1.C.n3 SARlogic_0.dffrs_1.nand3_1.C.n2 6.04952
R8631 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C.n0 5.13907
R8632 SARlogic_0.dffrs_1.nand3_0.Z SARlogic_0.dffrs_1.nand3_1.C.n4 4.72925
R8633 SARlogic_0.dffrs_1.nand3_1.C.n4 SARlogic_0.dffrs_1.nand3_1.C.n3 0.732092
R8634 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t2 0.7285
R8635 SARlogic_0.dffrs_1.nand3_1.C.n2 SARlogic_0.dffrs_1.nand3_1.C.t3 0.7285
R8636 SARlogic_0.dffrs_1.nand3_1.C.n1 SARlogic_0.dffrs_1.nand3_1.C 0.0455
R8637 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t3 41.0041
R8638 adc_PISO_0.2inmux_4.OUT.n0 adc_PISO_0.2inmux_4.OUT.t2 26.9438
R8639 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t0 9.6935
R8640 adc_PISO_0.dffrs_3.d adc_PISO_0.2inmux_4.OUT.n0 6.55979
R8641 adc_PISO_0.2inmux_4.OUT adc_PISO_0.dffrs_3.d 4.883
R8642 adc_PISO_0.2inmux_4.OUT.n1 adc_PISO_0.2inmux_4.OUT.t1 4.35383
R8643 adc_PISO_0.2inmux_4.OUT adc_PISO_0.2inmux_4.OUT.n1 0.350857
R8644 a_14313_31423.n1 a_14313_31423.t4 41.0041
R8645 a_14313_31423.n0 a_14313_31423.t6 40.8177
R8646 a_14313_31423.n2 a_14313_31423.t5 40.6313
R8647 a_14313_31423.n2 a_14313_31423.t8 27.3166
R8648 a_14313_31423.n0 a_14313_31423.t9 27.1302
R8649 a_14313_31423.n1 a_14313_31423.t7 26.9438
R8650 a_14313_31423.n3 a_14313_31423.n1 15.6312
R8651 a_14313_31423.n3 a_14313_31423.n2 15.046
R8652 a_14313_31423.n5 a_14313_31423.t1 10.0473
R8653 a_14313_31423.n6 a_14313_31423.t2 6.51042
R8654 a_14313_31423.n7 a_14313_31423.n6 6.04952
R8655 a_14313_31423.n4 a_14313_31423.n0 5.64619
R8656 a_14313_31423.n5 a_14313_31423.n4 5.17851
R8657 a_14313_31423.n4 a_14313_31423.n3 4.5005
R8658 a_14313_31423.n6 a_14313_31423.n5 0.732092
R8659 a_14313_31423.t0 a_14313_31423.n7 0.7285
R8660 a_14313_31423.n7 a_14313_31423.t3 0.7285
R8661 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t4 41.0041
R8662 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t7 40.6313
R8663 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t6 40.6313
R8664 SARlogic_0.dffrs_2.Qb SARlogic_0.dffrs_9.setb 28.021
R8665 SARlogic_0.dffrs_2.Qb.n4 SARlogic_0.dffrs_2.Qb.t9 27.3166
R8666 SARlogic_0.dffrs_2.Qb.n2 SARlogic_0.dffrs_2.Qb.t8 27.3166
R8667 SARlogic_0.dffrs_2.Qb.n0 SARlogic_0.dffrs_2.Qb.t5 26.9438
R8668 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.t0 10.0473
R8669 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb.n1 9.84255
R8670 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n3 9.22229
R8671 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.t1 6.51042
R8672 SARlogic_0.dffrs_2.Qb.n8 SARlogic_0.dffrs_2.Qb.n7 6.04952
R8673 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.Qb.n0 5.7305
R8674 SARlogic_0.dffrs_2.Qb.n5 SARlogic_0.dffrs_2.Qb.n4 5.14711
R8675 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_2.Qb.n2 5.13907
R8676 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n6 4.94976
R8677 SARlogic_0.dffrs_2.nand3_7.Z SARlogic_0.dffrs_2.Qb.n9 4.72925
R8678 SARlogic_0.dffrs_9.setb SARlogic_0.dffrs_9.nand3_0.C 0.784786
R8679 SARlogic_0.dffrs_2.Qb.n9 SARlogic_0.dffrs_2.Qb.n8 0.732092
R8680 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t2 0.7285
R8681 SARlogic_0.dffrs_2.Qb.n7 SARlogic_0.dffrs_2.Qb.t3 0.7285
R8682 SARlogic_0.dffrs_2.Qb.n6 SARlogic_0.dffrs_2.Qb 0.175225
R8683 SARlogic_0.dffrs_2.Qb.n1 SARlogic_0.dffrs_2.nand3_2.A 0.0455
R8684 SARlogic_0.dffrs_2.Qb.n3 SARlogic_0.dffrs_9.nand3_2.C 0.0455
R8685 SARlogic_0.dffrs_9.nand3_0.C SARlogic_0.dffrs_2.Qb.n5 0.0374643
.ends

