* NGSPICE file created from v2comp_SAR_final.ext - technology: (null)

.subckt comp_SAR_final Vdd Vss Clk Vin1 Vin2 Comp_out Reset SAR_in Clk_piso Load Piso_out
X0 a_n10869_517.t13 Clk.t0 Vdd.t31 Vdd.t30 pfet_03v3
**devattr s=14080,496 d=14080,496
X1 a_n9463_n751.t6 a_n10009_517.t9 a_n9733_n3007 Vss.t18 nfet_03v3
**devattr s=20800,504 d=20800,504
X2 a_n9429_n3007.t12 Vin1.t0 a_n10869_517.t9 Vss.t35 nfet_03v3
**devattr s=15600,404 d=15600,404
X3 Vdd.t7 a_n10831_3320 Comp_out.t3 Vdd.t6 pfet_03v3
**devattr s=18700,450 d=18700,450
X4 a_n10869_517.t3 a_n9463_n751.t9 a_n10009_517.t1 Vss.t31 nfet_03v3
**devattr s=20800,504 d=20800,504
X5 a_n9429_n3007.t18 Vin2.t0 a_n9733_n3007 Vss.t32 nfet_03v3
**devattr s=15600,404 d=15600,404
X6 a_n9733_n3007 Vin2.t1 a_n9429_n3007.t16 Vss.t24 nfet_03v3
**devattr s=15600,404 d=15600,404
X7 a_n9733_n3007 a_n9933_n3099 a_n10021_n3007 Vss.t20 nfet_03v3
**devattr s=26400,776 d=15600,404
X8 Vdd.t37 a_n10009_517.t10 a_n9463_n751.t3 Vdd.t36 pfet_03v3
**devattr s=10400,304 d=10400,304
X9 a_n9429_n3007.t19 Vin2.t2 a_n9733_n3007 Vss.t37 nfet_03v3
**devattr s=15600,404 d=15600,404
X10 a_n8351_n659 a_n8551_n751 a_n10009_517.t6 Vss.t40 nfet_03v3
**devattr s=20800,504 d=35200,976
X11 a_n9429_n3007.t17 Vin2.t3 a_n9733_n3007 Vss.t35 nfet_03v3
**devattr s=15600,404 d=15600,404
X12 a_n10211_3600 a_n8431_3575 Vdd.t17 Vdd.t16 pfet_03v3
**devattr s=17600,576 d=17600,576
X13 a_n10211_3600 a_n9321_1714 Vss.t22 Vss.t21 nfet_03v3
**devattr s=17600,576 d=17600,576
X14 a_n9733_n3007 a_n10009_517.t11 a_n9463_n751.t5 Vss.t17 nfet_03v3
**devattr s=20800,504 d=20800,504
X15 Comp_out.t7 a_n10831_3320 Vss.t7 Vss.t6 nfet_03v3
**devattr s=17000,540 d=9350,280
X16 a_n9321_1714 a_n10009_517.t12 Vss.t16 Vss.t15 nfet_03v3
**devattr s=35200,976 d=35200,976
X17 a_n10009_517.t3 a_n9463_n751.t10 Vdd.t19 Vdd.t18 pfet_03v3
**devattr s=10400,304 d=10400,304
X18 Vdd.t23 a_n9463_n751.t11 a_n10009_517.t4 Vdd.t22 pfet_03v3
**devattr s=10400,304 d=10400,304
X19 a_n10869_517.t5 Vin1.t1 a_n9429_n3007.t11 Vss.t24 nfet_03v3
**devattr s=15600,404 d=15600,404
X20 a_n10009_517.t2 a_n9463_n751.t12 Vdd.t15 Vdd.t14 pfet_03v3
**devattr s=10400,304 d=10400,304
X21 Vdd.t29 Clk.t1 a_n9733_n3007 Vdd.t28 pfet_03v3
**devattr s=14080,496 d=14080,496
X22 a_n6389_n2044 a_n6589_n2136 a_n9733_n3007 Vss.t19 nfet_03v3
**devattr s=15600,404 d=26400,776
X23 a_n10831_3320 a_n10211_3600 Vss.t11 Vss.t10 nfet_03v3
**devattr s=9350,280 d=17000,540
X24 a_n10869_517.t1 Vin1.t2 a_n9429_n3007.t10 Vss.t9 nfet_03v3
**devattr s=15600,404 d=15600,404
X25 a_n9429_n3007.t9 Vin1.t3 a_n10869_517.t11 Vss.t37 nfet_03v3
**devattr s=15600,404 d=15600,404
X26 Vdd.t27 Clk.t2 a_n9463_n751.t7 Vdd.t26 pfet_03v3
**devattr s=14080,496 d=14080,496
X27 Vss.t30 a_n9463_n751.t13 a_n7971_2755 Vss.t29 nfet_03v3
**devattr s=35200,976 d=35200,976
X28 Vdd.t43 a_n9629_405 a_n9717_497 Vdd.t42 pfet_03v3
**devattr s=17600,576 d=10400,304
X29 Comp_out.t2 a_n10831_3320 Vdd.t5 Vdd.t4 pfet_03v3
**devattr s=34000,880 d=18700,450
X30 Comp_out.t6 a_n10831_3320 Vss.t5 Vss.t4 nfet_03v3
**devattr s=9350,280 d=9350,280
X31 Vdd.t13 a_n9463_n751.t14 a_n10009_517.t0 Vdd.t12 pfet_03v3
**devattr s=10400,304 d=10400,304
X32 a_n10009_517.t7 a_n9463_n751.t15 a_n10869_517.t14 Vss.t28 nfet_03v3
**devattr s=20800,504 d=20800,504
X33 a_n9733_n3007 a_n10009_517.t13 a_n9463_n751.t4 Vss.t14 nfet_03v3
**devattr s=20800,504 d=20800,504
X34 a_n6389_n3007 a_n6589_n3099 a_n10869_517.t2 Vss.t19 nfet_03v3
**devattr s=15600,404 d=26400,776
X35 a_n10831_3320 a_n10211_3600 Vdd.t11 Vdd.t10 pfet_03v3
**devattr s=18700,450 d=34000,880
X36 a_n10009_517.t8 a_n9463_n751.t16 a_n10869_517.t16 Vss.t27 nfet_03v3
**devattr s=20800,504 d=20800,504
X37 a_n9429_n3007.t21 Vin2.t4 a_n9733_n3007 Vss.t34 nfet_03v3
**devattr s=15600,404 d=15600,404
X38 a_n9733_n3007 Vin2.t5 a_n9429_n3007.t20 Vss.t23 nfet_03v3
**devattr s=15600,404 d=15600,404
X39 a_n9733_n3007 Vin2.t6 a_n9429_n3007.t15 Vss.t36 nfet_03v3
**devattr s=15600,404 d=15600,404
X40 a_n9733_n3007 Vin2.t7 a_n9429_n3007.t2 Vss.t9 nfet_03v3
**devattr s=15600,404 d=15600,404
X41 Vss.t26 a_n8385_n3885 a_n8473_n3793 Vss.t25 nfet_03v3
**devattr s=14080,496 d=8320,264
X42 Comp_out.t1 a_n10831_3320 Vdd.t3 Vdd.t2 pfet_03v3
**devattr s=18700,450 d=18700,450
X43 a_n9463_n751.t2 a_n10009_517.t14 Vdd.t39 Vdd.t38 pfet_03v3
**devattr s=10400,304 d=10400,304
X44 a_n9429_n3007.t8 Vin1.t4 a_n10869_517.t7 Vss.t12 nfet_03v3
**devattr s=15600,404 d=15600,404
X45 a_n10869_517.t0 Vin1.t5 a_n9429_n3007.t7 Vss.t8 nfet_03v3
**devattr s=15600,404 d=15600,404
X46 a_n10009_517.t5 Clk.t3 Vdd.t25 Vdd.t24 pfet_03v3
**devattr s=14080,496 d=14080,496
X47 a_n9321_1714 a_n10009_517.t15 Vdd.t33 Vdd.t32 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X48 a_n9463_n751.t1 a_n10009_517.t16 Vdd.t41 Vdd.t40 pfet_03v3
**devattr s=10400,304 d=10400,304
X49 a_n6693_497 a_n6893_405 Vdd.t21 Vdd.t20 pfet_03v3
**devattr s=10400,304 d=17600,576
X50 a_n9463_n751.t8 a_n7971_n751 a_n8059_n659 Vss.t41 nfet_03v3
**devattr s=35200,976 d=20800,504
X51 a_n9429_n3007.t6 Vin1.t6 a_n10869_517.t8 Vss.t34 nfet_03v3
**devattr s=15600,404 d=15600,404
X52 Vss.t3 a_n10831_3320 Comp_out.t5 Vss.t2 nfet_03v3
**devattr s=9350,280 d=9350,280
X53 a_n10869_517.t4 Vin1.t7 a_n9429_n3007.t5 Vss.t23 nfet_03v3
**devattr s=15600,404 d=15600,404
X54 Vdd.t35 a_n10009_517.t17 a_n9463_n751.t0 Vdd.t34 pfet_03v3
**devattr s=10400,304 d=10400,304
X55 a_n10869_517.t15 a_n9767_n751 a_n9855_n659 Vss.t42 nfet_03v3
**devattr s=35200,976 d=20800,504
X56 a_n9429_n3007.t1 Vin2.t8 a_n9733_n3007 Vss.t12 nfet_03v3
**devattr s=15600,404 d=15600,404
X57 a_n10869_517.t10 Vin1.t8 a_n9429_n3007.t4 Vss.t36 nfet_03v3
**devattr s=15600,404 d=15600,404
X58 a_n9429_n3007.t14 Clk.t4 Vss.t39 Vss.t38 nfet_03v3
**devattr s=8320,264 d=8320,264
X59 Vdd.t45 a_n9463_n751.t17 a_n7971_2755 Vdd.t44 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X60 a_n9429_n3007.t3 Vin1.t9 a_n10869_517.t6 Vss.t32 nfet_03v3
**devattr s=15600,404 d=15600,404
X61 a_n9733_n3007 Vin2.t9 a_n9429_n3007.t0 Vss.t8 nfet_03v3
**devattr s=15600,404 d=15600,404
X62 Vss.t1 a_n10831_3320 Comp_out.t4 Vss.t0 nfet_03v3
**devattr s=9350,280 d=9350,280
X63 Vdd.t9 a_n10211_3600 a_n8431_3575 Vdd.t8 pfet_03v3
**devattr s=17600,576 d=17600,576
X64 a_n6555_n659 a_n6755_n751 a_n9733_n3007 Vss.t13 nfet_03v3
**devattr s=20800,504 d=35200,976
X65 a_n10869_517.t12 a_n9933_n2136 a_n10021_n2044 Vss.t20 nfet_03v3
**devattr s=26400,776 d=15600,404
X66 Vss.t44 a_n7971_2755 a_n8431_3575 Vss.t43 nfet_03v3
**devattr s=17600,576 d=17600,576
X67 Vdd.t1 a_n10831_3320 Comp_out.t0 Vdd.t0 pfet_03v3
**devattr s=18700,450 d=18700,450
X68 a_n7937_n3793 a_n8017_n3885 a_n9429_n3007.t13 Vss.t33 nfet_03v3
**devattr s=8320,264 d=14080,496
R0 Clk.n4 Clk.t0 21.1483
R1 Clk.n3 Clk.t3 21.1483
R2 Clk.n2 Clk.t2 21.1483
R3 Clk.n1 Clk.t1 21.1483
R4 Clk.n0 Clk.t4 20.5929
R5 Clk.n1 Clk.n0 19.1491
R6 Clk.n5 Clk.n4 15.5861
R7 Clk Clk.n5 7.2261
R8 Clk.n3 Clk.n2 4.47208
R9 Clk.n5 Clk.n0 3.56405
R10 Clk.n2 Clk.n1 1.01892
R11 Clk.n4 Clk.n3 1.01892
R12 Vdd.n11 Vdd.t32 869.717
R13 Vdd.n1 Vdd.t44 869.717
R14 Vdd.t22 Vdd.t20 490.324
R15 Vdd.t14 Vdd.t22 490.324
R16 Vdd.t36 Vdd.t14 490.324
R17 Vdd.t40 Vdd.t36 490.324
R18 Vdd.t12 Vdd.t40 490.324
R19 Vdd.t18 Vdd.t12 490.324
R20 Vdd.t34 Vdd.t18 490.324
R21 Vdd.t38 Vdd.t34 490.324
R22 Vdd.t42 Vdd.t38 490.324
R23 Vdd.t20 Vdd.n46 467.743
R24 Vdd.n48 Vdd.t42 467.743
R25 Vdd.n49 Vdd.t24 398.652
R26 Vdd.n31 Vdd.t26 398.652
R27 Vdd.t24 Vdd.n48 389.878
R28 Vdd.n46 Vdd.t26 389.878
R29 Vdd.t8 Vdd.n5 372.543
R30 Vdd.n8 Vdd.t16 372.543
R31 Vdd.n7 Vdd.t8 370.969
R32 Vdd.t16 Vdd.n7 370.969
R33 Vdd.n26 Vdd.n24 287.351
R34 Vdd.n27 Vdd.n25 287.351
R35 Vdd.t2 Vdd.t0 265.625
R36 Vdd.n17 Vdd.t10 242.189
R37 Vdd.t6 Vdd.n19 195.312
R38 Vdd.n53 Vdd.t30 190.464
R39 Vdd.n29 Vdd.t28 190.464
R40 Vdd.n20 Vdd.t6 179.689
R41 Vdd.t10 Vdd.n16 145.523
R42 Vdd.n20 Vdd.t2 85.938
R43 Vdd.n19 Vdd.t4 70.313
R44 Vdd.n5 Vdd.n3 58.9755
R45 Vdd.n8 Vdd.n3 58.9755
R46 Vdd.n8 Vdd.n4 58.9755
R47 Vdd.n5 Vdd.n4 58.9755
R48 Vdd.n49 Vdd.n24 54.0755
R49 Vdd.n31 Vdd.n26 54.0755
R50 Vdd.n31 Vdd.n27 54.0755
R51 Vdd.n49 Vdd.n25 54.0755
R52 Vdd.n53 Vdd.n52 29.3622
R53 Vdd.n30 Vdd.n29 29.3622
R54 Vdd.t0 Vdd.n17 23.438
R55 Vdd.n45 Vdd.n26 20.1255
R56 Vdd.n45 Vdd.n27 20.1255
R57 Vdd.n47 Vdd.n24 20.1255
R58 Vdd.n47 Vdd.n25 20.1255
R59 Vdd.n54 Vdd.n53 19.9167
R60 Vdd.n29 Vdd.n28 19.9167
R61 Vdd.n6 Vdd.n3 18.7255
R62 Vdd.n6 Vdd.n4 18.7255
R63 Vdd.n56 Vdd.n55 15.0415
R64 Vdd.n60 Vdd.n0 13.4987
R65 Vdd.n17 Vdd.n12 12.6005
R66 Vdd.n21 Vdd.n20 12.6005
R67 Vdd.n19 Vdd.n18 12.6005
R68 Vdd.n43 Vdd.n42 12.136
R69 Vdd.n41 Vdd.n40 12.136
R70 Vdd.n39 Vdd.n38 12.136
R71 Vdd.n37 Vdd.n36 12.136
R72 Vdd.n35 Vdd.n34 12.136
R73 Vdd.n47 Vdd.n23 11.111
R74 Vdd.n45 Vdd.n44 11.111
R75 Vdd.n28 Vdd.n0 9.86945
R76 Vdd.n33 Vdd.n32 9.536
R77 Vdd.n51 Vdd.n50 9.536
R78 Vdd.n55 Vdd.n54 9.536
R79 Vdd.n32 Vdd.t27 7.4755
R80 Vdd.n50 Vdd.t25 7.4755
R81 Vdd.n54 Vdd.t31 7.4755
R82 Vdd.n28 Vdd.t29 7.4755
R83 Vdd Vdd.n60 5.27311
R84 Vdd.n9 Vdd.t17 4.4205
R85 Vdd.n2 Vdd.t9 4.4205
R86 Vdd.n18 Vdd.t5 3.38176
R87 Vdd.n32 Vdd.n31 2.1905
R88 Vdd.n50 Vdd.n49 2.1905
R89 Vdd.n14 Vdd.n13 2.16583
R90 Vdd.n16 Vdd.n15 2.16583
R91 Vdd.n11 Vdd.t33 2.00711
R92 Vdd.n1 Vdd.t45 1.99236
R93 Vdd.n57 Vdd.n11 1.83762
R94 Vdd.n59 Vdd.n1 1.83762
R95 Vdd.n42 Vdd.t21 1.8205
R96 Vdd.n42 Vdd.t23 1.8205
R97 Vdd.n40 Vdd.t15 1.8205
R98 Vdd.n40 Vdd.t37 1.8205
R99 Vdd.n38 Vdd.t41 1.8205
R100 Vdd.n38 Vdd.t13 1.8205
R101 Vdd.n36 Vdd.t19 1.8205
R102 Vdd.n36 Vdd.t35 1.8205
R103 Vdd.n34 Vdd.t39 1.8205
R104 Vdd.n34 Vdd.t43 1.8205
R105 Vdd.n7 Vdd.n6 1.5755
R106 Vdd.n9 Vdd.n8 1.5755
R107 Vdd.n5 Vdd.n2 1.5755
R108 Vdd.n46 Vdd.n45 1.5755
R109 Vdd.n48 Vdd.n47 1.5755
R110 Vdd.n13 Vdd.t3 1.13285
R111 Vdd.n13 Vdd.t7 1.13285
R112 Vdd.n15 Vdd.t11 1.13285
R113 Vdd.n15 Vdd.t1 1.13285
R114 Vdd.n58 Vdd.n10 1.058
R115 Vdd.n10 Vdd.n2 1.01373
R116 Vdd.n10 Vdd.n9 0.979984
R117 Vdd.n56 Vdd.n22 0.750875
R118 Vdd.n37 Vdd.n35 0.667
R119 Vdd.n43 Vdd.n41 0.662
R120 Vdd.n39 Vdd.n37 0.643429
R121 Vdd.n41 Vdd.n39 0.638429
R122 Vdd.n52 Vdd.n51 0.58325
R123 Vdd.n33 Vdd.n30 0.58325
R124 Vdd.n35 Vdd.n23 0.47525
R125 Vdd.n44 Vdd.n43 0.47525
R126 Vdd.n55 Vdd.n52 0.34025
R127 Vdd.n51 Vdd.n23 0.34025
R128 Vdd.n44 Vdd.n33 0.34025
R129 Vdd.n60 Vdd.n59 0.313132
R130 Vdd.n59 Vdd.n58 0.289447
R131 Vdd.n58 Vdd.n57 0.279974
R132 Vdd.n57 Vdd.n56 0.256289
R133 Vdd.n18 Vdd.n14 0.1355
R134 Vdd.n22 Vdd.n12 0.103357
R135 Vdd.n22 Vdd.n21 0.0519286
R136 Vdd.n16 Vdd.n12 0.0455
R137 Vdd.n21 Vdd.n14 0.0197857
R138 Vdd.n30 Vdd.n0 0.0068
R139 a_n10869_517.n6 a_n10869_517.t13 19.5626
R140 a_n10869_517.n5 a_n10869_517.n3 11.9065
R141 a_n10869_517.n5 a_n10869_517.n4 11.2495
R142 a_n10869_517.n1 a_n10869_517.n0 11.243
R143 a_n10869_517.n12 a_n10869_517.n2 8.80104
R144 a_n10869_517.n16 a_n10869_517.n15 6.60725
R145 a_n10869_517.n11 a_n10869_517.n9 6.52262
R146 a_n10869_517.n15 a_n10869_517.n14 6.386
R147 a_n10869_517.n8 a_n10869_517.n6 5.44213
R148 a_n10869_517.n11 a_n10869_517.n10 4.36738
R149 a_n10869_517.n14 a_n10869_517.n13 4.36738
R150 a_n10869_517.n8 a_n10869_517.n7 4.3505
R151 a_n10869_517.n9 a_n10869_517.n8 2.2505
R152 a_n10869_517.n12 a_n10869_517.n11 2.14009
R153 a_n10869_517.n15 a_n10869_517.n1 1.50001
R154 a_n10869_517.n9 a_n10869_517.n1 1.49326
R155 a_n10869_517.n0 a_n10869_517.t6 1.0925
R156 a_n10869_517.n0 a_n10869_517.t1 1.0925
R157 a_n10869_517.n7 a_n10869_517.t7 1.0925
R158 a_n10869_517.n7 a_n10869_517.t12 1.0925
R159 a_n10869_517.n10 a_n10869_517.t8 1.0925
R160 a_n10869_517.n10 a_n10869_517.t5 1.0925
R161 a_n10869_517.n2 a_n10869_517.t2 1.0925
R162 a_n10869_517.n2 a_n10869_517.t10 1.0925
R163 a_n10869_517.n13 a_n10869_517.t11 1.0925
R164 a_n10869_517.n13 a_n10869_517.t4 1.0925
R165 a_n10869_517.n16 a_n10869_517.t9 1.0925
R166 a_n10869_517.t0 a_n10869_517.n16 1.0925
R167 a_n10869_517.n4 a_n10869_517.t16 0.8195
R168 a_n10869_517.n4 a_n10869_517.t15 0.8195
R169 a_n10869_517.n3 a_n10869_517.t14 0.8195
R170 a_n10869_517.n3 a_n10869_517.t3 0.8195
R171 a_n10869_517.n14 a_n10869_517.n12 0.314375
R172 a_n10869_517.n6 a_n10869_517.n5 0.16025
R173 a_n10009_517.n5 a_n10009_517.t15 49.7997
R174 a_n10009_517.n5 a_n10009_517.t12 31.5502
R175 a_n10009_517.t16 a_n10009_517.t10 19.735
R176 a_n10009_517.n12 a_n10009_517.n0 18.0852
R177 a_n10009_517.n6 a_n10009_517.t5 16.9998
R178 a_n10009_517.n3 a_n10009_517.t16 14.5537
R179 a_n10009_517.n3 a_n10009_517.n2 14.2885
R180 a_n10009_517.n1 a_n10009_517.t13 13.6729
R181 a_n10009_517.n2 a_n10009_517.t11 13.3844
R182 a_n10009_517.n1 a_n10009_517.t9 13.3445
R183 a_n10009_517.n6 a_n10009_517.n5 13.282
R184 a_n10009_517.n9 a_n10009_517.n8 11.24
R185 a_n10009_517.n13 a_n10009_517.n12 7.16477
R186 a_n10009_517.n10 a_n10009_517.n4 6.75194
R187 a_n10009_517.n7 a_n10009_517.t17 5.04666
R188 a_n10009_517.n7 a_n10009_517.t14 4.84137
R189 a_n10009_517.n10 a_n10009_517.n9 2.836
R190 a_n10009_517.n9 a_n10009_517.n7 2.75432
R191 a_n10009_517.n0 a_n10009_517.t4 1.8205
R192 a_n10009_517.n0 a_n10009_517.t2 1.8205
R193 a_n10009_517.t0 a_n10009_517.n13 1.8205
R194 a_n10009_517.n13 a_n10009_517.t3 1.8205
R195 a_n10009_517.n8 a_n10009_517.t1 0.8195
R196 a_n10009_517.n8 a_n10009_517.t8 0.8195
R197 a_n10009_517.n4 a_n10009_517.t6 0.8195
R198 a_n10009_517.n4 a_n10009_517.t7 0.8195
R199 a_n10009_517.n9 a_n10009_517.n6 0.733357
R200 a_n10009_517.n11 a_n10009_517.n3 0.440894
R201 a_n10009_517.n12 a_n10009_517.n11 0.426875
R202 a_n10009_517.n2 a_n10009_517.n1 0.289009
R203 a_n10009_517.n11 a_n10009_517.n10 0.0607115
R204 a_n9463_n751.n0 a_n9463_n751.t17 49.7997
R205 a_n9463_n751.n0 a_n9463_n751.t13 31.5502
R206 a_n9463_n751.t14 a_n9463_n751.t10 19.735
R207 a_n9463_n751.n11 a_n9463_n751.t14 18.9075
R208 a_n9463_n751.n1 a_n9463_n751.t7 16.9998
R209 a_n9463_n751.n8 a_n9463_n751.t16 13.6729
R210 a_n9463_n751.n9 a_n9463_n751.t15 13.3844
R211 a_n9463_n751.n8 a_n9463_n751.t9 13.3445
R212 a_n9463_n751.n1 a_n9463_n751.n0 13.2778
R213 a_n9463_n751.n10 a_n9463_n751.n7 12.247
R214 a_n9463_n751.n4 a_n9463_n751.n3 11.2403
R215 a_n9463_n751.n10 a_n9463_n751.n9 9.4181
R216 a_n9463_n751.n13 a_n9463_n751.n12 7.4449
R217 a_n9463_n751.n6 a_n9463_n751.n5 6.75194
R218 a_n9463_n751.n2 a_n9463_n751.t12 5.04666
R219 a_n9463_n751.n12 a_n9463_n751.n11 4.94262
R220 a_n9463_n751.n2 a_n9463_n751.t11 4.84137
R221 a_n9463_n751.n6 a_n9463_n751.n4 2.836
R222 a_n9463_n751.n4 a_n9463_n751.n2 2.75432
R223 a_n9463_n751.n7 a_n9463_n751.t0 1.8205
R224 a_n9463_n751.n7 a_n9463_n751.t2 1.8205
R225 a_n9463_n751.t3 a_n9463_n751.n13 1.8205
R226 a_n9463_n751.n13 a_n9463_n751.t1 1.8205
R227 a_n9463_n751.n5 a_n9463_n751.t5 0.8195
R228 a_n9463_n751.n5 a_n9463_n751.t8 0.8195
R229 a_n9463_n751.n3 a_n9463_n751.t4 0.8195
R230 a_n9463_n751.n3 a_n9463_n751.t6 0.8195
R231 a_n9463_n751.n4 a_n9463_n751.n1 0.733357
R232 a_n9463_n751.n11 a_n9463_n751.n10 0.5315
R233 a_n9463_n751.n9 a_n9463_n751.n8 0.289009
R234 a_n9463_n751.n12 a_n9463_n751.n6 0.184462
R235 Vss.n63 Vss.n62 259245
R236 Vss.n40 Vss.n4 148254
R237 Vss.n61 Vss.n2 59530.8
R238 Vss.n60 Vss.n59 25794.4
R239 Vss.n60 Vss.n4 23334.9
R240 Vss.n62 Vss.n61 18659
R241 Vss.n59 Vss.t10 10202.1
R242 Vss.n59 Vss.n16 5567.73
R243 Vss.n62 Vss.n3 2358.54
R244 Vss.n47 Vss.t15 1596.98
R245 Vss.n63 Vss.t29 1596.98
R246 Vss.t6 Vss.n4 1095.73
R247 Vss.n61 Vss.n60 924.742
R248 Vss.n48 Vss.n47 478.125
R249 Vss.n28 Vss.n18 414.478
R250 Vss.n9 Vss.n2 325
R251 Vss.n16 Vss.n15 325
R252 Vss.n9 Vss.t43 293.137
R253 Vss.t43 Vss.n8 293.137
R254 Vss.n8 Vss.t21 293.137
R255 Vss.n15 Vss.t21 293.137
R256 Vss.n63 Vss.n2 248.53
R257 Vss.n47 Vss.n16 248.53
R258 Vss.n30 Vss.n19 205.139
R259 Vss.n42 Vss.n19 205.139
R260 Vss.n42 Vss.n20 205.139
R261 Vss.n30 Vss.n20 205.139
R262 Vss.n41 Vss.n40 193.476
R263 Vss.n31 Vss.n3 192.703
R264 Vss.t2 Vss.t4 191.642
R265 Vss.t10 Vss.n58 174.732
R266 Vss.n26 Vss.n24 166.989
R267 Vss.n38 Vss.n21 166.989
R268 Vss.t0 Vss.n56 140.913
R269 Vss.n57 Vss.t0 129.641
R270 Vss.n35 Vss.n23 118.222
R271 Vss.t13 Vss.t19 108.138
R272 Vss.t14 Vss.t36 108.138
R273 Vss.t18 Vss.t35 108.138
R274 Vss.t17 Vss.t8 108.138
R275 Vss.t28 Vss.t34 108.138
R276 Vss.t31 Vss.t24 108.138
R277 Vss.t27 Vss.t12 108.138
R278 Vss.t42 Vss.t20 108.138
R279 Vss.t10 Vss.n48 105.561
R280 Vss.t38 Vss.t23 99.0183
R281 Vss.t32 Vss.t38 99.0183
R282 Vss.n47 Vss.n46 98.7258
R283 Vss.n64 Vss.n63 98.7258
R284 Vss.t36 Vss.t13 89.8983
R285 Vss.t35 Vss.t14 89.8983
R286 Vss.t8 Vss.t18 89.8983
R287 Vss.t37 Vss.t17 89.8983
R288 Vss.t9 Vss.t28 89.8983
R289 Vss.t34 Vss.t31 89.8983
R290 Vss.t24 Vss.t27 89.8983
R291 Vss.t12 Vss.t42 89.8983
R292 Vss.t41 Vss.n32 80.7782
R293 Vss.n34 Vss.t40 80.7782
R294 Vss.n41 Vss.t20 80.7782
R295 Vss.n24 Vss.n21 80.5005
R296 Vss.t33 Vss.t41 69.0524
R297 Vss.t40 Vss.t25 69.0524
R298 Vss.t19 Vss.n31 65.5624
R299 Vss.n10 Vss.n5 65.5283
R300 Vss.n14 Vss.n5 65.5283
R301 Vss.n14 Vss.n6 65.5283
R302 Vss.n10 Vss.n6 65.5283
R303 Vss.t4 Vss.n57 62.0024
R304 Vss.n56 Vss.t6 50.7294
R305 Vss.n33 Vss.n19 30.5283
R306 Vss.n33 Vss.n20 30.5283
R307 Vss.n32 Vss.t37 27.3607
R308 Vss.n34 Vss.t9 27.3607
R309 Vss.t23 Vss.t33 20.8464
R310 Vss.t25 Vss.t32 20.8464
R311 Vss.n7 Vss.n5 20.8061
R312 Vss.n7 Vss.n6 20.8061
R313 Vss.n35 Vss.n21 18.8616
R314 Vss.n24 Vss.n23 18.8616
R315 Vss.n45 Vss.n44 18.2476
R316 Vss.n66 Vss.n65 16.9448
R317 Vss.n58 Vss.t2 16.9105
R318 Vss.n57 Vss.n52 14.6641
R319 Vss.n56 Vss.n55 14.1923
R320 Vss.n58 Vss.n51 11.9681
R321 Vss.n36 Vss.n22 11.0305
R322 Vss.n50 Vss.n48 10.5098
R323 Vss Vss.n66 9.06952
R324 Vss.n55 Vss.t7 8.70131
R325 Vss.n44 Vss.n43 7.7564
R326 Vss.n29 Vss.n0 7.59387
R327 Vss.n26 Vss.n25 6.65104
R328 Vss.n50 Vss.n49 6.5795
R329 Vss.n54 Vss.n53 6.5795
R330 Vss.n43 Vss.n42 6.33584
R331 Vss.n30 Vss.n29 6.32806
R332 Vss.n36 Vss.n35 6.23383
R333 Vss.n11 Vss.t44 4.7885
R334 Vss.n13 Vss.t22 4.7885
R335 Vss.n38 Vss.n37 3.8722
R336 Vss.n29 Vss.n28 3.52248
R337 Vss.n43 Vss.n18 3.51469
R338 Vss.n45 Vss.t16 2.9111
R339 Vss.n65 Vss.t30 2.9111
R340 Vss.n22 Vss.t39 2.048
R341 Vss.n22 Vss.t26 2.048
R342 Vss.n49 Vss.t11 2.03874
R343 Vss.n49 Vss.t3 2.03874
R344 Vss.n53 Vss.t5 2.03874
R345 Vss.n53 Vss.t1 2.03874
R346 Vss.n35 Vss.n34 1.73383
R347 Vss.n32 Vss.n23 1.73383
R348 Vss.n64 Vss.n1 1.70279
R349 Vss.n46 Vss.n1 1.62925
R350 Vss.n11 Vss.n10 1.3005
R351 Vss.n10 Vss.n9 1.3005
R352 Vss.n8 Vss.n7 1.3005
R353 Vss.n14 Vss.n13 1.3005
R354 Vss.n15 Vss.n14 1.3005
R355 Vss.n12 Vss.n1 1.29323
R356 Vss.n12 Vss.n11 1.00923
R357 Vss.n28 Vss.n27 0.999917
R358 Vss.n27 Vss.n26 0.999917
R359 Vss.n39 Vss.n18 0.999917
R360 Vss.n39 Vss.n38 0.999917
R361 Vss.n13 Vss.n12 0.984484
R362 Vss.n37 Vss.n17 0.949529
R363 Vss.n25 Vss.n17 0.907842
R364 Vss.n31 Vss.n30 0.867167
R365 Vss.t38 Vss.n33 0.867167
R366 Vss.n42 Vss.n41 0.867167
R367 Vss.n37 Vss.n36 0.824071
R368 Vss.n66 Vss.n0 0.211763
R369 Vss.n44 Vss.n17 0.163684
R370 Vss.n52 Vss.n51 0.154786
R371 Vss.n55 Vss.n54 0.1355
R372 Vss.n65 Vss.n64 0.128901
R373 Vss.n46 Vss.n45 0.127885
R374 Vss.n25 Vss.n0 0.112526
R375 Vss.n51 Vss.n50 0.0455
R376 Vss.n27 Vss.n3 0.0215413
R377 Vss.n40 Vss.n39 0.0215413
R378 Vss.n54 Vss.n52 0.0197857
R379 Vin1.n7 Vin1.n6 23.1032
R380 Vin1.n3 Vin1.n2 23.1032
R381 Vin1.n0 Vin1.t8 22.5295
R382 Vin1.n2 Vin1.t3 16.3641
R383 Vin1.n6 Vin1.t6 16.3626
R384 Vin1.n2 Vin1.t7 16.0225
R385 Vin1.n6 Vin1.t1 16.021
R386 Vin1.n8 Vin1.t4 11.5195
R387 Vin1.n5 Vin1.t2 11.5195
R388 Vin1.n4 Vin1.t9 11.5195
R389 Vin1.n1 Vin1.t5 11.5195
R390 Vin1.n0 Vin1.t0 11.5195
R391 Vin1 Vin1.n8 9.6279
R392 Vin1.n1 Vin1.n0 4.00673
R393 Vin1.n7 Vin1.n5 3.16619
R394 Vin1.n3 Vin1.n1 0.650658
R395 Vin1.n8 Vin1.n7 0.280193
R396 Vin1.n4 Vin1.n3 0.279681
R397 Vin1.n5 Vin1.n4 0.231705
R398 a_n9429_n3007.n13 a_n9429_n3007.n5 11.2899
R399 a_n9429_n3007.n14 a_n9429_n3007.n13 8.49339
R400 a_n9429_n3007.n17 a_n9429_n3007.n16 4.89725
R401 a_n9429_n3007.n10 a_n9429_n3007.n6 4.89725
R402 a_n9429_n3007.n15 a_n9429_n3007.n3 4.89725
R403 a_n9429_n3007.n9 a_n9429_n3007.n7 4.89725
R404 a_n9429_n3007.n2 a_n9429_n3007.n0 4.89725
R405 a_n9429_n3007.n9 a_n9429_n3007.n8 4.88712
R406 a_n9429_n3007.n2 a_n9429_n3007.n1 4.88712
R407 a_n9429_n3007.n18 a_n9429_n3007.n17 4.88712
R408 a_n9429_n3007.n12 a_n9429_n3007.n11 4.4
R409 a_n9429_n3007.n14 a_n9429_n3007.n4 4.35275
R410 a_n9429_n3007.n5 a_n9429_n3007.t13 2.048
R411 a_n9429_n3007.n5 a_n9429_n3007.t14 2.048
R412 a_n9429_n3007.n13 a_n9429_n3007.n12 1.95895
R413 a_n9429_n3007.n16 a_n9429_n3007.t7 1.0925
R414 a_n9429_n3007.n16 a_n9429_n3007.t19 1.0925
R415 a_n9429_n3007.n6 a_n9429_n3007.t16 1.0925
R416 a_n9429_n3007.n6 a_n9429_n3007.t8 1.0925
R417 a_n9429_n3007.n11 a_n9429_n3007.t11 1.0925
R418 a_n9429_n3007.n11 a_n9429_n3007.t1 1.0925
R419 a_n9429_n3007.n3 a_n9429_n3007.t15 1.0925
R420 a_n9429_n3007.n3 a_n9429_n3007.t12 1.0925
R421 a_n9429_n3007.n4 a_n9429_n3007.t4 1.0925
R422 a_n9429_n3007.n4 a_n9429_n3007.t17 1.0925
R423 a_n9429_n3007.n7 a_n9429_n3007.t10 1.0925
R424 a_n9429_n3007.n7 a_n9429_n3007.t21 1.0925
R425 a_n9429_n3007.n8 a_n9429_n3007.t2 1.0925
R426 a_n9429_n3007.n8 a_n9429_n3007.t6 1.0925
R427 a_n9429_n3007.n0 a_n9429_n3007.t20 1.0925
R428 a_n9429_n3007.n0 a_n9429_n3007.t3 1.0925
R429 a_n9429_n3007.n1 a_n9429_n3007.t5 1.0925
R430 a_n9429_n3007.n1 a_n9429_n3007.t18 1.0925
R431 a_n9429_n3007.t0 a_n9429_n3007.n18 1.0925
R432 a_n9429_n3007.n18 a_n9429_n3007.t9 1.0925
R433 a_n9429_n3007.n10 a_n9429_n3007.n9 0.849071
R434 a_n9429_n3007.n9 a_n9429_n3007.n2 0.849071
R435 a_n9429_n3007.n17 a_n9429_n3007.n2 0.849071
R436 a_n9429_n3007.n17 a_n9429_n3007.n15 0.849071
R437 a_n9429_n3007.n15 a_n9429_n3007.n14 0.534875
R438 a_n9429_n3007.n12 a_n9429_n3007.n10 0.487625
R439 Comp_out Comp_out.n8 18.1644
R440 Comp_out.n5 Comp_out.n4 6.5435
R441 Comp_out.n2 Comp_out.n1 6.5435
R442 Comp_out.n6 Comp_out.n3 2.17483
R443 Comp_out.n4 Comp_out.t5 2.03874
R444 Comp_out.n4 Comp_out.t6 2.03874
R445 Comp_out.n1 Comp_out.t4 2.03874
R446 Comp_out.n1 Comp_out.t7 2.03874
R447 Comp_out.n8 Comp_out.n0 2.00383
R448 Comp_out.n0 Comp_out.t3 1.13285
R449 Comp_out.n0 Comp_out.t2 1.13285
R450 Comp_out.n3 Comp_out.t0 1.13285
R451 Comp_out.n3 Comp_out.t1 1.13285
R452 Comp_out.n5 Comp_out.n2 0.5105
R453 Comp_out.n7 Comp_out.n6 0.5105
R454 Comp_out.n7 Comp_out.n2 0.2165
R455 Comp_out.n6 Comp_out.n5 0.2165
R456 Comp_out.n8 Comp_out.n7 0.1175
R457 Vin2.n7 Vin2.n6 23.1032
R458 Vin2.n3 Vin2.n2 23.1032
R459 Vin2.n0 Vin2.t6 22.8502
R460 Vin2.n2 Vin2.t5 16.3656
R461 Vin2.n6 Vin2.t1 16.3641
R462 Vin2.n2 Vin2.t2 16.021
R463 Vin2.n6 Vin2.t4 16.0195
R464 Vin2.n8 Vin2.t8 11.5195
R465 Vin2.n5 Vin2.t7 11.5195
R466 Vin2.n4 Vin2.t0 11.5195
R467 Vin2.n1 Vin2.t9 11.5195
R468 Vin2.n0 Vin2.t3 11.5195
R469 Vin2 Vin2.n8 9.62695
R470 Vin2.n7 Vin2.n5 2.53166
R471 Vin2.n1 Vin2.n0 2.48408
R472 Vin2.n3 Vin2.n1 1.40666
R473 Vin2.n8 Vin2.n7 0.647658
R474 Vin2.n4 Vin2.n3 0.647132
R475 Vin2.n5 Vin2.n4 0.234605
R476 SARlogic_0.reset Reset 0.18425
R477 SARlogic_0.comp_in SAR_in 0.1775
.ends

