magic
tech gf180mcuD
magscale 1 10
timestamp 1757859636
<< error_p >>
rect -354 433 -343 479
rect -150 433 -139 479
rect 54 433 65 479
rect 258 433 269 479
rect -354 -479 -343 -433
rect -150 -479 -139 -433
rect 54 -479 65 -433
rect 258 -479 269 -433
<< nwell >>
rect -606 -610 606 610
<< pmos >>
rect -356 -400 -256 400
rect -152 -400 -52 400
rect 52 -400 152 400
rect 256 -400 356 400
<< pdiff >>
rect -444 387 -356 400
rect -444 -387 -431 387
rect -385 -387 -356 387
rect -444 -400 -356 -387
rect -256 387 -152 400
rect -256 -387 -227 387
rect -181 -387 -152 387
rect -256 -400 -152 -387
rect -52 387 52 400
rect -52 -387 -23 387
rect 23 -387 52 387
rect -52 -400 52 -387
rect 152 387 256 400
rect 152 -387 181 387
rect 227 -387 256 387
rect 152 -400 256 -387
rect 356 387 444 400
rect 356 -387 385 387
rect 431 -387 444 387
rect 356 -400 444 -387
<< pdiffc >>
rect -431 -387 -385 387
rect -227 -387 -181 387
rect -23 -387 23 387
rect 181 -387 227 387
rect 385 -387 431 387
<< nsubdiff >>
rect -582 514 582 586
rect -582 470 -510 514
rect -582 -470 -569 470
rect -523 -470 -510 470
rect 510 470 582 514
rect -582 -514 -510 -470
rect 510 -470 523 470
rect 569 -470 582 470
rect 510 -514 582 -470
rect -582 -586 582 -514
<< nsubdiffcont >>
rect -569 -470 -523 470
rect 523 -470 569 470
<< polysilicon >>
rect -356 479 -256 492
rect -356 433 -343 479
rect -269 433 -256 479
rect -356 400 -256 433
rect -152 479 -52 492
rect -152 433 -139 479
rect -65 433 -52 479
rect -152 400 -52 433
rect 52 479 152 492
rect 52 433 65 479
rect 139 433 152 479
rect 52 400 152 433
rect 256 479 356 492
rect 256 433 269 479
rect 343 433 356 479
rect 256 400 356 433
rect -356 -433 -256 -400
rect -356 -479 -343 -433
rect -269 -479 -256 -433
rect -356 -492 -256 -479
rect -152 -433 -52 -400
rect -152 -479 -139 -433
rect -65 -479 -52 -433
rect -152 -492 -52 -479
rect 52 -433 152 -400
rect 52 -479 65 -433
rect 139 -479 152 -433
rect 52 -492 152 -479
rect 256 -433 356 -400
rect 256 -479 269 -433
rect 343 -479 356 -433
rect 256 -492 356 -479
<< polycontact >>
rect -343 433 -269 479
rect -139 433 -65 479
rect 65 433 139 479
rect 269 433 343 479
rect -343 -479 -269 -433
rect -139 -479 -65 -433
rect 65 -479 139 -433
rect 269 -479 343 -433
<< metal1 >>
rect -569 527 569 573
rect -569 470 -523 527
rect -354 433 -343 479
rect -269 433 -258 479
rect -150 433 -139 479
rect -65 433 -54 479
rect 54 433 65 479
rect 139 433 150 479
rect 258 433 269 479
rect 343 433 354 479
rect 523 470 569 527
rect -431 387 -385 398
rect -431 -398 -385 -387
rect -227 387 -181 398
rect -227 -398 -181 -387
rect -23 387 23 398
rect -23 -398 23 -387
rect 181 387 227 398
rect 181 -398 227 -387
rect 385 387 431 398
rect 385 -398 431 -387
rect -569 -527 -523 -470
rect -354 -479 -343 -433
rect -269 -479 -258 -433
rect -150 -479 -139 -433
rect -65 -479 -54 -433
rect 54 -479 65 -433
rect 139 -479 150 -433
rect 258 -479 269 -433
rect 343 -479 354 -433
rect 523 -527 569 -470
rect -569 -573 569 -527
<< properties >>
string FIXED_BBOX -546 -550 546 550
string gencell pfet_03v3
string library gf180mcu
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
