magic
tech gf180mcuD
magscale 1 10
timestamp 1757285905
<< error_s >>
rect 783 -643 794 -597
rect 783 -1555 794 -1509
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 618 -2208 674 -2048
rect 615 -2877 671 -2717
use nfet_03v3_WAUSUP  XM3
timestamp 1757285905
transform 1 0 643 0 1 -2483
box -290 -410 290 410
use pfet_03v3_LSTY94  XM4
timestamp 1757285905
transform 1 0 821 0 1 -1076
box -290 -610 290 610
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 in
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 avss
port 3 nsew
<< end >>
