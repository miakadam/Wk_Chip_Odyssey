magic
tech gf180mcuD
magscale 1 10
timestamp 1758084968
<< nwell >>
rect 94 920 694 1940
rect 982 920 2062 1940
rect -800 -500 -200 520
rect 2322 -256 4290 764
rect 94 -1420 694 -400
rect 982 -1420 2062 -400
<< pwell >>
rect 1714 831 1800 911
rect 94 200 2062 820
rect 3942 -345 4028 -265
rect -548 -589 -462 -509
rect -800 -1220 -200 -600
rect 2322 -976 2922 -356
rect 3006 -446 3606 -356
rect 3006 -704 3652 -446
rect 3006 -976 3606 -704
rect 3690 -976 4290 -356
rect 1714 -1509 1800 -1429
rect 94 -2140 2062 -1520
<< nmos >>
rect 344 410 444 610
rect 548 410 648 610
rect 1028 410 1128 610
rect 1232 410 1332 610
rect 1712 410 1812 610
rect -550 -1010 -450 -810
rect 2572 -766 2672 -566
rect 3256 -766 3356 -566
rect 3940 -766 4040 -566
rect 344 -1930 444 -1730
rect 548 -1930 648 -1730
rect 1028 -1930 1128 -1730
rect 1232 -1930 1332 -1730
rect 1712 -1930 1812 -1730
<< pmos >>
rect 344 1130 444 1730
rect 1232 1130 1332 1730
rect 1712 1130 1812 1730
rect -550 -290 -450 310
rect 2572 -46 2672 554
rect 2776 -46 2876 554
rect 3256 -46 3356 554
rect 3460 -46 3560 554
rect 3940 -46 4040 554
rect 344 -1210 444 -610
rect 1232 -1210 1332 -610
rect 1712 -1210 1812 -610
<< ndiff >>
rect 256 597 344 610
rect 256 423 269 597
rect 315 423 344 597
rect 256 410 344 423
rect 444 597 548 610
rect 444 423 473 597
rect 519 423 548 597
rect 444 410 548 423
rect 648 597 736 610
rect 648 423 677 597
rect 723 423 736 597
rect 648 410 736 423
rect 940 597 1028 610
rect 940 423 953 597
rect 999 423 1028 597
rect 940 410 1028 423
rect 1128 597 1232 610
rect 1128 423 1157 597
rect 1203 423 1232 597
rect 1128 410 1232 423
rect 1332 597 1420 610
rect 1332 423 1361 597
rect 1407 423 1420 597
rect 1332 410 1420 423
rect 1624 597 1712 610
rect 1624 423 1637 597
rect 1683 423 1712 597
rect 1624 410 1712 423
rect 1812 597 1900 610
rect 1812 423 1841 597
rect 1887 423 1900 597
rect 1812 410 1900 423
rect -638 -823 -550 -810
rect -638 -997 -625 -823
rect -579 -997 -550 -823
rect -638 -1010 -550 -997
rect -450 -823 -362 -810
rect -450 -997 -421 -823
rect -375 -997 -362 -823
rect -450 -1010 -362 -997
rect 2484 -579 2572 -566
rect 2484 -753 2497 -579
rect 2543 -753 2572 -579
rect 2484 -766 2572 -753
rect 2672 -579 2760 -566
rect 2672 -753 2701 -579
rect 2747 -753 2760 -579
rect 2672 -766 2760 -753
rect 3168 -579 3256 -566
rect 3168 -753 3181 -579
rect 3227 -753 3256 -579
rect 3168 -766 3256 -753
rect 3356 -579 3444 -566
rect 3356 -753 3385 -579
rect 3431 -753 3444 -579
rect 3356 -766 3444 -753
rect 3852 -579 3940 -566
rect 3852 -753 3865 -579
rect 3911 -753 3940 -579
rect 3852 -766 3940 -753
rect 4040 -579 4128 -566
rect 4040 -753 4069 -579
rect 4115 -753 4128 -579
rect 4040 -766 4128 -753
rect 256 -1743 344 -1730
rect 256 -1917 269 -1743
rect 315 -1917 344 -1743
rect 256 -1930 344 -1917
rect 444 -1743 548 -1730
rect 444 -1917 473 -1743
rect 519 -1917 548 -1743
rect 444 -1930 548 -1917
rect 648 -1743 736 -1730
rect 648 -1917 677 -1743
rect 723 -1917 736 -1743
rect 648 -1930 736 -1917
rect 940 -1743 1028 -1730
rect 940 -1917 953 -1743
rect 999 -1917 1028 -1743
rect 940 -1930 1028 -1917
rect 1128 -1743 1232 -1730
rect 1128 -1917 1157 -1743
rect 1203 -1917 1232 -1743
rect 1128 -1930 1232 -1917
rect 1332 -1743 1420 -1730
rect 1332 -1917 1361 -1743
rect 1407 -1917 1420 -1743
rect 1332 -1930 1420 -1917
rect 1624 -1743 1712 -1730
rect 1624 -1917 1637 -1743
rect 1683 -1917 1712 -1743
rect 1624 -1930 1712 -1917
rect 1812 -1743 1900 -1730
rect 1812 -1917 1841 -1743
rect 1887 -1917 1900 -1743
rect 1812 -1930 1900 -1917
<< pdiff >>
rect 256 1717 344 1730
rect 256 1143 269 1717
rect 315 1143 344 1717
rect 256 1130 344 1143
rect 444 1717 532 1730
rect 444 1143 473 1717
rect 519 1143 532 1717
rect 444 1130 532 1143
rect 1144 1717 1232 1730
rect 1144 1143 1157 1717
rect 1203 1143 1232 1717
rect 1144 1130 1232 1143
rect 1332 1717 1420 1730
rect 1332 1143 1361 1717
rect 1407 1143 1420 1717
rect 1332 1130 1420 1143
rect 1624 1717 1712 1730
rect 1624 1143 1637 1717
rect 1683 1143 1712 1717
rect 1624 1130 1712 1143
rect 1812 1717 1900 1730
rect 1812 1143 1841 1717
rect 1887 1143 1900 1717
rect 1812 1130 1900 1143
rect -638 297 -550 310
rect -638 -277 -625 297
rect -579 -277 -550 297
rect -638 -290 -550 -277
rect -450 297 -362 310
rect -450 -277 -421 297
rect -375 -277 -362 297
rect -450 -290 -362 -277
rect 2484 541 2572 554
rect 2484 -33 2497 541
rect 2543 -33 2572 541
rect 2484 -46 2572 -33
rect 2672 541 2776 554
rect 2672 -33 2701 541
rect 2747 -33 2776 541
rect 2672 -46 2776 -33
rect 2876 541 2964 554
rect 2876 -33 2905 541
rect 2951 -33 2964 541
rect 2876 -46 2964 -33
rect 3168 541 3256 554
rect 3168 -33 3181 541
rect 3227 -33 3256 541
rect 3168 -46 3256 -33
rect 3356 541 3460 554
rect 3356 -33 3385 541
rect 3431 -33 3460 541
rect 3356 -46 3460 -33
rect 3560 541 3648 554
rect 3560 -33 3589 541
rect 3635 -33 3648 541
rect 3560 -46 3648 -33
rect 3852 541 3940 554
rect 3852 -33 3865 541
rect 3911 -33 3940 541
rect 3852 -46 3940 -33
rect 4040 541 4128 554
rect 4040 -33 4069 541
rect 4115 -33 4128 541
rect 4040 -46 4128 -33
rect 256 -623 344 -610
rect 256 -1197 269 -623
rect 315 -1197 344 -623
rect 256 -1210 344 -1197
rect 444 -623 532 -610
rect 444 -1197 473 -623
rect 519 -1197 532 -623
rect 444 -1210 532 -1197
rect 1144 -623 1232 -610
rect 1144 -1197 1157 -623
rect 1203 -1197 1232 -623
rect 1144 -1210 1232 -1197
rect 1332 -623 1420 -610
rect 1332 -1197 1361 -623
rect 1407 -1197 1420 -623
rect 1332 -1210 1420 -1197
rect 1624 -623 1712 -610
rect 1624 -1197 1637 -623
rect 1683 -1197 1712 -623
rect 1624 -1210 1712 -1197
rect 1812 -623 1900 -610
rect 1812 -1197 1841 -623
rect 1887 -1197 1900 -623
rect 1812 -1210 1900 -1197
<< ndiffc >>
rect 269 423 315 597
rect 473 423 519 597
rect 677 423 723 597
rect 953 423 999 597
rect 1157 423 1203 597
rect 1361 423 1407 597
rect 1637 423 1683 597
rect 1841 423 1887 597
rect -625 -997 -579 -823
rect -421 -997 -375 -823
rect 2497 -753 2543 -579
rect 2701 -753 2747 -579
rect 3181 -753 3227 -579
rect 3385 -753 3431 -579
rect 3865 -753 3911 -579
rect 4069 -753 4115 -579
rect 269 -1917 315 -1743
rect 473 -1917 519 -1743
rect 677 -1917 723 -1743
rect 953 -1917 999 -1743
rect 1157 -1917 1203 -1743
rect 1361 -1917 1407 -1743
rect 1637 -1917 1683 -1743
rect 1841 -1917 1887 -1743
<< pdiffc >>
rect 269 1143 315 1717
rect 473 1143 519 1717
rect 1157 1143 1203 1717
rect 1361 1143 1407 1717
rect 1637 1143 1683 1717
rect 1841 1143 1887 1717
rect -625 -277 -579 297
rect -421 -277 -375 297
rect 2497 -33 2543 541
rect 2701 -33 2747 541
rect 2905 -33 2951 541
rect 3181 -33 3227 541
rect 3385 -33 3431 541
rect 3589 -33 3635 541
rect 3865 -33 3911 541
rect 4069 -33 4115 541
rect 269 -1197 315 -623
rect 473 -1197 519 -623
rect 1157 -1197 1203 -623
rect 1361 -1197 1407 -623
rect 1637 -1197 1683 -623
rect 1841 -1197 1887 -623
<< psubdiff >>
rect 118 724 2038 796
rect 118 680 190 724
rect 118 340 131 680
rect 177 340 190 680
rect 802 680 874 724
rect 118 296 190 340
rect 802 340 815 680
rect 861 340 874 680
rect 1486 680 1558 724
rect 802 296 874 340
rect 1486 340 1499 680
rect 1545 340 1558 680
rect 1966 680 2038 724
rect 1486 296 1558 340
rect 1966 340 1979 680
rect 2025 340 2038 680
rect 1966 296 2038 340
rect 118 224 2038 296
rect -776 -696 -224 -624
rect -776 -740 -704 -696
rect -776 -1080 -763 -740
rect -717 -1080 -704 -740
rect -296 -740 -224 -696
rect -776 -1124 -704 -1080
rect -296 -1080 -283 -740
rect -237 -1080 -224 -740
rect -296 -1124 -224 -1080
rect -776 -1196 -224 -1124
rect 2346 -452 2898 -380
rect 2346 -496 2418 -452
rect 2346 -836 2359 -496
rect 2405 -836 2418 -496
rect 2826 -496 2898 -452
rect 2346 -880 2418 -836
rect 2826 -836 2839 -496
rect 2885 -836 2898 -496
rect 2826 -880 2898 -836
rect 2346 -952 2898 -880
rect 3030 -452 3582 -380
rect 3030 -496 3102 -452
rect 3030 -836 3043 -496
rect 3089 -836 3102 -496
rect 3510 -496 3582 -452
rect 3030 -880 3102 -836
rect 3510 -836 3523 -496
rect 3569 -836 3582 -496
rect 3510 -880 3582 -836
rect 3030 -952 3582 -880
rect 3714 -452 4266 -380
rect 3714 -496 3786 -452
rect 3714 -836 3727 -496
rect 3773 -836 3786 -496
rect 4194 -496 4266 -452
rect 3714 -880 3786 -836
rect 4194 -836 4207 -496
rect 4253 -836 4266 -496
rect 4194 -880 4266 -836
rect 3714 -952 4266 -880
rect 118 -1616 2038 -1544
rect 118 -1660 190 -1616
rect 118 -2000 131 -1660
rect 177 -2000 190 -1660
rect 802 -1660 874 -1616
rect 118 -2044 190 -2000
rect 802 -2000 815 -1660
rect 861 -2000 874 -1660
rect 1486 -1660 1558 -1616
rect 802 -2044 874 -2000
rect 1486 -2000 1499 -1660
rect 1545 -2000 1558 -1660
rect 1966 -1660 2038 -1616
rect 1486 -2044 1558 -2000
rect 1966 -2000 1979 -1660
rect 2025 -2000 2038 -1660
rect 1966 -2044 2038 -2000
rect 118 -2116 2038 -2044
<< nsubdiff >>
rect 118 1844 670 1916
rect 118 1800 190 1844
rect 118 1060 131 1800
rect 177 1060 190 1800
rect 598 1800 670 1844
rect 118 1016 190 1060
rect 598 1060 611 1800
rect 657 1060 670 1800
rect 598 1016 670 1060
rect 118 944 670 1016
rect 1006 1844 2038 1916
rect 1006 1800 1078 1844
rect 1006 1060 1019 1800
rect 1065 1060 1078 1800
rect 1486 1800 1558 1844
rect 1006 1016 1078 1060
rect 1486 1060 1499 1800
rect 1545 1060 1558 1800
rect 1966 1800 2038 1844
rect 1486 1016 1558 1060
rect 1966 1060 1979 1800
rect 2025 1060 2038 1800
rect 1966 1016 2038 1060
rect 1006 944 2038 1016
rect -776 424 -224 496
rect -776 380 -704 424
rect -776 -360 -763 380
rect -717 -360 -704 380
rect -296 380 -224 424
rect -776 -404 -704 -360
rect -296 -360 -283 380
rect -237 -360 -224 380
rect 2346 668 4266 740
rect 2346 624 2418 668
rect 2346 -116 2359 624
rect 2405 -116 2418 624
rect 3030 624 3102 668
rect 2346 -160 2418 -116
rect 3030 -116 3043 624
rect 3089 -116 3102 624
rect 3714 624 3786 668
rect 3030 -160 3102 -116
rect 3714 -116 3727 624
rect 3773 -116 3786 624
rect 4194 624 4266 668
rect 3714 -160 3786 -116
rect 4194 -116 4207 624
rect 4253 -116 4266 624
rect 4194 -160 4266 -116
rect 2346 -232 4266 -160
rect -296 -404 -224 -360
rect -776 -476 -224 -404
rect 118 -496 670 -424
rect 118 -540 190 -496
rect 118 -1280 131 -540
rect 177 -1280 190 -540
rect 598 -540 670 -496
rect 118 -1324 190 -1280
rect 598 -1280 611 -540
rect 657 -1280 670 -540
rect 598 -1324 670 -1280
rect 118 -1396 670 -1324
rect 1006 -496 2038 -424
rect 1006 -540 1078 -496
rect 1006 -1280 1019 -540
rect 1065 -1280 1078 -540
rect 1486 -540 1558 -496
rect 1006 -1324 1078 -1280
rect 1486 -1280 1499 -540
rect 1545 -1280 1558 -540
rect 1966 -540 2038 -496
rect 1486 -1324 1558 -1280
rect 1966 -1280 1979 -540
rect 2025 -1280 2038 -540
rect 1966 -1324 2038 -1280
rect 1006 -1396 2038 -1324
<< psubdiffcont >>
rect 131 340 177 680
rect 815 340 861 680
rect 1499 340 1545 680
rect 1979 340 2025 680
rect -763 -1080 -717 -740
rect -283 -1080 -237 -740
rect 2359 -836 2405 -496
rect 2839 -836 2885 -496
rect 3043 -836 3089 -496
rect 3523 -836 3569 -496
rect 3727 -836 3773 -496
rect 4207 -836 4253 -496
rect 131 -2000 177 -1660
rect 815 -2000 861 -1660
rect 1499 -2000 1545 -1660
rect 1979 -2000 2025 -1660
<< nsubdiffcont >>
rect 131 1060 177 1800
rect 611 1060 657 1800
rect 1019 1060 1065 1800
rect 1499 1060 1545 1800
rect 1979 1060 2025 1800
rect -763 -360 -717 380
rect -283 -360 -237 380
rect 2359 -116 2405 624
rect 3043 -116 3089 624
rect 3727 -116 3773 624
rect 4207 -116 4253 624
rect 131 -1280 177 -540
rect 611 -1280 657 -540
rect 1019 -1280 1065 -540
rect 1499 -1280 1545 -540
rect 1979 -1280 2025 -540
<< polysilicon >>
rect 344 1809 444 1822
rect 344 1763 357 1809
rect 431 1763 444 1809
rect 344 1730 444 1763
rect 344 1097 444 1130
rect 344 1051 357 1097
rect 431 1051 444 1097
rect 344 1038 444 1051
rect 1232 1809 1332 1822
rect 1232 1763 1245 1809
rect 1319 1763 1332 1809
rect 1232 1730 1332 1763
rect 1232 1097 1332 1130
rect 1232 1051 1245 1097
rect 1319 1051 1332 1097
rect 1232 1038 1332 1051
rect 1712 1809 1812 1822
rect 1712 1763 1725 1809
rect 1799 1763 1812 1809
rect 1712 1730 1812 1763
rect 1712 1097 1812 1130
rect 1712 1051 1725 1097
rect 1799 1051 1812 1097
rect 1712 1038 1812 1051
rect -550 389 -450 402
rect -550 343 -537 389
rect -463 343 -450 389
rect -550 310 -450 343
rect -550 -323 -450 -290
rect -550 -369 -537 -323
rect -463 -369 -450 -323
rect -550 -382 -450 -369
rect 344 689 444 702
rect 344 643 357 689
rect 431 643 444 689
rect 344 610 444 643
rect 548 689 648 702
rect 548 643 561 689
rect 635 643 648 689
rect 548 610 648 643
rect 344 377 444 410
rect 344 331 357 377
rect 431 331 444 377
rect 344 318 444 331
rect 548 377 648 410
rect 548 331 561 377
rect 635 331 648 377
rect 548 318 648 331
rect 1028 689 1128 702
rect 1028 643 1041 689
rect 1115 643 1128 689
rect 1028 610 1128 643
rect 1232 689 1332 702
rect 1232 643 1245 689
rect 1319 643 1332 689
rect 1232 610 1332 643
rect 1028 377 1128 410
rect 1028 331 1041 377
rect 1115 331 1128 377
rect 1028 318 1128 331
rect 1232 377 1332 410
rect 1232 331 1245 377
rect 1319 331 1332 377
rect 1232 318 1332 331
rect 1712 689 1812 702
rect 1712 643 1725 689
rect 1799 643 1812 689
rect 1712 610 1812 643
rect 1712 377 1812 410
rect 1712 331 1725 377
rect 1799 331 1812 377
rect 1712 318 1812 331
rect 2572 633 2672 646
rect 2572 587 2585 633
rect 2659 587 2672 633
rect 2572 554 2672 587
rect 2776 633 2876 646
rect 2776 587 2789 633
rect 2863 587 2876 633
rect 2776 554 2876 587
rect 2572 -79 2672 -46
rect 2572 -125 2585 -79
rect 2659 -125 2672 -79
rect 2572 -138 2672 -125
rect 2776 -79 2876 -46
rect 2776 -125 2789 -79
rect 2863 -125 2876 -79
rect 2776 -138 2876 -125
rect 3256 633 3356 646
rect 3256 587 3269 633
rect 3343 587 3356 633
rect 3256 554 3356 587
rect 3460 633 3560 646
rect 3460 587 3473 633
rect 3547 587 3560 633
rect 3460 554 3560 587
rect 3256 -79 3356 -46
rect 3256 -125 3269 -79
rect 3343 -125 3356 -79
rect 3256 -138 3356 -125
rect 3460 -79 3560 -46
rect 3460 -125 3473 -79
rect 3547 -125 3560 -79
rect 3460 -138 3560 -125
rect 3940 633 4040 646
rect 3940 587 3953 633
rect 4027 587 4040 633
rect 3940 554 4040 587
rect 3940 -79 4040 -46
rect 3940 -125 3953 -79
rect 4027 -125 4040 -79
rect 3940 -138 4040 -125
rect -550 -731 -450 -718
rect -550 -777 -537 -731
rect -463 -777 -450 -731
rect -550 -810 -450 -777
rect -550 -1043 -450 -1010
rect -550 -1089 -537 -1043
rect -463 -1089 -450 -1043
rect -550 -1102 -450 -1089
rect 344 -531 444 -518
rect 344 -577 357 -531
rect 431 -577 444 -531
rect 344 -610 444 -577
rect 344 -1243 444 -1210
rect 344 -1289 357 -1243
rect 431 -1289 444 -1243
rect 344 -1302 444 -1289
rect 1232 -531 1332 -518
rect 1232 -577 1245 -531
rect 1319 -577 1332 -531
rect 1232 -610 1332 -577
rect 1232 -1243 1332 -1210
rect 1232 -1289 1245 -1243
rect 1319 -1289 1332 -1243
rect 1232 -1302 1332 -1289
rect 1712 -531 1812 -518
rect 1712 -577 1725 -531
rect 1799 -577 1812 -531
rect 1712 -610 1812 -577
rect 1712 -1243 1812 -1210
rect 1712 -1289 1725 -1243
rect 1799 -1289 1812 -1243
rect 1712 -1302 1812 -1289
rect 2572 -487 2672 -474
rect 2572 -533 2585 -487
rect 2659 -533 2672 -487
rect 2572 -566 2672 -533
rect 2572 -799 2672 -766
rect 2572 -845 2585 -799
rect 2659 -845 2672 -799
rect 2572 -858 2672 -845
rect 3256 -487 3356 -474
rect 3256 -533 3269 -487
rect 3343 -533 3356 -487
rect 3256 -566 3356 -533
rect 3256 -799 3356 -766
rect 3256 -845 3269 -799
rect 3343 -845 3356 -799
rect 3256 -858 3356 -845
rect 3940 -487 4040 -474
rect 3940 -533 3953 -487
rect 4027 -533 4040 -487
rect 3940 -566 4040 -533
rect 3940 -799 4040 -766
rect 3940 -845 3953 -799
rect 4027 -845 4040 -799
rect 3940 -858 4040 -845
rect 344 -1651 444 -1638
rect 344 -1697 357 -1651
rect 431 -1697 444 -1651
rect 344 -1730 444 -1697
rect 548 -1651 648 -1638
rect 548 -1697 561 -1651
rect 635 -1697 648 -1651
rect 548 -1730 648 -1697
rect 344 -1963 444 -1930
rect 344 -2009 357 -1963
rect 431 -2009 444 -1963
rect 344 -2022 444 -2009
rect 548 -1963 648 -1930
rect 548 -2009 561 -1963
rect 635 -2009 648 -1963
rect 548 -2022 648 -2009
rect 1028 -1651 1128 -1638
rect 1028 -1697 1041 -1651
rect 1115 -1697 1128 -1651
rect 1028 -1730 1128 -1697
rect 1232 -1651 1332 -1638
rect 1232 -1697 1245 -1651
rect 1319 -1697 1332 -1651
rect 1232 -1730 1332 -1697
rect 1028 -1963 1128 -1930
rect 1028 -2009 1041 -1963
rect 1115 -2009 1128 -1963
rect 1028 -2022 1128 -2009
rect 1232 -1963 1332 -1930
rect 1232 -2009 1245 -1963
rect 1319 -2009 1332 -1963
rect 1232 -2022 1332 -2009
rect 1712 -1651 1812 -1638
rect 1712 -1697 1725 -1651
rect 1799 -1697 1812 -1651
rect 1712 -1730 1812 -1697
rect 1712 -1963 1812 -1930
rect 1712 -2009 1725 -1963
rect 1799 -2009 1812 -1963
rect 1712 -2022 1812 -2009
<< polycontact >>
rect 357 1763 431 1809
rect 357 1051 431 1097
rect 1245 1763 1319 1809
rect 1245 1051 1319 1097
rect 1725 1763 1799 1809
rect 1725 1051 1799 1097
rect -537 343 -463 389
rect -537 -369 -463 -323
rect 357 643 431 689
rect 561 643 635 689
rect 357 331 431 377
rect 561 331 635 377
rect 1041 643 1115 689
rect 1245 643 1319 689
rect 1041 331 1115 377
rect 1245 331 1319 377
rect 1725 643 1799 689
rect 1725 331 1799 377
rect 2585 587 2659 633
rect 2789 587 2863 633
rect 2585 -125 2659 -79
rect 2789 -125 2863 -79
rect 3269 587 3343 633
rect 3473 587 3547 633
rect 3269 -125 3343 -79
rect 3473 -125 3547 -79
rect 3953 587 4027 633
rect 3953 -125 4027 -79
rect -537 -777 -463 -731
rect -537 -1089 -463 -1043
rect 357 -577 431 -531
rect 357 -1289 431 -1243
rect 1245 -577 1319 -531
rect 1245 -1289 1319 -1243
rect 1725 -577 1799 -531
rect 1725 -1289 1799 -1243
rect 2585 -533 2659 -487
rect 2585 -845 2659 -799
rect 3269 -533 3343 -487
rect 3269 -845 3343 -799
rect 3953 -533 4027 -487
rect 3953 -845 4027 -799
rect 357 -1697 431 -1651
rect 561 -1697 635 -1651
rect 357 -2009 431 -1963
rect 561 -2009 635 -1963
rect 1041 -1697 1115 -1651
rect 1245 -1697 1319 -1651
rect 1041 -2009 1115 -1963
rect 1245 -2009 1319 -1963
rect 1725 -1697 1799 -1651
rect 1725 -2009 1799 -1963
<< metal1 >>
rect -800 1940 4290 2140
rect -800 520 -200 1940
rect 131 1800 177 1811
rect 346 1809 442 1840
rect 346 1763 357 1809
rect 431 1763 442 1809
rect 611 1800 1065 1940
rect 269 1717 315 1728
rect 252 1433 269 1443
rect 473 1717 611 1728
rect 315 1433 332 1443
rect 252 1193 264 1433
rect 320 1193 332 1433
rect 252 1183 269 1193
rect 315 1183 332 1193
rect 269 1132 315 1143
rect 519 1143 611 1717
rect 473 1132 611 1143
rect 131 1049 177 1060
rect 346 1051 357 1097
rect 431 1051 442 1097
rect 346 976 442 1051
rect 657 1132 1019 1800
rect 611 1049 657 1060
rect 1234 1809 1330 1840
rect 1234 1763 1245 1809
rect 1319 1763 1330 1809
rect 1499 1800 1545 1940
rect 1065 1717 1203 1728
rect 1065 1143 1157 1717
rect 1361 1717 1407 1728
rect 1344 1433 1361 1443
rect 1407 1433 1424 1443
rect 1344 1193 1356 1433
rect 1412 1193 1424 1433
rect 1344 1183 1361 1193
rect 1065 1132 1203 1143
rect 1407 1183 1424 1193
rect 1361 1132 1407 1143
rect 1019 1049 1065 1060
rect 1234 1051 1245 1097
rect 1319 1051 1330 1097
rect 346 920 366 976
rect 422 920 442 976
rect 346 702 442 920
rect 1234 832 1330 1051
rect 1714 1809 1810 1840
rect 1714 1763 1725 1809
rect 1799 1763 1810 1809
rect 1979 1800 2025 1940
rect 1545 1717 1683 1728
rect 1545 1143 1637 1717
rect 1841 1717 1887 1728
rect 1824 1433 1841 1443
rect 1887 1433 1904 1443
rect 1824 1193 1836 1433
rect 1892 1193 1904 1433
rect 1824 1183 1841 1193
rect 1545 1132 1683 1143
rect 1887 1183 1904 1193
rect 1841 1132 1887 1143
rect 1499 1049 1545 1060
rect 1714 1051 1725 1097
rect 1799 1051 1810 1097
rect 1714 910 1810 1051
rect 1979 1049 2025 1060
rect 1166 820 1330 832
rect 1646 898 1810 910
rect 1646 842 1658 898
rect 1714 842 1810 898
rect 1646 830 1810 842
rect 1166 764 1178 820
rect 1234 764 1330 820
rect 1166 752 1330 764
rect 1234 702 1330 752
rect 131 680 177 691
rect -763 380 -717 520
rect -548 389 -452 420
rect -548 343 -537 389
rect -463 343 -452 389
rect -283 380 -237 520
rect -717 297 -579 308
rect -717 -277 -625 297
rect -421 297 -375 308
rect -438 13 -421 23
rect -375 13 -358 23
rect -438 -227 -426 13
rect -370 -227 -358 13
rect -438 -237 -421 -227
rect -717 -288 -579 -277
rect -375 -237 -358 -227
rect -421 -288 -375 -277
rect -763 -371 -717 -360
rect -548 -369 -537 -323
rect -463 -369 -452 -323
rect -548 -510 -452 -369
rect 346 689 646 702
rect 346 643 357 689
rect 431 656 561 689
rect 431 643 442 656
rect 550 643 561 656
rect 635 643 646 689
rect 815 680 861 691
rect 177 597 315 608
rect 177 423 269 597
rect 473 597 519 608
rect 456 538 473 548
rect 677 597 815 608
rect 519 538 536 548
rect 456 482 468 538
rect 524 482 536 538
rect 456 472 473 482
rect 177 412 315 423
rect 519 472 536 482
rect 473 412 519 423
rect 723 423 815 597
rect 677 412 815 423
rect 131 200 177 340
rect 346 331 357 377
rect 431 331 442 377
rect 346 300 442 331
rect 550 331 561 377
rect 635 331 646 377
rect 550 300 646 331
rect 1030 689 1330 702
rect 1030 643 1041 689
rect 1115 656 1245 689
rect 1115 643 1126 656
rect 1234 643 1245 656
rect 1319 643 1330 689
rect 1499 680 1545 691
rect 953 597 999 608
rect 936 538 953 548
rect 1157 597 1203 608
rect 999 538 1016 548
rect 936 482 948 538
rect 1004 482 1016 538
rect 936 472 953 482
rect 999 472 1016 482
rect 1140 538 1157 548
rect 1361 597 1407 608
rect 1203 538 1220 548
rect 1140 482 1152 538
rect 1208 482 1220 538
rect 1140 472 1157 482
rect 953 412 999 423
rect 1203 472 1220 482
rect 1344 538 1361 548
rect 1407 538 1424 548
rect 1344 482 1356 538
rect 1412 482 1424 538
rect 1344 472 1361 482
rect 1157 412 1203 423
rect 1407 472 1424 482
rect 1361 412 1407 423
rect 815 200 861 340
rect 1030 331 1041 377
rect 1115 331 1126 377
rect 1030 300 1126 331
rect 1234 331 1245 377
rect 1319 331 1330 377
rect 1234 300 1330 331
rect 1714 689 1810 830
rect 2322 944 4290 1940
rect 2322 804 2422 944
rect 4190 804 4290 944
rect 2322 764 4290 804
rect 1714 643 1725 689
rect 1799 643 1810 689
rect 1979 680 2025 691
rect 1545 597 1683 608
rect 1545 423 1637 597
rect 1841 597 1887 608
rect 1824 538 1841 548
rect 1887 538 1904 548
rect 1824 482 1836 538
rect 1892 482 1904 538
rect 1824 472 1841 482
rect 1545 412 1683 423
rect 1887 472 1904 482
rect 1841 412 1887 423
rect 1499 200 1545 340
rect 1714 331 1725 377
rect 1799 331 1810 377
rect 1714 300 1810 331
rect 1979 200 2025 340
rect 2359 624 2405 764
rect 94 170 2062 200
rect 94 30 1362 170
rect 1962 30 2062 170
rect 94 0 2062 30
rect 2574 633 2670 664
rect 2574 587 2585 633
rect 2659 587 2670 633
rect 2778 633 2874 664
rect 2778 587 2789 633
rect 2863 587 2874 633
rect 3043 624 3089 764
rect 2405 541 2543 552
rect 2701 541 2747 552
rect 2905 541 3043 552
rect 2405 -33 2497 541
rect 2684 301 2696 541
rect 2752 301 2764 541
rect 2405 -44 2543 -33
rect 2701 -44 2747 -33
rect 2951 -33 3043 541
rect 2905 -44 3043 -33
rect 2359 -127 2405 -116
rect 2574 -125 2585 -79
rect 2659 -99 2670 -79
rect 2778 -99 2789 -79
rect 2659 -125 2789 -99
rect 2863 -125 2874 -79
rect 2574 -152 2874 -125
rect 3258 633 3354 664
rect 3258 587 3269 633
rect 3343 587 3354 633
rect 3462 633 3558 664
rect 3462 587 3473 633
rect 3547 587 3558 633
rect 3727 624 3773 764
rect 3181 541 3227 552
rect 3385 541 3431 552
rect 3589 541 3635 552
rect 3368 301 3380 541
rect 3436 301 3448 541
rect 3164 -33 3176 207
rect 3232 -33 3244 207
rect 3572 -33 3584 207
rect 3640 -33 3652 207
rect 3181 -44 3227 -33
rect 3385 -44 3431 -33
rect 3589 -44 3635 -33
rect 3043 -127 3089 -116
rect 3258 -125 3269 -79
rect 3343 -99 3354 -79
rect 3462 -99 3473 -79
rect 3343 -125 3473 -99
rect 3547 -125 3558 -79
rect 3258 -152 3558 -125
rect 3942 633 4038 664
rect 3942 587 3953 633
rect 4027 587 4038 633
rect 4207 624 4253 764
rect 3773 541 3911 552
rect 3773 -33 3865 541
rect 4069 541 4115 552
rect 4052 257 4069 267
rect 4115 257 4132 267
rect 4052 17 4064 257
rect 4120 17 4132 257
rect 4052 7 4069 17
rect 3773 -44 3911 -33
rect 4115 7 4132 17
rect 4069 -44 4115 -33
rect 3727 -127 3773 -116
rect 3942 -125 3953 -79
rect 4027 -125 4038 -79
rect 2574 -200 2670 -152
rect -283 -371 -237 -360
rect 94 -230 2062 -200
rect 94 -370 1362 -230
rect 1962 -370 2062 -230
rect 94 -400 2062 -370
rect 2574 -256 2594 -200
rect 2650 -256 2670 -200
rect -616 -522 -452 -510
rect -616 -578 -604 -522
rect -548 -578 -452 -522
rect -616 -590 -452 -578
rect -763 -740 -717 -729
rect -548 -731 -452 -590
rect 131 -540 177 -529
rect -548 -777 -537 -731
rect -463 -777 -452 -731
rect -283 -740 -237 -729
rect -717 -823 -579 -812
rect -717 -997 -625 -823
rect -421 -823 -375 -812
rect -438 -882 -421 -872
rect -375 -882 -358 -872
rect -438 -938 -426 -882
rect -370 -938 -358 -882
rect -438 -948 -421 -938
rect -717 -1008 -579 -997
rect -375 -948 -358 -938
rect -421 -1008 -375 -997
rect -763 -1220 -717 -1080
rect -548 -1089 -537 -1043
rect -463 -1089 -452 -1043
rect -548 -1120 -452 -1089
rect -283 -1220 -237 -1080
rect -800 -2140 -200 -1220
rect 346 -531 442 -500
rect 346 -577 357 -531
rect 431 -577 442 -531
rect 611 -540 1065 -400
rect 269 -623 315 -612
rect 252 -907 269 -897
rect 473 -623 611 -612
rect 315 -907 332 -897
rect 252 -1147 264 -907
rect 320 -1147 332 -907
rect 252 -1157 269 -1147
rect 315 -1157 332 -1147
rect 269 -1208 315 -1197
rect 519 -1197 611 -623
rect 473 -1208 611 -1197
rect 131 -1291 177 -1280
rect 346 -1289 357 -1243
rect 431 -1289 442 -1243
rect 346 -1364 442 -1289
rect 657 -1208 1019 -540
rect 611 -1291 657 -1280
rect 1234 -531 1330 -500
rect 1234 -577 1245 -531
rect 1319 -577 1330 -531
rect 1499 -540 1545 -400
rect 1065 -623 1203 -612
rect 1065 -1197 1157 -623
rect 1361 -623 1407 -612
rect 1344 -907 1361 -897
rect 1407 -907 1424 -897
rect 1344 -1147 1356 -907
rect 1412 -1147 1424 -907
rect 1344 -1157 1361 -1147
rect 1065 -1208 1203 -1197
rect 1407 -1157 1424 -1147
rect 1361 -1208 1407 -1197
rect 1019 -1291 1065 -1280
rect 1234 -1289 1245 -1243
rect 1319 -1289 1330 -1243
rect 346 -1420 366 -1364
rect 422 -1420 442 -1364
rect 346 -1638 442 -1420
rect 1234 -1508 1330 -1289
rect 1714 -531 1810 -500
rect 1714 -577 1725 -531
rect 1799 -577 1810 -531
rect 1979 -540 2025 -400
rect 1545 -623 1683 -612
rect 1545 -1197 1637 -623
rect 1841 -623 1887 -612
rect 1824 -907 1841 -897
rect 1887 -907 1904 -897
rect 1824 -1147 1836 -907
rect 1892 -1147 1904 -907
rect 1824 -1157 1841 -1147
rect 1545 -1208 1683 -1197
rect 1887 -1157 1904 -1147
rect 1841 -1208 1887 -1197
rect 1499 -1291 1545 -1280
rect 1714 -1289 1725 -1243
rect 1799 -1289 1810 -1243
rect 1714 -1430 1810 -1289
rect 2359 -496 2405 -485
rect 2574 -487 2670 -256
rect 3258 -356 3354 -152
rect 3942 -266 4038 -125
rect 4207 -127 4253 -116
rect 3874 -278 4038 -266
rect 3874 -334 3886 -278
rect 3942 -334 4038 -278
rect 3874 -346 4038 -334
rect 3258 -412 3278 -356
rect 3334 -412 3354 -356
rect 2574 -533 2585 -487
rect 2659 -533 2670 -487
rect 2839 -496 3089 -485
rect 2497 -579 2543 -568
rect 2480 -638 2497 -628
rect 2701 -579 2839 -568
rect 2543 -638 2560 -628
rect 2480 -694 2492 -638
rect 2548 -694 2560 -638
rect 2480 -704 2497 -694
rect 2543 -704 2560 -694
rect 2497 -764 2543 -753
rect 2747 -753 2839 -579
rect 2701 -764 2839 -753
rect 2359 -976 2405 -836
rect 2574 -845 2585 -799
rect 2659 -845 2670 -799
rect 2574 -876 2670 -845
rect 2885 -836 3043 -496
rect 3258 -487 3354 -412
rect 3258 -533 3269 -487
rect 3343 -533 3354 -487
rect 3523 -496 3569 -485
rect 3089 -579 3227 -568
rect 3089 -753 3181 -579
rect 3385 -579 3431 -568
rect 3368 -638 3385 -628
rect 3431 -638 3448 -628
rect 3368 -694 3380 -638
rect 3436 -694 3448 -638
rect 3368 -704 3385 -694
rect 3089 -764 3227 -753
rect 3431 -704 3448 -694
rect 3385 -764 3431 -753
rect 2839 -847 3089 -836
rect 3258 -845 3269 -799
rect 3343 -845 3354 -799
rect 2885 -976 3043 -847
rect 3258 -876 3354 -845
rect 3523 -976 3569 -836
rect 3727 -496 3773 -485
rect 3942 -487 4038 -346
rect 3942 -533 3953 -487
rect 4027 -533 4038 -487
rect 4207 -496 4253 -485
rect 3773 -579 3911 -568
rect 3773 -753 3865 -579
rect 4069 -579 4115 -568
rect 4052 -638 4069 -628
rect 4115 -638 4132 -628
rect 4052 -694 4064 -638
rect 4120 -694 4132 -638
rect 4052 -704 4069 -694
rect 3773 -764 3911 -753
rect 4115 -704 4132 -694
rect 4069 -764 4115 -753
rect 3727 -976 3773 -836
rect 3942 -845 3953 -799
rect 4027 -845 4038 -799
rect 3942 -876 4038 -845
rect 4207 -976 4253 -836
rect 1979 -1291 2025 -1280
rect 2322 -1016 4290 -976
rect 2322 -1156 2422 -1016
rect 4190 -1156 4290 -1016
rect 1166 -1520 1330 -1508
rect 1646 -1442 1810 -1430
rect 1646 -1498 1658 -1442
rect 1714 -1498 1810 -1442
rect 1646 -1510 1810 -1498
rect 1166 -1576 1178 -1520
rect 1234 -1576 1330 -1520
rect 1166 -1588 1330 -1576
rect 1234 -1638 1330 -1588
rect 131 -1660 177 -1649
rect 346 -1651 646 -1638
rect 346 -1697 357 -1651
rect 431 -1684 561 -1651
rect 431 -1697 442 -1684
rect 550 -1697 561 -1684
rect 635 -1697 646 -1651
rect 815 -1660 861 -1649
rect 177 -1743 315 -1732
rect 177 -1917 269 -1743
rect 473 -1743 519 -1732
rect 456 -1802 473 -1792
rect 677 -1743 815 -1732
rect 519 -1802 536 -1792
rect 456 -1858 468 -1802
rect 524 -1858 536 -1802
rect 456 -1868 473 -1858
rect 177 -1928 315 -1917
rect 519 -1868 536 -1858
rect 473 -1928 519 -1917
rect 723 -1917 815 -1743
rect 677 -1928 815 -1917
rect 131 -2140 177 -2000
rect 346 -2009 357 -1963
rect 431 -2009 442 -1963
rect 346 -2040 442 -2009
rect 550 -2009 561 -1963
rect 635 -2009 646 -1963
rect 550 -2040 646 -2009
rect 1030 -1651 1330 -1638
rect 1030 -1697 1041 -1651
rect 1115 -1684 1245 -1651
rect 1115 -1697 1126 -1684
rect 1234 -1697 1245 -1684
rect 1319 -1697 1330 -1651
rect 1499 -1660 1545 -1649
rect 953 -1743 999 -1732
rect 936 -1802 953 -1792
rect 1157 -1743 1203 -1732
rect 999 -1802 1016 -1792
rect 936 -1858 948 -1802
rect 1004 -1858 1016 -1802
rect 936 -1868 953 -1858
rect 999 -1868 1016 -1858
rect 1140 -1802 1157 -1792
rect 1361 -1743 1407 -1732
rect 1203 -1802 1220 -1792
rect 1140 -1858 1152 -1802
rect 1208 -1858 1220 -1802
rect 1140 -1868 1157 -1858
rect 953 -1928 999 -1917
rect 1203 -1868 1220 -1858
rect 1344 -1802 1361 -1792
rect 1407 -1802 1424 -1792
rect 1344 -1858 1356 -1802
rect 1412 -1858 1424 -1802
rect 1344 -1868 1361 -1858
rect 1157 -1928 1203 -1917
rect 1407 -1868 1424 -1858
rect 1361 -1928 1407 -1917
rect 815 -2140 861 -2000
rect 1030 -2009 1041 -1963
rect 1115 -2009 1126 -1963
rect 1030 -2040 1126 -2009
rect 1234 -2009 1245 -1963
rect 1319 -2009 1330 -1963
rect 1234 -2040 1330 -2009
rect 1714 -1651 1810 -1510
rect 1714 -1697 1725 -1651
rect 1799 -1697 1810 -1651
rect 1979 -1660 2025 -1649
rect 1545 -1743 1683 -1732
rect 1545 -1917 1637 -1743
rect 1841 -1743 1887 -1732
rect 1824 -1802 1841 -1792
rect 1887 -1802 1904 -1792
rect 1824 -1858 1836 -1802
rect 1892 -1858 1904 -1802
rect 1824 -1868 1841 -1858
rect 1545 -1928 1683 -1917
rect 1887 -1868 1904 -1858
rect 1841 -1928 1887 -1917
rect 1499 -2140 1545 -2000
rect 1714 -2009 1725 -1963
rect 1799 -2009 1810 -1963
rect 1714 -2040 1810 -2009
rect 1979 -2140 2025 -2000
rect 2322 -2140 4290 -1156
rect -800 -2340 4290 -2140
<< via1 >>
rect 264 1193 269 1433
rect 269 1193 315 1433
rect 315 1193 320 1433
rect 1356 1193 1361 1433
rect 1361 1193 1407 1433
rect 1407 1193 1412 1433
rect 366 920 422 976
rect 1836 1193 1841 1433
rect 1841 1193 1887 1433
rect 1887 1193 1892 1433
rect 1658 842 1714 898
rect 1178 764 1234 820
rect -426 -227 -421 13
rect -421 -227 -375 13
rect -375 -227 -370 13
rect 468 482 473 538
rect 473 482 519 538
rect 519 482 524 538
rect 948 482 953 538
rect 953 482 999 538
rect 999 482 1004 538
rect 1152 482 1157 538
rect 1157 482 1203 538
rect 1203 482 1208 538
rect 1356 482 1361 538
rect 1361 482 1407 538
rect 1407 482 1412 538
rect 2422 804 4190 944
rect 1836 482 1841 538
rect 1841 482 1887 538
rect 1887 482 1892 538
rect 1362 30 1962 170
rect 2696 301 2701 541
rect 2701 301 2747 541
rect 2747 301 2752 541
rect 3380 301 3385 541
rect 3385 301 3431 541
rect 3431 301 3436 541
rect 3176 -33 3181 207
rect 3181 -33 3227 207
rect 3227 -33 3232 207
rect 3584 -33 3589 207
rect 3589 -33 3635 207
rect 3635 -33 3640 207
rect 4064 17 4069 257
rect 4069 17 4115 257
rect 4115 17 4120 257
rect 1362 -370 1962 -230
rect 2594 -256 2650 -200
rect -604 -578 -548 -522
rect -426 -938 -421 -882
rect -421 -938 -375 -882
rect -375 -938 -370 -882
rect 264 -1147 269 -907
rect 269 -1147 315 -907
rect 315 -1147 320 -907
rect 1356 -1147 1361 -907
rect 1361 -1147 1407 -907
rect 1407 -1147 1412 -907
rect 366 -1420 422 -1364
rect 1836 -1147 1841 -907
rect 1841 -1147 1887 -907
rect 1887 -1147 1892 -907
rect 3886 -334 3942 -278
rect 3278 -412 3334 -356
rect 2492 -694 2497 -638
rect 2497 -694 2543 -638
rect 2543 -694 2548 -638
rect 3380 -694 3385 -638
rect 3385 -694 3431 -638
rect 3431 -694 3436 -638
rect 4064 -694 4069 -638
rect 4069 -694 4115 -638
rect 4115 -694 4120 -638
rect 2422 -1156 4190 -1016
rect 1658 -1498 1714 -1442
rect 1178 -1576 1234 -1520
rect 468 -1858 473 -1802
rect 473 -1858 519 -1802
rect 519 -1858 524 -1802
rect 948 -1858 953 -1802
rect 953 -1858 999 -1802
rect 999 -1858 1004 -1802
rect 1152 -1858 1157 -1802
rect 1157 -1858 1203 -1802
rect 1203 -1858 1208 -1802
rect 1356 -1858 1361 -1802
rect 1361 -1858 1407 -1802
rect 1407 -1858 1412 -1802
rect 1836 -1858 1841 -1802
rect 1841 -1858 1887 -1802
rect 1887 -1858 1892 -1802
<< metal2 >>
rect 252 1433 1424 1443
rect 252 1193 264 1433
rect 320 1193 1356 1433
rect 1412 1193 1424 1433
rect 252 1183 1424 1193
rect 346 976 424 988
rect -1024 920 366 976
rect 422 920 424 976
rect 346 908 424 920
rect 1344 898 1424 1183
rect 1824 1433 1904 1443
rect 1824 1193 1836 1433
rect 1892 1193 1904 1433
rect 1646 898 1716 910
rect 1344 842 1658 898
rect 1714 842 1716 898
rect 1166 820 1236 832
rect -1024 764 1178 820
rect 1234 764 1236 820
rect -912 -522 -856 764
rect 1166 752 1236 764
rect 456 538 536 548
rect 456 482 468 538
rect 524 482 536 538
rect 456 296 536 482
rect 936 538 1016 548
rect 936 482 948 538
rect 1004 482 1016 538
rect 936 472 1016 482
rect 1140 538 1220 548
rect 1140 482 1152 538
rect 1208 482 1220 538
rect 1140 296 1220 482
rect 1344 538 1424 842
rect 1646 830 1716 842
rect 1824 898 1904 1193
rect 2410 944 4202 956
rect 1824 842 2181 898
rect 1344 482 1356 538
rect 1412 482 1424 538
rect 1344 472 1424 482
rect 1824 538 1904 842
rect 1824 482 1836 538
rect 1892 482 1904 538
rect 1824 472 1904 482
rect 456 224 1220 296
rect 1350 170 1974 182
rect 1350 30 1362 170
rect 1962 30 1974 170
rect -438 13 -358 23
rect 1350 18 1974 30
rect -438 -227 -426 13
rect -370 -227 -358 13
rect 2125 -200 2181 842
rect 2410 804 2422 944
rect 4190 804 4202 944
rect 2410 792 4202 804
rect 2684 541 3448 551
rect 2684 301 2696 541
rect 2752 301 3380 541
rect 3436 301 3448 541
rect 2684 291 3448 301
rect 4052 257 4132 267
rect 3164 207 3652 217
rect 3164 -33 3176 207
rect 3232 -33 3584 207
rect 3640 -33 3652 207
rect 3164 -43 3652 -33
rect 2574 -200 2670 -188
rect -616 -522 -546 -510
rect -912 -578 -604 -522
rect -548 -578 -546 -522
rect -616 -590 -546 -578
rect -438 -522 -358 -227
rect 1350 -230 1974 -218
rect 1350 -370 1362 -230
rect 1962 -370 1974 -230
rect 2125 -256 2594 -200
rect 2650 -256 2670 -200
rect 2574 -268 2670 -256
rect 3572 -278 3652 -43
rect 4052 17 4064 257
rect 4120 17 4132 257
rect 3874 -278 3944 -266
rect 3572 -334 3886 -278
rect 3942 -334 3944 -278
rect 3258 -356 3354 -346
rect 1350 -382 1974 -370
rect 2125 -412 3278 -356
rect 3334 -412 3354 -356
rect -438 -578 0 -522
rect -438 -882 -358 -578
rect -438 -938 -426 -882
rect -370 -938 -358 -882
rect -438 -948 -358 -938
rect -56 -1364 0 -578
rect 252 -907 1424 -897
rect 252 -1147 264 -907
rect 320 -1147 1356 -907
rect 1412 -1147 1424 -907
rect 252 -1157 1424 -1147
rect 346 -1364 424 -1352
rect -56 -1420 366 -1364
rect 422 -1420 424 -1364
rect 346 -1432 424 -1420
rect 1344 -1442 1424 -1157
rect 1824 -907 1904 -897
rect 1824 -1147 1836 -907
rect 1892 -1147 1904 -907
rect 1646 -1442 1716 -1430
rect 1344 -1498 1658 -1442
rect 1714 -1498 1716 -1442
rect 1166 -1520 1236 -1508
rect -1024 -1576 1178 -1520
rect 1234 -1576 1236 -1520
rect 1166 -1588 1236 -1576
rect 456 -1802 536 -1792
rect 456 -1858 468 -1802
rect 524 -1858 536 -1802
rect 456 -2044 536 -1858
rect 936 -1802 1016 -1792
rect 936 -1858 948 -1802
rect 1004 -1858 1016 -1802
rect 936 -1868 1016 -1858
rect 1140 -1802 1220 -1792
rect 1140 -1858 1152 -1802
rect 1208 -1858 1220 -1802
rect 1140 -2044 1220 -1858
rect 1344 -1802 1424 -1498
rect 1646 -1510 1716 -1498
rect 1824 -1442 1904 -1147
rect 2125 -1442 2181 -412
rect 3258 -422 3354 -412
rect 3572 -628 3652 -334
rect 3874 -346 3944 -334
rect 4052 -278 4132 17
rect 4052 -334 4350 -278
rect 2480 -638 3652 -628
rect 2480 -694 2492 -638
rect 2548 -694 3380 -638
rect 3436 -694 3652 -638
rect 2480 -704 3652 -694
rect 4052 -638 4132 -334
rect 4052 -694 4064 -638
rect 4120 -694 4132 -638
rect 4052 -704 4132 -694
rect 2410 -1016 4202 -1004
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
rect 1824 -1498 2181 -1442
rect 1344 -1858 1356 -1802
rect 1412 -1858 1424 -1802
rect 1344 -1868 1424 -1858
rect 1824 -1802 1904 -1498
rect 1824 -1858 1836 -1802
rect 1892 -1858 1904 -1802
rect 1824 -1868 1904 -1858
rect 456 -2116 1220 -2044
<< via2 >>
rect 948 482 1004 538
rect 1356 482 1412 538
rect 1362 30 1962 170
rect 2422 804 4190 944
rect 1362 -370 1962 -230
rect 948 -1858 1004 -1802
rect 2422 -1156 4190 -1016
rect 1356 -1858 1412 -1802
<< metal3 >>
rect 2410 944 4202 956
rect 2410 804 2422 944
rect 4190 804 4202 944
rect 936 538 1424 548
rect 936 482 948 538
rect 1004 482 1356 538
rect 1412 482 1424 538
rect 936 472 1424 482
rect 1350 170 1974 182
rect 1350 30 1362 170
rect 1962 30 1974 170
rect 1350 18 1974 30
rect 2410 -218 4202 804
rect 1350 -230 4202 -218
rect 1350 -370 1362 -230
rect 1962 -370 4202 -230
rect 1350 -382 4202 -370
rect 2410 -1016 4202 -1004
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
rect 936 -1802 1424 -1792
rect 936 -1858 948 -1802
rect 1004 -1858 1356 -1802
rect 1412 -1858 1424 -1802
rect 936 -1868 1424 -1858
<< via3 >>
rect 1362 30 1962 170
rect 2422 -1156 4190 -1016
<< metal4 >>
rect 1350 170 4202 182
rect 1350 30 1362 170
rect 1962 30 4202 170
rect 1350 18 4202 30
rect 2410 -1016 4202 18
rect 2410 -1156 2422 -1016
rect 4190 -1156 4202 -1016
rect 2410 -1168 4202 -1156
<< labels >>
rlabel metal2 -1024 947 -1024 947 7 Bit
port 0 w
rlabel metal2 -1024 791 -1024 791 7 Load
port 1 w
rlabel metal1 -469 2140 -469 2140 1 VDD
port 2 n
rlabel metal2 4350 -306 4350 -306 3 OUT
port 3 e
rlabel metal1 -500 -2340 -500 -2340 5 VSS
port 4 s
rlabel metal2 -1024 -1549 -1024 -1549 7 In
port 5 w
<< end >>
