magic
tech gf180mcuD
magscale 1 10
timestamp 1758085300
<< nwell >>
rect -222 1780 726 2700
rect -222 -425 726 495
rect 1264 -425 2212 495
rect -222 -2630 726 -1710
rect 1264 -2629 2212 -1709
rect -222 -4835 726 -3915
<< pwell >>
rect 541 1540 609 1780
rect -222 920 726 1540
rect 541 -665 609 -425
rect 2027 -665 2095 -425
rect -222 -1285 726 -665
rect 1264 -1285 2212 -665
rect 541 -2870 609 -2630
rect 2027 -2869 2095 -2629
rect -222 -3490 726 -2870
rect 1264 -3489 2212 -2869
rect 541 -5075 609 -4835
rect -222 -5695 726 -5075
<< nmos >>
rect 28 1130 108 1330
rect 212 1130 292 1330
rect 396 1130 476 1330
rect 28 -1075 108 -875
rect 212 -1075 292 -875
rect 396 -1075 476 -875
rect 1514 -1075 1594 -875
rect 1698 -1075 1778 -875
rect 1882 -1075 1962 -875
rect 28 -3280 108 -3080
rect 212 -3280 292 -3080
rect 396 -3280 476 -3080
rect 1514 -3279 1594 -3079
rect 1698 -3279 1778 -3079
rect 1882 -3279 1962 -3079
rect 28 -5485 108 -5285
rect 212 -5485 292 -5285
rect 396 -5485 476 -5285
<< pmos >>
rect 28 1990 108 2490
rect 212 1990 292 2490
rect 396 1990 476 2490
rect 28 -215 108 285
rect 212 -215 292 285
rect 396 -215 476 285
rect 1514 -215 1594 285
rect 1698 -215 1778 285
rect 1882 -215 1962 285
rect 28 -2420 108 -1920
rect 212 -2420 292 -1920
rect 396 -2420 476 -1920
rect 1514 -2419 1594 -1919
rect 1698 -2419 1778 -1919
rect 1882 -2419 1962 -1919
rect 28 -4625 108 -4125
rect 212 -4625 292 -4125
rect 396 -4625 476 -4125
<< ndiff >>
rect -60 1317 28 1330
rect -60 1143 -47 1317
rect -1 1143 28 1317
rect -60 1130 28 1143
rect 108 1317 212 1330
rect 108 1143 137 1317
rect 183 1143 212 1317
rect 108 1130 212 1143
rect 292 1317 396 1330
rect 292 1143 321 1317
rect 367 1143 396 1317
rect 292 1130 396 1143
rect 476 1317 564 1330
rect 476 1143 505 1317
rect 551 1143 564 1317
rect 476 1130 564 1143
rect -60 -888 28 -875
rect -60 -1062 -47 -888
rect -1 -1062 28 -888
rect -60 -1075 28 -1062
rect 108 -888 212 -875
rect 108 -1062 137 -888
rect 183 -1062 212 -888
rect 108 -1075 212 -1062
rect 292 -888 396 -875
rect 292 -1062 321 -888
rect 367 -1062 396 -888
rect 292 -1075 396 -1062
rect 476 -888 564 -875
rect 476 -1062 505 -888
rect 551 -1062 564 -888
rect 476 -1075 564 -1062
rect 1426 -888 1514 -875
rect 1426 -1062 1439 -888
rect 1485 -1062 1514 -888
rect 1426 -1075 1514 -1062
rect 1594 -888 1698 -875
rect 1594 -1062 1623 -888
rect 1669 -1062 1698 -888
rect 1594 -1075 1698 -1062
rect 1778 -888 1882 -875
rect 1778 -1062 1807 -888
rect 1853 -1062 1882 -888
rect 1778 -1075 1882 -1062
rect 1962 -888 2050 -875
rect 1962 -1062 1991 -888
rect 2037 -1062 2050 -888
rect 1962 -1075 2050 -1062
rect -60 -3093 28 -3080
rect -60 -3267 -47 -3093
rect -1 -3267 28 -3093
rect -60 -3280 28 -3267
rect 108 -3093 212 -3080
rect 108 -3267 137 -3093
rect 183 -3267 212 -3093
rect 108 -3280 212 -3267
rect 292 -3093 396 -3080
rect 292 -3267 321 -3093
rect 367 -3267 396 -3093
rect 292 -3280 396 -3267
rect 476 -3093 564 -3080
rect 476 -3267 505 -3093
rect 551 -3267 564 -3093
rect 476 -3280 564 -3267
rect 1426 -3092 1514 -3079
rect 1426 -3266 1439 -3092
rect 1485 -3266 1514 -3092
rect 1426 -3279 1514 -3266
rect 1594 -3092 1698 -3079
rect 1594 -3266 1623 -3092
rect 1669 -3266 1698 -3092
rect 1594 -3279 1698 -3266
rect 1778 -3092 1882 -3079
rect 1778 -3266 1807 -3092
rect 1853 -3266 1882 -3092
rect 1778 -3279 1882 -3266
rect 1962 -3092 2050 -3079
rect 1962 -3266 1991 -3092
rect 2037 -3266 2050 -3092
rect 1962 -3279 2050 -3266
rect -60 -5298 28 -5285
rect -60 -5472 -47 -5298
rect -1 -5472 28 -5298
rect -60 -5485 28 -5472
rect 108 -5298 212 -5285
rect 108 -5472 137 -5298
rect 183 -5472 212 -5298
rect 108 -5485 212 -5472
rect 292 -5298 396 -5285
rect 292 -5472 321 -5298
rect 367 -5472 396 -5298
rect 292 -5485 396 -5472
rect 476 -5298 564 -5285
rect 476 -5472 505 -5298
rect 551 -5472 564 -5298
rect 476 -5485 564 -5472
<< pdiff >>
rect -60 2477 28 2490
rect -60 2003 -47 2477
rect -1 2003 28 2477
rect -60 1990 28 2003
rect 108 2477 212 2490
rect 108 2003 137 2477
rect 183 2003 212 2477
rect 108 1990 212 2003
rect 292 2477 396 2490
rect 292 2003 321 2477
rect 367 2003 396 2477
rect 292 1990 396 2003
rect 476 2477 564 2490
rect 476 2003 505 2477
rect 551 2003 564 2477
rect 476 1990 564 2003
rect -60 272 28 285
rect -60 -202 -47 272
rect -1 -202 28 272
rect -60 -215 28 -202
rect 108 272 212 285
rect 108 -202 137 272
rect 183 -202 212 272
rect 108 -215 212 -202
rect 292 272 396 285
rect 292 -202 321 272
rect 367 -202 396 272
rect 292 -215 396 -202
rect 476 272 564 285
rect 476 -202 505 272
rect 551 -202 564 272
rect 476 -215 564 -202
rect 1426 272 1514 285
rect 1426 -202 1439 272
rect 1485 -202 1514 272
rect 1426 -215 1514 -202
rect 1594 272 1698 285
rect 1594 -202 1623 272
rect 1669 -202 1698 272
rect 1594 -215 1698 -202
rect 1778 272 1882 285
rect 1778 -202 1807 272
rect 1853 -202 1882 272
rect 1778 -215 1882 -202
rect 1962 272 2050 285
rect 1962 -202 1991 272
rect 2037 -202 2050 272
rect 1962 -215 2050 -202
rect -60 -1933 28 -1920
rect -60 -2407 -47 -1933
rect -1 -2407 28 -1933
rect -60 -2420 28 -2407
rect 108 -1933 212 -1920
rect 108 -2407 137 -1933
rect 183 -2407 212 -1933
rect 108 -2420 212 -2407
rect 292 -1933 396 -1920
rect 292 -2407 321 -1933
rect 367 -2407 396 -1933
rect 292 -2420 396 -2407
rect 476 -1933 564 -1920
rect 476 -2407 505 -1933
rect 551 -2407 564 -1933
rect 476 -2420 564 -2407
rect 1426 -1932 1514 -1919
rect 1426 -2406 1439 -1932
rect 1485 -2406 1514 -1932
rect 1426 -2419 1514 -2406
rect 1594 -1932 1698 -1919
rect 1594 -2406 1623 -1932
rect 1669 -2406 1698 -1932
rect 1594 -2419 1698 -2406
rect 1778 -1932 1882 -1919
rect 1778 -2406 1807 -1932
rect 1853 -2406 1882 -1932
rect 1778 -2419 1882 -2406
rect 1962 -1932 2050 -1919
rect 1962 -2406 1991 -1932
rect 2037 -2406 2050 -1932
rect 1962 -2419 2050 -2406
rect -60 -4138 28 -4125
rect -60 -4612 -47 -4138
rect -1 -4612 28 -4138
rect -60 -4625 28 -4612
rect 108 -4138 212 -4125
rect 108 -4612 137 -4138
rect 183 -4612 212 -4138
rect 108 -4625 212 -4612
rect 292 -4138 396 -4125
rect 292 -4612 321 -4138
rect 367 -4612 396 -4138
rect 292 -4625 396 -4612
rect 476 -4138 564 -4125
rect 476 -4612 505 -4138
rect 551 -4612 564 -4138
rect 476 -4625 564 -4612
<< ndiffc >>
rect -47 1143 -1 1317
rect 137 1143 183 1317
rect 321 1143 367 1317
rect 505 1143 551 1317
rect -47 -1062 -1 -888
rect 137 -1062 183 -888
rect 321 -1062 367 -888
rect 505 -1062 551 -888
rect 1439 -1062 1485 -888
rect 1623 -1062 1669 -888
rect 1807 -1062 1853 -888
rect 1991 -1062 2037 -888
rect -47 -3267 -1 -3093
rect 137 -3267 183 -3093
rect 321 -3267 367 -3093
rect 505 -3267 551 -3093
rect 1439 -3266 1485 -3092
rect 1623 -3266 1669 -3092
rect 1807 -3266 1853 -3092
rect 1991 -3266 2037 -3092
rect -47 -5472 -1 -5298
rect 137 -5472 183 -5298
rect 321 -5472 367 -5298
rect 505 -5472 551 -5298
<< pdiffc >>
rect -47 2003 -1 2477
rect 137 2003 183 2477
rect 321 2003 367 2477
rect 505 2003 551 2477
rect -47 -202 -1 272
rect 137 -202 183 272
rect 321 -202 367 272
rect 505 -202 551 272
rect 1439 -202 1485 272
rect 1623 -202 1669 272
rect 1807 -202 1853 272
rect 1991 -202 2037 272
rect -47 -2407 -1 -1933
rect 137 -2407 183 -1933
rect 321 -2407 367 -1933
rect 505 -2407 551 -1933
rect 1439 -2406 1485 -1932
rect 1623 -2406 1669 -1932
rect 1807 -2406 1853 -1932
rect 1991 -2406 2037 -1932
rect -47 -4612 -1 -4138
rect 137 -4612 183 -4138
rect 321 -4612 367 -4138
rect 505 -4612 551 -4138
<< psubdiff >>
rect -198 1444 702 1516
rect -198 1400 -126 1444
rect -198 1060 -185 1400
rect -139 1060 -126 1400
rect 630 1400 702 1444
rect -198 1016 -126 1060
rect 630 1060 643 1400
rect 689 1060 702 1400
rect 630 1016 702 1060
rect -198 944 702 1016
rect -198 -761 702 -689
rect -198 -805 -126 -761
rect -198 -1145 -185 -805
rect -139 -1145 -126 -805
rect 630 -805 702 -761
rect -198 -1189 -126 -1145
rect 630 -1145 643 -805
rect 689 -1145 702 -805
rect 630 -1189 702 -1145
rect -198 -1261 702 -1189
rect 1288 -761 2188 -689
rect 1288 -805 1360 -761
rect 1288 -1145 1301 -805
rect 1347 -1145 1360 -805
rect 2116 -805 2188 -761
rect 1288 -1189 1360 -1145
rect 2116 -1145 2129 -805
rect 2175 -1145 2188 -805
rect 2116 -1189 2188 -1145
rect 1288 -1261 2188 -1189
rect -198 -2966 702 -2894
rect -198 -3010 -126 -2966
rect -198 -3350 -185 -3010
rect -139 -3350 -126 -3010
rect 630 -3010 702 -2966
rect -198 -3394 -126 -3350
rect 630 -3350 643 -3010
rect 689 -3350 702 -3010
rect 630 -3394 702 -3350
rect -198 -3466 702 -3394
rect 1288 -2965 2188 -2893
rect 1288 -3009 1360 -2965
rect 1288 -3349 1301 -3009
rect 1347 -3349 1360 -3009
rect 2116 -3009 2188 -2965
rect 1288 -3393 1360 -3349
rect 2116 -3349 2129 -3009
rect 2175 -3349 2188 -3009
rect 2116 -3393 2188 -3349
rect 1288 -3465 2188 -3393
rect -198 -5171 702 -5099
rect -198 -5215 -126 -5171
rect -198 -5555 -185 -5215
rect -139 -5555 -126 -5215
rect 630 -5215 702 -5171
rect -198 -5599 -126 -5555
rect 630 -5555 643 -5215
rect 689 -5555 702 -5215
rect 630 -5599 702 -5555
rect -198 -5671 702 -5599
<< nsubdiff >>
rect -198 2604 702 2676
rect -198 2560 -126 2604
rect -198 1920 -185 2560
rect -139 1920 -126 2560
rect 630 2560 702 2604
rect -198 1876 -126 1920
rect 630 1920 643 2560
rect 689 1920 702 2560
rect 630 1876 702 1920
rect -198 1804 702 1876
rect -198 399 702 471
rect -198 355 -126 399
rect -198 -285 -185 355
rect -139 -285 -126 355
rect 630 355 702 399
rect -198 -329 -126 -285
rect 630 -285 643 355
rect 689 -285 702 355
rect 630 -329 702 -285
rect -198 -401 702 -329
rect 1288 399 2188 471
rect 1288 355 1360 399
rect 1288 -285 1301 355
rect 1347 -285 1360 355
rect 2116 355 2188 399
rect 1288 -329 1360 -285
rect 2116 -285 2129 355
rect 2175 -285 2188 355
rect 2116 -329 2188 -285
rect 1288 -401 2188 -329
rect -198 -1806 702 -1734
rect -198 -1850 -126 -1806
rect -198 -2490 -185 -1850
rect -139 -2490 -126 -1850
rect 630 -1850 702 -1806
rect -198 -2534 -126 -2490
rect 630 -2490 643 -1850
rect 689 -2490 702 -1850
rect 630 -2534 702 -2490
rect -198 -2606 702 -2534
rect 1288 -1805 2188 -1733
rect 1288 -1849 1360 -1805
rect 1288 -2489 1301 -1849
rect 1347 -2489 1360 -1849
rect 2116 -1849 2188 -1805
rect 1288 -2533 1360 -2489
rect 2116 -2489 2129 -1849
rect 2175 -2489 2188 -1849
rect 2116 -2533 2188 -2489
rect 1288 -2605 2188 -2533
rect -198 -4011 702 -3939
rect -198 -4055 -126 -4011
rect -198 -4695 -185 -4055
rect -139 -4695 -126 -4055
rect 630 -4055 702 -4011
rect -198 -4739 -126 -4695
rect 630 -4695 643 -4055
rect 689 -4695 702 -4055
rect 630 -4739 702 -4695
rect -198 -4811 702 -4739
<< psubdiffcont >>
rect -185 1060 -139 1400
rect 643 1060 689 1400
rect -185 -1145 -139 -805
rect 643 -1145 689 -805
rect 1301 -1145 1347 -805
rect 2129 -1145 2175 -805
rect -185 -3350 -139 -3010
rect 643 -3350 689 -3010
rect 1301 -3349 1347 -3009
rect 2129 -3349 2175 -3009
rect -185 -5555 -139 -5215
rect 643 -5555 689 -5215
<< nsubdiffcont >>
rect -185 1920 -139 2560
rect 643 1920 689 2560
rect -185 -285 -139 355
rect 643 -285 689 355
rect 1301 -285 1347 355
rect 2129 -285 2175 355
rect -185 -2490 -139 -1850
rect 643 -2490 689 -1850
rect 1301 -2489 1347 -1849
rect 2129 -2489 2175 -1849
rect -185 -4695 -139 -4055
rect 643 -4695 689 -4055
<< polysilicon >>
rect 28 2569 108 2582
rect 28 2523 41 2569
rect 95 2523 108 2569
rect 28 2490 108 2523
rect 212 2569 292 2582
rect 212 2523 225 2569
rect 279 2523 292 2569
rect 212 2490 292 2523
rect 396 2569 476 2582
rect 396 2523 409 2569
rect 463 2523 476 2569
rect 396 2490 476 2523
rect 28 1957 108 1990
rect 28 1911 41 1957
rect 95 1911 108 1957
rect 28 1898 108 1911
rect 212 1957 292 1990
rect 212 1911 225 1957
rect 279 1911 292 1957
rect 212 1898 292 1911
rect 396 1957 476 1990
rect 396 1911 409 1957
rect 463 1911 476 1957
rect 396 1898 476 1911
rect 28 1409 108 1422
rect 28 1363 41 1409
rect 95 1363 108 1409
rect 28 1330 108 1363
rect 212 1409 292 1422
rect 212 1363 225 1409
rect 279 1363 292 1409
rect 212 1330 292 1363
rect 396 1409 476 1422
rect 396 1363 409 1409
rect 463 1363 476 1409
rect 396 1330 476 1363
rect 28 1097 108 1130
rect 28 1051 41 1097
rect 95 1051 108 1097
rect 28 1038 108 1051
rect 212 1097 292 1130
rect 212 1051 225 1097
rect 279 1051 292 1097
rect 212 1038 292 1051
rect 396 1097 476 1130
rect 396 1051 409 1097
rect 463 1051 476 1097
rect 396 1038 476 1051
rect 28 364 108 377
rect 28 318 41 364
rect 95 318 108 364
rect 28 285 108 318
rect 212 364 292 377
rect 212 318 225 364
rect 279 318 292 364
rect 212 285 292 318
rect 396 364 476 377
rect 396 318 409 364
rect 463 318 476 364
rect 396 285 476 318
rect 28 -248 108 -215
rect 28 -294 41 -248
rect 95 -294 108 -248
rect 28 -307 108 -294
rect 212 -248 292 -215
rect 212 -294 225 -248
rect 279 -294 292 -248
rect 212 -307 292 -294
rect 396 -248 476 -215
rect 396 -294 409 -248
rect 463 -294 476 -248
rect 396 -307 476 -294
rect 1514 364 1594 377
rect 1514 318 1527 364
rect 1581 318 1594 364
rect 1514 285 1594 318
rect 1698 364 1778 377
rect 1698 318 1711 364
rect 1765 318 1778 364
rect 1698 285 1778 318
rect 1882 364 1962 377
rect 1882 318 1895 364
rect 1949 318 1962 364
rect 1882 285 1962 318
rect 1514 -248 1594 -215
rect 1514 -294 1527 -248
rect 1581 -294 1594 -248
rect 1514 -307 1594 -294
rect 1698 -248 1778 -215
rect 1698 -294 1711 -248
rect 1765 -294 1778 -248
rect 1698 -307 1778 -294
rect 1882 -248 1962 -215
rect 1882 -294 1895 -248
rect 1949 -294 1962 -248
rect 1882 -307 1962 -294
rect 28 -796 108 -783
rect 28 -842 41 -796
rect 95 -842 108 -796
rect 28 -875 108 -842
rect 212 -796 292 -783
rect 212 -842 225 -796
rect 279 -842 292 -796
rect 212 -875 292 -842
rect 396 -796 476 -783
rect 396 -842 409 -796
rect 463 -842 476 -796
rect 396 -875 476 -842
rect 28 -1108 108 -1075
rect 28 -1154 41 -1108
rect 95 -1154 108 -1108
rect 28 -1167 108 -1154
rect 212 -1108 292 -1075
rect 212 -1154 225 -1108
rect 279 -1154 292 -1108
rect 212 -1167 292 -1154
rect 396 -1108 476 -1075
rect 396 -1154 409 -1108
rect 463 -1154 476 -1108
rect 396 -1167 476 -1154
rect 1514 -796 1594 -783
rect 1514 -842 1527 -796
rect 1581 -842 1594 -796
rect 1514 -875 1594 -842
rect 1698 -796 1778 -783
rect 1698 -842 1711 -796
rect 1765 -842 1778 -796
rect 1698 -875 1778 -842
rect 1882 -796 1962 -783
rect 1882 -842 1895 -796
rect 1949 -842 1962 -796
rect 1882 -875 1962 -842
rect 1514 -1108 1594 -1075
rect 1514 -1154 1527 -1108
rect 1581 -1154 1594 -1108
rect 1514 -1167 1594 -1154
rect 1698 -1108 1778 -1075
rect 1698 -1154 1711 -1108
rect 1765 -1154 1778 -1108
rect 1698 -1167 1778 -1154
rect 1882 -1108 1962 -1075
rect 1882 -1154 1895 -1108
rect 1949 -1154 1962 -1108
rect 1882 -1167 1962 -1154
rect 28 -1841 108 -1828
rect 28 -1887 41 -1841
rect 95 -1887 108 -1841
rect 28 -1920 108 -1887
rect 212 -1841 292 -1828
rect 212 -1887 225 -1841
rect 279 -1887 292 -1841
rect 212 -1920 292 -1887
rect 396 -1841 476 -1828
rect 396 -1887 409 -1841
rect 463 -1887 476 -1841
rect 396 -1920 476 -1887
rect 28 -2453 108 -2420
rect 28 -2499 41 -2453
rect 95 -2499 108 -2453
rect 28 -2512 108 -2499
rect 212 -2453 292 -2420
rect 212 -2499 225 -2453
rect 279 -2499 292 -2453
rect 212 -2512 292 -2499
rect 396 -2453 476 -2420
rect 396 -2499 409 -2453
rect 463 -2499 476 -2453
rect 396 -2512 476 -2499
rect 1514 -1840 1594 -1827
rect 1514 -1886 1527 -1840
rect 1581 -1886 1594 -1840
rect 1514 -1919 1594 -1886
rect 1698 -1840 1778 -1827
rect 1698 -1886 1711 -1840
rect 1765 -1886 1778 -1840
rect 1698 -1919 1778 -1886
rect 1882 -1840 1962 -1827
rect 1882 -1886 1895 -1840
rect 1949 -1886 1962 -1840
rect 1882 -1919 1962 -1886
rect 1514 -2452 1594 -2419
rect 1514 -2498 1527 -2452
rect 1581 -2498 1594 -2452
rect 1514 -2511 1594 -2498
rect 1698 -2452 1778 -2419
rect 1698 -2498 1711 -2452
rect 1765 -2498 1778 -2452
rect 1698 -2511 1778 -2498
rect 1882 -2452 1962 -2419
rect 1882 -2498 1895 -2452
rect 1949 -2498 1962 -2452
rect 1882 -2511 1962 -2498
rect 28 -3001 108 -2988
rect 28 -3047 41 -3001
rect 95 -3047 108 -3001
rect 28 -3080 108 -3047
rect 212 -3001 292 -2988
rect 212 -3047 225 -3001
rect 279 -3047 292 -3001
rect 212 -3080 292 -3047
rect 396 -3001 476 -2988
rect 396 -3047 409 -3001
rect 463 -3047 476 -3001
rect 396 -3080 476 -3047
rect 28 -3313 108 -3280
rect 28 -3359 41 -3313
rect 95 -3359 108 -3313
rect 28 -3372 108 -3359
rect 212 -3313 292 -3280
rect 212 -3359 225 -3313
rect 279 -3359 292 -3313
rect 212 -3372 292 -3359
rect 396 -3313 476 -3280
rect 396 -3359 409 -3313
rect 463 -3359 476 -3313
rect 396 -3372 476 -3359
rect 1514 -3000 1594 -2987
rect 1514 -3046 1527 -3000
rect 1581 -3046 1594 -3000
rect 1514 -3079 1594 -3046
rect 1698 -3000 1778 -2987
rect 1698 -3046 1711 -3000
rect 1765 -3046 1778 -3000
rect 1698 -3079 1778 -3046
rect 1882 -3000 1962 -2987
rect 1882 -3046 1895 -3000
rect 1949 -3046 1962 -3000
rect 1882 -3079 1962 -3046
rect 1514 -3312 1594 -3279
rect 1514 -3358 1527 -3312
rect 1581 -3358 1594 -3312
rect 1514 -3371 1594 -3358
rect 1698 -3312 1778 -3279
rect 1698 -3358 1711 -3312
rect 1765 -3358 1778 -3312
rect 1698 -3371 1778 -3358
rect 1882 -3312 1962 -3279
rect 1882 -3358 1895 -3312
rect 1949 -3358 1962 -3312
rect 1882 -3371 1962 -3358
rect 28 -4046 108 -4033
rect 28 -4092 41 -4046
rect 95 -4092 108 -4046
rect 28 -4125 108 -4092
rect 212 -4046 292 -4033
rect 212 -4092 225 -4046
rect 279 -4092 292 -4046
rect 212 -4125 292 -4092
rect 396 -4046 476 -4033
rect 396 -4092 409 -4046
rect 463 -4092 476 -4046
rect 396 -4125 476 -4092
rect 28 -4658 108 -4625
rect 28 -4704 41 -4658
rect 95 -4704 108 -4658
rect 28 -4717 108 -4704
rect 212 -4658 292 -4625
rect 212 -4704 225 -4658
rect 279 -4704 292 -4658
rect 212 -4717 292 -4704
rect 396 -4658 476 -4625
rect 396 -4704 409 -4658
rect 463 -4704 476 -4658
rect 396 -4717 476 -4704
rect 28 -5206 108 -5193
rect 28 -5252 41 -5206
rect 95 -5252 108 -5206
rect 28 -5285 108 -5252
rect 212 -5206 292 -5193
rect 212 -5252 225 -5206
rect 279 -5252 292 -5206
rect 212 -5285 292 -5252
rect 396 -5206 476 -5193
rect 396 -5252 409 -5206
rect 463 -5252 476 -5206
rect 396 -5285 476 -5252
rect 28 -5518 108 -5485
rect 28 -5564 41 -5518
rect 95 -5564 108 -5518
rect 28 -5577 108 -5564
rect 212 -5518 292 -5485
rect 212 -5564 225 -5518
rect 279 -5564 292 -5518
rect 212 -5577 292 -5564
rect 396 -5518 476 -5485
rect 396 -5564 409 -5518
rect 463 -5564 476 -5518
rect 396 -5577 476 -5564
<< polycontact >>
rect 41 2523 95 2569
rect 225 2523 279 2569
rect 409 2523 463 2569
rect 41 1911 95 1957
rect 225 1911 279 1957
rect 409 1911 463 1957
rect 41 1363 95 1409
rect 225 1363 279 1409
rect 409 1363 463 1409
rect 41 1051 95 1097
rect 225 1051 279 1097
rect 409 1051 463 1097
rect 41 318 95 364
rect 225 318 279 364
rect 409 318 463 364
rect 41 -294 95 -248
rect 225 -294 279 -248
rect 409 -294 463 -248
rect 1527 318 1581 364
rect 1711 318 1765 364
rect 1895 318 1949 364
rect 1527 -294 1581 -248
rect 1711 -294 1765 -248
rect 1895 -294 1949 -248
rect 41 -842 95 -796
rect 225 -842 279 -796
rect 409 -842 463 -796
rect 41 -1154 95 -1108
rect 225 -1154 279 -1108
rect 409 -1154 463 -1108
rect 1527 -842 1581 -796
rect 1711 -842 1765 -796
rect 1895 -842 1949 -796
rect 1527 -1154 1581 -1108
rect 1711 -1154 1765 -1108
rect 1895 -1154 1949 -1108
rect 41 -1887 95 -1841
rect 225 -1887 279 -1841
rect 409 -1887 463 -1841
rect 41 -2499 95 -2453
rect 225 -2499 279 -2453
rect 409 -2499 463 -2453
rect 1527 -1886 1581 -1840
rect 1711 -1886 1765 -1840
rect 1895 -1886 1949 -1840
rect 1527 -2498 1581 -2452
rect 1711 -2498 1765 -2452
rect 1895 -2498 1949 -2452
rect 41 -3047 95 -3001
rect 225 -3047 279 -3001
rect 409 -3047 463 -3001
rect 41 -3359 95 -3313
rect 225 -3359 279 -3313
rect 409 -3359 463 -3313
rect 1527 -3046 1581 -3000
rect 1711 -3046 1765 -3000
rect 1895 -3046 1949 -3000
rect 1527 -3358 1581 -3312
rect 1711 -3358 1765 -3312
rect 1895 -3358 1949 -3312
rect 41 -4092 95 -4046
rect 225 -4092 279 -4046
rect 409 -4092 463 -4046
rect 41 -4704 95 -4658
rect 225 -4704 279 -4658
rect 409 -4704 463 -4658
rect 41 -5252 95 -5206
rect 225 -5252 279 -5206
rect 409 -5252 463 -5206
rect 41 -5564 95 -5518
rect 225 -5564 279 -5518
rect 409 -5564 463 -5518
<< metal1 >>
rect -365 2825 1182 2881
rect -365 1804 -309 2825
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -185 2560 -139 2571
rect 30 2569 106 2602
rect 30 2523 41 2569
rect 95 2523 106 2569
rect 214 2569 290 2602
rect 214 2523 225 2569
rect 279 2523 290 2569
rect 398 2569 474 2602
rect 398 2523 409 2569
rect 463 2523 474 2569
rect 643 2560 689 2571
rect -47 2477 -1 2488
rect -64 2450 -47 2452
rect 137 2477 183 2488
rect -1 2450 16 2452
rect -139 2330 -52 2450
rect 4 2330 16 2450
rect -64 2328 -47 2330
rect -139 2030 -47 2150
rect -1 2328 16 2330
rect 120 2150 137 2152
rect 321 2477 367 2488
rect 304 2450 321 2452
rect 505 2477 551 2488
rect 367 2450 384 2452
rect 304 2330 316 2450
rect 372 2330 384 2450
rect 304 2328 321 2330
rect 183 2150 200 2152
rect 120 2030 132 2150
rect 188 2030 200 2150
rect 120 2028 137 2030
rect -47 1992 -1 2003
rect 183 2028 200 2030
rect 137 1992 183 2003
rect 367 2328 384 2330
rect 488 2150 505 2152
rect 626 2450 643 2452
rect 689 2450 706 2452
rect 626 2329 638 2450
rect 694 2329 706 2450
rect 626 2327 643 2329
rect 551 2150 568 2152
rect 488 2030 500 2150
rect 556 2030 568 2150
rect 488 2028 505 2030
rect 321 1992 367 2003
rect 551 2028 568 2030
rect 505 1992 551 2003
rect 30 1954 41 1957
rect 95 1954 106 1957
rect 214 1954 225 1957
rect 279 1954 290 1957
rect 398 1954 409 1957
rect 463 1954 474 1957
rect -185 1909 -139 1920
rect 28 1898 40 1954
rect 96 1898 108 1954
rect 28 1884 108 1898
rect 212 1898 224 1954
rect 280 1898 292 1954
rect 212 1884 292 1898
rect 396 1898 408 1954
rect 464 1898 476 1954
rect 689 2327 706 2329
rect 643 1909 689 1920
rect 396 1884 476 1898
rect 28 1804 108 1806
rect -848 1748 40 1804
rect 96 1748 108 1804
rect 28 1746 108 1748
rect -644 1688 -574 1700
rect 212 1688 292 1690
rect -644 1632 -632 1688
rect -576 1632 224 1688
rect 280 1632 292 1688
rect -644 1620 -574 1632
rect 212 1630 292 1632
rect 541 1688 621 1690
rect 808 1688 878 1700
rect 541 1632 553 1688
rect 609 1632 810 1688
rect 866 1632 878 1688
rect 541 1630 621 1632
rect 808 1622 878 1632
rect 396 1572 476 1574
rect -360 1516 408 1572
rect 464 1516 476 1572
rect -360 785 -304 1516
rect 396 1514 476 1516
rect 28 1422 108 1436
rect -185 1400 -139 1411
rect 28 1366 40 1422
rect 96 1366 108 1422
rect 212 1422 292 1436
rect 212 1366 224 1422
rect 280 1366 292 1422
rect 396 1422 476 1436
rect 396 1366 408 1422
rect 464 1366 476 1422
rect 643 1400 689 1411
rect 30 1363 41 1366
rect 95 1363 106 1366
rect 214 1363 225 1366
rect 279 1363 290 1366
rect 398 1363 409 1366
rect 463 1363 474 1366
rect -47 1317 -1 1328
rect -139 1143 -47 1317
rect -47 1132 -1 1143
rect 137 1317 183 1328
rect 137 1132 183 1143
rect 321 1317 367 1328
rect 505 1317 551 1328
rect 488 1290 505 1292
rect 551 1290 568 1292
rect 488 1170 500 1290
rect 556 1170 568 1290
rect 488 1168 505 1170
rect 321 1132 367 1143
rect 551 1168 568 1170
rect 505 1132 551 1143
rect -185 915 -139 1060
rect 30 1051 41 1097
rect 95 1051 106 1097
rect 30 1018 106 1051
rect 214 1051 225 1097
rect 279 1051 290 1097
rect 214 1018 290 1051
rect 398 1051 409 1097
rect 463 1051 474 1097
rect 398 1018 474 1051
rect 643 915 689 1060
rect -197 903 -117 915
rect -197 847 -185 903
rect -129 847 -117 903
rect -197 835 -117 847
rect 621 903 701 915
rect 621 847 633 903
rect 689 847 701 903
rect 621 835 701 847
rect 974 785 1054 795
rect -360 729 986 785
rect 1042 729 1054 785
rect 974 727 1054 729
rect 808 676 878 678
rect -360 675 878 676
rect -360 621 810 675
rect 866 621 878 675
rect -360 620 878 621
rect -360 -401 -304 620
rect 808 612 878 620
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect -185 355 -139 366
rect 30 364 106 397
rect 30 318 41 364
rect 95 318 106 364
rect 214 364 290 397
rect 214 318 225 364
rect 279 318 290 364
rect 398 364 474 397
rect 398 318 409 364
rect 463 318 474 364
rect 643 355 689 366
rect -47 272 -1 283
rect -64 245 -47 247
rect 137 272 183 283
rect -1 245 16 247
rect -139 125 -52 245
rect 4 125 16 245
rect -64 123 -47 125
rect -139 -175 -47 -55
rect -1 123 16 125
rect 120 -55 137 -53
rect 321 272 367 283
rect 304 245 321 247
rect 505 272 551 283
rect 367 245 384 247
rect 304 125 316 245
rect 372 125 384 245
rect 304 123 321 125
rect 183 -55 200 -53
rect 120 -175 132 -55
rect 188 -175 200 -55
rect 120 -177 137 -175
rect -47 -213 -1 -202
rect 183 -177 200 -175
rect 137 -213 183 -202
rect 367 123 384 125
rect 488 -55 505 -53
rect 626 245 643 247
rect 689 245 706 247
rect 626 124 638 245
rect 694 124 706 245
rect 626 122 643 124
rect 551 -55 568 -53
rect 488 -175 500 -55
rect 556 -175 568 -55
rect 488 -177 505 -175
rect 321 -213 367 -202
rect 551 -177 568 -175
rect 505 -213 551 -202
rect 30 -251 41 -248
rect 95 -251 106 -248
rect 214 -251 225 -248
rect 279 -251 290 -248
rect 398 -251 409 -248
rect 463 -251 474 -248
rect -185 -296 -139 -285
rect 28 -307 40 -251
rect 96 -307 108 -251
rect 28 -321 108 -307
rect 212 -307 224 -251
rect 280 -307 292 -251
rect 212 -321 292 -307
rect 396 -307 408 -251
rect 464 -307 476 -251
rect 689 122 706 124
rect 643 -296 689 -285
rect 396 -321 476 -307
rect 28 -401 108 -399
rect -360 -457 40 -401
rect 96 -457 108 -401
rect 1126 -401 1182 2825
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect 1301 355 1347 366
rect 1516 364 1592 397
rect 1516 318 1527 364
rect 1581 318 1592 364
rect 1700 364 1776 397
rect 1700 318 1711 364
rect 1765 318 1776 364
rect 1884 364 1960 397
rect 1884 318 1895 364
rect 1949 318 1960 364
rect 2129 355 2175 366
rect 1439 272 1485 283
rect 1422 245 1439 247
rect 1623 272 1669 283
rect 1485 245 1502 247
rect 1347 125 1434 245
rect 1490 125 1502 245
rect 1422 123 1439 125
rect 1347 -175 1439 -55
rect 1485 123 1502 125
rect 1606 -55 1623 -53
rect 1807 272 1853 283
rect 1790 245 1807 247
rect 1991 272 2037 283
rect 1853 245 1870 247
rect 1790 125 1802 245
rect 1858 125 1870 245
rect 1790 123 1807 125
rect 1669 -55 1686 -53
rect 1606 -175 1618 -55
rect 1674 -175 1686 -55
rect 1606 -177 1623 -175
rect 1439 -213 1485 -202
rect 1669 -177 1686 -175
rect 1623 -213 1669 -202
rect 1853 123 1870 125
rect 1974 -55 1991 -53
rect 2112 245 2129 247
rect 2175 245 2192 247
rect 2112 124 2124 245
rect 2180 124 2192 245
rect 2112 122 2129 124
rect 2037 -55 2054 -53
rect 1974 -175 1986 -55
rect 2042 -175 2054 -55
rect 1974 -177 1991 -175
rect 1807 -213 1853 -202
rect 2037 -177 2054 -175
rect 1991 -213 2037 -202
rect 1516 -251 1527 -248
rect 1581 -251 1592 -248
rect 1700 -251 1711 -248
rect 1765 -251 1776 -248
rect 1884 -251 1895 -248
rect 1949 -251 1960 -248
rect 1301 -296 1347 -285
rect 1514 -307 1526 -251
rect 1582 -307 1594 -251
rect 1514 -321 1594 -307
rect 1698 -307 1710 -251
rect 1766 -307 1778 -251
rect 1698 -321 1778 -307
rect 1882 -307 1894 -251
rect 1950 -307 1962 -251
rect 2175 122 2192 124
rect 2129 -296 2175 -285
rect 1882 -321 1962 -307
rect 1514 -401 1594 -399
rect 1126 -457 1526 -401
rect 1582 -457 1594 -401
rect 28 -459 108 -457
rect 1514 -459 1594 -457
rect -780 -517 -710 -503
rect 212 -517 292 -515
rect -780 -573 -768 -517
rect -712 -573 224 -517
rect 280 -573 292 -517
rect -780 -585 -710 -573
rect 212 -575 292 -573
rect 541 -517 621 -515
rect 984 -517 1044 -507
rect 1698 -517 1778 -515
rect 541 -573 553 -517
rect 609 -573 986 -517
rect 1042 -573 1710 -517
rect 1766 -573 1778 -517
rect 541 -575 621 -573
rect 984 -585 1044 -573
rect 1698 -575 1778 -573
rect 2027 -517 2107 -515
rect 2294 -517 2364 -505
rect 2027 -573 2039 -517
rect 2095 -573 2296 -517
rect 2352 -573 2364 -517
rect 2027 -575 2107 -573
rect 2294 -583 2364 -573
rect 396 -633 476 -631
rect 1882 -633 1962 -631
rect -496 -689 408 -633
rect 464 -689 476 -633
rect -496 -1419 -440 -689
rect 396 -691 476 -689
rect 1126 -689 1894 -633
rect 1950 -689 1962 -633
rect 28 -783 108 -769
rect -185 -805 -139 -794
rect 28 -839 40 -783
rect 96 -839 108 -783
rect 212 -783 292 -769
rect 212 -839 224 -783
rect 280 -839 292 -783
rect 396 -783 476 -769
rect 396 -839 408 -783
rect 464 -839 476 -783
rect 643 -805 689 -794
rect 30 -842 41 -839
rect 95 -842 106 -839
rect 214 -842 225 -839
rect 279 -842 290 -839
rect 398 -842 409 -839
rect 463 -842 474 -839
rect -47 -888 -1 -877
rect -139 -1062 -47 -888
rect -47 -1073 -1 -1062
rect 137 -888 183 -877
rect 137 -1073 183 -1062
rect 321 -888 367 -877
rect 505 -888 551 -877
rect 488 -915 505 -913
rect 551 -915 568 -913
rect 488 -1035 500 -915
rect 556 -1035 568 -915
rect 488 -1037 505 -1035
rect 321 -1073 367 -1062
rect 551 -1037 568 -1035
rect 505 -1073 551 -1062
rect -185 -1290 -139 -1145
rect 30 -1154 41 -1108
rect 95 -1154 106 -1108
rect 30 -1187 106 -1154
rect 214 -1154 225 -1108
rect 279 -1154 290 -1108
rect 214 -1187 290 -1154
rect 398 -1154 409 -1108
rect 463 -1154 474 -1108
rect 398 -1187 474 -1154
rect 643 -1290 689 -1145
rect -197 -1302 -117 -1290
rect -197 -1358 -185 -1302
rect -129 -1358 -117 -1302
rect -197 -1370 -117 -1358
rect 621 -1302 699 -1290
rect 621 -1358 633 -1302
rect 689 -1358 699 -1302
rect 621 -1370 699 -1358
rect -848 -1475 -440 -1419
rect 1126 -1419 1182 -689
rect 1882 -691 1962 -689
rect 1514 -783 1594 -769
rect 1301 -805 1347 -794
rect 1514 -839 1526 -783
rect 1582 -839 1594 -783
rect 1698 -783 1778 -769
rect 1698 -839 1710 -783
rect 1766 -839 1778 -783
rect 1882 -783 1962 -769
rect 1882 -839 1894 -783
rect 1950 -839 1962 -783
rect 2129 -805 2175 -794
rect 1516 -842 1527 -839
rect 1581 -842 1592 -839
rect 1700 -842 1711 -839
rect 1765 -842 1776 -839
rect 1884 -842 1895 -839
rect 1949 -842 1960 -839
rect 1439 -888 1485 -877
rect 1347 -1062 1439 -888
rect 1439 -1073 1485 -1062
rect 1623 -888 1669 -877
rect 1623 -1073 1669 -1062
rect 1807 -888 1853 -877
rect 1991 -888 2037 -877
rect 1974 -915 1991 -913
rect 2037 -915 2054 -913
rect 1974 -1035 1986 -915
rect 2042 -1035 2054 -915
rect 1974 -1037 1991 -1035
rect 1807 -1073 1853 -1062
rect 2037 -1037 2054 -1035
rect 1991 -1073 2037 -1062
rect 1301 -1290 1347 -1145
rect 1516 -1154 1527 -1108
rect 1581 -1154 1592 -1108
rect 1516 -1187 1592 -1154
rect 1700 -1154 1711 -1108
rect 1765 -1154 1776 -1108
rect 1700 -1187 1776 -1154
rect 1884 -1154 1895 -1108
rect 1949 -1154 1960 -1108
rect 1884 -1187 1960 -1154
rect 2129 -1290 2175 -1145
rect 1289 -1302 1369 -1290
rect 1289 -1358 1301 -1302
rect 1357 -1358 1369 -1302
rect 1289 -1370 1369 -1358
rect 2107 -1302 2185 -1290
rect 2107 -1358 2119 -1302
rect 2175 -1358 2185 -1302
rect 2107 -1370 2185 -1358
rect 2460 -1419 2540 -1409
rect 1126 -1475 2472 -1419
rect 2528 -1475 2540 -1419
rect -496 -2722 -440 -1475
rect 2460 -1477 2540 -1475
rect 984 -1530 1054 -1528
rect 2284 -1529 2364 -1527
rect -360 -1586 986 -1530
rect 1042 -1586 1054 -1530
rect -360 -2606 -304 -1586
rect 984 -1598 1054 -1586
rect 1126 -1585 2296 -1529
rect 2352 -1585 2364 -1529
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect -185 -1850 -139 -1839
rect 30 -1841 106 -1808
rect 30 -1887 41 -1841
rect 95 -1887 106 -1841
rect 214 -1841 290 -1808
rect 214 -1887 225 -1841
rect 279 -1887 290 -1841
rect 398 -1841 474 -1808
rect 398 -1887 409 -1841
rect 463 -1887 474 -1841
rect 643 -1850 689 -1839
rect -47 -1933 -1 -1922
rect -64 -1960 -47 -1958
rect 137 -1933 183 -1922
rect -1 -1960 16 -1958
rect -139 -2080 -52 -1960
rect 4 -2080 16 -1960
rect -64 -2082 -47 -2080
rect -139 -2380 -47 -2260
rect -1 -2082 16 -2080
rect 120 -2260 137 -2258
rect 321 -1933 367 -1922
rect 304 -1960 321 -1958
rect 505 -1933 551 -1922
rect 367 -1960 384 -1958
rect 304 -2080 316 -1960
rect 372 -2080 384 -1960
rect 304 -2082 321 -2080
rect 183 -2260 200 -2258
rect 120 -2380 132 -2260
rect 188 -2380 200 -2260
rect 120 -2382 137 -2380
rect -47 -2418 -1 -2407
rect 183 -2382 200 -2380
rect 137 -2418 183 -2407
rect 367 -2082 384 -2080
rect 488 -2260 505 -2258
rect 626 -1960 643 -1958
rect 689 -1960 706 -1958
rect 626 -2081 638 -1960
rect 694 -2081 706 -1960
rect 626 -2083 643 -2081
rect 551 -2260 568 -2258
rect 488 -2380 500 -2260
rect 556 -2380 568 -2260
rect 488 -2382 505 -2380
rect 321 -2418 367 -2407
rect 551 -2382 568 -2380
rect 505 -2418 551 -2407
rect 30 -2456 41 -2453
rect 95 -2456 106 -2453
rect 214 -2456 225 -2453
rect 279 -2456 290 -2453
rect 398 -2456 409 -2453
rect 463 -2456 474 -2453
rect -185 -2501 -139 -2490
rect 28 -2512 40 -2456
rect 96 -2512 108 -2456
rect 28 -2526 108 -2512
rect 212 -2512 224 -2456
rect 280 -2512 292 -2456
rect 212 -2526 292 -2512
rect 396 -2512 408 -2456
rect 464 -2512 476 -2456
rect 689 -2083 706 -2081
rect 643 -2501 689 -2490
rect 396 -2526 476 -2512
rect 28 -2606 108 -2604
rect -360 -2662 40 -2606
rect 96 -2662 108 -2606
rect 1126 -2605 1182 -1585
rect 2284 -1597 2364 -1585
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect 1301 -1849 1347 -1838
rect 1516 -1840 1592 -1807
rect 1516 -1886 1527 -1840
rect 1581 -1886 1592 -1840
rect 1700 -1840 1776 -1807
rect 1700 -1886 1711 -1840
rect 1765 -1886 1776 -1840
rect 1884 -1840 1960 -1807
rect 1884 -1886 1895 -1840
rect 1949 -1886 1960 -1840
rect 2129 -1849 2175 -1838
rect 1439 -1932 1485 -1921
rect 1422 -1959 1439 -1957
rect 1623 -1932 1669 -1921
rect 1485 -1959 1502 -1957
rect 1347 -2079 1434 -1959
rect 1490 -2079 1502 -1959
rect 1422 -2081 1439 -2079
rect 1347 -2379 1439 -2259
rect 1485 -2081 1502 -2079
rect 1606 -2259 1623 -2257
rect 1807 -1932 1853 -1921
rect 1790 -1959 1807 -1957
rect 1991 -1932 2037 -1921
rect 1853 -1959 1870 -1957
rect 1790 -2079 1802 -1959
rect 1858 -2079 1870 -1959
rect 1790 -2081 1807 -2079
rect 1669 -2259 1686 -2257
rect 1606 -2379 1618 -2259
rect 1674 -2379 1686 -2259
rect 1606 -2381 1623 -2379
rect 1439 -2417 1485 -2406
rect 1669 -2381 1686 -2379
rect 1623 -2417 1669 -2406
rect 1853 -2081 1870 -2079
rect 1974 -2259 1991 -2257
rect 2112 -1959 2129 -1957
rect 2175 -1959 2192 -1957
rect 2112 -2080 2124 -1959
rect 2180 -2080 2192 -1959
rect 2112 -2082 2129 -2080
rect 2037 -2259 2054 -2257
rect 1974 -2379 1986 -2259
rect 2042 -2379 2054 -2259
rect 1974 -2381 1991 -2379
rect 1807 -2417 1853 -2406
rect 2037 -2381 2054 -2379
rect 1991 -2417 2037 -2406
rect 1516 -2455 1527 -2452
rect 1581 -2455 1592 -2452
rect 1700 -2455 1711 -2452
rect 1765 -2455 1776 -2452
rect 1884 -2455 1895 -2452
rect 1949 -2455 1960 -2452
rect 1301 -2500 1347 -2489
rect 1514 -2511 1526 -2455
rect 1582 -2511 1594 -2455
rect 1514 -2525 1594 -2511
rect 1698 -2511 1710 -2455
rect 1766 -2511 1778 -2455
rect 1698 -2525 1778 -2511
rect 1882 -2511 1894 -2455
rect 1950 -2511 1962 -2455
rect 2175 -2082 2192 -2080
rect 2129 -2500 2175 -2489
rect 1882 -2525 1962 -2511
rect 1514 -2605 1594 -2603
rect 1126 -2661 1526 -2605
rect 1582 -2661 1594 -2605
rect 28 -2664 108 -2662
rect 1514 -2663 1594 -2661
rect 212 -2722 292 -2720
rect -496 -2778 224 -2722
rect 280 -2778 292 -2722
rect 212 -2780 292 -2778
rect 541 -2722 621 -2720
rect 808 -2721 878 -2710
rect 1698 -2721 1778 -2719
rect 808 -2722 1710 -2721
rect 541 -2778 553 -2722
rect 609 -2778 810 -2722
rect 866 -2777 1710 -2722
rect 1766 -2777 1778 -2721
rect 866 -2778 1126 -2777
rect 541 -2780 621 -2778
rect 808 -2788 878 -2778
rect 1698 -2779 1778 -2777
rect 2027 -2721 2107 -2719
rect 2470 -2721 2540 -2711
rect 2027 -2777 2039 -2721
rect 2095 -2777 2472 -2721
rect 2528 -2777 2540 -2721
rect 2027 -2779 2107 -2777
rect 2470 -2789 2540 -2777
rect -644 -2838 -574 -2826
rect 396 -2838 476 -2836
rect 1882 -2837 1962 -2835
rect -644 -2894 -632 -2838
rect -576 -2894 408 -2838
rect 464 -2894 476 -2838
rect -644 -2906 -574 -2894
rect -360 -3625 -304 -2894
rect 396 -2896 476 -2894
rect 1126 -2893 1894 -2837
rect 1950 -2893 1962 -2837
rect 28 -2988 108 -2974
rect -185 -3010 -139 -2999
rect 28 -3044 40 -2988
rect 96 -3044 108 -2988
rect 212 -2988 292 -2974
rect 212 -3044 224 -2988
rect 280 -3044 292 -2988
rect 396 -2988 476 -2974
rect 396 -3044 408 -2988
rect 464 -3044 476 -2988
rect 643 -3010 689 -2999
rect 30 -3047 41 -3044
rect 95 -3047 106 -3044
rect 214 -3047 225 -3044
rect 279 -3047 290 -3044
rect 398 -3047 409 -3044
rect 463 -3047 474 -3044
rect -47 -3093 -1 -3082
rect -139 -3267 -47 -3093
rect -47 -3278 -1 -3267
rect 137 -3093 183 -3082
rect 137 -3278 183 -3267
rect 321 -3093 367 -3082
rect 505 -3093 551 -3082
rect 488 -3120 505 -3118
rect 551 -3120 568 -3118
rect 488 -3240 500 -3120
rect 556 -3240 568 -3120
rect 488 -3242 505 -3240
rect 321 -3278 367 -3267
rect 551 -3242 568 -3240
rect 505 -3278 551 -3267
rect -185 -3495 -139 -3350
rect 30 -3359 41 -3313
rect 95 -3359 106 -3313
rect 30 -3392 106 -3359
rect 214 -3359 225 -3313
rect 279 -3359 290 -3313
rect 214 -3392 290 -3359
rect 398 -3359 409 -3313
rect 463 -3359 474 -3313
rect 398 -3392 474 -3359
rect 643 -3495 689 -3350
rect -197 -3507 -117 -3495
rect -197 -3563 -185 -3507
rect -129 -3563 -117 -3507
rect -197 -3575 -117 -3563
rect 621 -3507 699 -3495
rect 621 -3563 633 -3507
rect 689 -3563 699 -3507
rect 621 -3575 699 -3563
rect 974 -3625 1054 -3615
rect -360 -3681 986 -3625
rect 1042 -3681 1054 -3625
rect 974 -3683 1054 -3681
rect 808 -3734 878 -3732
rect -360 -3735 878 -3734
rect -360 -3789 810 -3735
rect 866 -3789 878 -3735
rect -360 -3790 878 -3789
rect -360 -4811 -304 -3790
rect 808 -3798 878 -3790
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect -185 -4055 -139 -4044
rect 30 -4046 106 -4013
rect 30 -4092 41 -4046
rect 95 -4092 106 -4046
rect 214 -4046 290 -4013
rect 214 -4092 225 -4046
rect 279 -4092 290 -4046
rect 398 -4046 474 -4013
rect 398 -4092 409 -4046
rect 463 -4092 474 -4046
rect 643 -4055 689 -4044
rect -47 -4138 -1 -4127
rect -64 -4165 -47 -4163
rect 137 -4138 183 -4127
rect -1 -4165 16 -4163
rect -139 -4285 -52 -4165
rect 4 -4285 16 -4165
rect -64 -4287 -47 -4285
rect -139 -4585 -47 -4465
rect -1 -4287 16 -4285
rect 120 -4465 137 -4463
rect 321 -4138 367 -4127
rect 304 -4165 321 -4163
rect 505 -4138 551 -4127
rect 367 -4165 384 -4163
rect 304 -4285 316 -4165
rect 372 -4285 384 -4165
rect 304 -4287 321 -4285
rect 183 -4465 200 -4463
rect 120 -4585 132 -4465
rect 188 -4585 200 -4465
rect 120 -4587 137 -4585
rect -47 -4623 -1 -4612
rect 183 -4587 200 -4585
rect 137 -4623 183 -4612
rect 367 -4287 384 -4285
rect 488 -4465 505 -4463
rect 626 -4165 643 -4163
rect 689 -4165 706 -4163
rect 626 -4286 638 -4165
rect 694 -4286 706 -4165
rect 626 -4288 643 -4286
rect 551 -4465 568 -4463
rect 488 -4585 500 -4465
rect 556 -4585 568 -4465
rect 488 -4587 505 -4585
rect 321 -4623 367 -4612
rect 551 -4587 568 -4585
rect 505 -4623 551 -4612
rect 30 -4661 41 -4658
rect 95 -4661 106 -4658
rect 214 -4661 225 -4658
rect 279 -4661 290 -4658
rect 398 -4661 409 -4658
rect 463 -4661 474 -4658
rect -185 -4706 -139 -4695
rect 28 -4717 40 -4661
rect 96 -4717 108 -4661
rect 28 -4731 108 -4717
rect 212 -4717 224 -4661
rect 280 -4717 292 -4661
rect 212 -4731 292 -4717
rect 396 -4717 408 -4661
rect 464 -4717 476 -4661
rect 689 -4288 706 -4286
rect 643 -4706 689 -4695
rect 396 -4731 476 -4717
rect 28 -4811 108 -4809
rect -360 -4867 40 -4811
rect 96 -4867 108 -4811
rect 28 -4869 108 -4867
rect -780 -4927 -710 -4913
rect 212 -4927 292 -4925
rect -780 -4983 -768 -4927
rect -712 -4983 224 -4927
rect 280 -4983 292 -4927
rect -780 -4995 -710 -4983
rect 212 -4985 292 -4983
rect 541 -4927 621 -4925
rect 984 -4927 1044 -4915
rect 541 -4983 553 -4927
rect 609 -4983 986 -4927
rect 1042 -4983 1044 -4927
rect 541 -4985 621 -4983
rect 984 -4995 1044 -4983
rect 396 -5043 476 -5041
rect -848 -5099 408 -5043
rect 464 -5099 476 -5043
rect 396 -5101 476 -5099
rect 28 -5193 108 -5179
rect -185 -5215 -139 -5204
rect 28 -5249 40 -5193
rect 96 -5249 108 -5193
rect 212 -5193 292 -5179
rect 212 -5249 224 -5193
rect 280 -5249 292 -5193
rect 396 -5193 476 -5179
rect 396 -5249 408 -5193
rect 464 -5249 476 -5193
rect 643 -5215 689 -5204
rect 30 -5252 41 -5249
rect 95 -5252 106 -5249
rect 214 -5252 225 -5249
rect 279 -5252 290 -5249
rect 398 -5252 409 -5249
rect 463 -5252 474 -5249
rect -47 -5298 -1 -5287
rect -139 -5472 -47 -5298
rect -47 -5483 -1 -5472
rect 137 -5298 183 -5287
rect 137 -5483 183 -5472
rect 321 -5298 367 -5287
rect 505 -5298 551 -5287
rect 488 -5325 505 -5323
rect 551 -5325 568 -5323
rect 488 -5445 500 -5325
rect 556 -5445 568 -5325
rect 488 -5447 505 -5445
rect 321 -5483 367 -5472
rect 551 -5447 568 -5445
rect 505 -5483 551 -5472
rect -185 -5700 -139 -5555
rect 30 -5564 41 -5518
rect 95 -5564 106 -5518
rect 30 -5597 106 -5564
rect 214 -5564 225 -5518
rect 279 -5564 290 -5518
rect 214 -5597 290 -5564
rect 398 -5564 409 -5518
rect 463 -5564 474 -5518
rect 398 -5597 474 -5564
rect 643 -5700 689 -5555
rect -197 -5712 -117 -5700
rect -197 -5768 -185 -5712
rect -129 -5768 -117 -5712
rect -197 -5780 -117 -5768
rect 621 -5712 701 -5700
rect 621 -5768 633 -5712
rect 689 -5768 701 -5712
rect 621 -5780 701 -5768
rect -770 -5830 -710 -5826
rect 1126 -5830 1182 -2893
rect 1882 -2895 1962 -2893
rect 1514 -2987 1594 -2973
rect 1301 -3009 1347 -2998
rect 1514 -3043 1526 -2987
rect 1582 -3043 1594 -2987
rect 1698 -2987 1778 -2973
rect 1698 -3043 1710 -2987
rect 1766 -3043 1778 -2987
rect 1882 -2987 1962 -2973
rect 1882 -3043 1894 -2987
rect 1950 -3043 1962 -2987
rect 2129 -3009 2175 -2998
rect 1516 -3046 1527 -3043
rect 1581 -3046 1592 -3043
rect 1700 -3046 1711 -3043
rect 1765 -3046 1776 -3043
rect 1884 -3046 1895 -3043
rect 1949 -3046 1960 -3043
rect 1439 -3092 1485 -3081
rect 1347 -3266 1439 -3092
rect 1439 -3277 1485 -3266
rect 1623 -3092 1669 -3081
rect 1623 -3277 1669 -3266
rect 1807 -3092 1853 -3081
rect 1991 -3092 2037 -3081
rect 1974 -3119 1991 -3117
rect 2037 -3119 2054 -3117
rect 1974 -3239 1986 -3119
rect 2042 -3239 2054 -3119
rect 1974 -3241 1991 -3239
rect 1807 -3277 1853 -3266
rect 2037 -3241 2054 -3239
rect 1991 -3277 2037 -3266
rect 1301 -3494 1347 -3349
rect 1516 -3358 1527 -3312
rect 1581 -3358 1592 -3312
rect 1516 -3391 1592 -3358
rect 1700 -3358 1711 -3312
rect 1765 -3358 1776 -3312
rect 1700 -3391 1776 -3358
rect 1884 -3358 1895 -3312
rect 1949 -3358 1960 -3312
rect 1884 -3391 1960 -3358
rect 2129 -3494 2175 -3349
rect 1289 -3506 1369 -3494
rect 1289 -3562 1301 -3506
rect 1357 -3562 1369 -3506
rect 1289 -3574 1369 -3562
rect 2107 -3506 2185 -3494
rect 2107 -3562 2119 -3506
rect 2175 -3562 2185 -3506
rect 2107 -3574 2185 -3562
rect -831 -5886 -768 -5830
rect -712 -5886 1182 -5830
rect -770 -5898 -710 -5886
<< via1 >>
rect 316 2717 372 2773
rect -52 2330 -47 2450
rect -47 2330 -1 2450
rect -1 2330 4 2450
rect 316 2330 321 2450
rect 321 2330 367 2450
rect 367 2330 372 2450
rect 132 2030 137 2150
rect 137 2030 183 2150
rect 183 2030 188 2150
rect 638 2329 643 2450
rect 643 2329 689 2450
rect 689 2329 694 2450
rect 500 2030 505 2150
rect 505 2030 551 2150
rect 551 2030 556 2150
rect 40 1911 41 1954
rect 41 1911 95 1954
rect 95 1911 96 1954
rect 40 1898 96 1911
rect 224 1911 225 1954
rect 225 1911 279 1954
rect 279 1911 280 1954
rect 224 1898 280 1911
rect 408 1911 409 1954
rect 409 1911 463 1954
rect 463 1911 464 1954
rect 408 1898 464 1911
rect 40 1748 96 1804
rect -632 1632 -576 1688
rect 224 1632 280 1688
rect 553 1632 609 1688
rect 810 1632 866 1688
rect 408 1516 464 1572
rect 40 1409 96 1422
rect 40 1366 41 1409
rect 41 1366 95 1409
rect 95 1366 96 1409
rect 224 1409 280 1422
rect 224 1366 225 1409
rect 225 1366 279 1409
rect 279 1366 280 1409
rect 408 1409 464 1422
rect 408 1366 409 1409
rect 409 1366 463 1409
rect 463 1366 464 1409
rect 500 1170 505 1290
rect 505 1170 551 1290
rect 551 1170 556 1290
rect -185 847 -129 903
rect 633 847 689 903
rect 986 729 1042 785
rect 810 621 866 675
rect 316 512 372 568
rect -52 125 -47 245
rect -47 125 -1 245
rect -1 125 4 245
rect 316 125 321 245
rect 321 125 367 245
rect 367 125 372 245
rect 132 -175 137 -55
rect 137 -175 183 -55
rect 183 -175 188 -55
rect 638 124 643 245
rect 643 124 689 245
rect 689 124 694 245
rect 500 -175 505 -55
rect 505 -175 551 -55
rect 551 -175 556 -55
rect 40 -294 41 -251
rect 41 -294 95 -251
rect 95 -294 96 -251
rect 40 -307 96 -294
rect 224 -294 225 -251
rect 225 -294 279 -251
rect 279 -294 280 -251
rect 224 -307 280 -294
rect 408 -294 409 -251
rect 409 -294 463 -251
rect 463 -294 464 -251
rect 408 -307 464 -294
rect 40 -457 96 -401
rect 1802 512 1858 568
rect 1434 125 1439 245
rect 1439 125 1485 245
rect 1485 125 1490 245
rect 1802 125 1807 245
rect 1807 125 1853 245
rect 1853 125 1858 245
rect 1618 -175 1623 -55
rect 1623 -175 1669 -55
rect 1669 -175 1674 -55
rect 2124 124 2129 245
rect 2129 124 2175 245
rect 2175 124 2180 245
rect 1986 -175 1991 -55
rect 1991 -175 2037 -55
rect 2037 -175 2042 -55
rect 1526 -294 1527 -251
rect 1527 -294 1581 -251
rect 1581 -294 1582 -251
rect 1526 -307 1582 -294
rect 1710 -294 1711 -251
rect 1711 -294 1765 -251
rect 1765 -294 1766 -251
rect 1710 -307 1766 -294
rect 1894 -294 1895 -251
rect 1895 -294 1949 -251
rect 1949 -294 1950 -251
rect 1894 -307 1950 -294
rect 1526 -457 1582 -401
rect -768 -573 -712 -517
rect 224 -573 280 -517
rect 553 -573 609 -517
rect 986 -573 1042 -517
rect 1710 -573 1766 -517
rect 2039 -573 2095 -517
rect 2296 -573 2352 -517
rect 408 -689 464 -633
rect 1894 -689 1950 -633
rect 40 -796 96 -783
rect 40 -839 41 -796
rect 41 -839 95 -796
rect 95 -839 96 -796
rect 224 -796 280 -783
rect 224 -839 225 -796
rect 225 -839 279 -796
rect 279 -839 280 -796
rect 408 -796 464 -783
rect 408 -839 409 -796
rect 409 -839 463 -796
rect 463 -839 464 -796
rect 500 -1035 505 -915
rect 505 -1035 551 -915
rect 551 -1035 556 -915
rect -185 -1358 -129 -1302
rect 633 -1358 689 -1302
rect 1526 -796 1582 -783
rect 1526 -839 1527 -796
rect 1527 -839 1581 -796
rect 1581 -839 1582 -796
rect 1710 -796 1766 -783
rect 1710 -839 1711 -796
rect 1711 -839 1765 -796
rect 1765 -839 1766 -796
rect 1894 -796 1950 -783
rect 1894 -839 1895 -796
rect 1895 -839 1949 -796
rect 1949 -839 1950 -796
rect 1986 -1035 1991 -915
rect 1991 -1035 2037 -915
rect 2037 -1035 2042 -915
rect 1301 -1358 1357 -1302
rect 2119 -1358 2175 -1302
rect 2472 -1475 2528 -1419
rect 986 -1586 1042 -1530
rect 2296 -1585 2352 -1529
rect 316 -1693 372 -1637
rect -52 -2080 -47 -1960
rect -47 -2080 -1 -1960
rect -1 -2080 4 -1960
rect 316 -2080 321 -1960
rect 321 -2080 367 -1960
rect 367 -2080 372 -1960
rect 132 -2380 137 -2260
rect 137 -2380 183 -2260
rect 183 -2380 188 -2260
rect 638 -2081 643 -1960
rect 643 -2081 689 -1960
rect 689 -2081 694 -1960
rect 500 -2380 505 -2260
rect 505 -2380 551 -2260
rect 551 -2380 556 -2260
rect 40 -2499 41 -2456
rect 41 -2499 95 -2456
rect 95 -2499 96 -2456
rect 40 -2512 96 -2499
rect 224 -2499 225 -2456
rect 225 -2499 279 -2456
rect 279 -2499 280 -2456
rect 224 -2512 280 -2499
rect 408 -2499 409 -2456
rect 409 -2499 463 -2456
rect 463 -2499 464 -2456
rect 408 -2512 464 -2499
rect 40 -2662 96 -2606
rect 1802 -1692 1858 -1636
rect 1434 -2079 1439 -1959
rect 1439 -2079 1485 -1959
rect 1485 -2079 1490 -1959
rect 1802 -2079 1807 -1959
rect 1807 -2079 1853 -1959
rect 1853 -2079 1858 -1959
rect 1618 -2379 1623 -2259
rect 1623 -2379 1669 -2259
rect 1669 -2379 1674 -2259
rect 2124 -2080 2129 -1959
rect 2129 -2080 2175 -1959
rect 2175 -2080 2180 -1959
rect 1986 -2379 1991 -2259
rect 1991 -2379 2037 -2259
rect 2037 -2379 2042 -2259
rect 1526 -2498 1527 -2455
rect 1527 -2498 1581 -2455
rect 1581 -2498 1582 -2455
rect 1526 -2511 1582 -2498
rect 1710 -2498 1711 -2455
rect 1711 -2498 1765 -2455
rect 1765 -2498 1766 -2455
rect 1710 -2511 1766 -2498
rect 1894 -2498 1895 -2455
rect 1895 -2498 1949 -2455
rect 1949 -2498 1950 -2455
rect 1894 -2511 1950 -2498
rect 1526 -2661 1582 -2605
rect 224 -2778 280 -2722
rect 553 -2778 609 -2722
rect 810 -2778 866 -2722
rect 1710 -2777 1766 -2721
rect 2039 -2777 2095 -2721
rect 2472 -2777 2528 -2721
rect -632 -2894 -576 -2838
rect 408 -2894 464 -2838
rect 1894 -2893 1950 -2837
rect 40 -3001 96 -2988
rect 40 -3044 41 -3001
rect 41 -3044 95 -3001
rect 95 -3044 96 -3001
rect 224 -3001 280 -2988
rect 224 -3044 225 -3001
rect 225 -3044 279 -3001
rect 279 -3044 280 -3001
rect 408 -3001 464 -2988
rect 408 -3044 409 -3001
rect 409 -3044 463 -3001
rect 463 -3044 464 -3001
rect 500 -3240 505 -3120
rect 505 -3240 551 -3120
rect 551 -3240 556 -3120
rect -185 -3563 -129 -3507
rect 633 -3563 689 -3507
rect 986 -3681 1042 -3625
rect 810 -3789 866 -3735
rect 316 -3898 372 -3842
rect -52 -4285 -47 -4165
rect -47 -4285 -1 -4165
rect -1 -4285 4 -4165
rect 316 -4285 321 -4165
rect 321 -4285 367 -4165
rect 367 -4285 372 -4165
rect 132 -4585 137 -4465
rect 137 -4585 183 -4465
rect 183 -4585 188 -4465
rect 638 -4286 643 -4165
rect 643 -4286 689 -4165
rect 689 -4286 694 -4165
rect 500 -4585 505 -4465
rect 505 -4585 551 -4465
rect 551 -4585 556 -4465
rect 40 -4704 41 -4661
rect 41 -4704 95 -4661
rect 95 -4704 96 -4661
rect 40 -4717 96 -4704
rect 224 -4704 225 -4661
rect 225 -4704 279 -4661
rect 279 -4704 280 -4661
rect 224 -4717 280 -4704
rect 408 -4704 409 -4661
rect 409 -4704 463 -4661
rect 463 -4704 464 -4661
rect 408 -4717 464 -4704
rect 40 -4867 96 -4811
rect -768 -4983 -712 -4927
rect 224 -4983 280 -4927
rect 553 -4983 609 -4927
rect 986 -4983 1042 -4927
rect 408 -5099 464 -5043
rect 40 -5206 96 -5193
rect 40 -5249 41 -5206
rect 41 -5249 95 -5206
rect 95 -5249 96 -5206
rect 224 -5206 280 -5193
rect 224 -5249 225 -5206
rect 225 -5249 279 -5206
rect 279 -5249 280 -5206
rect 408 -5206 464 -5193
rect 408 -5249 409 -5206
rect 409 -5249 463 -5206
rect 463 -5249 464 -5206
rect 500 -5445 505 -5325
rect 505 -5445 551 -5325
rect 551 -5445 556 -5325
rect -185 -5768 -129 -5712
rect 633 -5768 689 -5712
rect 1526 -3000 1582 -2987
rect 1526 -3043 1527 -3000
rect 1527 -3043 1581 -3000
rect 1581 -3043 1582 -3000
rect 1710 -3000 1766 -2987
rect 1710 -3043 1711 -3000
rect 1711 -3043 1765 -3000
rect 1765 -3043 1766 -3000
rect 1894 -3000 1950 -2987
rect 1894 -3043 1895 -3000
rect 1895 -3043 1949 -3000
rect 1949 -3043 1950 -3000
rect 1986 -3239 1991 -3119
rect 1991 -3239 2037 -3119
rect 2037 -3239 2042 -3119
rect 1301 -3562 1357 -3506
rect 2119 -3562 2175 -3506
rect -768 -5886 -712 -5830
<< metal2 >>
rect -52 2773 694 2785
rect -52 2717 316 2773
rect 372 2717 694 2773
rect -52 2705 694 2717
rect -52 2452 4 2705
rect 316 2452 372 2705
rect 638 2452 694 2705
rect -64 2450 16 2452
rect -64 2330 -52 2450
rect 4 2330 16 2450
rect -64 2328 16 2330
rect 304 2450 384 2452
rect 304 2330 316 2450
rect 372 2330 384 2450
rect 304 2328 384 2330
rect 626 2450 706 2452
rect 626 2329 638 2450
rect 694 2329 706 2450
rect -52 2320 4 2328
rect 316 2320 372 2328
rect 626 2327 706 2329
rect 638 2319 694 2327
rect 132 2152 188 2160
rect 500 2152 556 2160
rect 120 2150 609 2152
rect 120 2030 132 2150
rect 188 2030 500 2150
rect 556 2030 609 2150
rect 120 2028 609 2030
rect 132 2020 188 2028
rect 500 2020 609 2028
rect 28 1954 108 1964
rect 28 1898 40 1954
rect 96 1898 108 1954
rect 28 1888 108 1898
rect 212 1954 292 1964
rect 212 1898 224 1954
rect 280 1898 292 1954
rect 212 1888 292 1898
rect 396 1954 476 1964
rect 396 1898 408 1954
rect 464 1898 476 1954
rect 396 1888 476 1898
rect 40 1806 96 1888
rect 28 1804 108 1806
rect 28 1748 40 1804
rect 96 1748 108 1804
rect 28 1746 108 1748
rect -644 1688 -574 1700
rect -644 1632 -632 1688
rect -576 1632 -574 1688
rect -644 1620 -574 1632
rect -780 -517 -710 -503
rect -780 -573 -768 -517
rect -712 -573 -710 -517
rect -780 -585 -710 -573
rect -768 -4913 -712 -585
rect -632 -2826 -576 1620
rect 40 1432 96 1746
rect 224 1690 280 1888
rect 212 1688 292 1690
rect 212 1632 224 1688
rect 280 1632 292 1688
rect 212 1630 292 1632
rect 224 1432 280 1630
rect 408 1574 464 1888
rect 541 1690 609 2020
rect 541 1688 621 1690
rect 541 1632 553 1688
rect 609 1632 621 1688
rect 541 1630 621 1632
rect 808 1688 878 1700
rect 808 1632 810 1688
rect 866 1632 878 1688
rect 396 1572 476 1574
rect 396 1516 408 1572
rect 464 1516 476 1572
rect 396 1514 476 1516
rect 408 1432 464 1514
rect 28 1422 108 1432
rect 28 1366 40 1422
rect 96 1366 108 1422
rect 28 1356 108 1366
rect 212 1422 292 1432
rect 212 1366 224 1422
rect 280 1366 292 1422
rect 212 1356 292 1366
rect 396 1422 476 1432
rect 396 1366 408 1422
rect 464 1366 476 1422
rect 396 1356 476 1366
rect 541 1300 609 1630
rect 808 1622 878 1632
rect 500 1292 609 1300
rect 488 1290 609 1292
rect 488 1170 500 1290
rect 556 1170 609 1290
rect 488 1168 609 1170
rect 500 1160 556 1168
rect -197 903 701 915
rect -197 847 -185 903
rect -129 847 633 903
rect 689 847 701 903
rect -197 835 701 847
rect 810 678 866 1622
rect 974 785 1054 795
rect 974 729 986 785
rect 1042 729 1054 785
rect 974 727 1054 729
rect 808 675 878 678
rect 808 621 810 675
rect 866 621 878 675
rect 808 609 878 621
rect -52 568 694 580
rect -52 512 316 568
rect 372 512 694 568
rect -52 500 694 512
rect -52 247 4 500
rect 316 247 372 500
rect 638 247 694 500
rect -64 245 16 247
rect -64 125 -52 245
rect 4 125 16 245
rect -64 123 16 125
rect 304 245 384 247
rect 304 125 316 245
rect 372 125 384 245
rect 304 123 384 125
rect 626 245 706 247
rect 626 124 638 245
rect 694 124 706 245
rect -52 115 4 123
rect 316 115 372 123
rect 626 122 706 124
rect 638 114 694 122
rect 132 -53 188 -45
rect 500 -53 556 -45
rect 120 -55 609 -53
rect 120 -175 132 -55
rect 188 -175 500 -55
rect 556 -175 609 -55
rect 120 -177 609 -175
rect 132 -185 188 -177
rect 500 -185 609 -177
rect 28 -251 108 -241
rect 28 -307 40 -251
rect 96 -307 108 -251
rect 28 -317 108 -307
rect 212 -251 292 -241
rect 212 -307 224 -251
rect 280 -307 292 -251
rect 212 -317 292 -307
rect 396 -251 476 -241
rect 396 -307 408 -251
rect 464 -307 476 -251
rect 396 -317 476 -307
rect 40 -399 96 -317
rect 28 -401 108 -399
rect 28 -457 40 -401
rect 96 -457 108 -401
rect 28 -459 108 -457
rect 40 -773 96 -459
rect 224 -515 280 -317
rect 212 -517 292 -515
rect 212 -573 224 -517
rect 280 -573 292 -517
rect 212 -575 292 -573
rect 224 -773 280 -575
rect 408 -631 464 -317
rect 541 -515 609 -185
rect 986 -507 1042 727
rect 1434 568 2180 580
rect 1434 512 1802 568
rect 1858 512 2180 568
rect 1434 500 2180 512
rect 1434 247 1490 500
rect 1802 247 1858 500
rect 2124 247 2180 500
rect 1422 245 1502 247
rect 1422 125 1434 245
rect 1490 125 1502 245
rect 1422 123 1502 125
rect 1790 245 1870 247
rect 1790 125 1802 245
rect 1858 125 1870 245
rect 1790 123 1870 125
rect 2112 245 2192 247
rect 2112 124 2124 245
rect 2180 124 2192 245
rect 1434 115 1490 123
rect 1802 115 1858 123
rect 2112 122 2192 124
rect 2124 114 2180 122
rect 1618 -53 1674 -45
rect 1986 -53 2042 -45
rect 1606 -55 2095 -53
rect 1606 -175 1618 -55
rect 1674 -175 1986 -55
rect 2042 -175 2095 -55
rect 1606 -177 2095 -175
rect 1618 -185 1674 -177
rect 1986 -185 2095 -177
rect 1514 -251 1594 -241
rect 1514 -307 1526 -251
rect 1582 -307 1594 -251
rect 1514 -317 1594 -307
rect 1698 -251 1778 -241
rect 1698 -307 1710 -251
rect 1766 -307 1778 -251
rect 1698 -317 1778 -307
rect 1882 -251 1962 -241
rect 1882 -307 1894 -251
rect 1950 -307 1962 -251
rect 1882 -317 1962 -307
rect 1526 -399 1582 -317
rect 1514 -401 1594 -399
rect 1514 -457 1526 -401
rect 1582 -457 1594 -401
rect 1514 -459 1594 -457
rect 541 -517 621 -515
rect 541 -573 553 -517
rect 609 -573 621 -517
rect 541 -575 621 -573
rect 984 -517 1044 -507
rect 984 -573 986 -517
rect 1042 -573 1044 -517
rect 396 -633 476 -631
rect 396 -689 408 -633
rect 464 -689 476 -633
rect 396 -691 476 -689
rect 408 -773 464 -691
rect 28 -783 108 -773
rect 28 -839 40 -783
rect 96 -839 108 -783
rect 28 -849 108 -839
rect 212 -783 292 -773
rect 212 -839 224 -783
rect 280 -839 292 -783
rect 212 -849 292 -839
rect 396 -783 476 -773
rect 396 -839 408 -783
rect 464 -839 476 -783
rect 396 -849 476 -839
rect 541 -905 609 -575
rect 984 -585 1044 -573
rect 500 -913 609 -905
rect 488 -915 609 -913
rect 488 -1035 500 -915
rect 556 -1035 609 -915
rect 488 -1037 609 -1035
rect 500 -1045 556 -1037
rect -197 -1302 699 -1290
rect -197 -1358 -185 -1302
rect -129 -1358 633 -1302
rect 689 -1358 699 -1302
rect -197 -1370 699 -1358
rect 986 -1528 1042 -585
rect 1526 -773 1582 -459
rect 1710 -515 1766 -317
rect 1698 -517 1778 -515
rect 1698 -573 1710 -517
rect 1766 -573 1778 -517
rect 1698 -575 1778 -573
rect 1710 -773 1766 -575
rect 1894 -631 1950 -317
rect 2027 -515 2095 -185
rect 2027 -517 2107 -515
rect 2027 -573 2039 -517
rect 2095 -573 2107 -517
rect 2027 -575 2107 -573
rect 2294 -517 2364 -505
rect 2294 -573 2296 -517
rect 2352 -573 2620 -517
rect 1882 -633 1962 -631
rect 1882 -689 1894 -633
rect 1950 -689 1962 -633
rect 1882 -691 1962 -689
rect 1894 -773 1950 -691
rect 1514 -783 1594 -773
rect 1514 -839 1526 -783
rect 1582 -839 1594 -783
rect 1514 -849 1594 -839
rect 1698 -783 1778 -773
rect 1698 -839 1710 -783
rect 1766 -839 1778 -783
rect 1698 -849 1778 -839
rect 1882 -783 1962 -773
rect 1882 -839 1894 -783
rect 1950 -839 1962 -783
rect 1882 -849 1962 -839
rect 2027 -905 2095 -575
rect 2294 -583 2364 -573
rect 1986 -913 2095 -905
rect 1974 -915 2095 -913
rect 1974 -1035 1986 -915
rect 2042 -1035 2095 -915
rect 1974 -1037 2095 -1035
rect 1986 -1045 2042 -1037
rect 1289 -1302 2185 -1290
rect 1289 -1358 1301 -1302
rect 1357 -1358 2119 -1302
rect 2175 -1358 2185 -1302
rect 1289 -1370 2185 -1358
rect 2296 -1527 2352 -583
rect 2460 -1419 2540 -1409
rect 2460 -1475 2472 -1419
rect 2528 -1475 2540 -1419
rect 2460 -1477 2540 -1475
rect 984 -1530 1054 -1528
rect 984 -1586 986 -1530
rect 1042 -1586 1054 -1530
rect 984 -1598 1054 -1586
rect 2284 -1529 2364 -1527
rect 2284 -1585 2296 -1529
rect 2352 -1585 2364 -1529
rect 2284 -1597 2364 -1585
rect -52 -1637 694 -1625
rect -52 -1693 316 -1637
rect 372 -1693 694 -1637
rect -52 -1705 694 -1693
rect -52 -1958 4 -1705
rect 316 -1958 372 -1705
rect 638 -1958 694 -1705
rect 1434 -1636 2180 -1624
rect 1434 -1692 1802 -1636
rect 1858 -1692 2180 -1636
rect 1434 -1704 2180 -1692
rect 1434 -1957 1490 -1704
rect 1802 -1957 1858 -1704
rect 2124 -1957 2180 -1704
rect -64 -1960 16 -1958
rect -64 -2080 -52 -1960
rect 4 -2080 16 -1960
rect -64 -2082 16 -2080
rect 304 -1960 384 -1958
rect 304 -2080 316 -1960
rect 372 -2080 384 -1960
rect 304 -2082 384 -2080
rect 626 -1960 706 -1958
rect 626 -2081 638 -1960
rect 694 -2081 706 -1960
rect 1422 -1959 1502 -1957
rect 1422 -2079 1434 -1959
rect 1490 -2079 1502 -1959
rect 1422 -2081 1502 -2079
rect 1790 -1959 1870 -1957
rect 1790 -2079 1802 -1959
rect 1858 -2079 1870 -1959
rect 1790 -2081 1870 -2079
rect 2112 -1959 2192 -1957
rect 2112 -2080 2124 -1959
rect 2180 -2080 2192 -1959
rect -52 -2090 4 -2082
rect 316 -2090 372 -2082
rect 626 -2083 706 -2081
rect 638 -2091 694 -2083
rect 1434 -2089 1490 -2081
rect 1802 -2089 1858 -2081
rect 2112 -2082 2192 -2080
rect 2124 -2090 2180 -2082
rect 132 -2258 188 -2250
rect 500 -2258 556 -2250
rect 1618 -2257 1674 -2249
rect 1986 -2257 2042 -2249
rect 120 -2260 609 -2258
rect 120 -2380 132 -2260
rect 188 -2380 500 -2260
rect 556 -2380 609 -2260
rect 120 -2382 609 -2380
rect 1606 -2259 2095 -2257
rect 1606 -2379 1618 -2259
rect 1674 -2379 1986 -2259
rect 2042 -2379 2095 -2259
rect 1606 -2381 2095 -2379
rect 132 -2390 188 -2382
rect 500 -2390 609 -2382
rect 1618 -2389 1674 -2381
rect 1986 -2389 2095 -2381
rect 28 -2456 108 -2446
rect 28 -2512 40 -2456
rect 96 -2512 108 -2456
rect 28 -2522 108 -2512
rect 212 -2456 292 -2446
rect 212 -2512 224 -2456
rect 280 -2512 292 -2456
rect 212 -2522 292 -2512
rect 396 -2456 476 -2446
rect 396 -2512 408 -2456
rect 464 -2512 476 -2456
rect 396 -2522 476 -2512
rect 40 -2604 96 -2522
rect 28 -2606 108 -2604
rect 28 -2662 40 -2606
rect 96 -2662 108 -2606
rect 28 -2664 108 -2662
rect -644 -2838 -574 -2826
rect -644 -2894 -632 -2838
rect -576 -2894 -574 -2838
rect -644 -2906 -574 -2894
rect 40 -2978 96 -2664
rect 224 -2720 280 -2522
rect 212 -2722 292 -2720
rect 212 -2778 224 -2722
rect 280 -2778 292 -2722
rect 212 -2780 292 -2778
rect 224 -2978 280 -2780
rect 408 -2836 464 -2522
rect 541 -2720 609 -2390
rect 1514 -2455 1594 -2445
rect 1514 -2511 1526 -2455
rect 1582 -2511 1594 -2455
rect 1514 -2521 1594 -2511
rect 1698 -2455 1778 -2445
rect 1698 -2511 1710 -2455
rect 1766 -2511 1778 -2455
rect 1698 -2521 1778 -2511
rect 1882 -2455 1962 -2445
rect 1882 -2511 1894 -2455
rect 1950 -2511 1962 -2455
rect 1882 -2521 1962 -2511
rect 1526 -2603 1582 -2521
rect 1514 -2605 1594 -2603
rect 1514 -2661 1526 -2605
rect 1582 -2661 1594 -2605
rect 1514 -2663 1594 -2661
rect 541 -2722 621 -2720
rect 541 -2778 553 -2722
rect 609 -2778 621 -2722
rect 541 -2780 621 -2778
rect 808 -2722 878 -2710
rect 808 -2778 810 -2722
rect 866 -2778 878 -2722
rect 396 -2838 476 -2836
rect 396 -2894 408 -2838
rect 464 -2894 476 -2838
rect 396 -2896 476 -2894
rect 408 -2978 464 -2896
rect 28 -2988 108 -2978
rect 28 -3044 40 -2988
rect 96 -3044 108 -2988
rect 28 -3054 108 -3044
rect 212 -2988 292 -2978
rect 212 -3044 224 -2988
rect 280 -3044 292 -2988
rect 212 -3054 292 -3044
rect 396 -2988 476 -2978
rect 396 -3044 408 -2988
rect 464 -3044 476 -2988
rect 396 -3054 476 -3044
rect 541 -3110 609 -2780
rect 808 -2788 878 -2778
rect 500 -3118 609 -3110
rect 488 -3120 609 -3118
rect 488 -3240 500 -3120
rect 556 -3240 609 -3120
rect 488 -3242 609 -3240
rect 500 -3250 556 -3242
rect -197 -3507 699 -3495
rect -197 -3563 -185 -3507
rect -129 -3563 633 -3507
rect 689 -3563 699 -3507
rect -197 -3575 699 -3563
rect 810 -3732 866 -2788
rect 1526 -2977 1582 -2663
rect 1710 -2719 1766 -2521
rect 1698 -2721 1778 -2719
rect 1698 -2777 1710 -2721
rect 1766 -2777 1778 -2721
rect 1698 -2779 1778 -2777
rect 1710 -2977 1766 -2779
rect 1894 -2835 1950 -2521
rect 2027 -2719 2095 -2389
rect 2472 -2711 2528 -1477
rect 2027 -2721 2107 -2719
rect 2027 -2777 2039 -2721
rect 2095 -2777 2107 -2721
rect 2027 -2779 2107 -2777
rect 2470 -2721 2540 -2711
rect 2470 -2777 2472 -2721
rect 2528 -2777 2620 -2721
rect 1882 -2837 1962 -2835
rect 1882 -2893 1894 -2837
rect 1950 -2893 1962 -2837
rect 1882 -2895 1962 -2893
rect 1894 -2977 1950 -2895
rect 1514 -2987 1594 -2977
rect 1514 -3043 1526 -2987
rect 1582 -3043 1594 -2987
rect 1514 -3053 1594 -3043
rect 1698 -2987 1778 -2977
rect 1698 -3043 1710 -2987
rect 1766 -3043 1778 -2987
rect 1698 -3053 1778 -3043
rect 1882 -2987 1962 -2977
rect 1882 -3043 1894 -2987
rect 1950 -3043 1962 -2987
rect 1882 -3053 1962 -3043
rect 2027 -3109 2095 -2779
rect 2470 -2789 2540 -2777
rect 1986 -3117 2095 -3109
rect 1974 -3119 2095 -3117
rect 1974 -3239 1986 -3119
rect 2042 -3239 2095 -3119
rect 1974 -3241 2095 -3239
rect 1986 -3249 2042 -3241
rect 1289 -3506 2185 -3494
rect 1289 -3562 1301 -3506
rect 1357 -3562 2119 -3506
rect 2175 -3562 2185 -3506
rect 1289 -3574 2185 -3562
rect 974 -3625 1054 -3615
rect 974 -3681 986 -3625
rect 1042 -3681 1054 -3625
rect 974 -3683 1054 -3681
rect 808 -3735 878 -3732
rect 808 -3789 810 -3735
rect 866 -3789 878 -3735
rect 808 -3801 878 -3789
rect -52 -3842 694 -3830
rect -52 -3898 316 -3842
rect 372 -3898 694 -3842
rect -52 -3910 694 -3898
rect -52 -4163 4 -3910
rect 316 -4163 372 -3910
rect 638 -4163 694 -3910
rect -64 -4165 16 -4163
rect -64 -4285 -52 -4165
rect 4 -4285 16 -4165
rect -64 -4287 16 -4285
rect 304 -4165 384 -4163
rect 304 -4285 316 -4165
rect 372 -4285 384 -4165
rect 304 -4287 384 -4285
rect 626 -4165 706 -4163
rect 626 -4286 638 -4165
rect 694 -4286 706 -4165
rect -52 -4295 4 -4287
rect 316 -4295 372 -4287
rect 626 -4288 706 -4286
rect 638 -4296 694 -4288
rect 132 -4463 188 -4455
rect 500 -4463 556 -4455
rect 120 -4465 609 -4463
rect 120 -4585 132 -4465
rect 188 -4585 500 -4465
rect 556 -4585 609 -4465
rect 120 -4587 609 -4585
rect 132 -4595 188 -4587
rect 500 -4595 609 -4587
rect 28 -4661 108 -4651
rect 28 -4717 40 -4661
rect 96 -4717 108 -4661
rect 28 -4727 108 -4717
rect 212 -4661 292 -4651
rect 212 -4717 224 -4661
rect 280 -4717 292 -4661
rect 212 -4727 292 -4717
rect 396 -4661 476 -4651
rect 396 -4717 408 -4661
rect 464 -4717 476 -4661
rect 396 -4727 476 -4717
rect 40 -4809 96 -4727
rect 28 -4811 108 -4809
rect 28 -4867 40 -4811
rect 96 -4867 108 -4811
rect 28 -4869 108 -4867
rect -780 -4927 -710 -4913
rect -780 -4983 -768 -4927
rect -712 -4983 -710 -4927
rect -780 -4995 -710 -4983
rect -768 -5826 -712 -4995
rect 40 -5183 96 -4869
rect 224 -4925 280 -4727
rect 212 -4927 292 -4925
rect 212 -4983 224 -4927
rect 280 -4983 292 -4927
rect 212 -4985 292 -4983
rect 224 -5183 280 -4985
rect 408 -5041 464 -4727
rect 541 -4925 609 -4595
rect 986 -4915 1042 -3683
rect 541 -4927 621 -4925
rect 541 -4983 553 -4927
rect 609 -4983 621 -4927
rect 541 -4985 621 -4983
rect 984 -4927 1044 -4915
rect 984 -4983 986 -4927
rect 1042 -4983 1044 -4927
rect 396 -5043 476 -5041
rect 396 -5099 408 -5043
rect 464 -5099 476 -5043
rect 396 -5101 476 -5099
rect 408 -5183 464 -5101
rect 28 -5193 108 -5183
rect 28 -5249 40 -5193
rect 96 -5249 108 -5193
rect 28 -5259 108 -5249
rect 212 -5193 292 -5183
rect 212 -5249 224 -5193
rect 280 -5249 292 -5193
rect 212 -5259 292 -5249
rect 396 -5193 476 -5183
rect 396 -5249 408 -5193
rect 464 -5249 476 -5193
rect 396 -5259 476 -5249
rect 541 -5315 609 -4985
rect 984 -4995 1044 -4983
rect 500 -5323 609 -5315
rect 488 -5325 609 -5323
rect 488 -5445 500 -5325
rect 556 -5445 609 -5325
rect 488 -5447 609 -5445
rect 500 -5455 556 -5447
rect -197 -5712 701 -5700
rect -197 -5768 -185 -5712
rect -129 -5768 633 -5712
rect 689 -5768 701 -5712
rect -197 -5780 701 -5768
rect -770 -5830 -710 -5826
rect -770 -5886 -768 -5830
rect -712 -5886 -710 -5830
rect -770 -5898 -710 -5886
<< via2 >>
rect 316 2717 372 2773
rect -185 847 -129 903
rect 633 847 689 903
rect 316 512 372 568
rect 1802 512 1858 568
rect -185 -1358 -129 -1302
rect 633 -1358 689 -1302
rect 1301 -1358 1357 -1302
rect 2119 -1358 2175 -1302
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect -185 -3563 -129 -3507
rect 633 -3563 689 -3507
rect 1301 -3562 1357 -3506
rect 2119 -3562 2175 -3506
rect 316 -3898 372 -3842
rect -185 -5768 -129 -5712
rect 633 -5768 689 -5712
<< metal3 >>
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -197 903 -117 915
rect -197 847 -185 903
rect -129 847 -117 903
rect -197 835 -117 847
rect 621 903 701 915
rect 621 847 633 903
rect 689 847 701 903
rect 621 835 701 847
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect -197 -1302 -117 -1290
rect -197 -1358 -185 -1302
rect -129 -1358 -117 -1302
rect -197 -1370 -117 -1358
rect 621 -1302 701 -1290
rect 621 -1358 633 -1302
rect 689 -1358 701 -1302
rect 621 -1370 701 -1358
rect 1289 -1302 1369 -1290
rect 1289 -1358 1301 -1302
rect 1357 -1358 1369 -1302
rect 1289 -1370 1369 -1358
rect 2107 -1302 2187 -1290
rect 2107 -1358 2119 -1302
rect 2175 -1358 2187 -1302
rect 2107 -1370 2187 -1358
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect -197 -3507 -117 -3495
rect -197 -3563 -185 -3507
rect -129 -3563 -117 -3507
rect -197 -3575 -117 -3563
rect 621 -3507 701 -3495
rect 621 -3563 633 -3507
rect 689 -3563 701 -3507
rect 621 -3575 701 -3563
rect 1289 -3506 1369 -3494
rect 1289 -3562 1301 -3506
rect 1357 -3562 1369 -3506
rect 1289 -3574 1369 -3562
rect 2107 -3506 2187 -3494
rect 2107 -3562 2119 -3506
rect 2175 -3562 2187 -3506
rect 2107 -3574 2187 -3562
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect -197 -5712 -117 -5700
rect -197 -5768 -185 -5712
rect -129 -5768 -117 -5712
rect -197 -5780 -117 -5768
rect 621 -5712 701 -5700
rect 621 -5768 633 -5712
rect 689 -5768 701 -5712
rect 621 -5780 701 -5768
<< via3 >>
rect 316 2717 372 2773
rect -185 847 -129 903
rect 633 847 689 903
rect 316 512 372 568
rect 1802 512 1858 568
rect -185 -1358 -129 -1302
rect 633 -1358 689 -1302
rect 1301 -1358 1357 -1302
rect 2119 -1358 2175 -1302
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect -185 -3563 -129 -3507
rect 633 -3563 689 -3507
rect 1301 -3562 1357 -3506
rect 2119 -3562 2175 -3506
rect 316 -3898 372 -3842
rect -185 -5768 -129 -5712
rect 633 -5768 689 -5712
<< metal4 >>
rect 304 2773 390 2777
rect 304 2717 316 2773
rect 372 2717 390 2773
rect 304 2705 390 2717
rect -710 903 2590 2569
rect -710 847 -185 903
rect -129 847 633 903
rect 689 847 2590 903
rect -710 729 2590 847
rect -710 364 122 729
rect 304 568 390 572
rect 304 512 316 568
rect 372 512 390 568
rect 304 500 390 512
rect 572 364 1608 729
rect 1790 568 1876 572
rect 1790 512 1802 568
rect 1858 512 1876 568
rect 1790 500 1876 512
rect 2058 364 2590 729
rect -710 -1302 2590 364
rect -710 -1358 -185 -1302
rect -129 -1358 633 -1302
rect 689 -1358 1301 -1302
rect 1357 -1358 2119 -1302
rect 2175 -1358 2590 -1302
rect -710 -1476 2590 -1358
rect -710 -1841 122 -1476
rect 304 -1637 390 -1633
rect 304 -1693 316 -1637
rect 372 -1693 390 -1637
rect 304 -1705 390 -1693
rect 572 -1841 1608 -1476
rect 1790 -1636 1876 -1632
rect 1790 -1692 1802 -1636
rect 1858 -1692 1876 -1636
rect 1790 -1704 1876 -1692
rect 2058 -1841 2590 -1476
rect -710 -3506 2590 -1841
rect -710 -3507 1301 -3506
rect -710 -3563 -185 -3507
rect -129 -3563 633 -3507
rect 689 -3562 1301 -3507
rect 1357 -3562 2119 -3506
rect 2175 -3562 2590 -3506
rect 689 -3563 2590 -3562
rect -710 -3681 2590 -3563
rect -710 -4046 122 -3681
rect 304 -3842 390 -3838
rect 304 -3898 316 -3842
rect 372 -3898 390 -3842
rect 304 -3910 390 -3898
rect 572 -4046 2590 -3681
rect -710 -5712 2590 -4046
rect -710 -5768 -185 -5712
rect -129 -5768 633 -5712
rect 689 -5768 2590 -5712
rect -710 -5898 2590 -5768
<< via4 >>
rect 316 2717 372 2773
rect 316 512 372 568
rect 1802 512 1858 568
rect 316 -1693 372 -1637
rect 1802 -1692 1858 -1636
rect 316 -3898 372 -3842
<< metal5 >>
rect -710 2773 2590 2881
rect -710 2717 316 2773
rect 372 2717 2590 2773
rect -710 568 2590 2717
rect -710 512 316 568
rect 372 512 1802 568
rect 1858 512 2590 568
rect -710 -1636 2590 512
rect -710 -1637 1802 -1636
rect -710 -1693 316 -1637
rect 372 -1692 1802 -1637
rect 1858 -1692 2590 -1636
rect 372 -1693 2590 -1692
rect -710 -3842 2590 -1693
rect -710 -3898 316 -3842
rect 372 -3898 2590 -3842
rect -710 -5898 2590 -3898
<< labels >>
rlabel metal1 -848 1776 -848 1776 7 setb
port 4 w
rlabel metal1 -848 -1447 -848 -1447 7 clk
port 3 w
rlabel metal1 -848 -5072 -848 -5072 7 d
port 2 w
rlabel metal1 -831 -5859 -831 -5859 7 resetb
port 5 w
rlabel metal2 2620 -545 2620 -545 3 Q
port 6 e
rlabel metal2 2620 -2750 2620 -2750 3 Qb
port 7 e
rlabel metal5 1260 2881 1260 2881 1 vdd
port 0 n
rlabel metal4 1219 -5898 1219 -5898 5 vss
port 1 s
<< end >>
