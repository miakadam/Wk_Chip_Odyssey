magic
tech gf180mcuD
magscale 1 10
timestamp 1757591539
<< nwell >>
rect 0 630 780 1270
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
rect 440 210 500 380
<< pmos >>
rect 190 720 250 1060
rect 360 720 420 1060
rect 530 720 590 1060
<< ndiff >>
rect 120 290 220 380
rect 120 230 140 290
rect 190 230 220 290
rect 120 210 220 230
rect 280 210 330 380
rect 390 210 440 380
rect 500 360 600 380
rect 500 230 530 360
rect 580 230 600 360
rect 500 210 600 230
<< pdiff >>
rect 90 1040 190 1060
rect 90 740 110 1040
rect 160 740 190 1040
rect 90 720 190 740
rect 250 1040 360 1060
rect 250 790 280 1040
rect 330 790 360 1040
rect 250 720 360 790
rect 420 1040 530 1060
rect 420 740 450 1040
rect 500 740 530 1040
rect 420 720 530 740
rect 590 1040 690 1060
rect 590 790 620 1040
rect 670 790 690 1040
rect 590 720 690 790
<< ndiffc >>
rect 140 230 190 290
rect 530 230 580 360
<< pdiffc >>
rect 110 740 160 1040
rect 280 790 330 1040
rect 450 740 500 1040
rect 620 790 670 1040
<< psubdiff >>
rect 60 120 210 140
rect 60 70 110 120
rect 160 70 210 120
rect 60 50 210 70
rect 300 120 450 140
rect 300 70 350 120
rect 400 70 450 120
rect 300 50 450 70
rect 540 120 690 140
rect 540 70 590 120
rect 640 70 690 120
rect 540 50 690 70
<< nsubdiff >>
rect 60 1200 210 1220
rect 60 1150 110 1200
rect 160 1150 210 1200
rect 60 1130 210 1150
rect 300 1200 450 1220
rect 300 1150 350 1200
rect 400 1150 450 1200
rect 300 1130 450 1150
rect 540 1200 690 1220
rect 540 1150 590 1200
rect 640 1150 690 1200
rect 540 1130 690 1150
<< psubdiffcont >>
rect 110 70 160 120
rect 350 70 400 120
rect 590 70 640 120
<< nsubdiffcont >>
rect 110 1150 160 1200
rect 350 1150 400 1200
rect 590 1150 640 1200
<< polysilicon >>
rect 190 1060 250 1110
rect 360 1060 420 1110
rect 530 1060 590 1110
rect 190 660 250 720
rect 360 660 420 720
rect 190 549 280 660
rect 110 529 280 549
rect 110 469 140 529
rect 200 469 280 529
rect 110 449 280 469
rect 220 380 280 449
rect 330 653 420 660
rect 330 633 477 653
rect 330 573 397 633
rect 457 573 477 633
rect 330 553 477 573
rect 330 486 420 553
rect 530 509 590 720
rect 530 501 670 509
rect 475 489 670 501
rect 330 380 390 486
rect 475 440 590 489
rect 440 429 590 440
rect 650 429 670 489
rect 440 409 670 429
rect 440 404 590 409
rect 440 380 500 404
rect 220 160 280 210
rect 330 160 390 210
rect 440 160 500 210
<< polycontact >>
rect 140 469 200 529
rect 397 573 457 633
rect 590 429 650 489
<< metal1 >>
rect 0 1200 780 1270
rect 0 1150 110 1200
rect 160 1150 350 1200
rect 400 1150 590 1200
rect 640 1150 780 1200
rect 0 1130 780 1150
rect 110 1040 160 1130
rect 280 1040 330 1060
rect 280 780 330 790
rect 450 1040 500 1130
rect 110 720 160 740
rect 260 720 280 780
rect 340 720 360 780
rect 620 1040 670 1060
rect 450 720 500 740
rect 598 780 682 790
rect 598 720 610 780
rect 670 720 682 780
rect 120 469 140 529
rect 200 469 220 529
rect 280 370 330 720
rect 377 573 397 633
rect 457 573 477 633
rect 570 429 590 489
rect 650 429 670 489
rect 140 320 330 370
rect 530 360 580 380
rect 140 290 190 320
rect 140 210 190 230
rect 530 140 580 230
rect 0 120 780 140
rect 0 70 110 120
rect 160 70 350 120
rect 400 70 590 120
rect 640 70 780 120
rect 0 0 780 70
<< via1 >>
rect 280 720 340 780
rect 610 720 670 780
rect 140 469 200 529
rect 397 573 457 633
rect 590 429 650 489
<< metal2 >>
rect 260 780 360 790
rect 598 780 682 790
rect 260 720 280 780
rect 340 720 610 780
rect 670 720 682 780
rect 260 710 360 720
rect 598 710 682 720
rect 377 633 477 643
rect 377 573 397 633
rect 457 573 477 633
rect 377 563 477 573
rect 120 529 220 539
rect 120 469 140 529
rect 200 469 220 529
rect 120 459 220 469
rect 570 489 670 499
rect 570 429 590 489
rect 650 429 670 489
rect 570 419 670 429
<< labels >>
rlabel metal2 310 750 310 750 1 Y
port 3 n
rlabel metal1 130 1180 130 1180 1 VDD
port 4 n
rlabel metal1 130 90 130 90 1 VSS
port 5 n
rlabel via1 170 499 170 499 1 A
port 1 n
rlabel via1 427 603 427 603 1 B
port 2 n
rlabel via1 620 459 620 459 1 C
port 6 n
<< end >>
