* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__buf_2 A Y VDD VSS
X0 VSS A a_90_210# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 VDD A a_90_210# VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 Y a_90_210# VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 Y a_90_210# VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X4 VSS a_90_210# Y VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X5 VDD a_90_210# Y VDD pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
.ends
