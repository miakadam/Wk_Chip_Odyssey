* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_2.ext - technology: (null)

.subckt gf180mcu_osu_sc_gp9t3v3__buf_2 A Y VDD VSS
X0 VSS.t1 A.t0 a_90_210# VSS.t0 nfet_03v3
**devattr s=17000,540 d=9350,280
X1 VDD.t1 A.t1 a_90_210# VDD.t0 pfet_03v3
**devattr s=34000,880 d=18700,450
X2 Y.t3 a_90_210# VSS.t5 VSS.t4 nfet_03v3
**devattr s=9350,280 d=9350,280
X3 Y.t1 a_90_210# VDD.t5 VDD.t4 pfet_03v3
**devattr s=18700,450 d=18700,450
X4 VSS.t3 a_90_210# Y.t2 VSS.t2 nfet_03v3
**devattr s=9350,280 d=17000,540
X5 VDD.t3 a_90_210# Y.t0 VDD.t2 pfet_03v3
**devattr s=18700,450 d=34000,880
R0 A.n0 A.t1 45.6255
R1 A.n0 A.t0 20.6838
R2 A A.n0 12.5005
R3 VSS.t2 VSS.t4 876.985
R4 VSS.t0 VSS.n4 799.604
R5 VSS.n5 VSS.t0 448.892
R6 VSS.n2 VSS.t2 294.13
R7 VSS.n4 VSS.t4 77.3815
R8 VSS.n4 VSS.n3 10.4005
R9 VSS.n2 VSS.t3 8.63702
R10 VSS.n1 VSS.n0 6.5795
R11 VSS.n0 VSS.t5 2.03874
R12 VSS.n0 VSS.t1 2.03874
R13 VSS.n3 VSS.n2 0.154786
R14 VSS.n5 VSS.n1 0.109786
R15 VSS.n3 VSS.n1 0.0455
R16 VSS VSS.n5 0.00371429
R17 VDD.t2 VDD.t4 265.625
R18 VDD.t0 VDD.n4 242.189
R19 VDD.n5 VDD.t0 145.413
R20 VDD.n2 VDD.t2 98.538
R21 VDD.n4 VDD.t4 23.438
R22 VDD.n4 VDD.n3 12.6005
R23 VDD.n2 VDD.t3 3.31747
R24 VDD.n1 VDD.n0 2.16583
R25 VDD.n0 VDD.t5 1.13285
R26 VDD.n0 VDD.t1 1.13285
R27 VDD.n3 VDD.n2 0.154786
R28 VDD.n5 VDD.n1 0.109786
R29 VDD.n3 VDD.n1 0.0455
R30 VDD VDD.n5 0.00371429
R31 Y.n2 Y.n1 7.0925
R32 Y Y.n2 4.5005
R33 Y.n1 Y.t2 2.03874
R34 Y.n1 Y.t3 2.03874
R35 Y.n2 Y.n0 2.00383
R36 Y.n0 Y.t0 1.13285
R37 Y.n0 Y.t1 1.13285
.ends

