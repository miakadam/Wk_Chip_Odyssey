magic
tech gf180mcuD
magscale 1 10
timestamp 1757668849
<< nwell >>
rect 1854 414 1880 435
rect 2146 191 2241 217
rect 2120 160 2250 191
rect 2118 132 2250 160
rect 2118 129 2248 132
rect 2118 101 2271 129
rect 2141 70 2271 101
<< pwell >>
rect 2146 -74 2224 70
rect 1910 -130 2224 -74
rect 2146 -231 2224 -130
rect 2146 -277 2241 -231
<< metal1 >>
rect 1962 699 2038 730
rect 2146 699 2222 730
rect 2330 699 2406 730
rect 2483 435 2578 607
rect 1854 433 1948 435
rect 1854 313 1880 433
rect 1936 313 1948 433
rect 1854 311 1948 313
rect 2052 433 2132 435
rect 2052 313 2064 433
rect 2120 313 2132 433
rect 2052 311 2132 313
rect 2236 433 2316 435
rect 2236 313 2248 433
rect 2304 313 2316 433
rect 2236 311 2316 313
rect 2420 433 2578 435
rect 2420 313 2432 433
rect 2488 313 2578 433
rect 2420 311 2578 313
rect 1854 -74 1910 311
rect 2483 293 2578 311
rect 1960 227 2040 229
rect 1960 171 1972 227
rect 2028 171 2040 227
rect 1960 169 2040 171
rect 2146 201 2334 217
rect 2146 171 2406 201
rect 2146 -74 2224 171
rect 1854 -130 2224 -74
rect 1854 -363 1910 -130
rect 1960 -231 2040 -229
rect 1960 -287 1972 -231
rect 2028 -287 2040 -231
rect 2146 -231 2224 -130
rect 2146 -261 2406 -231
rect 2146 -277 2341 -261
rect 1960 -289 2040 -287
rect 2330 -307 2341 -277
rect 2395 -307 2406 -261
rect 1854 -365 1948 -363
rect 1854 -485 1880 -365
rect 1936 -485 1948 -365
rect 1854 -487 1948 -485
rect 2052 -365 2132 -363
rect 2052 -485 2064 -365
rect 2120 -485 2132 -365
rect 2052 -487 2132 -485
rect 2236 -365 2316 -363
rect 2236 -485 2248 -365
rect 2304 -485 2316 -365
rect 2236 -487 2316 -485
rect 2420 -365 2588 -363
rect 2420 -485 2432 -365
rect 2488 -485 2588 -365
rect 2420 -487 2588 -485
rect 1962 -620 2038 -589
rect 2146 -620 2222 -589
rect 2330 -620 2406 -589
<< via1 >>
rect 1880 313 1936 433
rect 2064 313 2120 433
rect 2248 313 2304 433
rect 2432 313 2488 433
rect 1972 171 2028 227
rect 1972 -287 2028 -231
rect 1880 -485 1936 -365
rect 2064 -485 2120 -365
rect 2248 -485 2304 -365
rect 2432 -485 2488 -365
<< metal2 >>
rect 1710 830 2657 930
rect 1880 435 1936 443
rect 2064 435 2120 830
rect 2248 435 2304 443
rect 2432 435 2488 830
rect 1868 433 1948 435
rect 1868 313 1880 433
rect 1936 313 1948 433
rect 1868 311 1948 313
rect 2052 433 2132 435
rect 2052 313 2064 433
rect 2120 313 2132 433
rect 2052 311 2132 313
rect 2236 433 2316 435
rect 2236 313 2248 433
rect 2304 313 2316 433
rect 2236 311 2316 313
rect 2420 433 2500 435
rect 2420 313 2432 433
rect 2488 313 2500 433
rect 2420 311 2500 313
rect 1880 303 1936 311
rect 2064 303 2120 311
rect 1972 229 2028 237
rect 1960 227 2040 229
rect 1960 171 1972 227
rect 2028 171 2040 227
rect 1960 169 2040 171
rect 1972 26 2028 169
rect 1628 -30 2028 26
rect 1972 -229 2028 -30
rect 2248 26 2304 311
rect 2432 303 2488 311
rect 2248 -30 2740 26
rect 1960 -231 2040 -229
rect 1960 -287 1972 -231
rect 2028 -287 2040 -231
rect 1960 -289 2040 -287
rect 1972 -297 2028 -289
rect 1880 -363 1936 -355
rect 2064 -363 2120 -355
rect 2248 -363 2304 -30
rect 2432 -363 2488 -355
rect 1868 -365 1948 -363
rect 1868 -485 1880 -365
rect 1936 -485 1948 -365
rect 1868 -487 1948 -485
rect 2052 -365 2132 -363
rect 2052 -485 2064 -365
rect 2120 -485 2132 -365
rect 2052 -487 2132 -485
rect 2236 -365 2316 -363
rect 2236 -485 2248 -365
rect 2304 -485 2316 -365
rect 2236 -487 2316 -485
rect 2420 -365 2500 -363
rect 2420 -485 2432 -365
rect 2488 -485 2500 -365
rect 2420 -487 2500 -485
rect 1880 -495 1936 -487
rect 2064 -720 2120 -487
rect 2248 -495 2304 -487
rect 2432 -720 2488 -487
rect 1710 -820 2657 -720
use pfet_03v3_FUEB84  M3
timestamp 1757668360
transform 1 0 2184 0 1 450
box -474 -380 474 380
use nfet_03v3_5ZFFTM  M4
timestamp 1757668360
transform 1 0 2184 0 1 -425
box -474 -295 474 295
<< labels >>
rlabel metal2 2190 930 2190 930 1 VDD
port 0 n
rlabel metal2 2180 -820 2180 -820 5 VSS
port 3 s
rlabel metal2 1628 -1 1628 -1 7 A
port 1 w
rlabel metal2 2740 -4 2740 -4 3 Y
port 2 e
<< end >>
