magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 73 -23 119
rect 23 73 34 84
rect -103 -38 -57 38
rect 57 -38 103 38
rect -34 -119 -23 -73
<< pwell >>
rect -278 -250 278 250
<< nmos >>
rect -28 -40 28 40
<< ndiff >>
rect -116 27 -28 40
rect -116 -27 -103 27
rect -57 -27 -28 27
rect -116 -40 -28 -27
rect 28 27 116 40
rect 28 -27 57 27
rect 103 -27 116 27
rect 28 -40 116 -27
<< ndiffc >>
rect -103 -27 -57 27
rect 57 -27 103 27
<< psubdiff >>
rect -254 154 254 226
rect -254 110 -182 154
rect -254 -110 -241 110
rect -195 -110 -182 110
rect 182 110 254 154
rect -254 -154 -182 -110
rect 182 -110 195 110
rect 241 -110 254 110
rect 182 -154 254 -110
rect -254 -226 254 -154
<< psubdiffcont >>
rect -241 -110 -195 110
rect 195 -110 241 110
<< polysilicon >>
rect -36 119 36 132
rect -36 73 -23 119
rect 23 73 36 119
rect -36 60 36 73
rect -28 40 28 60
rect -28 -60 28 -40
rect -36 -73 36 -60
rect -36 -119 -23 -73
rect 23 -119 36 -73
rect -36 -132 36 -119
<< polycontact >>
rect -23 73 23 119
rect -23 -119 23 -73
<< metal1 >>
rect -241 167 241 213
rect -241 110 -195 167
rect -34 73 -23 119
rect 23 73 34 119
rect 195 110 241 167
rect -103 27 -57 38
rect -103 -38 -57 -27
rect 57 27 103 38
rect 57 -38 103 -27
rect -241 -167 -195 -110
rect -34 -119 -23 -73
rect 23 -119 34 -73
rect 195 -167 241 -110
rect -241 -213 241 -167
<< properties >>
string FIXED_BBOX -218 -190 218 190
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.4 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
