magic
tech gf180mcuD
magscale 1 10
timestamp 1758101161
<< nwell >>
rect 6270 8915 7218 9835
rect 15742 8915 16690 9835
rect 25214 8916 26162 9836
rect 34686 8916 35634 9836
rect 44158 8916 45106 9836
rect 53630 8916 54578 9836
rect 6270 6710 7218 7630
rect 7756 6710 8704 7630
rect 15742 6710 16690 7630
rect 17228 6710 18176 7630
rect 25214 6711 26162 7631
rect 26700 6711 27648 7631
rect 34686 6711 35634 7631
rect 36172 6711 37120 7631
rect 44158 6711 45106 7631
rect 45644 6711 46592 7631
rect 53630 6711 54578 7631
rect 55116 6711 56064 7631
rect 6270 4505 7218 5425
rect 7756 4506 8704 5426
rect 1128 3290 1728 4310
rect 2016 3290 3096 4310
rect 15742 4505 16690 5425
rect 17228 4506 18176 5426
rect 25214 4506 26162 5426
rect 26700 4507 27648 5427
rect 10600 3290 11200 4310
rect 11488 3290 12568 4310
rect 20072 3291 20672 4311
rect 20960 3291 22040 4311
rect 34686 4506 35634 5426
rect 36172 4507 37120 5427
rect 29544 3291 30144 4311
rect 30432 3291 31512 4311
rect 44158 4506 45106 5426
rect 45644 4507 46592 5427
rect 39016 3291 39616 4311
rect 39904 3291 40984 4311
rect 53630 4506 54578 5426
rect 55116 4507 56064 5427
rect 48488 3291 49088 4311
rect 49376 3291 50456 4311
rect 234 1870 834 2890
rect 3356 2114 5324 3134
rect 6270 2300 7218 3220
rect 1128 950 1728 1970
rect 2016 950 3096 1970
rect 9706 1870 10306 2890
rect 12828 2114 14796 3134
rect 15742 2300 16690 3220
rect 10600 950 11200 1970
rect 11488 950 12568 1970
rect 19178 1871 19778 2891
rect 22300 2115 24268 3135
rect 25214 2301 26162 3221
rect 20072 951 20672 1971
rect 20960 951 22040 1971
rect 28650 1871 29250 2891
rect 31772 2115 33740 3135
rect 34686 2301 35634 3221
rect 29544 951 30144 1971
rect 30432 951 31512 1971
rect 38122 1871 38722 2891
rect 41244 2115 43212 3135
rect 44158 2301 45106 3221
rect 39016 951 39616 1971
rect 39904 951 40984 1971
rect 47594 1871 48194 2891
rect 50716 2115 52684 3135
rect 53630 2301 54578 3221
rect 48488 951 49088 1971
rect 49376 951 50456 1971
<< pwell >>
rect 7033 8675 7101 8915
rect 16505 8675 16573 8915
rect 25977 8676 26045 8916
rect 35449 8676 35517 8916
rect 44921 8676 44989 8916
rect 54393 8676 54461 8916
rect 6270 8055 7218 8675
rect 15742 8055 16690 8675
rect 25214 8056 26162 8676
rect 34686 8056 35634 8676
rect 44158 8056 45106 8676
rect 53630 8056 54578 8676
rect 7033 6470 7101 6710
rect 8519 6470 8587 6710
rect 16505 6470 16573 6710
rect 17991 6470 18059 6710
rect 25977 6471 26045 6711
rect 27463 6471 27531 6711
rect 35449 6471 35517 6711
rect 36935 6471 37003 6711
rect 44921 6471 44989 6711
rect 46407 6471 46475 6711
rect 54393 6471 54461 6711
rect 55879 6471 55947 6711
rect 6270 5850 7218 6470
rect 7756 5850 8704 6470
rect 15742 5850 16690 6470
rect 17228 5850 18176 6470
rect 25214 5851 26162 6471
rect 26700 5851 27648 6471
rect 34686 5851 35634 6471
rect 36172 5851 37120 6471
rect 44158 5851 45106 6471
rect 45644 5851 46592 6471
rect 53630 5851 54578 6471
rect 55116 5851 56064 6471
rect 7033 4265 7101 4505
rect 8519 4266 8587 4506
rect 6270 3645 7218 4265
rect 7756 3646 8704 4266
rect 16505 4265 16573 4505
rect 17991 4266 18059 4506
rect 15742 3645 16690 4265
rect 17228 3646 18176 4266
rect 25977 4266 26045 4506
rect 27463 4267 27531 4507
rect 25214 3646 26162 4266
rect 26700 3647 27648 4267
rect 35449 4266 35517 4506
rect 36935 4267 37003 4507
rect 34686 3646 35634 4266
rect 36172 3647 37120 4267
rect 44921 4266 44989 4506
rect 46407 4267 46475 4507
rect 44158 3646 45106 4266
rect 45644 3647 46592 4267
rect 54393 4266 54461 4506
rect 55879 4267 55947 4507
rect 53630 3646 54578 4266
rect 55116 3647 56064 4267
rect 2748 3201 2834 3281
rect 1128 2570 3096 3190
rect 12220 3201 12306 3281
rect 4976 2025 5062 2105
rect 7033 2060 7101 2300
rect 486 1781 572 1861
rect 234 1150 834 1770
rect 3356 1394 3956 2014
rect 4040 1924 4640 2014
rect 4040 1666 4686 1924
rect 4040 1394 4640 1666
rect 4724 1394 5324 2014
rect 6270 1440 7218 2060
rect 10600 2570 12568 3190
rect 21692 3202 21778 3282
rect 14448 2025 14534 2105
rect 16505 2060 16573 2300
rect 9958 1781 10044 1861
rect 9706 1150 10306 1770
rect 12828 1394 13428 2014
rect 13512 1924 14112 2014
rect 13512 1666 14158 1924
rect 13512 1394 14112 1666
rect 14196 1394 14796 2014
rect 15742 1440 16690 2060
rect 20072 2571 22040 3191
rect 31164 3202 31250 3282
rect 23920 2026 24006 2106
rect 25977 2061 26045 2301
rect 19430 1782 19516 1862
rect 19178 1151 19778 1771
rect 22300 1395 22900 2015
rect 22984 1925 23584 2015
rect 22984 1667 23630 1925
rect 22984 1395 23584 1667
rect 23668 1395 24268 2015
rect 25214 1441 26162 2061
rect 29544 2571 31512 3191
rect 40636 3202 40722 3282
rect 33392 2026 33478 2106
rect 35449 2061 35517 2301
rect 28902 1782 28988 1862
rect 28650 1151 29250 1771
rect 31772 1395 32372 2015
rect 32456 1925 33056 2015
rect 32456 1667 33102 1925
rect 32456 1395 33056 1667
rect 33140 1395 33740 2015
rect 34686 1441 35634 2061
rect 39016 2571 40984 3191
rect 50108 3202 50194 3282
rect 42864 2026 42950 2106
rect 44921 2061 44989 2301
rect 38374 1782 38460 1862
rect 38122 1151 38722 1771
rect 41244 1395 41844 2015
rect 41928 1925 42528 2015
rect 41928 1667 42574 1925
rect 41928 1395 42528 1667
rect 42612 1395 43212 2015
rect 44158 1441 45106 2061
rect 48488 2571 50456 3191
rect 52336 2026 52422 2106
rect 54393 2061 54461 2301
rect 47846 1782 47932 1862
rect 47594 1151 48194 1771
rect 50716 1395 51316 2015
rect 51400 1925 52000 2015
rect 51400 1667 52046 1925
rect 51400 1395 52000 1667
rect 52084 1395 52684 2015
rect 53630 1441 54578 2061
rect 2748 861 2834 941
rect 12220 861 12306 941
rect 21692 862 21778 942
rect 31164 862 31250 942
rect 40636 862 40722 942
rect 50108 862 50194 942
rect 1128 230 3096 850
rect 10600 230 12568 850
rect 20072 231 22040 851
rect 29544 231 31512 851
rect 39016 231 40984 851
rect 48488 231 50456 851
<< nmos >>
rect 6520 8265 6600 8465
rect 6704 8265 6784 8465
rect 6888 8265 6968 8465
rect 15992 8265 16072 8465
rect 16176 8265 16256 8465
rect 16360 8265 16440 8465
rect 25464 8266 25544 8466
rect 25648 8266 25728 8466
rect 25832 8266 25912 8466
rect 34936 8266 35016 8466
rect 35120 8266 35200 8466
rect 35304 8266 35384 8466
rect 44408 8266 44488 8466
rect 44592 8266 44672 8466
rect 44776 8266 44856 8466
rect 53880 8266 53960 8466
rect 54064 8266 54144 8466
rect 54248 8266 54328 8466
rect 6520 6060 6600 6260
rect 6704 6060 6784 6260
rect 6888 6060 6968 6260
rect 8006 6060 8086 6260
rect 8190 6060 8270 6260
rect 8374 6060 8454 6260
rect 15992 6060 16072 6260
rect 16176 6060 16256 6260
rect 16360 6060 16440 6260
rect 17478 6060 17558 6260
rect 17662 6060 17742 6260
rect 17846 6060 17926 6260
rect 25464 6061 25544 6261
rect 25648 6061 25728 6261
rect 25832 6061 25912 6261
rect 26950 6061 27030 6261
rect 27134 6061 27214 6261
rect 27318 6061 27398 6261
rect 34936 6061 35016 6261
rect 35120 6061 35200 6261
rect 35304 6061 35384 6261
rect 36422 6061 36502 6261
rect 36606 6061 36686 6261
rect 36790 6061 36870 6261
rect 44408 6061 44488 6261
rect 44592 6061 44672 6261
rect 44776 6061 44856 6261
rect 45894 6061 45974 6261
rect 46078 6061 46158 6261
rect 46262 6061 46342 6261
rect 53880 6061 53960 6261
rect 54064 6061 54144 6261
rect 54248 6061 54328 6261
rect 55366 6061 55446 6261
rect 55550 6061 55630 6261
rect 55734 6061 55814 6261
rect 6520 3855 6600 4055
rect 6704 3855 6784 4055
rect 6888 3855 6968 4055
rect 8006 3856 8086 4056
rect 8190 3856 8270 4056
rect 8374 3856 8454 4056
rect 15992 3855 16072 4055
rect 16176 3855 16256 4055
rect 16360 3855 16440 4055
rect 17478 3856 17558 4056
rect 17662 3856 17742 4056
rect 17846 3856 17926 4056
rect 25464 3856 25544 4056
rect 25648 3856 25728 4056
rect 25832 3856 25912 4056
rect 26950 3857 27030 4057
rect 27134 3857 27214 4057
rect 27318 3857 27398 4057
rect 34936 3856 35016 4056
rect 35120 3856 35200 4056
rect 35304 3856 35384 4056
rect 36422 3857 36502 4057
rect 36606 3857 36686 4057
rect 36790 3857 36870 4057
rect 44408 3856 44488 4056
rect 44592 3856 44672 4056
rect 44776 3856 44856 4056
rect 45894 3857 45974 4057
rect 46078 3857 46158 4057
rect 46262 3857 46342 4057
rect 53880 3856 53960 4056
rect 54064 3856 54144 4056
rect 54248 3856 54328 4056
rect 55366 3857 55446 4057
rect 55550 3857 55630 4057
rect 55734 3857 55814 4057
rect 1378 2780 1478 2980
rect 1582 2780 1682 2980
rect 2062 2780 2162 2980
rect 2266 2780 2366 2980
rect 2746 2780 2846 2980
rect 484 1360 584 1560
rect 3606 1604 3706 1804
rect 4290 1604 4390 1804
rect 4974 1604 5074 1804
rect 6520 1650 6600 1850
rect 6704 1650 6784 1850
rect 6888 1650 6968 1850
rect 10850 2780 10950 2980
rect 11054 2780 11154 2980
rect 11534 2780 11634 2980
rect 11738 2780 11838 2980
rect 12218 2780 12318 2980
rect 9956 1360 10056 1560
rect 13078 1604 13178 1804
rect 13762 1604 13862 1804
rect 14446 1604 14546 1804
rect 15992 1650 16072 1850
rect 16176 1650 16256 1850
rect 16360 1650 16440 1850
rect 20322 2781 20422 2981
rect 20526 2781 20626 2981
rect 21006 2781 21106 2981
rect 21210 2781 21310 2981
rect 21690 2781 21790 2981
rect 19428 1361 19528 1561
rect 22550 1605 22650 1805
rect 23234 1605 23334 1805
rect 23918 1605 24018 1805
rect 25464 1651 25544 1851
rect 25648 1651 25728 1851
rect 25832 1651 25912 1851
rect 29794 2781 29894 2981
rect 29998 2781 30098 2981
rect 30478 2781 30578 2981
rect 30682 2781 30782 2981
rect 31162 2781 31262 2981
rect 28900 1361 29000 1561
rect 32022 1605 32122 1805
rect 32706 1605 32806 1805
rect 33390 1605 33490 1805
rect 34936 1651 35016 1851
rect 35120 1651 35200 1851
rect 35304 1651 35384 1851
rect 39266 2781 39366 2981
rect 39470 2781 39570 2981
rect 39950 2781 40050 2981
rect 40154 2781 40254 2981
rect 40634 2781 40734 2981
rect 38372 1361 38472 1561
rect 41494 1605 41594 1805
rect 42178 1605 42278 1805
rect 42862 1605 42962 1805
rect 44408 1651 44488 1851
rect 44592 1651 44672 1851
rect 44776 1651 44856 1851
rect 48738 2781 48838 2981
rect 48942 2781 49042 2981
rect 49422 2781 49522 2981
rect 49626 2781 49726 2981
rect 50106 2781 50206 2981
rect 47844 1361 47944 1561
rect 50966 1605 51066 1805
rect 51650 1605 51750 1805
rect 52334 1605 52434 1805
rect 53880 1651 53960 1851
rect 54064 1651 54144 1851
rect 54248 1651 54328 1851
rect 1378 440 1478 640
rect 1582 440 1682 640
rect 2062 440 2162 640
rect 2266 440 2366 640
rect 2746 440 2846 640
rect 10850 440 10950 640
rect 11054 440 11154 640
rect 11534 440 11634 640
rect 11738 440 11838 640
rect 12218 440 12318 640
rect 20322 441 20422 641
rect 20526 441 20626 641
rect 21006 441 21106 641
rect 21210 441 21310 641
rect 21690 441 21790 641
rect 29794 441 29894 641
rect 29998 441 30098 641
rect 30478 441 30578 641
rect 30682 441 30782 641
rect 31162 441 31262 641
rect 39266 441 39366 641
rect 39470 441 39570 641
rect 39950 441 40050 641
rect 40154 441 40254 641
rect 40634 441 40734 641
rect 48738 441 48838 641
rect 48942 441 49042 641
rect 49422 441 49522 641
rect 49626 441 49726 641
rect 50106 441 50206 641
<< pmos >>
rect 6520 9125 6600 9625
rect 6704 9125 6784 9625
rect 6888 9125 6968 9625
rect 15992 9125 16072 9625
rect 16176 9125 16256 9625
rect 16360 9125 16440 9625
rect 25464 9126 25544 9626
rect 25648 9126 25728 9626
rect 25832 9126 25912 9626
rect 34936 9126 35016 9626
rect 35120 9126 35200 9626
rect 35304 9126 35384 9626
rect 44408 9126 44488 9626
rect 44592 9126 44672 9626
rect 44776 9126 44856 9626
rect 53880 9126 53960 9626
rect 54064 9126 54144 9626
rect 54248 9126 54328 9626
rect 6520 6920 6600 7420
rect 6704 6920 6784 7420
rect 6888 6920 6968 7420
rect 8006 6920 8086 7420
rect 8190 6920 8270 7420
rect 8374 6920 8454 7420
rect 15992 6920 16072 7420
rect 16176 6920 16256 7420
rect 16360 6920 16440 7420
rect 17478 6920 17558 7420
rect 17662 6920 17742 7420
rect 17846 6920 17926 7420
rect 25464 6921 25544 7421
rect 25648 6921 25728 7421
rect 25832 6921 25912 7421
rect 26950 6921 27030 7421
rect 27134 6921 27214 7421
rect 27318 6921 27398 7421
rect 34936 6921 35016 7421
rect 35120 6921 35200 7421
rect 35304 6921 35384 7421
rect 36422 6921 36502 7421
rect 36606 6921 36686 7421
rect 36790 6921 36870 7421
rect 44408 6921 44488 7421
rect 44592 6921 44672 7421
rect 44776 6921 44856 7421
rect 45894 6921 45974 7421
rect 46078 6921 46158 7421
rect 46262 6921 46342 7421
rect 53880 6921 53960 7421
rect 54064 6921 54144 7421
rect 54248 6921 54328 7421
rect 55366 6921 55446 7421
rect 55550 6921 55630 7421
rect 55734 6921 55814 7421
rect 6520 4715 6600 5215
rect 6704 4715 6784 5215
rect 6888 4715 6968 5215
rect 8006 4716 8086 5216
rect 8190 4716 8270 5216
rect 8374 4716 8454 5216
rect 15992 4715 16072 5215
rect 16176 4715 16256 5215
rect 16360 4715 16440 5215
rect 17478 4716 17558 5216
rect 17662 4716 17742 5216
rect 17846 4716 17926 5216
rect 25464 4716 25544 5216
rect 25648 4716 25728 5216
rect 25832 4716 25912 5216
rect 26950 4717 27030 5217
rect 27134 4717 27214 5217
rect 27318 4717 27398 5217
rect 34936 4716 35016 5216
rect 35120 4716 35200 5216
rect 35304 4716 35384 5216
rect 36422 4717 36502 5217
rect 36606 4717 36686 5217
rect 36790 4717 36870 5217
rect 44408 4716 44488 5216
rect 44592 4716 44672 5216
rect 44776 4716 44856 5216
rect 45894 4717 45974 5217
rect 46078 4717 46158 5217
rect 46262 4717 46342 5217
rect 53880 4716 53960 5216
rect 54064 4716 54144 5216
rect 54248 4716 54328 5216
rect 55366 4717 55446 5217
rect 55550 4717 55630 5217
rect 55734 4717 55814 5217
rect 1378 3500 1478 4100
rect 2266 3500 2366 4100
rect 2746 3500 2846 4100
rect 10850 3500 10950 4100
rect 11738 3500 11838 4100
rect 12218 3500 12318 4100
rect 20322 3501 20422 4101
rect 21210 3501 21310 4101
rect 21690 3501 21790 4101
rect 29794 3501 29894 4101
rect 30682 3501 30782 4101
rect 31162 3501 31262 4101
rect 39266 3501 39366 4101
rect 40154 3501 40254 4101
rect 40634 3501 40734 4101
rect 48738 3501 48838 4101
rect 49626 3501 49726 4101
rect 50106 3501 50206 4101
rect 484 2080 584 2680
rect 3606 2324 3706 2924
rect 3810 2324 3910 2924
rect 4290 2324 4390 2924
rect 4494 2324 4594 2924
rect 4974 2324 5074 2924
rect 6520 2510 6600 3010
rect 6704 2510 6784 3010
rect 6888 2510 6968 3010
rect 1378 1160 1478 1760
rect 2266 1160 2366 1760
rect 2746 1160 2846 1760
rect 9956 2080 10056 2680
rect 13078 2324 13178 2924
rect 13282 2324 13382 2924
rect 13762 2324 13862 2924
rect 13966 2324 14066 2924
rect 14446 2324 14546 2924
rect 15992 2510 16072 3010
rect 16176 2510 16256 3010
rect 16360 2510 16440 3010
rect 10850 1160 10950 1760
rect 11738 1160 11838 1760
rect 12218 1160 12318 1760
rect 19428 2081 19528 2681
rect 22550 2325 22650 2925
rect 22754 2325 22854 2925
rect 23234 2325 23334 2925
rect 23438 2325 23538 2925
rect 23918 2325 24018 2925
rect 25464 2511 25544 3011
rect 25648 2511 25728 3011
rect 25832 2511 25912 3011
rect 20322 1161 20422 1761
rect 21210 1161 21310 1761
rect 21690 1161 21790 1761
rect 28900 2081 29000 2681
rect 32022 2325 32122 2925
rect 32226 2325 32326 2925
rect 32706 2325 32806 2925
rect 32910 2325 33010 2925
rect 33390 2325 33490 2925
rect 34936 2511 35016 3011
rect 35120 2511 35200 3011
rect 35304 2511 35384 3011
rect 29794 1161 29894 1761
rect 30682 1161 30782 1761
rect 31162 1161 31262 1761
rect 38372 2081 38472 2681
rect 41494 2325 41594 2925
rect 41698 2325 41798 2925
rect 42178 2325 42278 2925
rect 42382 2325 42482 2925
rect 42862 2325 42962 2925
rect 44408 2511 44488 3011
rect 44592 2511 44672 3011
rect 44776 2511 44856 3011
rect 39266 1161 39366 1761
rect 40154 1161 40254 1761
rect 40634 1161 40734 1761
rect 47844 2081 47944 2681
rect 50966 2325 51066 2925
rect 51170 2325 51270 2925
rect 51650 2325 51750 2925
rect 51854 2325 51954 2925
rect 52334 2325 52434 2925
rect 53880 2511 53960 3011
rect 54064 2511 54144 3011
rect 54248 2511 54328 3011
rect 48738 1161 48838 1761
rect 49626 1161 49726 1761
rect 50106 1161 50206 1761
<< ndiff >>
rect 6432 8452 6520 8465
rect 6432 8278 6445 8452
rect 6491 8278 6520 8452
rect 6432 8265 6520 8278
rect 6600 8452 6704 8465
rect 6600 8278 6629 8452
rect 6675 8278 6704 8452
rect 6600 8265 6704 8278
rect 6784 8452 6888 8465
rect 6784 8278 6813 8452
rect 6859 8278 6888 8452
rect 6784 8265 6888 8278
rect 6968 8452 7056 8465
rect 6968 8278 6997 8452
rect 7043 8278 7056 8452
rect 6968 8265 7056 8278
rect 15904 8452 15992 8465
rect 15904 8278 15917 8452
rect 15963 8278 15992 8452
rect 15904 8265 15992 8278
rect 16072 8452 16176 8465
rect 16072 8278 16101 8452
rect 16147 8278 16176 8452
rect 16072 8265 16176 8278
rect 16256 8452 16360 8465
rect 16256 8278 16285 8452
rect 16331 8278 16360 8452
rect 16256 8265 16360 8278
rect 16440 8452 16528 8465
rect 16440 8278 16469 8452
rect 16515 8278 16528 8452
rect 16440 8265 16528 8278
rect 25376 8453 25464 8466
rect 25376 8279 25389 8453
rect 25435 8279 25464 8453
rect 25376 8266 25464 8279
rect 25544 8453 25648 8466
rect 25544 8279 25573 8453
rect 25619 8279 25648 8453
rect 25544 8266 25648 8279
rect 25728 8453 25832 8466
rect 25728 8279 25757 8453
rect 25803 8279 25832 8453
rect 25728 8266 25832 8279
rect 25912 8453 26000 8466
rect 25912 8279 25941 8453
rect 25987 8279 26000 8453
rect 25912 8266 26000 8279
rect 34848 8453 34936 8466
rect 34848 8279 34861 8453
rect 34907 8279 34936 8453
rect 34848 8266 34936 8279
rect 35016 8453 35120 8466
rect 35016 8279 35045 8453
rect 35091 8279 35120 8453
rect 35016 8266 35120 8279
rect 35200 8453 35304 8466
rect 35200 8279 35229 8453
rect 35275 8279 35304 8453
rect 35200 8266 35304 8279
rect 35384 8453 35472 8466
rect 35384 8279 35413 8453
rect 35459 8279 35472 8453
rect 35384 8266 35472 8279
rect 44320 8453 44408 8466
rect 44320 8279 44333 8453
rect 44379 8279 44408 8453
rect 44320 8266 44408 8279
rect 44488 8453 44592 8466
rect 44488 8279 44517 8453
rect 44563 8279 44592 8453
rect 44488 8266 44592 8279
rect 44672 8453 44776 8466
rect 44672 8279 44701 8453
rect 44747 8279 44776 8453
rect 44672 8266 44776 8279
rect 44856 8453 44944 8466
rect 44856 8279 44885 8453
rect 44931 8279 44944 8453
rect 44856 8266 44944 8279
rect 53792 8453 53880 8466
rect 53792 8279 53805 8453
rect 53851 8279 53880 8453
rect 53792 8266 53880 8279
rect 53960 8453 54064 8466
rect 53960 8279 53989 8453
rect 54035 8279 54064 8453
rect 53960 8266 54064 8279
rect 54144 8453 54248 8466
rect 54144 8279 54173 8453
rect 54219 8279 54248 8453
rect 54144 8266 54248 8279
rect 54328 8453 54416 8466
rect 54328 8279 54357 8453
rect 54403 8279 54416 8453
rect 54328 8266 54416 8279
rect 6432 6247 6520 6260
rect 6432 6073 6445 6247
rect 6491 6073 6520 6247
rect 6432 6060 6520 6073
rect 6600 6247 6704 6260
rect 6600 6073 6629 6247
rect 6675 6073 6704 6247
rect 6600 6060 6704 6073
rect 6784 6247 6888 6260
rect 6784 6073 6813 6247
rect 6859 6073 6888 6247
rect 6784 6060 6888 6073
rect 6968 6247 7056 6260
rect 6968 6073 6997 6247
rect 7043 6073 7056 6247
rect 6968 6060 7056 6073
rect 7918 6247 8006 6260
rect 7918 6073 7931 6247
rect 7977 6073 8006 6247
rect 7918 6060 8006 6073
rect 8086 6247 8190 6260
rect 8086 6073 8115 6247
rect 8161 6073 8190 6247
rect 8086 6060 8190 6073
rect 8270 6247 8374 6260
rect 8270 6073 8299 6247
rect 8345 6073 8374 6247
rect 8270 6060 8374 6073
rect 8454 6247 8542 6260
rect 8454 6073 8483 6247
rect 8529 6073 8542 6247
rect 8454 6060 8542 6073
rect 15904 6247 15992 6260
rect 15904 6073 15917 6247
rect 15963 6073 15992 6247
rect 15904 6060 15992 6073
rect 16072 6247 16176 6260
rect 16072 6073 16101 6247
rect 16147 6073 16176 6247
rect 16072 6060 16176 6073
rect 16256 6247 16360 6260
rect 16256 6073 16285 6247
rect 16331 6073 16360 6247
rect 16256 6060 16360 6073
rect 16440 6247 16528 6260
rect 16440 6073 16469 6247
rect 16515 6073 16528 6247
rect 16440 6060 16528 6073
rect 17390 6247 17478 6260
rect 17390 6073 17403 6247
rect 17449 6073 17478 6247
rect 17390 6060 17478 6073
rect 17558 6247 17662 6260
rect 17558 6073 17587 6247
rect 17633 6073 17662 6247
rect 17558 6060 17662 6073
rect 17742 6247 17846 6260
rect 17742 6073 17771 6247
rect 17817 6073 17846 6247
rect 17742 6060 17846 6073
rect 17926 6247 18014 6260
rect 17926 6073 17955 6247
rect 18001 6073 18014 6247
rect 17926 6060 18014 6073
rect 25376 6248 25464 6261
rect 25376 6074 25389 6248
rect 25435 6074 25464 6248
rect 25376 6061 25464 6074
rect 25544 6248 25648 6261
rect 25544 6074 25573 6248
rect 25619 6074 25648 6248
rect 25544 6061 25648 6074
rect 25728 6248 25832 6261
rect 25728 6074 25757 6248
rect 25803 6074 25832 6248
rect 25728 6061 25832 6074
rect 25912 6248 26000 6261
rect 25912 6074 25941 6248
rect 25987 6074 26000 6248
rect 25912 6061 26000 6074
rect 26862 6248 26950 6261
rect 26862 6074 26875 6248
rect 26921 6074 26950 6248
rect 26862 6061 26950 6074
rect 27030 6248 27134 6261
rect 27030 6074 27059 6248
rect 27105 6074 27134 6248
rect 27030 6061 27134 6074
rect 27214 6248 27318 6261
rect 27214 6074 27243 6248
rect 27289 6074 27318 6248
rect 27214 6061 27318 6074
rect 27398 6248 27486 6261
rect 27398 6074 27427 6248
rect 27473 6074 27486 6248
rect 27398 6061 27486 6074
rect 34848 6248 34936 6261
rect 34848 6074 34861 6248
rect 34907 6074 34936 6248
rect 34848 6061 34936 6074
rect 35016 6248 35120 6261
rect 35016 6074 35045 6248
rect 35091 6074 35120 6248
rect 35016 6061 35120 6074
rect 35200 6248 35304 6261
rect 35200 6074 35229 6248
rect 35275 6074 35304 6248
rect 35200 6061 35304 6074
rect 35384 6248 35472 6261
rect 35384 6074 35413 6248
rect 35459 6074 35472 6248
rect 35384 6061 35472 6074
rect 36334 6248 36422 6261
rect 36334 6074 36347 6248
rect 36393 6074 36422 6248
rect 36334 6061 36422 6074
rect 36502 6248 36606 6261
rect 36502 6074 36531 6248
rect 36577 6074 36606 6248
rect 36502 6061 36606 6074
rect 36686 6248 36790 6261
rect 36686 6074 36715 6248
rect 36761 6074 36790 6248
rect 36686 6061 36790 6074
rect 36870 6248 36958 6261
rect 36870 6074 36899 6248
rect 36945 6074 36958 6248
rect 36870 6061 36958 6074
rect 44320 6248 44408 6261
rect 44320 6074 44333 6248
rect 44379 6074 44408 6248
rect 44320 6061 44408 6074
rect 44488 6248 44592 6261
rect 44488 6074 44517 6248
rect 44563 6074 44592 6248
rect 44488 6061 44592 6074
rect 44672 6248 44776 6261
rect 44672 6074 44701 6248
rect 44747 6074 44776 6248
rect 44672 6061 44776 6074
rect 44856 6248 44944 6261
rect 44856 6074 44885 6248
rect 44931 6074 44944 6248
rect 44856 6061 44944 6074
rect 45806 6248 45894 6261
rect 45806 6074 45819 6248
rect 45865 6074 45894 6248
rect 45806 6061 45894 6074
rect 45974 6248 46078 6261
rect 45974 6074 46003 6248
rect 46049 6074 46078 6248
rect 45974 6061 46078 6074
rect 46158 6248 46262 6261
rect 46158 6074 46187 6248
rect 46233 6074 46262 6248
rect 46158 6061 46262 6074
rect 46342 6248 46430 6261
rect 46342 6074 46371 6248
rect 46417 6074 46430 6248
rect 46342 6061 46430 6074
rect 53792 6248 53880 6261
rect 53792 6074 53805 6248
rect 53851 6074 53880 6248
rect 53792 6061 53880 6074
rect 53960 6248 54064 6261
rect 53960 6074 53989 6248
rect 54035 6074 54064 6248
rect 53960 6061 54064 6074
rect 54144 6248 54248 6261
rect 54144 6074 54173 6248
rect 54219 6074 54248 6248
rect 54144 6061 54248 6074
rect 54328 6248 54416 6261
rect 54328 6074 54357 6248
rect 54403 6074 54416 6248
rect 54328 6061 54416 6074
rect 55278 6248 55366 6261
rect 55278 6074 55291 6248
rect 55337 6074 55366 6248
rect 55278 6061 55366 6074
rect 55446 6248 55550 6261
rect 55446 6074 55475 6248
rect 55521 6074 55550 6248
rect 55446 6061 55550 6074
rect 55630 6248 55734 6261
rect 55630 6074 55659 6248
rect 55705 6074 55734 6248
rect 55630 6061 55734 6074
rect 55814 6248 55902 6261
rect 55814 6074 55843 6248
rect 55889 6074 55902 6248
rect 55814 6061 55902 6074
rect 6432 4042 6520 4055
rect 6432 3868 6445 4042
rect 6491 3868 6520 4042
rect 6432 3855 6520 3868
rect 6600 4042 6704 4055
rect 6600 3868 6629 4042
rect 6675 3868 6704 4042
rect 6600 3855 6704 3868
rect 6784 4042 6888 4055
rect 6784 3868 6813 4042
rect 6859 3868 6888 4042
rect 6784 3855 6888 3868
rect 6968 4042 7056 4055
rect 6968 3868 6997 4042
rect 7043 3868 7056 4042
rect 6968 3855 7056 3868
rect 7918 4043 8006 4056
rect 7918 3869 7931 4043
rect 7977 3869 8006 4043
rect 7918 3856 8006 3869
rect 8086 4043 8190 4056
rect 8086 3869 8115 4043
rect 8161 3869 8190 4043
rect 8086 3856 8190 3869
rect 8270 4043 8374 4056
rect 8270 3869 8299 4043
rect 8345 3869 8374 4043
rect 8270 3856 8374 3869
rect 8454 4043 8542 4056
rect 8454 3869 8483 4043
rect 8529 3869 8542 4043
rect 8454 3856 8542 3869
rect 15904 4042 15992 4055
rect 15904 3868 15917 4042
rect 15963 3868 15992 4042
rect 15904 3855 15992 3868
rect 16072 4042 16176 4055
rect 16072 3868 16101 4042
rect 16147 3868 16176 4042
rect 16072 3855 16176 3868
rect 16256 4042 16360 4055
rect 16256 3868 16285 4042
rect 16331 3868 16360 4042
rect 16256 3855 16360 3868
rect 16440 4042 16528 4055
rect 16440 3868 16469 4042
rect 16515 3868 16528 4042
rect 16440 3855 16528 3868
rect 17390 4043 17478 4056
rect 17390 3869 17403 4043
rect 17449 3869 17478 4043
rect 17390 3856 17478 3869
rect 17558 4043 17662 4056
rect 17558 3869 17587 4043
rect 17633 3869 17662 4043
rect 17558 3856 17662 3869
rect 17742 4043 17846 4056
rect 17742 3869 17771 4043
rect 17817 3869 17846 4043
rect 17742 3856 17846 3869
rect 17926 4043 18014 4056
rect 17926 3869 17955 4043
rect 18001 3869 18014 4043
rect 17926 3856 18014 3869
rect 25376 4043 25464 4056
rect 25376 3869 25389 4043
rect 25435 3869 25464 4043
rect 25376 3856 25464 3869
rect 25544 4043 25648 4056
rect 25544 3869 25573 4043
rect 25619 3869 25648 4043
rect 25544 3856 25648 3869
rect 25728 4043 25832 4056
rect 25728 3869 25757 4043
rect 25803 3869 25832 4043
rect 25728 3856 25832 3869
rect 25912 4043 26000 4056
rect 25912 3869 25941 4043
rect 25987 3869 26000 4043
rect 25912 3856 26000 3869
rect 26862 4044 26950 4057
rect 26862 3870 26875 4044
rect 26921 3870 26950 4044
rect 26862 3857 26950 3870
rect 27030 4044 27134 4057
rect 27030 3870 27059 4044
rect 27105 3870 27134 4044
rect 27030 3857 27134 3870
rect 27214 4044 27318 4057
rect 27214 3870 27243 4044
rect 27289 3870 27318 4044
rect 27214 3857 27318 3870
rect 27398 4044 27486 4057
rect 27398 3870 27427 4044
rect 27473 3870 27486 4044
rect 27398 3857 27486 3870
rect 34848 4043 34936 4056
rect 34848 3869 34861 4043
rect 34907 3869 34936 4043
rect 34848 3856 34936 3869
rect 35016 4043 35120 4056
rect 35016 3869 35045 4043
rect 35091 3869 35120 4043
rect 35016 3856 35120 3869
rect 35200 4043 35304 4056
rect 35200 3869 35229 4043
rect 35275 3869 35304 4043
rect 35200 3856 35304 3869
rect 35384 4043 35472 4056
rect 35384 3869 35413 4043
rect 35459 3869 35472 4043
rect 35384 3856 35472 3869
rect 36334 4044 36422 4057
rect 36334 3870 36347 4044
rect 36393 3870 36422 4044
rect 36334 3857 36422 3870
rect 36502 4044 36606 4057
rect 36502 3870 36531 4044
rect 36577 3870 36606 4044
rect 36502 3857 36606 3870
rect 36686 4044 36790 4057
rect 36686 3870 36715 4044
rect 36761 3870 36790 4044
rect 36686 3857 36790 3870
rect 36870 4044 36958 4057
rect 36870 3870 36899 4044
rect 36945 3870 36958 4044
rect 36870 3857 36958 3870
rect 44320 4043 44408 4056
rect 44320 3869 44333 4043
rect 44379 3869 44408 4043
rect 44320 3856 44408 3869
rect 44488 4043 44592 4056
rect 44488 3869 44517 4043
rect 44563 3869 44592 4043
rect 44488 3856 44592 3869
rect 44672 4043 44776 4056
rect 44672 3869 44701 4043
rect 44747 3869 44776 4043
rect 44672 3856 44776 3869
rect 44856 4043 44944 4056
rect 44856 3869 44885 4043
rect 44931 3869 44944 4043
rect 44856 3856 44944 3869
rect 45806 4044 45894 4057
rect 45806 3870 45819 4044
rect 45865 3870 45894 4044
rect 45806 3857 45894 3870
rect 45974 4044 46078 4057
rect 45974 3870 46003 4044
rect 46049 3870 46078 4044
rect 45974 3857 46078 3870
rect 46158 4044 46262 4057
rect 46158 3870 46187 4044
rect 46233 3870 46262 4044
rect 46158 3857 46262 3870
rect 46342 4044 46430 4057
rect 46342 3870 46371 4044
rect 46417 3870 46430 4044
rect 46342 3857 46430 3870
rect 53792 4043 53880 4056
rect 53792 3869 53805 4043
rect 53851 3869 53880 4043
rect 53792 3856 53880 3869
rect 53960 4043 54064 4056
rect 53960 3869 53989 4043
rect 54035 3869 54064 4043
rect 53960 3856 54064 3869
rect 54144 4043 54248 4056
rect 54144 3869 54173 4043
rect 54219 3869 54248 4043
rect 54144 3856 54248 3869
rect 54328 4043 54416 4056
rect 54328 3869 54357 4043
rect 54403 3869 54416 4043
rect 54328 3856 54416 3869
rect 55278 4044 55366 4057
rect 55278 3870 55291 4044
rect 55337 3870 55366 4044
rect 55278 3857 55366 3870
rect 55446 4044 55550 4057
rect 55446 3870 55475 4044
rect 55521 3870 55550 4044
rect 55446 3857 55550 3870
rect 55630 4044 55734 4057
rect 55630 3870 55659 4044
rect 55705 3870 55734 4044
rect 55630 3857 55734 3870
rect 55814 4044 55902 4057
rect 55814 3870 55843 4044
rect 55889 3870 55902 4044
rect 55814 3857 55902 3870
rect 1290 2967 1378 2980
rect 1290 2793 1303 2967
rect 1349 2793 1378 2967
rect 1290 2780 1378 2793
rect 1478 2967 1582 2980
rect 1478 2793 1507 2967
rect 1553 2793 1582 2967
rect 1478 2780 1582 2793
rect 1682 2967 1770 2980
rect 1682 2793 1711 2967
rect 1757 2793 1770 2967
rect 1682 2780 1770 2793
rect 1974 2967 2062 2980
rect 1974 2793 1987 2967
rect 2033 2793 2062 2967
rect 1974 2780 2062 2793
rect 2162 2967 2266 2980
rect 2162 2793 2191 2967
rect 2237 2793 2266 2967
rect 2162 2780 2266 2793
rect 2366 2967 2454 2980
rect 2366 2793 2395 2967
rect 2441 2793 2454 2967
rect 2366 2780 2454 2793
rect 2658 2967 2746 2980
rect 2658 2793 2671 2967
rect 2717 2793 2746 2967
rect 2658 2780 2746 2793
rect 2846 2967 2934 2980
rect 2846 2793 2875 2967
rect 2921 2793 2934 2967
rect 2846 2780 2934 2793
rect 396 1547 484 1560
rect 396 1373 409 1547
rect 455 1373 484 1547
rect 396 1360 484 1373
rect 584 1547 672 1560
rect 584 1373 613 1547
rect 659 1373 672 1547
rect 584 1360 672 1373
rect 3518 1791 3606 1804
rect 3518 1617 3531 1791
rect 3577 1617 3606 1791
rect 3518 1604 3606 1617
rect 3706 1791 3794 1804
rect 3706 1617 3735 1791
rect 3781 1617 3794 1791
rect 3706 1604 3794 1617
rect 4202 1791 4290 1804
rect 4202 1617 4215 1791
rect 4261 1617 4290 1791
rect 4202 1604 4290 1617
rect 4390 1791 4478 1804
rect 4390 1617 4419 1791
rect 4465 1617 4478 1791
rect 4390 1604 4478 1617
rect 4886 1791 4974 1804
rect 4886 1617 4899 1791
rect 4945 1617 4974 1791
rect 4886 1604 4974 1617
rect 5074 1791 5162 1804
rect 5074 1617 5103 1791
rect 5149 1617 5162 1791
rect 5074 1604 5162 1617
rect 6432 1837 6520 1850
rect 6432 1663 6445 1837
rect 6491 1663 6520 1837
rect 6432 1650 6520 1663
rect 6600 1837 6704 1850
rect 6600 1663 6629 1837
rect 6675 1663 6704 1837
rect 6600 1650 6704 1663
rect 6784 1837 6888 1850
rect 6784 1663 6813 1837
rect 6859 1663 6888 1837
rect 6784 1650 6888 1663
rect 6968 1837 7056 1850
rect 6968 1663 6997 1837
rect 7043 1663 7056 1837
rect 6968 1650 7056 1663
rect 10762 2967 10850 2980
rect 10762 2793 10775 2967
rect 10821 2793 10850 2967
rect 10762 2780 10850 2793
rect 10950 2967 11054 2980
rect 10950 2793 10979 2967
rect 11025 2793 11054 2967
rect 10950 2780 11054 2793
rect 11154 2967 11242 2980
rect 11154 2793 11183 2967
rect 11229 2793 11242 2967
rect 11154 2780 11242 2793
rect 11446 2967 11534 2980
rect 11446 2793 11459 2967
rect 11505 2793 11534 2967
rect 11446 2780 11534 2793
rect 11634 2967 11738 2980
rect 11634 2793 11663 2967
rect 11709 2793 11738 2967
rect 11634 2780 11738 2793
rect 11838 2967 11926 2980
rect 11838 2793 11867 2967
rect 11913 2793 11926 2967
rect 11838 2780 11926 2793
rect 12130 2967 12218 2980
rect 12130 2793 12143 2967
rect 12189 2793 12218 2967
rect 12130 2780 12218 2793
rect 12318 2967 12406 2980
rect 12318 2793 12347 2967
rect 12393 2793 12406 2967
rect 12318 2780 12406 2793
rect 9868 1547 9956 1560
rect 9868 1373 9881 1547
rect 9927 1373 9956 1547
rect 9868 1360 9956 1373
rect 10056 1547 10144 1560
rect 10056 1373 10085 1547
rect 10131 1373 10144 1547
rect 10056 1360 10144 1373
rect 12990 1791 13078 1804
rect 12990 1617 13003 1791
rect 13049 1617 13078 1791
rect 12990 1604 13078 1617
rect 13178 1791 13266 1804
rect 13178 1617 13207 1791
rect 13253 1617 13266 1791
rect 13178 1604 13266 1617
rect 13674 1791 13762 1804
rect 13674 1617 13687 1791
rect 13733 1617 13762 1791
rect 13674 1604 13762 1617
rect 13862 1791 13950 1804
rect 13862 1617 13891 1791
rect 13937 1617 13950 1791
rect 13862 1604 13950 1617
rect 14358 1791 14446 1804
rect 14358 1617 14371 1791
rect 14417 1617 14446 1791
rect 14358 1604 14446 1617
rect 14546 1791 14634 1804
rect 14546 1617 14575 1791
rect 14621 1617 14634 1791
rect 14546 1604 14634 1617
rect 15904 1837 15992 1850
rect 15904 1663 15917 1837
rect 15963 1663 15992 1837
rect 15904 1650 15992 1663
rect 16072 1837 16176 1850
rect 16072 1663 16101 1837
rect 16147 1663 16176 1837
rect 16072 1650 16176 1663
rect 16256 1837 16360 1850
rect 16256 1663 16285 1837
rect 16331 1663 16360 1837
rect 16256 1650 16360 1663
rect 16440 1837 16528 1850
rect 16440 1663 16469 1837
rect 16515 1663 16528 1837
rect 16440 1650 16528 1663
rect 20234 2968 20322 2981
rect 20234 2794 20247 2968
rect 20293 2794 20322 2968
rect 20234 2781 20322 2794
rect 20422 2968 20526 2981
rect 20422 2794 20451 2968
rect 20497 2794 20526 2968
rect 20422 2781 20526 2794
rect 20626 2968 20714 2981
rect 20626 2794 20655 2968
rect 20701 2794 20714 2968
rect 20626 2781 20714 2794
rect 20918 2968 21006 2981
rect 20918 2794 20931 2968
rect 20977 2794 21006 2968
rect 20918 2781 21006 2794
rect 21106 2968 21210 2981
rect 21106 2794 21135 2968
rect 21181 2794 21210 2968
rect 21106 2781 21210 2794
rect 21310 2968 21398 2981
rect 21310 2794 21339 2968
rect 21385 2794 21398 2968
rect 21310 2781 21398 2794
rect 21602 2968 21690 2981
rect 21602 2794 21615 2968
rect 21661 2794 21690 2968
rect 21602 2781 21690 2794
rect 21790 2968 21878 2981
rect 21790 2794 21819 2968
rect 21865 2794 21878 2968
rect 21790 2781 21878 2794
rect 19340 1548 19428 1561
rect 19340 1374 19353 1548
rect 19399 1374 19428 1548
rect 19340 1361 19428 1374
rect 19528 1548 19616 1561
rect 19528 1374 19557 1548
rect 19603 1374 19616 1548
rect 19528 1361 19616 1374
rect 22462 1792 22550 1805
rect 22462 1618 22475 1792
rect 22521 1618 22550 1792
rect 22462 1605 22550 1618
rect 22650 1792 22738 1805
rect 22650 1618 22679 1792
rect 22725 1618 22738 1792
rect 22650 1605 22738 1618
rect 23146 1792 23234 1805
rect 23146 1618 23159 1792
rect 23205 1618 23234 1792
rect 23146 1605 23234 1618
rect 23334 1792 23422 1805
rect 23334 1618 23363 1792
rect 23409 1618 23422 1792
rect 23334 1605 23422 1618
rect 23830 1792 23918 1805
rect 23830 1618 23843 1792
rect 23889 1618 23918 1792
rect 23830 1605 23918 1618
rect 24018 1792 24106 1805
rect 24018 1618 24047 1792
rect 24093 1618 24106 1792
rect 24018 1605 24106 1618
rect 25376 1838 25464 1851
rect 25376 1664 25389 1838
rect 25435 1664 25464 1838
rect 25376 1651 25464 1664
rect 25544 1838 25648 1851
rect 25544 1664 25573 1838
rect 25619 1664 25648 1838
rect 25544 1651 25648 1664
rect 25728 1838 25832 1851
rect 25728 1664 25757 1838
rect 25803 1664 25832 1838
rect 25728 1651 25832 1664
rect 25912 1838 26000 1851
rect 25912 1664 25941 1838
rect 25987 1664 26000 1838
rect 25912 1651 26000 1664
rect 29706 2968 29794 2981
rect 29706 2794 29719 2968
rect 29765 2794 29794 2968
rect 29706 2781 29794 2794
rect 29894 2968 29998 2981
rect 29894 2794 29923 2968
rect 29969 2794 29998 2968
rect 29894 2781 29998 2794
rect 30098 2968 30186 2981
rect 30098 2794 30127 2968
rect 30173 2794 30186 2968
rect 30098 2781 30186 2794
rect 30390 2968 30478 2981
rect 30390 2794 30403 2968
rect 30449 2794 30478 2968
rect 30390 2781 30478 2794
rect 30578 2968 30682 2981
rect 30578 2794 30607 2968
rect 30653 2794 30682 2968
rect 30578 2781 30682 2794
rect 30782 2968 30870 2981
rect 30782 2794 30811 2968
rect 30857 2794 30870 2968
rect 30782 2781 30870 2794
rect 31074 2968 31162 2981
rect 31074 2794 31087 2968
rect 31133 2794 31162 2968
rect 31074 2781 31162 2794
rect 31262 2968 31350 2981
rect 31262 2794 31291 2968
rect 31337 2794 31350 2968
rect 31262 2781 31350 2794
rect 28812 1548 28900 1561
rect 28812 1374 28825 1548
rect 28871 1374 28900 1548
rect 28812 1361 28900 1374
rect 29000 1548 29088 1561
rect 29000 1374 29029 1548
rect 29075 1374 29088 1548
rect 29000 1361 29088 1374
rect 31934 1792 32022 1805
rect 31934 1618 31947 1792
rect 31993 1618 32022 1792
rect 31934 1605 32022 1618
rect 32122 1792 32210 1805
rect 32122 1618 32151 1792
rect 32197 1618 32210 1792
rect 32122 1605 32210 1618
rect 32618 1792 32706 1805
rect 32618 1618 32631 1792
rect 32677 1618 32706 1792
rect 32618 1605 32706 1618
rect 32806 1792 32894 1805
rect 32806 1618 32835 1792
rect 32881 1618 32894 1792
rect 32806 1605 32894 1618
rect 33302 1792 33390 1805
rect 33302 1618 33315 1792
rect 33361 1618 33390 1792
rect 33302 1605 33390 1618
rect 33490 1792 33578 1805
rect 33490 1618 33519 1792
rect 33565 1618 33578 1792
rect 33490 1605 33578 1618
rect 34848 1838 34936 1851
rect 34848 1664 34861 1838
rect 34907 1664 34936 1838
rect 34848 1651 34936 1664
rect 35016 1838 35120 1851
rect 35016 1664 35045 1838
rect 35091 1664 35120 1838
rect 35016 1651 35120 1664
rect 35200 1838 35304 1851
rect 35200 1664 35229 1838
rect 35275 1664 35304 1838
rect 35200 1651 35304 1664
rect 35384 1838 35472 1851
rect 35384 1664 35413 1838
rect 35459 1664 35472 1838
rect 35384 1651 35472 1664
rect 39178 2968 39266 2981
rect 39178 2794 39191 2968
rect 39237 2794 39266 2968
rect 39178 2781 39266 2794
rect 39366 2968 39470 2981
rect 39366 2794 39395 2968
rect 39441 2794 39470 2968
rect 39366 2781 39470 2794
rect 39570 2968 39658 2981
rect 39570 2794 39599 2968
rect 39645 2794 39658 2968
rect 39570 2781 39658 2794
rect 39862 2968 39950 2981
rect 39862 2794 39875 2968
rect 39921 2794 39950 2968
rect 39862 2781 39950 2794
rect 40050 2968 40154 2981
rect 40050 2794 40079 2968
rect 40125 2794 40154 2968
rect 40050 2781 40154 2794
rect 40254 2968 40342 2981
rect 40254 2794 40283 2968
rect 40329 2794 40342 2968
rect 40254 2781 40342 2794
rect 40546 2968 40634 2981
rect 40546 2794 40559 2968
rect 40605 2794 40634 2968
rect 40546 2781 40634 2794
rect 40734 2968 40822 2981
rect 40734 2794 40763 2968
rect 40809 2794 40822 2968
rect 40734 2781 40822 2794
rect 38284 1548 38372 1561
rect 38284 1374 38297 1548
rect 38343 1374 38372 1548
rect 38284 1361 38372 1374
rect 38472 1548 38560 1561
rect 38472 1374 38501 1548
rect 38547 1374 38560 1548
rect 38472 1361 38560 1374
rect 41406 1792 41494 1805
rect 41406 1618 41419 1792
rect 41465 1618 41494 1792
rect 41406 1605 41494 1618
rect 41594 1792 41682 1805
rect 41594 1618 41623 1792
rect 41669 1618 41682 1792
rect 41594 1605 41682 1618
rect 42090 1792 42178 1805
rect 42090 1618 42103 1792
rect 42149 1618 42178 1792
rect 42090 1605 42178 1618
rect 42278 1792 42366 1805
rect 42278 1618 42307 1792
rect 42353 1618 42366 1792
rect 42278 1605 42366 1618
rect 42774 1792 42862 1805
rect 42774 1618 42787 1792
rect 42833 1618 42862 1792
rect 42774 1605 42862 1618
rect 42962 1792 43050 1805
rect 42962 1618 42991 1792
rect 43037 1618 43050 1792
rect 42962 1605 43050 1618
rect 44320 1838 44408 1851
rect 44320 1664 44333 1838
rect 44379 1664 44408 1838
rect 44320 1651 44408 1664
rect 44488 1838 44592 1851
rect 44488 1664 44517 1838
rect 44563 1664 44592 1838
rect 44488 1651 44592 1664
rect 44672 1838 44776 1851
rect 44672 1664 44701 1838
rect 44747 1664 44776 1838
rect 44672 1651 44776 1664
rect 44856 1838 44944 1851
rect 44856 1664 44885 1838
rect 44931 1664 44944 1838
rect 44856 1651 44944 1664
rect 48650 2968 48738 2981
rect 48650 2794 48663 2968
rect 48709 2794 48738 2968
rect 48650 2781 48738 2794
rect 48838 2968 48942 2981
rect 48838 2794 48867 2968
rect 48913 2794 48942 2968
rect 48838 2781 48942 2794
rect 49042 2968 49130 2981
rect 49042 2794 49071 2968
rect 49117 2794 49130 2968
rect 49042 2781 49130 2794
rect 49334 2968 49422 2981
rect 49334 2794 49347 2968
rect 49393 2794 49422 2968
rect 49334 2781 49422 2794
rect 49522 2968 49626 2981
rect 49522 2794 49551 2968
rect 49597 2794 49626 2968
rect 49522 2781 49626 2794
rect 49726 2968 49814 2981
rect 49726 2794 49755 2968
rect 49801 2794 49814 2968
rect 49726 2781 49814 2794
rect 50018 2968 50106 2981
rect 50018 2794 50031 2968
rect 50077 2794 50106 2968
rect 50018 2781 50106 2794
rect 50206 2968 50294 2981
rect 50206 2794 50235 2968
rect 50281 2794 50294 2968
rect 50206 2781 50294 2794
rect 47756 1548 47844 1561
rect 47756 1374 47769 1548
rect 47815 1374 47844 1548
rect 47756 1361 47844 1374
rect 47944 1548 48032 1561
rect 47944 1374 47973 1548
rect 48019 1374 48032 1548
rect 47944 1361 48032 1374
rect 50878 1792 50966 1805
rect 50878 1618 50891 1792
rect 50937 1618 50966 1792
rect 50878 1605 50966 1618
rect 51066 1792 51154 1805
rect 51066 1618 51095 1792
rect 51141 1618 51154 1792
rect 51066 1605 51154 1618
rect 51562 1792 51650 1805
rect 51562 1618 51575 1792
rect 51621 1618 51650 1792
rect 51562 1605 51650 1618
rect 51750 1792 51838 1805
rect 51750 1618 51779 1792
rect 51825 1618 51838 1792
rect 51750 1605 51838 1618
rect 52246 1792 52334 1805
rect 52246 1618 52259 1792
rect 52305 1618 52334 1792
rect 52246 1605 52334 1618
rect 52434 1792 52522 1805
rect 52434 1618 52463 1792
rect 52509 1618 52522 1792
rect 52434 1605 52522 1618
rect 53792 1838 53880 1851
rect 53792 1664 53805 1838
rect 53851 1664 53880 1838
rect 53792 1651 53880 1664
rect 53960 1838 54064 1851
rect 53960 1664 53989 1838
rect 54035 1664 54064 1838
rect 53960 1651 54064 1664
rect 54144 1838 54248 1851
rect 54144 1664 54173 1838
rect 54219 1664 54248 1838
rect 54144 1651 54248 1664
rect 54328 1838 54416 1851
rect 54328 1664 54357 1838
rect 54403 1664 54416 1838
rect 54328 1651 54416 1664
rect 1290 627 1378 640
rect 1290 453 1303 627
rect 1349 453 1378 627
rect 1290 440 1378 453
rect 1478 627 1582 640
rect 1478 453 1507 627
rect 1553 453 1582 627
rect 1478 440 1582 453
rect 1682 627 1770 640
rect 1682 453 1711 627
rect 1757 453 1770 627
rect 1682 440 1770 453
rect 1974 627 2062 640
rect 1974 453 1987 627
rect 2033 453 2062 627
rect 1974 440 2062 453
rect 2162 627 2266 640
rect 2162 453 2191 627
rect 2237 453 2266 627
rect 2162 440 2266 453
rect 2366 627 2454 640
rect 2366 453 2395 627
rect 2441 453 2454 627
rect 2366 440 2454 453
rect 2658 627 2746 640
rect 2658 453 2671 627
rect 2717 453 2746 627
rect 2658 440 2746 453
rect 2846 627 2934 640
rect 2846 453 2875 627
rect 2921 453 2934 627
rect 2846 440 2934 453
rect 10762 627 10850 640
rect 10762 453 10775 627
rect 10821 453 10850 627
rect 10762 440 10850 453
rect 10950 627 11054 640
rect 10950 453 10979 627
rect 11025 453 11054 627
rect 10950 440 11054 453
rect 11154 627 11242 640
rect 11154 453 11183 627
rect 11229 453 11242 627
rect 11154 440 11242 453
rect 11446 627 11534 640
rect 11446 453 11459 627
rect 11505 453 11534 627
rect 11446 440 11534 453
rect 11634 627 11738 640
rect 11634 453 11663 627
rect 11709 453 11738 627
rect 11634 440 11738 453
rect 11838 627 11926 640
rect 11838 453 11867 627
rect 11913 453 11926 627
rect 11838 440 11926 453
rect 12130 627 12218 640
rect 12130 453 12143 627
rect 12189 453 12218 627
rect 12130 440 12218 453
rect 12318 627 12406 640
rect 12318 453 12347 627
rect 12393 453 12406 627
rect 12318 440 12406 453
rect 20234 628 20322 641
rect 20234 454 20247 628
rect 20293 454 20322 628
rect 20234 441 20322 454
rect 20422 628 20526 641
rect 20422 454 20451 628
rect 20497 454 20526 628
rect 20422 441 20526 454
rect 20626 628 20714 641
rect 20626 454 20655 628
rect 20701 454 20714 628
rect 20626 441 20714 454
rect 20918 628 21006 641
rect 20918 454 20931 628
rect 20977 454 21006 628
rect 20918 441 21006 454
rect 21106 628 21210 641
rect 21106 454 21135 628
rect 21181 454 21210 628
rect 21106 441 21210 454
rect 21310 628 21398 641
rect 21310 454 21339 628
rect 21385 454 21398 628
rect 21310 441 21398 454
rect 21602 628 21690 641
rect 21602 454 21615 628
rect 21661 454 21690 628
rect 21602 441 21690 454
rect 21790 628 21878 641
rect 21790 454 21819 628
rect 21865 454 21878 628
rect 21790 441 21878 454
rect 29706 628 29794 641
rect 29706 454 29719 628
rect 29765 454 29794 628
rect 29706 441 29794 454
rect 29894 628 29998 641
rect 29894 454 29923 628
rect 29969 454 29998 628
rect 29894 441 29998 454
rect 30098 628 30186 641
rect 30098 454 30127 628
rect 30173 454 30186 628
rect 30098 441 30186 454
rect 30390 628 30478 641
rect 30390 454 30403 628
rect 30449 454 30478 628
rect 30390 441 30478 454
rect 30578 628 30682 641
rect 30578 454 30607 628
rect 30653 454 30682 628
rect 30578 441 30682 454
rect 30782 628 30870 641
rect 30782 454 30811 628
rect 30857 454 30870 628
rect 30782 441 30870 454
rect 31074 628 31162 641
rect 31074 454 31087 628
rect 31133 454 31162 628
rect 31074 441 31162 454
rect 31262 628 31350 641
rect 31262 454 31291 628
rect 31337 454 31350 628
rect 31262 441 31350 454
rect 39178 628 39266 641
rect 39178 454 39191 628
rect 39237 454 39266 628
rect 39178 441 39266 454
rect 39366 628 39470 641
rect 39366 454 39395 628
rect 39441 454 39470 628
rect 39366 441 39470 454
rect 39570 628 39658 641
rect 39570 454 39599 628
rect 39645 454 39658 628
rect 39570 441 39658 454
rect 39862 628 39950 641
rect 39862 454 39875 628
rect 39921 454 39950 628
rect 39862 441 39950 454
rect 40050 628 40154 641
rect 40050 454 40079 628
rect 40125 454 40154 628
rect 40050 441 40154 454
rect 40254 628 40342 641
rect 40254 454 40283 628
rect 40329 454 40342 628
rect 40254 441 40342 454
rect 40546 628 40634 641
rect 40546 454 40559 628
rect 40605 454 40634 628
rect 40546 441 40634 454
rect 40734 628 40822 641
rect 40734 454 40763 628
rect 40809 454 40822 628
rect 40734 441 40822 454
rect 48650 628 48738 641
rect 48650 454 48663 628
rect 48709 454 48738 628
rect 48650 441 48738 454
rect 48838 628 48942 641
rect 48838 454 48867 628
rect 48913 454 48942 628
rect 48838 441 48942 454
rect 49042 628 49130 641
rect 49042 454 49071 628
rect 49117 454 49130 628
rect 49042 441 49130 454
rect 49334 628 49422 641
rect 49334 454 49347 628
rect 49393 454 49422 628
rect 49334 441 49422 454
rect 49522 628 49626 641
rect 49522 454 49551 628
rect 49597 454 49626 628
rect 49522 441 49626 454
rect 49726 628 49814 641
rect 49726 454 49755 628
rect 49801 454 49814 628
rect 49726 441 49814 454
rect 50018 628 50106 641
rect 50018 454 50031 628
rect 50077 454 50106 628
rect 50018 441 50106 454
rect 50206 628 50294 641
rect 50206 454 50235 628
rect 50281 454 50294 628
rect 50206 441 50294 454
<< pdiff >>
rect 6432 9612 6520 9625
rect 6432 9138 6445 9612
rect 6491 9138 6520 9612
rect 6432 9125 6520 9138
rect 6600 9612 6704 9625
rect 6600 9138 6629 9612
rect 6675 9138 6704 9612
rect 6600 9125 6704 9138
rect 6784 9612 6888 9625
rect 6784 9138 6813 9612
rect 6859 9138 6888 9612
rect 6784 9125 6888 9138
rect 6968 9612 7056 9625
rect 6968 9138 6997 9612
rect 7043 9138 7056 9612
rect 6968 9125 7056 9138
rect 15904 9612 15992 9625
rect 15904 9138 15917 9612
rect 15963 9138 15992 9612
rect 15904 9125 15992 9138
rect 16072 9612 16176 9625
rect 16072 9138 16101 9612
rect 16147 9138 16176 9612
rect 16072 9125 16176 9138
rect 16256 9612 16360 9625
rect 16256 9138 16285 9612
rect 16331 9138 16360 9612
rect 16256 9125 16360 9138
rect 16440 9612 16528 9625
rect 16440 9138 16469 9612
rect 16515 9138 16528 9612
rect 16440 9125 16528 9138
rect 25376 9613 25464 9626
rect 25376 9139 25389 9613
rect 25435 9139 25464 9613
rect 25376 9126 25464 9139
rect 25544 9613 25648 9626
rect 25544 9139 25573 9613
rect 25619 9139 25648 9613
rect 25544 9126 25648 9139
rect 25728 9613 25832 9626
rect 25728 9139 25757 9613
rect 25803 9139 25832 9613
rect 25728 9126 25832 9139
rect 25912 9613 26000 9626
rect 25912 9139 25941 9613
rect 25987 9139 26000 9613
rect 25912 9126 26000 9139
rect 34848 9613 34936 9626
rect 34848 9139 34861 9613
rect 34907 9139 34936 9613
rect 34848 9126 34936 9139
rect 35016 9613 35120 9626
rect 35016 9139 35045 9613
rect 35091 9139 35120 9613
rect 35016 9126 35120 9139
rect 35200 9613 35304 9626
rect 35200 9139 35229 9613
rect 35275 9139 35304 9613
rect 35200 9126 35304 9139
rect 35384 9613 35472 9626
rect 35384 9139 35413 9613
rect 35459 9139 35472 9613
rect 35384 9126 35472 9139
rect 44320 9613 44408 9626
rect 44320 9139 44333 9613
rect 44379 9139 44408 9613
rect 44320 9126 44408 9139
rect 44488 9613 44592 9626
rect 44488 9139 44517 9613
rect 44563 9139 44592 9613
rect 44488 9126 44592 9139
rect 44672 9613 44776 9626
rect 44672 9139 44701 9613
rect 44747 9139 44776 9613
rect 44672 9126 44776 9139
rect 44856 9613 44944 9626
rect 44856 9139 44885 9613
rect 44931 9139 44944 9613
rect 44856 9126 44944 9139
rect 53792 9613 53880 9626
rect 53792 9139 53805 9613
rect 53851 9139 53880 9613
rect 53792 9126 53880 9139
rect 53960 9613 54064 9626
rect 53960 9139 53989 9613
rect 54035 9139 54064 9613
rect 53960 9126 54064 9139
rect 54144 9613 54248 9626
rect 54144 9139 54173 9613
rect 54219 9139 54248 9613
rect 54144 9126 54248 9139
rect 54328 9613 54416 9626
rect 54328 9139 54357 9613
rect 54403 9139 54416 9613
rect 54328 9126 54416 9139
rect 6432 7407 6520 7420
rect 6432 6933 6445 7407
rect 6491 6933 6520 7407
rect 6432 6920 6520 6933
rect 6600 7407 6704 7420
rect 6600 6933 6629 7407
rect 6675 6933 6704 7407
rect 6600 6920 6704 6933
rect 6784 7407 6888 7420
rect 6784 6933 6813 7407
rect 6859 6933 6888 7407
rect 6784 6920 6888 6933
rect 6968 7407 7056 7420
rect 6968 6933 6997 7407
rect 7043 6933 7056 7407
rect 6968 6920 7056 6933
rect 7918 7407 8006 7420
rect 7918 6933 7931 7407
rect 7977 6933 8006 7407
rect 7918 6920 8006 6933
rect 8086 7407 8190 7420
rect 8086 6933 8115 7407
rect 8161 6933 8190 7407
rect 8086 6920 8190 6933
rect 8270 7407 8374 7420
rect 8270 6933 8299 7407
rect 8345 6933 8374 7407
rect 8270 6920 8374 6933
rect 8454 7407 8542 7420
rect 8454 6933 8483 7407
rect 8529 6933 8542 7407
rect 8454 6920 8542 6933
rect 15904 7407 15992 7420
rect 15904 6933 15917 7407
rect 15963 6933 15992 7407
rect 15904 6920 15992 6933
rect 16072 7407 16176 7420
rect 16072 6933 16101 7407
rect 16147 6933 16176 7407
rect 16072 6920 16176 6933
rect 16256 7407 16360 7420
rect 16256 6933 16285 7407
rect 16331 6933 16360 7407
rect 16256 6920 16360 6933
rect 16440 7407 16528 7420
rect 16440 6933 16469 7407
rect 16515 6933 16528 7407
rect 16440 6920 16528 6933
rect 17390 7407 17478 7420
rect 17390 6933 17403 7407
rect 17449 6933 17478 7407
rect 17390 6920 17478 6933
rect 17558 7407 17662 7420
rect 17558 6933 17587 7407
rect 17633 6933 17662 7407
rect 17558 6920 17662 6933
rect 17742 7407 17846 7420
rect 17742 6933 17771 7407
rect 17817 6933 17846 7407
rect 17742 6920 17846 6933
rect 17926 7407 18014 7420
rect 17926 6933 17955 7407
rect 18001 6933 18014 7407
rect 17926 6920 18014 6933
rect 25376 7408 25464 7421
rect 25376 6934 25389 7408
rect 25435 6934 25464 7408
rect 25376 6921 25464 6934
rect 25544 7408 25648 7421
rect 25544 6934 25573 7408
rect 25619 6934 25648 7408
rect 25544 6921 25648 6934
rect 25728 7408 25832 7421
rect 25728 6934 25757 7408
rect 25803 6934 25832 7408
rect 25728 6921 25832 6934
rect 25912 7408 26000 7421
rect 25912 6934 25941 7408
rect 25987 6934 26000 7408
rect 25912 6921 26000 6934
rect 26862 7408 26950 7421
rect 26862 6934 26875 7408
rect 26921 6934 26950 7408
rect 26862 6921 26950 6934
rect 27030 7408 27134 7421
rect 27030 6934 27059 7408
rect 27105 6934 27134 7408
rect 27030 6921 27134 6934
rect 27214 7408 27318 7421
rect 27214 6934 27243 7408
rect 27289 6934 27318 7408
rect 27214 6921 27318 6934
rect 27398 7408 27486 7421
rect 27398 6934 27427 7408
rect 27473 6934 27486 7408
rect 27398 6921 27486 6934
rect 34848 7408 34936 7421
rect 34848 6934 34861 7408
rect 34907 6934 34936 7408
rect 34848 6921 34936 6934
rect 35016 7408 35120 7421
rect 35016 6934 35045 7408
rect 35091 6934 35120 7408
rect 35016 6921 35120 6934
rect 35200 7408 35304 7421
rect 35200 6934 35229 7408
rect 35275 6934 35304 7408
rect 35200 6921 35304 6934
rect 35384 7408 35472 7421
rect 35384 6934 35413 7408
rect 35459 6934 35472 7408
rect 35384 6921 35472 6934
rect 36334 7408 36422 7421
rect 36334 6934 36347 7408
rect 36393 6934 36422 7408
rect 36334 6921 36422 6934
rect 36502 7408 36606 7421
rect 36502 6934 36531 7408
rect 36577 6934 36606 7408
rect 36502 6921 36606 6934
rect 36686 7408 36790 7421
rect 36686 6934 36715 7408
rect 36761 6934 36790 7408
rect 36686 6921 36790 6934
rect 36870 7408 36958 7421
rect 36870 6934 36899 7408
rect 36945 6934 36958 7408
rect 36870 6921 36958 6934
rect 44320 7408 44408 7421
rect 44320 6934 44333 7408
rect 44379 6934 44408 7408
rect 44320 6921 44408 6934
rect 44488 7408 44592 7421
rect 44488 6934 44517 7408
rect 44563 6934 44592 7408
rect 44488 6921 44592 6934
rect 44672 7408 44776 7421
rect 44672 6934 44701 7408
rect 44747 6934 44776 7408
rect 44672 6921 44776 6934
rect 44856 7408 44944 7421
rect 44856 6934 44885 7408
rect 44931 6934 44944 7408
rect 44856 6921 44944 6934
rect 45806 7408 45894 7421
rect 45806 6934 45819 7408
rect 45865 6934 45894 7408
rect 45806 6921 45894 6934
rect 45974 7408 46078 7421
rect 45974 6934 46003 7408
rect 46049 6934 46078 7408
rect 45974 6921 46078 6934
rect 46158 7408 46262 7421
rect 46158 6934 46187 7408
rect 46233 6934 46262 7408
rect 46158 6921 46262 6934
rect 46342 7408 46430 7421
rect 46342 6934 46371 7408
rect 46417 6934 46430 7408
rect 46342 6921 46430 6934
rect 53792 7408 53880 7421
rect 53792 6934 53805 7408
rect 53851 6934 53880 7408
rect 53792 6921 53880 6934
rect 53960 7408 54064 7421
rect 53960 6934 53989 7408
rect 54035 6934 54064 7408
rect 53960 6921 54064 6934
rect 54144 7408 54248 7421
rect 54144 6934 54173 7408
rect 54219 6934 54248 7408
rect 54144 6921 54248 6934
rect 54328 7408 54416 7421
rect 54328 6934 54357 7408
rect 54403 6934 54416 7408
rect 54328 6921 54416 6934
rect 55278 7408 55366 7421
rect 55278 6934 55291 7408
rect 55337 6934 55366 7408
rect 55278 6921 55366 6934
rect 55446 7408 55550 7421
rect 55446 6934 55475 7408
rect 55521 6934 55550 7408
rect 55446 6921 55550 6934
rect 55630 7408 55734 7421
rect 55630 6934 55659 7408
rect 55705 6934 55734 7408
rect 55630 6921 55734 6934
rect 55814 7408 55902 7421
rect 55814 6934 55843 7408
rect 55889 6934 55902 7408
rect 55814 6921 55902 6934
rect 6432 5202 6520 5215
rect 6432 4728 6445 5202
rect 6491 4728 6520 5202
rect 6432 4715 6520 4728
rect 6600 5202 6704 5215
rect 6600 4728 6629 5202
rect 6675 4728 6704 5202
rect 6600 4715 6704 4728
rect 6784 5202 6888 5215
rect 6784 4728 6813 5202
rect 6859 4728 6888 5202
rect 6784 4715 6888 4728
rect 6968 5202 7056 5215
rect 6968 4728 6997 5202
rect 7043 4728 7056 5202
rect 6968 4715 7056 4728
rect 7918 5203 8006 5216
rect 7918 4729 7931 5203
rect 7977 4729 8006 5203
rect 7918 4716 8006 4729
rect 8086 5203 8190 5216
rect 8086 4729 8115 5203
rect 8161 4729 8190 5203
rect 8086 4716 8190 4729
rect 8270 5203 8374 5216
rect 8270 4729 8299 5203
rect 8345 4729 8374 5203
rect 8270 4716 8374 4729
rect 8454 5203 8542 5216
rect 8454 4729 8483 5203
rect 8529 4729 8542 5203
rect 8454 4716 8542 4729
rect 15904 5202 15992 5215
rect 15904 4728 15917 5202
rect 15963 4728 15992 5202
rect 15904 4715 15992 4728
rect 16072 5202 16176 5215
rect 16072 4728 16101 5202
rect 16147 4728 16176 5202
rect 16072 4715 16176 4728
rect 16256 5202 16360 5215
rect 16256 4728 16285 5202
rect 16331 4728 16360 5202
rect 16256 4715 16360 4728
rect 16440 5202 16528 5215
rect 16440 4728 16469 5202
rect 16515 4728 16528 5202
rect 16440 4715 16528 4728
rect 17390 5203 17478 5216
rect 17390 4729 17403 5203
rect 17449 4729 17478 5203
rect 17390 4716 17478 4729
rect 17558 5203 17662 5216
rect 17558 4729 17587 5203
rect 17633 4729 17662 5203
rect 17558 4716 17662 4729
rect 17742 5203 17846 5216
rect 17742 4729 17771 5203
rect 17817 4729 17846 5203
rect 17742 4716 17846 4729
rect 17926 5203 18014 5216
rect 17926 4729 17955 5203
rect 18001 4729 18014 5203
rect 17926 4716 18014 4729
rect 25376 5203 25464 5216
rect 25376 4729 25389 5203
rect 25435 4729 25464 5203
rect 25376 4716 25464 4729
rect 25544 5203 25648 5216
rect 25544 4729 25573 5203
rect 25619 4729 25648 5203
rect 25544 4716 25648 4729
rect 25728 5203 25832 5216
rect 25728 4729 25757 5203
rect 25803 4729 25832 5203
rect 25728 4716 25832 4729
rect 25912 5203 26000 5216
rect 25912 4729 25941 5203
rect 25987 4729 26000 5203
rect 25912 4716 26000 4729
rect 26862 5204 26950 5217
rect 26862 4730 26875 5204
rect 26921 4730 26950 5204
rect 26862 4717 26950 4730
rect 27030 5204 27134 5217
rect 27030 4730 27059 5204
rect 27105 4730 27134 5204
rect 27030 4717 27134 4730
rect 27214 5204 27318 5217
rect 27214 4730 27243 5204
rect 27289 4730 27318 5204
rect 27214 4717 27318 4730
rect 27398 5204 27486 5217
rect 27398 4730 27427 5204
rect 27473 4730 27486 5204
rect 27398 4717 27486 4730
rect 34848 5203 34936 5216
rect 34848 4729 34861 5203
rect 34907 4729 34936 5203
rect 34848 4716 34936 4729
rect 35016 5203 35120 5216
rect 35016 4729 35045 5203
rect 35091 4729 35120 5203
rect 35016 4716 35120 4729
rect 35200 5203 35304 5216
rect 35200 4729 35229 5203
rect 35275 4729 35304 5203
rect 35200 4716 35304 4729
rect 35384 5203 35472 5216
rect 35384 4729 35413 5203
rect 35459 4729 35472 5203
rect 35384 4716 35472 4729
rect 36334 5204 36422 5217
rect 36334 4730 36347 5204
rect 36393 4730 36422 5204
rect 36334 4717 36422 4730
rect 36502 5204 36606 5217
rect 36502 4730 36531 5204
rect 36577 4730 36606 5204
rect 36502 4717 36606 4730
rect 36686 5204 36790 5217
rect 36686 4730 36715 5204
rect 36761 4730 36790 5204
rect 36686 4717 36790 4730
rect 36870 5204 36958 5217
rect 36870 4730 36899 5204
rect 36945 4730 36958 5204
rect 36870 4717 36958 4730
rect 44320 5203 44408 5216
rect 44320 4729 44333 5203
rect 44379 4729 44408 5203
rect 44320 4716 44408 4729
rect 44488 5203 44592 5216
rect 44488 4729 44517 5203
rect 44563 4729 44592 5203
rect 44488 4716 44592 4729
rect 44672 5203 44776 5216
rect 44672 4729 44701 5203
rect 44747 4729 44776 5203
rect 44672 4716 44776 4729
rect 44856 5203 44944 5216
rect 44856 4729 44885 5203
rect 44931 4729 44944 5203
rect 44856 4716 44944 4729
rect 45806 5204 45894 5217
rect 45806 4730 45819 5204
rect 45865 4730 45894 5204
rect 45806 4717 45894 4730
rect 45974 5204 46078 5217
rect 45974 4730 46003 5204
rect 46049 4730 46078 5204
rect 45974 4717 46078 4730
rect 46158 5204 46262 5217
rect 46158 4730 46187 5204
rect 46233 4730 46262 5204
rect 46158 4717 46262 4730
rect 46342 5204 46430 5217
rect 46342 4730 46371 5204
rect 46417 4730 46430 5204
rect 46342 4717 46430 4730
rect 53792 5203 53880 5216
rect 53792 4729 53805 5203
rect 53851 4729 53880 5203
rect 53792 4716 53880 4729
rect 53960 5203 54064 5216
rect 53960 4729 53989 5203
rect 54035 4729 54064 5203
rect 53960 4716 54064 4729
rect 54144 5203 54248 5216
rect 54144 4729 54173 5203
rect 54219 4729 54248 5203
rect 54144 4716 54248 4729
rect 54328 5203 54416 5216
rect 54328 4729 54357 5203
rect 54403 4729 54416 5203
rect 54328 4716 54416 4729
rect 55278 5204 55366 5217
rect 55278 4730 55291 5204
rect 55337 4730 55366 5204
rect 55278 4717 55366 4730
rect 55446 5204 55550 5217
rect 55446 4730 55475 5204
rect 55521 4730 55550 5204
rect 55446 4717 55550 4730
rect 55630 5204 55734 5217
rect 55630 4730 55659 5204
rect 55705 4730 55734 5204
rect 55630 4717 55734 4730
rect 55814 5204 55902 5217
rect 55814 4730 55843 5204
rect 55889 4730 55902 5204
rect 55814 4717 55902 4730
rect 1290 4087 1378 4100
rect 1290 3513 1303 4087
rect 1349 3513 1378 4087
rect 1290 3500 1378 3513
rect 1478 4087 1566 4100
rect 1478 3513 1507 4087
rect 1553 3513 1566 4087
rect 1478 3500 1566 3513
rect 2178 4087 2266 4100
rect 2178 3513 2191 4087
rect 2237 3513 2266 4087
rect 2178 3500 2266 3513
rect 2366 4087 2454 4100
rect 2366 3513 2395 4087
rect 2441 3513 2454 4087
rect 2366 3500 2454 3513
rect 2658 4087 2746 4100
rect 2658 3513 2671 4087
rect 2717 3513 2746 4087
rect 2658 3500 2746 3513
rect 2846 4087 2934 4100
rect 2846 3513 2875 4087
rect 2921 3513 2934 4087
rect 2846 3500 2934 3513
rect 10762 4087 10850 4100
rect 10762 3513 10775 4087
rect 10821 3513 10850 4087
rect 10762 3500 10850 3513
rect 10950 4087 11038 4100
rect 10950 3513 10979 4087
rect 11025 3513 11038 4087
rect 10950 3500 11038 3513
rect 11650 4087 11738 4100
rect 11650 3513 11663 4087
rect 11709 3513 11738 4087
rect 11650 3500 11738 3513
rect 11838 4087 11926 4100
rect 11838 3513 11867 4087
rect 11913 3513 11926 4087
rect 11838 3500 11926 3513
rect 12130 4087 12218 4100
rect 12130 3513 12143 4087
rect 12189 3513 12218 4087
rect 12130 3500 12218 3513
rect 12318 4087 12406 4100
rect 12318 3513 12347 4087
rect 12393 3513 12406 4087
rect 12318 3500 12406 3513
rect 20234 4088 20322 4101
rect 20234 3514 20247 4088
rect 20293 3514 20322 4088
rect 20234 3501 20322 3514
rect 20422 4088 20510 4101
rect 20422 3514 20451 4088
rect 20497 3514 20510 4088
rect 20422 3501 20510 3514
rect 21122 4088 21210 4101
rect 21122 3514 21135 4088
rect 21181 3514 21210 4088
rect 21122 3501 21210 3514
rect 21310 4088 21398 4101
rect 21310 3514 21339 4088
rect 21385 3514 21398 4088
rect 21310 3501 21398 3514
rect 21602 4088 21690 4101
rect 21602 3514 21615 4088
rect 21661 3514 21690 4088
rect 21602 3501 21690 3514
rect 21790 4088 21878 4101
rect 21790 3514 21819 4088
rect 21865 3514 21878 4088
rect 21790 3501 21878 3514
rect 29706 4088 29794 4101
rect 29706 3514 29719 4088
rect 29765 3514 29794 4088
rect 29706 3501 29794 3514
rect 29894 4088 29982 4101
rect 29894 3514 29923 4088
rect 29969 3514 29982 4088
rect 29894 3501 29982 3514
rect 30594 4088 30682 4101
rect 30594 3514 30607 4088
rect 30653 3514 30682 4088
rect 30594 3501 30682 3514
rect 30782 4088 30870 4101
rect 30782 3514 30811 4088
rect 30857 3514 30870 4088
rect 30782 3501 30870 3514
rect 31074 4088 31162 4101
rect 31074 3514 31087 4088
rect 31133 3514 31162 4088
rect 31074 3501 31162 3514
rect 31262 4088 31350 4101
rect 31262 3514 31291 4088
rect 31337 3514 31350 4088
rect 31262 3501 31350 3514
rect 39178 4088 39266 4101
rect 39178 3514 39191 4088
rect 39237 3514 39266 4088
rect 39178 3501 39266 3514
rect 39366 4088 39454 4101
rect 39366 3514 39395 4088
rect 39441 3514 39454 4088
rect 39366 3501 39454 3514
rect 40066 4088 40154 4101
rect 40066 3514 40079 4088
rect 40125 3514 40154 4088
rect 40066 3501 40154 3514
rect 40254 4088 40342 4101
rect 40254 3514 40283 4088
rect 40329 3514 40342 4088
rect 40254 3501 40342 3514
rect 40546 4088 40634 4101
rect 40546 3514 40559 4088
rect 40605 3514 40634 4088
rect 40546 3501 40634 3514
rect 40734 4088 40822 4101
rect 40734 3514 40763 4088
rect 40809 3514 40822 4088
rect 40734 3501 40822 3514
rect 48650 4088 48738 4101
rect 48650 3514 48663 4088
rect 48709 3514 48738 4088
rect 48650 3501 48738 3514
rect 48838 4088 48926 4101
rect 48838 3514 48867 4088
rect 48913 3514 48926 4088
rect 48838 3501 48926 3514
rect 49538 4088 49626 4101
rect 49538 3514 49551 4088
rect 49597 3514 49626 4088
rect 49538 3501 49626 3514
rect 49726 4088 49814 4101
rect 49726 3514 49755 4088
rect 49801 3514 49814 4088
rect 49726 3501 49814 3514
rect 50018 4088 50106 4101
rect 50018 3514 50031 4088
rect 50077 3514 50106 4088
rect 50018 3501 50106 3514
rect 50206 4088 50294 4101
rect 50206 3514 50235 4088
rect 50281 3514 50294 4088
rect 50206 3501 50294 3514
rect 396 2667 484 2680
rect 396 2093 409 2667
rect 455 2093 484 2667
rect 396 2080 484 2093
rect 584 2667 672 2680
rect 584 2093 613 2667
rect 659 2093 672 2667
rect 584 2080 672 2093
rect 3518 2911 3606 2924
rect 3518 2337 3531 2911
rect 3577 2337 3606 2911
rect 3518 2324 3606 2337
rect 3706 2911 3810 2924
rect 3706 2337 3735 2911
rect 3781 2337 3810 2911
rect 3706 2324 3810 2337
rect 3910 2911 3998 2924
rect 3910 2337 3939 2911
rect 3985 2337 3998 2911
rect 3910 2324 3998 2337
rect 4202 2911 4290 2924
rect 4202 2337 4215 2911
rect 4261 2337 4290 2911
rect 4202 2324 4290 2337
rect 4390 2911 4494 2924
rect 4390 2337 4419 2911
rect 4465 2337 4494 2911
rect 4390 2324 4494 2337
rect 4594 2911 4682 2924
rect 4594 2337 4623 2911
rect 4669 2337 4682 2911
rect 4594 2324 4682 2337
rect 4886 2911 4974 2924
rect 4886 2337 4899 2911
rect 4945 2337 4974 2911
rect 4886 2324 4974 2337
rect 5074 2911 5162 2924
rect 5074 2337 5103 2911
rect 5149 2337 5162 2911
rect 5074 2324 5162 2337
rect 6432 2997 6520 3010
rect 6432 2523 6445 2997
rect 6491 2523 6520 2997
rect 6432 2510 6520 2523
rect 6600 2997 6704 3010
rect 6600 2523 6629 2997
rect 6675 2523 6704 2997
rect 6600 2510 6704 2523
rect 6784 2997 6888 3010
rect 6784 2523 6813 2997
rect 6859 2523 6888 2997
rect 6784 2510 6888 2523
rect 6968 2997 7056 3010
rect 6968 2523 6997 2997
rect 7043 2523 7056 2997
rect 6968 2510 7056 2523
rect 1290 1747 1378 1760
rect 1290 1173 1303 1747
rect 1349 1173 1378 1747
rect 1290 1160 1378 1173
rect 1478 1747 1566 1760
rect 1478 1173 1507 1747
rect 1553 1173 1566 1747
rect 1478 1160 1566 1173
rect 2178 1747 2266 1760
rect 2178 1173 2191 1747
rect 2237 1173 2266 1747
rect 2178 1160 2266 1173
rect 2366 1747 2454 1760
rect 2366 1173 2395 1747
rect 2441 1173 2454 1747
rect 2366 1160 2454 1173
rect 2658 1747 2746 1760
rect 2658 1173 2671 1747
rect 2717 1173 2746 1747
rect 2658 1160 2746 1173
rect 2846 1747 2934 1760
rect 2846 1173 2875 1747
rect 2921 1173 2934 1747
rect 2846 1160 2934 1173
rect 9868 2667 9956 2680
rect 9868 2093 9881 2667
rect 9927 2093 9956 2667
rect 9868 2080 9956 2093
rect 10056 2667 10144 2680
rect 10056 2093 10085 2667
rect 10131 2093 10144 2667
rect 10056 2080 10144 2093
rect 12990 2911 13078 2924
rect 12990 2337 13003 2911
rect 13049 2337 13078 2911
rect 12990 2324 13078 2337
rect 13178 2911 13282 2924
rect 13178 2337 13207 2911
rect 13253 2337 13282 2911
rect 13178 2324 13282 2337
rect 13382 2911 13470 2924
rect 13382 2337 13411 2911
rect 13457 2337 13470 2911
rect 13382 2324 13470 2337
rect 13674 2911 13762 2924
rect 13674 2337 13687 2911
rect 13733 2337 13762 2911
rect 13674 2324 13762 2337
rect 13862 2911 13966 2924
rect 13862 2337 13891 2911
rect 13937 2337 13966 2911
rect 13862 2324 13966 2337
rect 14066 2911 14154 2924
rect 14066 2337 14095 2911
rect 14141 2337 14154 2911
rect 14066 2324 14154 2337
rect 14358 2911 14446 2924
rect 14358 2337 14371 2911
rect 14417 2337 14446 2911
rect 14358 2324 14446 2337
rect 14546 2911 14634 2924
rect 14546 2337 14575 2911
rect 14621 2337 14634 2911
rect 14546 2324 14634 2337
rect 15904 2997 15992 3010
rect 15904 2523 15917 2997
rect 15963 2523 15992 2997
rect 15904 2510 15992 2523
rect 16072 2997 16176 3010
rect 16072 2523 16101 2997
rect 16147 2523 16176 2997
rect 16072 2510 16176 2523
rect 16256 2997 16360 3010
rect 16256 2523 16285 2997
rect 16331 2523 16360 2997
rect 16256 2510 16360 2523
rect 16440 2997 16528 3010
rect 16440 2523 16469 2997
rect 16515 2523 16528 2997
rect 16440 2510 16528 2523
rect 10762 1747 10850 1760
rect 10762 1173 10775 1747
rect 10821 1173 10850 1747
rect 10762 1160 10850 1173
rect 10950 1747 11038 1760
rect 10950 1173 10979 1747
rect 11025 1173 11038 1747
rect 10950 1160 11038 1173
rect 11650 1747 11738 1760
rect 11650 1173 11663 1747
rect 11709 1173 11738 1747
rect 11650 1160 11738 1173
rect 11838 1747 11926 1760
rect 11838 1173 11867 1747
rect 11913 1173 11926 1747
rect 11838 1160 11926 1173
rect 12130 1747 12218 1760
rect 12130 1173 12143 1747
rect 12189 1173 12218 1747
rect 12130 1160 12218 1173
rect 12318 1747 12406 1760
rect 12318 1173 12347 1747
rect 12393 1173 12406 1747
rect 12318 1160 12406 1173
rect 19340 2668 19428 2681
rect 19340 2094 19353 2668
rect 19399 2094 19428 2668
rect 19340 2081 19428 2094
rect 19528 2668 19616 2681
rect 19528 2094 19557 2668
rect 19603 2094 19616 2668
rect 19528 2081 19616 2094
rect 22462 2912 22550 2925
rect 22462 2338 22475 2912
rect 22521 2338 22550 2912
rect 22462 2325 22550 2338
rect 22650 2912 22754 2925
rect 22650 2338 22679 2912
rect 22725 2338 22754 2912
rect 22650 2325 22754 2338
rect 22854 2912 22942 2925
rect 22854 2338 22883 2912
rect 22929 2338 22942 2912
rect 22854 2325 22942 2338
rect 23146 2912 23234 2925
rect 23146 2338 23159 2912
rect 23205 2338 23234 2912
rect 23146 2325 23234 2338
rect 23334 2912 23438 2925
rect 23334 2338 23363 2912
rect 23409 2338 23438 2912
rect 23334 2325 23438 2338
rect 23538 2912 23626 2925
rect 23538 2338 23567 2912
rect 23613 2338 23626 2912
rect 23538 2325 23626 2338
rect 23830 2912 23918 2925
rect 23830 2338 23843 2912
rect 23889 2338 23918 2912
rect 23830 2325 23918 2338
rect 24018 2912 24106 2925
rect 24018 2338 24047 2912
rect 24093 2338 24106 2912
rect 24018 2325 24106 2338
rect 25376 2998 25464 3011
rect 25376 2524 25389 2998
rect 25435 2524 25464 2998
rect 25376 2511 25464 2524
rect 25544 2998 25648 3011
rect 25544 2524 25573 2998
rect 25619 2524 25648 2998
rect 25544 2511 25648 2524
rect 25728 2998 25832 3011
rect 25728 2524 25757 2998
rect 25803 2524 25832 2998
rect 25728 2511 25832 2524
rect 25912 2998 26000 3011
rect 25912 2524 25941 2998
rect 25987 2524 26000 2998
rect 25912 2511 26000 2524
rect 20234 1748 20322 1761
rect 20234 1174 20247 1748
rect 20293 1174 20322 1748
rect 20234 1161 20322 1174
rect 20422 1748 20510 1761
rect 20422 1174 20451 1748
rect 20497 1174 20510 1748
rect 20422 1161 20510 1174
rect 21122 1748 21210 1761
rect 21122 1174 21135 1748
rect 21181 1174 21210 1748
rect 21122 1161 21210 1174
rect 21310 1748 21398 1761
rect 21310 1174 21339 1748
rect 21385 1174 21398 1748
rect 21310 1161 21398 1174
rect 21602 1748 21690 1761
rect 21602 1174 21615 1748
rect 21661 1174 21690 1748
rect 21602 1161 21690 1174
rect 21790 1748 21878 1761
rect 21790 1174 21819 1748
rect 21865 1174 21878 1748
rect 21790 1161 21878 1174
rect 28812 2668 28900 2681
rect 28812 2094 28825 2668
rect 28871 2094 28900 2668
rect 28812 2081 28900 2094
rect 29000 2668 29088 2681
rect 29000 2094 29029 2668
rect 29075 2094 29088 2668
rect 29000 2081 29088 2094
rect 31934 2912 32022 2925
rect 31934 2338 31947 2912
rect 31993 2338 32022 2912
rect 31934 2325 32022 2338
rect 32122 2912 32226 2925
rect 32122 2338 32151 2912
rect 32197 2338 32226 2912
rect 32122 2325 32226 2338
rect 32326 2912 32414 2925
rect 32326 2338 32355 2912
rect 32401 2338 32414 2912
rect 32326 2325 32414 2338
rect 32618 2912 32706 2925
rect 32618 2338 32631 2912
rect 32677 2338 32706 2912
rect 32618 2325 32706 2338
rect 32806 2912 32910 2925
rect 32806 2338 32835 2912
rect 32881 2338 32910 2912
rect 32806 2325 32910 2338
rect 33010 2912 33098 2925
rect 33010 2338 33039 2912
rect 33085 2338 33098 2912
rect 33010 2325 33098 2338
rect 33302 2912 33390 2925
rect 33302 2338 33315 2912
rect 33361 2338 33390 2912
rect 33302 2325 33390 2338
rect 33490 2912 33578 2925
rect 33490 2338 33519 2912
rect 33565 2338 33578 2912
rect 33490 2325 33578 2338
rect 34848 2998 34936 3011
rect 34848 2524 34861 2998
rect 34907 2524 34936 2998
rect 34848 2511 34936 2524
rect 35016 2998 35120 3011
rect 35016 2524 35045 2998
rect 35091 2524 35120 2998
rect 35016 2511 35120 2524
rect 35200 2998 35304 3011
rect 35200 2524 35229 2998
rect 35275 2524 35304 2998
rect 35200 2511 35304 2524
rect 35384 2998 35472 3011
rect 35384 2524 35413 2998
rect 35459 2524 35472 2998
rect 35384 2511 35472 2524
rect 29706 1748 29794 1761
rect 29706 1174 29719 1748
rect 29765 1174 29794 1748
rect 29706 1161 29794 1174
rect 29894 1748 29982 1761
rect 29894 1174 29923 1748
rect 29969 1174 29982 1748
rect 29894 1161 29982 1174
rect 30594 1748 30682 1761
rect 30594 1174 30607 1748
rect 30653 1174 30682 1748
rect 30594 1161 30682 1174
rect 30782 1748 30870 1761
rect 30782 1174 30811 1748
rect 30857 1174 30870 1748
rect 30782 1161 30870 1174
rect 31074 1748 31162 1761
rect 31074 1174 31087 1748
rect 31133 1174 31162 1748
rect 31074 1161 31162 1174
rect 31262 1748 31350 1761
rect 31262 1174 31291 1748
rect 31337 1174 31350 1748
rect 31262 1161 31350 1174
rect 38284 2668 38372 2681
rect 38284 2094 38297 2668
rect 38343 2094 38372 2668
rect 38284 2081 38372 2094
rect 38472 2668 38560 2681
rect 38472 2094 38501 2668
rect 38547 2094 38560 2668
rect 38472 2081 38560 2094
rect 41406 2912 41494 2925
rect 41406 2338 41419 2912
rect 41465 2338 41494 2912
rect 41406 2325 41494 2338
rect 41594 2912 41698 2925
rect 41594 2338 41623 2912
rect 41669 2338 41698 2912
rect 41594 2325 41698 2338
rect 41798 2912 41886 2925
rect 41798 2338 41827 2912
rect 41873 2338 41886 2912
rect 41798 2325 41886 2338
rect 42090 2912 42178 2925
rect 42090 2338 42103 2912
rect 42149 2338 42178 2912
rect 42090 2325 42178 2338
rect 42278 2912 42382 2925
rect 42278 2338 42307 2912
rect 42353 2338 42382 2912
rect 42278 2325 42382 2338
rect 42482 2912 42570 2925
rect 42482 2338 42511 2912
rect 42557 2338 42570 2912
rect 42482 2325 42570 2338
rect 42774 2912 42862 2925
rect 42774 2338 42787 2912
rect 42833 2338 42862 2912
rect 42774 2325 42862 2338
rect 42962 2912 43050 2925
rect 42962 2338 42991 2912
rect 43037 2338 43050 2912
rect 42962 2325 43050 2338
rect 44320 2998 44408 3011
rect 44320 2524 44333 2998
rect 44379 2524 44408 2998
rect 44320 2511 44408 2524
rect 44488 2998 44592 3011
rect 44488 2524 44517 2998
rect 44563 2524 44592 2998
rect 44488 2511 44592 2524
rect 44672 2998 44776 3011
rect 44672 2524 44701 2998
rect 44747 2524 44776 2998
rect 44672 2511 44776 2524
rect 44856 2998 44944 3011
rect 44856 2524 44885 2998
rect 44931 2524 44944 2998
rect 44856 2511 44944 2524
rect 39178 1748 39266 1761
rect 39178 1174 39191 1748
rect 39237 1174 39266 1748
rect 39178 1161 39266 1174
rect 39366 1748 39454 1761
rect 39366 1174 39395 1748
rect 39441 1174 39454 1748
rect 39366 1161 39454 1174
rect 40066 1748 40154 1761
rect 40066 1174 40079 1748
rect 40125 1174 40154 1748
rect 40066 1161 40154 1174
rect 40254 1748 40342 1761
rect 40254 1174 40283 1748
rect 40329 1174 40342 1748
rect 40254 1161 40342 1174
rect 40546 1748 40634 1761
rect 40546 1174 40559 1748
rect 40605 1174 40634 1748
rect 40546 1161 40634 1174
rect 40734 1748 40822 1761
rect 40734 1174 40763 1748
rect 40809 1174 40822 1748
rect 40734 1161 40822 1174
rect 47756 2668 47844 2681
rect 47756 2094 47769 2668
rect 47815 2094 47844 2668
rect 47756 2081 47844 2094
rect 47944 2668 48032 2681
rect 47944 2094 47973 2668
rect 48019 2094 48032 2668
rect 47944 2081 48032 2094
rect 50878 2912 50966 2925
rect 50878 2338 50891 2912
rect 50937 2338 50966 2912
rect 50878 2325 50966 2338
rect 51066 2912 51170 2925
rect 51066 2338 51095 2912
rect 51141 2338 51170 2912
rect 51066 2325 51170 2338
rect 51270 2912 51358 2925
rect 51270 2338 51299 2912
rect 51345 2338 51358 2912
rect 51270 2325 51358 2338
rect 51562 2912 51650 2925
rect 51562 2338 51575 2912
rect 51621 2338 51650 2912
rect 51562 2325 51650 2338
rect 51750 2912 51854 2925
rect 51750 2338 51779 2912
rect 51825 2338 51854 2912
rect 51750 2325 51854 2338
rect 51954 2912 52042 2925
rect 51954 2338 51983 2912
rect 52029 2338 52042 2912
rect 51954 2325 52042 2338
rect 52246 2912 52334 2925
rect 52246 2338 52259 2912
rect 52305 2338 52334 2912
rect 52246 2325 52334 2338
rect 52434 2912 52522 2925
rect 52434 2338 52463 2912
rect 52509 2338 52522 2912
rect 52434 2325 52522 2338
rect 53792 2998 53880 3011
rect 53792 2524 53805 2998
rect 53851 2524 53880 2998
rect 53792 2511 53880 2524
rect 53960 2998 54064 3011
rect 53960 2524 53989 2998
rect 54035 2524 54064 2998
rect 53960 2511 54064 2524
rect 54144 2998 54248 3011
rect 54144 2524 54173 2998
rect 54219 2524 54248 2998
rect 54144 2511 54248 2524
rect 54328 2998 54416 3011
rect 54328 2524 54357 2998
rect 54403 2524 54416 2998
rect 54328 2511 54416 2524
rect 48650 1748 48738 1761
rect 48650 1174 48663 1748
rect 48709 1174 48738 1748
rect 48650 1161 48738 1174
rect 48838 1748 48926 1761
rect 48838 1174 48867 1748
rect 48913 1174 48926 1748
rect 48838 1161 48926 1174
rect 49538 1748 49626 1761
rect 49538 1174 49551 1748
rect 49597 1174 49626 1748
rect 49538 1161 49626 1174
rect 49726 1748 49814 1761
rect 49726 1174 49755 1748
rect 49801 1174 49814 1748
rect 49726 1161 49814 1174
rect 50018 1748 50106 1761
rect 50018 1174 50031 1748
rect 50077 1174 50106 1748
rect 50018 1161 50106 1174
rect 50206 1748 50294 1761
rect 50206 1174 50235 1748
rect 50281 1174 50294 1748
rect 50206 1161 50294 1174
<< ndiffc >>
rect 6445 8278 6491 8452
rect 6629 8278 6675 8452
rect 6813 8278 6859 8452
rect 6997 8278 7043 8452
rect 15917 8278 15963 8452
rect 16101 8278 16147 8452
rect 16285 8278 16331 8452
rect 16469 8278 16515 8452
rect 25389 8279 25435 8453
rect 25573 8279 25619 8453
rect 25757 8279 25803 8453
rect 25941 8279 25987 8453
rect 34861 8279 34907 8453
rect 35045 8279 35091 8453
rect 35229 8279 35275 8453
rect 35413 8279 35459 8453
rect 44333 8279 44379 8453
rect 44517 8279 44563 8453
rect 44701 8279 44747 8453
rect 44885 8279 44931 8453
rect 53805 8279 53851 8453
rect 53989 8279 54035 8453
rect 54173 8279 54219 8453
rect 54357 8279 54403 8453
rect 6445 6073 6491 6247
rect 6629 6073 6675 6247
rect 6813 6073 6859 6247
rect 6997 6073 7043 6247
rect 7931 6073 7977 6247
rect 8115 6073 8161 6247
rect 8299 6073 8345 6247
rect 8483 6073 8529 6247
rect 15917 6073 15963 6247
rect 16101 6073 16147 6247
rect 16285 6073 16331 6247
rect 16469 6073 16515 6247
rect 17403 6073 17449 6247
rect 17587 6073 17633 6247
rect 17771 6073 17817 6247
rect 17955 6073 18001 6247
rect 25389 6074 25435 6248
rect 25573 6074 25619 6248
rect 25757 6074 25803 6248
rect 25941 6074 25987 6248
rect 26875 6074 26921 6248
rect 27059 6074 27105 6248
rect 27243 6074 27289 6248
rect 27427 6074 27473 6248
rect 34861 6074 34907 6248
rect 35045 6074 35091 6248
rect 35229 6074 35275 6248
rect 35413 6074 35459 6248
rect 36347 6074 36393 6248
rect 36531 6074 36577 6248
rect 36715 6074 36761 6248
rect 36899 6074 36945 6248
rect 44333 6074 44379 6248
rect 44517 6074 44563 6248
rect 44701 6074 44747 6248
rect 44885 6074 44931 6248
rect 45819 6074 45865 6248
rect 46003 6074 46049 6248
rect 46187 6074 46233 6248
rect 46371 6074 46417 6248
rect 53805 6074 53851 6248
rect 53989 6074 54035 6248
rect 54173 6074 54219 6248
rect 54357 6074 54403 6248
rect 55291 6074 55337 6248
rect 55475 6074 55521 6248
rect 55659 6074 55705 6248
rect 55843 6074 55889 6248
rect 6445 3868 6491 4042
rect 6629 3868 6675 4042
rect 6813 3868 6859 4042
rect 6997 3868 7043 4042
rect 7931 3869 7977 4043
rect 8115 3869 8161 4043
rect 8299 3869 8345 4043
rect 8483 3869 8529 4043
rect 15917 3868 15963 4042
rect 16101 3868 16147 4042
rect 16285 3868 16331 4042
rect 16469 3868 16515 4042
rect 17403 3869 17449 4043
rect 17587 3869 17633 4043
rect 17771 3869 17817 4043
rect 17955 3869 18001 4043
rect 25389 3869 25435 4043
rect 25573 3869 25619 4043
rect 25757 3869 25803 4043
rect 25941 3869 25987 4043
rect 26875 3870 26921 4044
rect 27059 3870 27105 4044
rect 27243 3870 27289 4044
rect 27427 3870 27473 4044
rect 34861 3869 34907 4043
rect 35045 3869 35091 4043
rect 35229 3869 35275 4043
rect 35413 3869 35459 4043
rect 36347 3870 36393 4044
rect 36531 3870 36577 4044
rect 36715 3870 36761 4044
rect 36899 3870 36945 4044
rect 44333 3869 44379 4043
rect 44517 3869 44563 4043
rect 44701 3869 44747 4043
rect 44885 3869 44931 4043
rect 45819 3870 45865 4044
rect 46003 3870 46049 4044
rect 46187 3870 46233 4044
rect 46371 3870 46417 4044
rect 53805 3869 53851 4043
rect 53989 3869 54035 4043
rect 54173 3869 54219 4043
rect 54357 3869 54403 4043
rect 55291 3870 55337 4044
rect 55475 3870 55521 4044
rect 55659 3870 55705 4044
rect 55843 3870 55889 4044
rect 1303 2793 1349 2967
rect 1507 2793 1553 2967
rect 1711 2793 1757 2967
rect 1987 2793 2033 2967
rect 2191 2793 2237 2967
rect 2395 2793 2441 2967
rect 2671 2793 2717 2967
rect 2875 2793 2921 2967
rect 409 1373 455 1547
rect 613 1373 659 1547
rect 3531 1617 3577 1791
rect 3735 1617 3781 1791
rect 4215 1617 4261 1791
rect 4419 1617 4465 1791
rect 4899 1617 4945 1791
rect 5103 1617 5149 1791
rect 6445 1663 6491 1837
rect 6629 1663 6675 1837
rect 6813 1663 6859 1837
rect 6997 1663 7043 1837
rect 10775 2793 10821 2967
rect 10979 2793 11025 2967
rect 11183 2793 11229 2967
rect 11459 2793 11505 2967
rect 11663 2793 11709 2967
rect 11867 2793 11913 2967
rect 12143 2793 12189 2967
rect 12347 2793 12393 2967
rect 9881 1373 9927 1547
rect 10085 1373 10131 1547
rect 13003 1617 13049 1791
rect 13207 1617 13253 1791
rect 13687 1617 13733 1791
rect 13891 1617 13937 1791
rect 14371 1617 14417 1791
rect 14575 1617 14621 1791
rect 15917 1663 15963 1837
rect 16101 1663 16147 1837
rect 16285 1663 16331 1837
rect 16469 1663 16515 1837
rect 20247 2794 20293 2968
rect 20451 2794 20497 2968
rect 20655 2794 20701 2968
rect 20931 2794 20977 2968
rect 21135 2794 21181 2968
rect 21339 2794 21385 2968
rect 21615 2794 21661 2968
rect 21819 2794 21865 2968
rect 19353 1374 19399 1548
rect 19557 1374 19603 1548
rect 22475 1618 22521 1792
rect 22679 1618 22725 1792
rect 23159 1618 23205 1792
rect 23363 1618 23409 1792
rect 23843 1618 23889 1792
rect 24047 1618 24093 1792
rect 25389 1664 25435 1838
rect 25573 1664 25619 1838
rect 25757 1664 25803 1838
rect 25941 1664 25987 1838
rect 29719 2794 29765 2968
rect 29923 2794 29969 2968
rect 30127 2794 30173 2968
rect 30403 2794 30449 2968
rect 30607 2794 30653 2968
rect 30811 2794 30857 2968
rect 31087 2794 31133 2968
rect 31291 2794 31337 2968
rect 28825 1374 28871 1548
rect 29029 1374 29075 1548
rect 31947 1618 31993 1792
rect 32151 1618 32197 1792
rect 32631 1618 32677 1792
rect 32835 1618 32881 1792
rect 33315 1618 33361 1792
rect 33519 1618 33565 1792
rect 34861 1664 34907 1838
rect 35045 1664 35091 1838
rect 35229 1664 35275 1838
rect 35413 1664 35459 1838
rect 39191 2794 39237 2968
rect 39395 2794 39441 2968
rect 39599 2794 39645 2968
rect 39875 2794 39921 2968
rect 40079 2794 40125 2968
rect 40283 2794 40329 2968
rect 40559 2794 40605 2968
rect 40763 2794 40809 2968
rect 38297 1374 38343 1548
rect 38501 1374 38547 1548
rect 41419 1618 41465 1792
rect 41623 1618 41669 1792
rect 42103 1618 42149 1792
rect 42307 1618 42353 1792
rect 42787 1618 42833 1792
rect 42991 1618 43037 1792
rect 44333 1664 44379 1838
rect 44517 1664 44563 1838
rect 44701 1664 44747 1838
rect 44885 1664 44931 1838
rect 48663 2794 48709 2968
rect 48867 2794 48913 2968
rect 49071 2794 49117 2968
rect 49347 2794 49393 2968
rect 49551 2794 49597 2968
rect 49755 2794 49801 2968
rect 50031 2794 50077 2968
rect 50235 2794 50281 2968
rect 47769 1374 47815 1548
rect 47973 1374 48019 1548
rect 50891 1618 50937 1792
rect 51095 1618 51141 1792
rect 51575 1618 51621 1792
rect 51779 1618 51825 1792
rect 52259 1618 52305 1792
rect 52463 1618 52509 1792
rect 53805 1664 53851 1838
rect 53989 1664 54035 1838
rect 54173 1664 54219 1838
rect 54357 1664 54403 1838
rect 1303 453 1349 627
rect 1507 453 1553 627
rect 1711 453 1757 627
rect 1987 453 2033 627
rect 2191 453 2237 627
rect 2395 453 2441 627
rect 2671 453 2717 627
rect 2875 453 2921 627
rect 10775 453 10821 627
rect 10979 453 11025 627
rect 11183 453 11229 627
rect 11459 453 11505 627
rect 11663 453 11709 627
rect 11867 453 11913 627
rect 12143 453 12189 627
rect 12347 453 12393 627
rect 20247 454 20293 628
rect 20451 454 20497 628
rect 20655 454 20701 628
rect 20931 454 20977 628
rect 21135 454 21181 628
rect 21339 454 21385 628
rect 21615 454 21661 628
rect 21819 454 21865 628
rect 29719 454 29765 628
rect 29923 454 29969 628
rect 30127 454 30173 628
rect 30403 454 30449 628
rect 30607 454 30653 628
rect 30811 454 30857 628
rect 31087 454 31133 628
rect 31291 454 31337 628
rect 39191 454 39237 628
rect 39395 454 39441 628
rect 39599 454 39645 628
rect 39875 454 39921 628
rect 40079 454 40125 628
rect 40283 454 40329 628
rect 40559 454 40605 628
rect 40763 454 40809 628
rect 48663 454 48709 628
rect 48867 454 48913 628
rect 49071 454 49117 628
rect 49347 454 49393 628
rect 49551 454 49597 628
rect 49755 454 49801 628
rect 50031 454 50077 628
rect 50235 454 50281 628
<< pdiffc >>
rect 6445 9138 6491 9612
rect 6629 9138 6675 9612
rect 6813 9138 6859 9612
rect 6997 9138 7043 9612
rect 15917 9138 15963 9612
rect 16101 9138 16147 9612
rect 16285 9138 16331 9612
rect 16469 9138 16515 9612
rect 25389 9139 25435 9613
rect 25573 9139 25619 9613
rect 25757 9139 25803 9613
rect 25941 9139 25987 9613
rect 34861 9139 34907 9613
rect 35045 9139 35091 9613
rect 35229 9139 35275 9613
rect 35413 9139 35459 9613
rect 44333 9139 44379 9613
rect 44517 9139 44563 9613
rect 44701 9139 44747 9613
rect 44885 9139 44931 9613
rect 53805 9139 53851 9613
rect 53989 9139 54035 9613
rect 54173 9139 54219 9613
rect 54357 9139 54403 9613
rect 6445 6933 6491 7407
rect 6629 6933 6675 7407
rect 6813 6933 6859 7407
rect 6997 6933 7043 7407
rect 7931 6933 7977 7407
rect 8115 6933 8161 7407
rect 8299 6933 8345 7407
rect 8483 6933 8529 7407
rect 15917 6933 15963 7407
rect 16101 6933 16147 7407
rect 16285 6933 16331 7407
rect 16469 6933 16515 7407
rect 17403 6933 17449 7407
rect 17587 6933 17633 7407
rect 17771 6933 17817 7407
rect 17955 6933 18001 7407
rect 25389 6934 25435 7408
rect 25573 6934 25619 7408
rect 25757 6934 25803 7408
rect 25941 6934 25987 7408
rect 26875 6934 26921 7408
rect 27059 6934 27105 7408
rect 27243 6934 27289 7408
rect 27427 6934 27473 7408
rect 34861 6934 34907 7408
rect 35045 6934 35091 7408
rect 35229 6934 35275 7408
rect 35413 6934 35459 7408
rect 36347 6934 36393 7408
rect 36531 6934 36577 7408
rect 36715 6934 36761 7408
rect 36899 6934 36945 7408
rect 44333 6934 44379 7408
rect 44517 6934 44563 7408
rect 44701 6934 44747 7408
rect 44885 6934 44931 7408
rect 45819 6934 45865 7408
rect 46003 6934 46049 7408
rect 46187 6934 46233 7408
rect 46371 6934 46417 7408
rect 53805 6934 53851 7408
rect 53989 6934 54035 7408
rect 54173 6934 54219 7408
rect 54357 6934 54403 7408
rect 55291 6934 55337 7408
rect 55475 6934 55521 7408
rect 55659 6934 55705 7408
rect 55843 6934 55889 7408
rect 6445 4728 6491 5202
rect 6629 4728 6675 5202
rect 6813 4728 6859 5202
rect 6997 4728 7043 5202
rect 7931 4729 7977 5203
rect 8115 4729 8161 5203
rect 8299 4729 8345 5203
rect 8483 4729 8529 5203
rect 15917 4728 15963 5202
rect 16101 4728 16147 5202
rect 16285 4728 16331 5202
rect 16469 4728 16515 5202
rect 17403 4729 17449 5203
rect 17587 4729 17633 5203
rect 17771 4729 17817 5203
rect 17955 4729 18001 5203
rect 25389 4729 25435 5203
rect 25573 4729 25619 5203
rect 25757 4729 25803 5203
rect 25941 4729 25987 5203
rect 26875 4730 26921 5204
rect 27059 4730 27105 5204
rect 27243 4730 27289 5204
rect 27427 4730 27473 5204
rect 34861 4729 34907 5203
rect 35045 4729 35091 5203
rect 35229 4729 35275 5203
rect 35413 4729 35459 5203
rect 36347 4730 36393 5204
rect 36531 4730 36577 5204
rect 36715 4730 36761 5204
rect 36899 4730 36945 5204
rect 44333 4729 44379 5203
rect 44517 4729 44563 5203
rect 44701 4729 44747 5203
rect 44885 4729 44931 5203
rect 45819 4730 45865 5204
rect 46003 4730 46049 5204
rect 46187 4730 46233 5204
rect 46371 4730 46417 5204
rect 53805 4729 53851 5203
rect 53989 4729 54035 5203
rect 54173 4729 54219 5203
rect 54357 4729 54403 5203
rect 55291 4730 55337 5204
rect 55475 4730 55521 5204
rect 55659 4730 55705 5204
rect 55843 4730 55889 5204
rect 1303 3513 1349 4087
rect 1507 3513 1553 4087
rect 2191 3513 2237 4087
rect 2395 3513 2441 4087
rect 2671 3513 2717 4087
rect 2875 3513 2921 4087
rect 10775 3513 10821 4087
rect 10979 3513 11025 4087
rect 11663 3513 11709 4087
rect 11867 3513 11913 4087
rect 12143 3513 12189 4087
rect 12347 3513 12393 4087
rect 20247 3514 20293 4088
rect 20451 3514 20497 4088
rect 21135 3514 21181 4088
rect 21339 3514 21385 4088
rect 21615 3514 21661 4088
rect 21819 3514 21865 4088
rect 29719 3514 29765 4088
rect 29923 3514 29969 4088
rect 30607 3514 30653 4088
rect 30811 3514 30857 4088
rect 31087 3514 31133 4088
rect 31291 3514 31337 4088
rect 39191 3514 39237 4088
rect 39395 3514 39441 4088
rect 40079 3514 40125 4088
rect 40283 3514 40329 4088
rect 40559 3514 40605 4088
rect 40763 3514 40809 4088
rect 48663 3514 48709 4088
rect 48867 3514 48913 4088
rect 49551 3514 49597 4088
rect 49755 3514 49801 4088
rect 50031 3514 50077 4088
rect 50235 3514 50281 4088
rect 409 2093 455 2667
rect 613 2093 659 2667
rect 3531 2337 3577 2911
rect 3735 2337 3781 2911
rect 3939 2337 3985 2911
rect 4215 2337 4261 2911
rect 4419 2337 4465 2911
rect 4623 2337 4669 2911
rect 4899 2337 4945 2911
rect 5103 2337 5149 2911
rect 6445 2523 6491 2997
rect 6629 2523 6675 2997
rect 6813 2523 6859 2997
rect 6997 2523 7043 2997
rect 1303 1173 1349 1747
rect 1507 1173 1553 1747
rect 2191 1173 2237 1747
rect 2395 1173 2441 1747
rect 2671 1173 2717 1747
rect 2875 1173 2921 1747
rect 9881 2093 9927 2667
rect 10085 2093 10131 2667
rect 13003 2337 13049 2911
rect 13207 2337 13253 2911
rect 13411 2337 13457 2911
rect 13687 2337 13733 2911
rect 13891 2337 13937 2911
rect 14095 2337 14141 2911
rect 14371 2337 14417 2911
rect 14575 2337 14621 2911
rect 15917 2523 15963 2997
rect 16101 2523 16147 2997
rect 16285 2523 16331 2997
rect 16469 2523 16515 2997
rect 10775 1173 10821 1747
rect 10979 1173 11025 1747
rect 11663 1173 11709 1747
rect 11867 1173 11913 1747
rect 12143 1173 12189 1747
rect 12347 1173 12393 1747
rect 19353 2094 19399 2668
rect 19557 2094 19603 2668
rect 22475 2338 22521 2912
rect 22679 2338 22725 2912
rect 22883 2338 22929 2912
rect 23159 2338 23205 2912
rect 23363 2338 23409 2912
rect 23567 2338 23613 2912
rect 23843 2338 23889 2912
rect 24047 2338 24093 2912
rect 25389 2524 25435 2998
rect 25573 2524 25619 2998
rect 25757 2524 25803 2998
rect 25941 2524 25987 2998
rect 20247 1174 20293 1748
rect 20451 1174 20497 1748
rect 21135 1174 21181 1748
rect 21339 1174 21385 1748
rect 21615 1174 21661 1748
rect 21819 1174 21865 1748
rect 28825 2094 28871 2668
rect 29029 2094 29075 2668
rect 31947 2338 31993 2912
rect 32151 2338 32197 2912
rect 32355 2338 32401 2912
rect 32631 2338 32677 2912
rect 32835 2338 32881 2912
rect 33039 2338 33085 2912
rect 33315 2338 33361 2912
rect 33519 2338 33565 2912
rect 34861 2524 34907 2998
rect 35045 2524 35091 2998
rect 35229 2524 35275 2998
rect 35413 2524 35459 2998
rect 29719 1174 29765 1748
rect 29923 1174 29969 1748
rect 30607 1174 30653 1748
rect 30811 1174 30857 1748
rect 31087 1174 31133 1748
rect 31291 1174 31337 1748
rect 38297 2094 38343 2668
rect 38501 2094 38547 2668
rect 41419 2338 41465 2912
rect 41623 2338 41669 2912
rect 41827 2338 41873 2912
rect 42103 2338 42149 2912
rect 42307 2338 42353 2912
rect 42511 2338 42557 2912
rect 42787 2338 42833 2912
rect 42991 2338 43037 2912
rect 44333 2524 44379 2998
rect 44517 2524 44563 2998
rect 44701 2524 44747 2998
rect 44885 2524 44931 2998
rect 39191 1174 39237 1748
rect 39395 1174 39441 1748
rect 40079 1174 40125 1748
rect 40283 1174 40329 1748
rect 40559 1174 40605 1748
rect 40763 1174 40809 1748
rect 47769 2094 47815 2668
rect 47973 2094 48019 2668
rect 50891 2338 50937 2912
rect 51095 2338 51141 2912
rect 51299 2338 51345 2912
rect 51575 2338 51621 2912
rect 51779 2338 51825 2912
rect 51983 2338 52029 2912
rect 52259 2338 52305 2912
rect 52463 2338 52509 2912
rect 53805 2524 53851 2998
rect 53989 2524 54035 2998
rect 54173 2524 54219 2998
rect 54357 2524 54403 2998
rect 48663 1174 48709 1748
rect 48867 1174 48913 1748
rect 49551 1174 49597 1748
rect 49755 1174 49801 1748
rect 50031 1174 50077 1748
rect 50235 1174 50281 1748
<< psubdiff >>
rect 6294 8579 7194 8651
rect 6294 8535 6366 8579
rect 6294 8195 6307 8535
rect 6353 8195 6366 8535
rect 7122 8535 7194 8579
rect 6294 8151 6366 8195
rect 7122 8195 7135 8535
rect 7181 8195 7194 8535
rect 7122 8151 7194 8195
rect 6294 8079 7194 8151
rect 15766 8579 16666 8651
rect 15766 8535 15838 8579
rect 15766 8195 15779 8535
rect 15825 8195 15838 8535
rect 16594 8535 16666 8579
rect 15766 8151 15838 8195
rect 16594 8195 16607 8535
rect 16653 8195 16666 8535
rect 16594 8151 16666 8195
rect 15766 8079 16666 8151
rect 25238 8580 26138 8652
rect 25238 8536 25310 8580
rect 25238 8196 25251 8536
rect 25297 8196 25310 8536
rect 26066 8536 26138 8580
rect 25238 8152 25310 8196
rect 26066 8196 26079 8536
rect 26125 8196 26138 8536
rect 26066 8152 26138 8196
rect 25238 8080 26138 8152
rect 34710 8580 35610 8652
rect 34710 8536 34782 8580
rect 34710 8196 34723 8536
rect 34769 8196 34782 8536
rect 35538 8536 35610 8580
rect 34710 8152 34782 8196
rect 35538 8196 35551 8536
rect 35597 8196 35610 8536
rect 35538 8152 35610 8196
rect 34710 8080 35610 8152
rect 44182 8580 45082 8652
rect 44182 8536 44254 8580
rect 44182 8196 44195 8536
rect 44241 8196 44254 8536
rect 45010 8536 45082 8580
rect 44182 8152 44254 8196
rect 45010 8196 45023 8536
rect 45069 8196 45082 8536
rect 45010 8152 45082 8196
rect 44182 8080 45082 8152
rect 53654 8580 54554 8652
rect 53654 8536 53726 8580
rect 53654 8196 53667 8536
rect 53713 8196 53726 8536
rect 54482 8536 54554 8580
rect 53654 8152 53726 8196
rect 54482 8196 54495 8536
rect 54541 8196 54554 8536
rect 54482 8152 54554 8196
rect 53654 8080 54554 8152
rect 6294 6374 7194 6446
rect 6294 6330 6366 6374
rect 6294 5990 6307 6330
rect 6353 5990 6366 6330
rect 7122 6330 7194 6374
rect 6294 5946 6366 5990
rect 7122 5990 7135 6330
rect 7181 5990 7194 6330
rect 7122 5946 7194 5990
rect 6294 5874 7194 5946
rect 7780 6374 8680 6446
rect 7780 6330 7852 6374
rect 7780 5990 7793 6330
rect 7839 5990 7852 6330
rect 8608 6330 8680 6374
rect 7780 5946 7852 5990
rect 8608 5990 8621 6330
rect 8667 5990 8680 6330
rect 8608 5946 8680 5990
rect 7780 5874 8680 5946
rect 15766 6374 16666 6446
rect 15766 6330 15838 6374
rect 15766 5990 15779 6330
rect 15825 5990 15838 6330
rect 16594 6330 16666 6374
rect 15766 5946 15838 5990
rect 16594 5990 16607 6330
rect 16653 5990 16666 6330
rect 16594 5946 16666 5990
rect 15766 5874 16666 5946
rect 17252 6374 18152 6446
rect 17252 6330 17324 6374
rect 17252 5990 17265 6330
rect 17311 5990 17324 6330
rect 18080 6330 18152 6374
rect 17252 5946 17324 5990
rect 18080 5990 18093 6330
rect 18139 5990 18152 6330
rect 18080 5946 18152 5990
rect 17252 5874 18152 5946
rect 25238 6375 26138 6447
rect 25238 6331 25310 6375
rect 25238 5991 25251 6331
rect 25297 5991 25310 6331
rect 26066 6331 26138 6375
rect 25238 5947 25310 5991
rect 26066 5991 26079 6331
rect 26125 5991 26138 6331
rect 26066 5947 26138 5991
rect 25238 5875 26138 5947
rect 26724 6375 27624 6447
rect 26724 6331 26796 6375
rect 26724 5991 26737 6331
rect 26783 5991 26796 6331
rect 27552 6331 27624 6375
rect 26724 5947 26796 5991
rect 27552 5991 27565 6331
rect 27611 5991 27624 6331
rect 27552 5947 27624 5991
rect 26724 5875 27624 5947
rect 34710 6375 35610 6447
rect 34710 6331 34782 6375
rect 34710 5991 34723 6331
rect 34769 5991 34782 6331
rect 35538 6331 35610 6375
rect 34710 5947 34782 5991
rect 35538 5991 35551 6331
rect 35597 5991 35610 6331
rect 35538 5947 35610 5991
rect 34710 5875 35610 5947
rect 36196 6375 37096 6447
rect 36196 6331 36268 6375
rect 36196 5991 36209 6331
rect 36255 5991 36268 6331
rect 37024 6331 37096 6375
rect 36196 5947 36268 5991
rect 37024 5991 37037 6331
rect 37083 5991 37096 6331
rect 37024 5947 37096 5991
rect 36196 5875 37096 5947
rect 44182 6375 45082 6447
rect 44182 6331 44254 6375
rect 44182 5991 44195 6331
rect 44241 5991 44254 6331
rect 45010 6331 45082 6375
rect 44182 5947 44254 5991
rect 45010 5991 45023 6331
rect 45069 5991 45082 6331
rect 45010 5947 45082 5991
rect 44182 5875 45082 5947
rect 45668 6375 46568 6447
rect 45668 6331 45740 6375
rect 45668 5991 45681 6331
rect 45727 5991 45740 6331
rect 46496 6331 46568 6375
rect 45668 5947 45740 5991
rect 46496 5991 46509 6331
rect 46555 5991 46568 6331
rect 46496 5947 46568 5991
rect 45668 5875 46568 5947
rect 53654 6375 54554 6447
rect 53654 6331 53726 6375
rect 53654 5991 53667 6331
rect 53713 5991 53726 6331
rect 54482 6331 54554 6375
rect 53654 5947 53726 5991
rect 54482 5991 54495 6331
rect 54541 5991 54554 6331
rect 54482 5947 54554 5991
rect 53654 5875 54554 5947
rect 55140 6375 56040 6447
rect 55140 6331 55212 6375
rect 55140 5991 55153 6331
rect 55199 5991 55212 6331
rect 55968 6331 56040 6375
rect 55140 5947 55212 5991
rect 55968 5991 55981 6331
rect 56027 5991 56040 6331
rect 55968 5947 56040 5991
rect 55140 5875 56040 5947
rect 6294 4169 7194 4241
rect 6294 4125 6366 4169
rect 6294 3785 6307 4125
rect 6353 3785 6366 4125
rect 7122 4125 7194 4169
rect 6294 3741 6366 3785
rect 7122 3785 7135 4125
rect 7181 3785 7194 4125
rect 7122 3741 7194 3785
rect 6294 3669 7194 3741
rect 7780 4170 8680 4242
rect 7780 4126 7852 4170
rect 7780 3786 7793 4126
rect 7839 3786 7852 4126
rect 8608 4126 8680 4170
rect 7780 3742 7852 3786
rect 8608 3786 8621 4126
rect 8667 3786 8680 4126
rect 8608 3742 8680 3786
rect 7780 3670 8680 3742
rect 15766 4169 16666 4241
rect 15766 4125 15838 4169
rect 15766 3785 15779 4125
rect 15825 3785 15838 4125
rect 16594 4125 16666 4169
rect 15766 3741 15838 3785
rect 16594 3785 16607 4125
rect 16653 3785 16666 4125
rect 16594 3741 16666 3785
rect 15766 3669 16666 3741
rect 17252 4170 18152 4242
rect 17252 4126 17324 4170
rect 17252 3786 17265 4126
rect 17311 3786 17324 4126
rect 18080 4126 18152 4170
rect 17252 3742 17324 3786
rect 18080 3786 18093 4126
rect 18139 3786 18152 4126
rect 18080 3742 18152 3786
rect 17252 3670 18152 3742
rect 25238 4170 26138 4242
rect 25238 4126 25310 4170
rect 25238 3786 25251 4126
rect 25297 3786 25310 4126
rect 26066 4126 26138 4170
rect 25238 3742 25310 3786
rect 26066 3786 26079 4126
rect 26125 3786 26138 4126
rect 26066 3742 26138 3786
rect 25238 3670 26138 3742
rect 26724 4171 27624 4243
rect 26724 4127 26796 4171
rect 26724 3787 26737 4127
rect 26783 3787 26796 4127
rect 27552 4127 27624 4171
rect 26724 3743 26796 3787
rect 27552 3787 27565 4127
rect 27611 3787 27624 4127
rect 27552 3743 27624 3787
rect 26724 3671 27624 3743
rect 34710 4170 35610 4242
rect 34710 4126 34782 4170
rect 34710 3786 34723 4126
rect 34769 3786 34782 4126
rect 35538 4126 35610 4170
rect 34710 3742 34782 3786
rect 35538 3786 35551 4126
rect 35597 3786 35610 4126
rect 35538 3742 35610 3786
rect 34710 3670 35610 3742
rect 36196 4171 37096 4243
rect 36196 4127 36268 4171
rect 36196 3787 36209 4127
rect 36255 3787 36268 4127
rect 37024 4127 37096 4171
rect 36196 3743 36268 3787
rect 37024 3787 37037 4127
rect 37083 3787 37096 4127
rect 37024 3743 37096 3787
rect 36196 3671 37096 3743
rect 44182 4170 45082 4242
rect 44182 4126 44254 4170
rect 44182 3786 44195 4126
rect 44241 3786 44254 4126
rect 45010 4126 45082 4170
rect 44182 3742 44254 3786
rect 45010 3786 45023 4126
rect 45069 3786 45082 4126
rect 45010 3742 45082 3786
rect 44182 3670 45082 3742
rect 45668 4171 46568 4243
rect 45668 4127 45740 4171
rect 45668 3787 45681 4127
rect 45727 3787 45740 4127
rect 46496 4127 46568 4171
rect 45668 3743 45740 3787
rect 46496 3787 46509 4127
rect 46555 3787 46568 4127
rect 46496 3743 46568 3787
rect 45668 3671 46568 3743
rect 53654 4170 54554 4242
rect 53654 4126 53726 4170
rect 53654 3786 53667 4126
rect 53713 3786 53726 4126
rect 54482 4126 54554 4170
rect 53654 3742 53726 3786
rect 54482 3786 54495 4126
rect 54541 3786 54554 4126
rect 54482 3742 54554 3786
rect 53654 3670 54554 3742
rect 55140 4171 56040 4243
rect 55140 4127 55212 4171
rect 55140 3787 55153 4127
rect 55199 3787 55212 4127
rect 55968 4127 56040 4171
rect 55140 3743 55212 3787
rect 55968 3787 55981 4127
rect 56027 3787 56040 4127
rect 55968 3743 56040 3787
rect 55140 3671 56040 3743
rect 1152 3094 3072 3166
rect 1152 3050 1224 3094
rect 1152 2710 1165 3050
rect 1211 2710 1224 3050
rect 1836 3050 1908 3094
rect 1152 2666 1224 2710
rect 1836 2710 1849 3050
rect 1895 2710 1908 3050
rect 2520 3050 2592 3094
rect 1836 2666 1908 2710
rect 2520 2710 2533 3050
rect 2579 2710 2592 3050
rect 3000 3050 3072 3094
rect 2520 2666 2592 2710
rect 3000 2710 3013 3050
rect 3059 2710 3072 3050
rect 3000 2666 3072 2710
rect 1152 2594 3072 2666
rect 10624 3094 12544 3166
rect 10624 3050 10696 3094
rect 258 1674 810 1746
rect 258 1630 330 1674
rect 258 1290 271 1630
rect 317 1290 330 1630
rect 738 1630 810 1674
rect 258 1246 330 1290
rect 738 1290 751 1630
rect 797 1290 810 1630
rect 738 1246 810 1290
rect 258 1174 810 1246
rect 3380 1918 3932 1990
rect 3380 1874 3452 1918
rect 3380 1534 3393 1874
rect 3439 1534 3452 1874
rect 3860 1874 3932 1918
rect 3380 1490 3452 1534
rect 3860 1534 3873 1874
rect 3919 1534 3932 1874
rect 3860 1490 3932 1534
rect 3380 1418 3932 1490
rect 4064 1918 4616 1990
rect 4064 1874 4136 1918
rect 4064 1534 4077 1874
rect 4123 1534 4136 1874
rect 4544 1874 4616 1918
rect 4064 1490 4136 1534
rect 4544 1534 4557 1874
rect 4603 1534 4616 1874
rect 4544 1490 4616 1534
rect 4064 1418 4616 1490
rect 4748 1918 5300 1990
rect 4748 1874 4820 1918
rect 4748 1534 4761 1874
rect 4807 1534 4820 1874
rect 5228 1874 5300 1918
rect 4748 1490 4820 1534
rect 5228 1534 5241 1874
rect 5287 1534 5300 1874
rect 5228 1490 5300 1534
rect 4748 1418 5300 1490
rect 6294 1964 7194 2036
rect 6294 1920 6366 1964
rect 6294 1580 6307 1920
rect 6353 1580 6366 1920
rect 7122 1920 7194 1964
rect 6294 1536 6366 1580
rect 7122 1580 7135 1920
rect 7181 1580 7194 1920
rect 10624 2710 10637 3050
rect 10683 2710 10696 3050
rect 11308 3050 11380 3094
rect 10624 2666 10696 2710
rect 11308 2710 11321 3050
rect 11367 2710 11380 3050
rect 11992 3050 12064 3094
rect 11308 2666 11380 2710
rect 11992 2710 12005 3050
rect 12051 2710 12064 3050
rect 12472 3050 12544 3094
rect 11992 2666 12064 2710
rect 12472 2710 12485 3050
rect 12531 2710 12544 3050
rect 12472 2666 12544 2710
rect 10624 2594 12544 2666
rect 20096 3095 22016 3167
rect 20096 3051 20168 3095
rect 7122 1536 7194 1580
rect 6294 1464 7194 1536
rect 9730 1674 10282 1746
rect 9730 1630 9802 1674
rect 9730 1290 9743 1630
rect 9789 1290 9802 1630
rect 10210 1630 10282 1674
rect 9730 1246 9802 1290
rect 10210 1290 10223 1630
rect 10269 1290 10282 1630
rect 10210 1246 10282 1290
rect 9730 1174 10282 1246
rect 12852 1918 13404 1990
rect 12852 1874 12924 1918
rect 12852 1534 12865 1874
rect 12911 1534 12924 1874
rect 13332 1874 13404 1918
rect 12852 1490 12924 1534
rect 13332 1534 13345 1874
rect 13391 1534 13404 1874
rect 13332 1490 13404 1534
rect 12852 1418 13404 1490
rect 13536 1918 14088 1990
rect 13536 1874 13608 1918
rect 13536 1534 13549 1874
rect 13595 1534 13608 1874
rect 14016 1874 14088 1918
rect 13536 1490 13608 1534
rect 14016 1534 14029 1874
rect 14075 1534 14088 1874
rect 14016 1490 14088 1534
rect 13536 1418 14088 1490
rect 14220 1918 14772 1990
rect 14220 1874 14292 1918
rect 14220 1534 14233 1874
rect 14279 1534 14292 1874
rect 14700 1874 14772 1918
rect 14220 1490 14292 1534
rect 14700 1534 14713 1874
rect 14759 1534 14772 1874
rect 14700 1490 14772 1534
rect 14220 1418 14772 1490
rect 15766 1964 16666 2036
rect 15766 1920 15838 1964
rect 15766 1580 15779 1920
rect 15825 1580 15838 1920
rect 16594 1920 16666 1964
rect 15766 1536 15838 1580
rect 16594 1580 16607 1920
rect 16653 1580 16666 1920
rect 20096 2711 20109 3051
rect 20155 2711 20168 3051
rect 20780 3051 20852 3095
rect 20096 2667 20168 2711
rect 20780 2711 20793 3051
rect 20839 2711 20852 3051
rect 21464 3051 21536 3095
rect 20780 2667 20852 2711
rect 21464 2711 21477 3051
rect 21523 2711 21536 3051
rect 21944 3051 22016 3095
rect 21464 2667 21536 2711
rect 21944 2711 21957 3051
rect 22003 2711 22016 3051
rect 21944 2667 22016 2711
rect 20096 2595 22016 2667
rect 29568 3095 31488 3167
rect 29568 3051 29640 3095
rect 16594 1536 16666 1580
rect 15766 1464 16666 1536
rect 19202 1675 19754 1747
rect 19202 1631 19274 1675
rect 19202 1291 19215 1631
rect 19261 1291 19274 1631
rect 19682 1631 19754 1675
rect 19202 1247 19274 1291
rect 19682 1291 19695 1631
rect 19741 1291 19754 1631
rect 19682 1247 19754 1291
rect 19202 1175 19754 1247
rect 22324 1919 22876 1991
rect 22324 1875 22396 1919
rect 22324 1535 22337 1875
rect 22383 1535 22396 1875
rect 22804 1875 22876 1919
rect 22324 1491 22396 1535
rect 22804 1535 22817 1875
rect 22863 1535 22876 1875
rect 22804 1491 22876 1535
rect 22324 1419 22876 1491
rect 23008 1919 23560 1991
rect 23008 1875 23080 1919
rect 23008 1535 23021 1875
rect 23067 1535 23080 1875
rect 23488 1875 23560 1919
rect 23008 1491 23080 1535
rect 23488 1535 23501 1875
rect 23547 1535 23560 1875
rect 23488 1491 23560 1535
rect 23008 1419 23560 1491
rect 23692 1919 24244 1991
rect 23692 1875 23764 1919
rect 23692 1535 23705 1875
rect 23751 1535 23764 1875
rect 24172 1875 24244 1919
rect 23692 1491 23764 1535
rect 24172 1535 24185 1875
rect 24231 1535 24244 1875
rect 24172 1491 24244 1535
rect 23692 1419 24244 1491
rect 25238 1965 26138 2037
rect 25238 1921 25310 1965
rect 25238 1581 25251 1921
rect 25297 1581 25310 1921
rect 26066 1921 26138 1965
rect 25238 1537 25310 1581
rect 26066 1581 26079 1921
rect 26125 1581 26138 1921
rect 29568 2711 29581 3051
rect 29627 2711 29640 3051
rect 30252 3051 30324 3095
rect 29568 2667 29640 2711
rect 30252 2711 30265 3051
rect 30311 2711 30324 3051
rect 30936 3051 31008 3095
rect 30252 2667 30324 2711
rect 30936 2711 30949 3051
rect 30995 2711 31008 3051
rect 31416 3051 31488 3095
rect 30936 2667 31008 2711
rect 31416 2711 31429 3051
rect 31475 2711 31488 3051
rect 31416 2667 31488 2711
rect 29568 2595 31488 2667
rect 39040 3095 40960 3167
rect 39040 3051 39112 3095
rect 26066 1537 26138 1581
rect 25238 1465 26138 1537
rect 28674 1675 29226 1747
rect 28674 1631 28746 1675
rect 28674 1291 28687 1631
rect 28733 1291 28746 1631
rect 29154 1631 29226 1675
rect 28674 1247 28746 1291
rect 29154 1291 29167 1631
rect 29213 1291 29226 1631
rect 29154 1247 29226 1291
rect 28674 1175 29226 1247
rect 31796 1919 32348 1991
rect 31796 1875 31868 1919
rect 31796 1535 31809 1875
rect 31855 1535 31868 1875
rect 32276 1875 32348 1919
rect 31796 1491 31868 1535
rect 32276 1535 32289 1875
rect 32335 1535 32348 1875
rect 32276 1491 32348 1535
rect 31796 1419 32348 1491
rect 32480 1919 33032 1991
rect 32480 1875 32552 1919
rect 32480 1535 32493 1875
rect 32539 1535 32552 1875
rect 32960 1875 33032 1919
rect 32480 1491 32552 1535
rect 32960 1535 32973 1875
rect 33019 1535 33032 1875
rect 32960 1491 33032 1535
rect 32480 1419 33032 1491
rect 33164 1919 33716 1991
rect 33164 1875 33236 1919
rect 33164 1535 33177 1875
rect 33223 1535 33236 1875
rect 33644 1875 33716 1919
rect 33164 1491 33236 1535
rect 33644 1535 33657 1875
rect 33703 1535 33716 1875
rect 33644 1491 33716 1535
rect 33164 1419 33716 1491
rect 34710 1965 35610 2037
rect 34710 1921 34782 1965
rect 34710 1581 34723 1921
rect 34769 1581 34782 1921
rect 35538 1921 35610 1965
rect 34710 1537 34782 1581
rect 35538 1581 35551 1921
rect 35597 1581 35610 1921
rect 39040 2711 39053 3051
rect 39099 2711 39112 3051
rect 39724 3051 39796 3095
rect 39040 2667 39112 2711
rect 39724 2711 39737 3051
rect 39783 2711 39796 3051
rect 40408 3051 40480 3095
rect 39724 2667 39796 2711
rect 40408 2711 40421 3051
rect 40467 2711 40480 3051
rect 40888 3051 40960 3095
rect 40408 2667 40480 2711
rect 40888 2711 40901 3051
rect 40947 2711 40960 3051
rect 40888 2667 40960 2711
rect 39040 2595 40960 2667
rect 48512 3095 50432 3167
rect 48512 3051 48584 3095
rect 35538 1537 35610 1581
rect 34710 1465 35610 1537
rect 38146 1675 38698 1747
rect 38146 1631 38218 1675
rect 38146 1291 38159 1631
rect 38205 1291 38218 1631
rect 38626 1631 38698 1675
rect 38146 1247 38218 1291
rect 38626 1291 38639 1631
rect 38685 1291 38698 1631
rect 38626 1247 38698 1291
rect 38146 1175 38698 1247
rect 41268 1919 41820 1991
rect 41268 1875 41340 1919
rect 41268 1535 41281 1875
rect 41327 1535 41340 1875
rect 41748 1875 41820 1919
rect 41268 1491 41340 1535
rect 41748 1535 41761 1875
rect 41807 1535 41820 1875
rect 41748 1491 41820 1535
rect 41268 1419 41820 1491
rect 41952 1919 42504 1991
rect 41952 1875 42024 1919
rect 41952 1535 41965 1875
rect 42011 1535 42024 1875
rect 42432 1875 42504 1919
rect 41952 1491 42024 1535
rect 42432 1535 42445 1875
rect 42491 1535 42504 1875
rect 42432 1491 42504 1535
rect 41952 1419 42504 1491
rect 42636 1919 43188 1991
rect 42636 1875 42708 1919
rect 42636 1535 42649 1875
rect 42695 1535 42708 1875
rect 43116 1875 43188 1919
rect 42636 1491 42708 1535
rect 43116 1535 43129 1875
rect 43175 1535 43188 1875
rect 43116 1491 43188 1535
rect 42636 1419 43188 1491
rect 44182 1965 45082 2037
rect 44182 1921 44254 1965
rect 44182 1581 44195 1921
rect 44241 1581 44254 1921
rect 45010 1921 45082 1965
rect 44182 1537 44254 1581
rect 45010 1581 45023 1921
rect 45069 1581 45082 1921
rect 48512 2711 48525 3051
rect 48571 2711 48584 3051
rect 49196 3051 49268 3095
rect 48512 2667 48584 2711
rect 49196 2711 49209 3051
rect 49255 2711 49268 3051
rect 49880 3051 49952 3095
rect 49196 2667 49268 2711
rect 49880 2711 49893 3051
rect 49939 2711 49952 3051
rect 50360 3051 50432 3095
rect 49880 2667 49952 2711
rect 50360 2711 50373 3051
rect 50419 2711 50432 3051
rect 50360 2667 50432 2711
rect 48512 2595 50432 2667
rect 45010 1537 45082 1581
rect 44182 1465 45082 1537
rect 47618 1675 48170 1747
rect 47618 1631 47690 1675
rect 47618 1291 47631 1631
rect 47677 1291 47690 1631
rect 48098 1631 48170 1675
rect 47618 1247 47690 1291
rect 48098 1291 48111 1631
rect 48157 1291 48170 1631
rect 48098 1247 48170 1291
rect 47618 1175 48170 1247
rect 50740 1919 51292 1991
rect 50740 1875 50812 1919
rect 50740 1535 50753 1875
rect 50799 1535 50812 1875
rect 51220 1875 51292 1919
rect 50740 1491 50812 1535
rect 51220 1535 51233 1875
rect 51279 1535 51292 1875
rect 51220 1491 51292 1535
rect 50740 1419 51292 1491
rect 51424 1919 51976 1991
rect 51424 1875 51496 1919
rect 51424 1535 51437 1875
rect 51483 1535 51496 1875
rect 51904 1875 51976 1919
rect 51424 1491 51496 1535
rect 51904 1535 51917 1875
rect 51963 1535 51976 1875
rect 51904 1491 51976 1535
rect 51424 1419 51976 1491
rect 52108 1919 52660 1991
rect 52108 1875 52180 1919
rect 52108 1535 52121 1875
rect 52167 1535 52180 1875
rect 52588 1875 52660 1919
rect 52108 1491 52180 1535
rect 52588 1535 52601 1875
rect 52647 1535 52660 1875
rect 52588 1491 52660 1535
rect 52108 1419 52660 1491
rect 53654 1965 54554 2037
rect 53654 1921 53726 1965
rect 53654 1581 53667 1921
rect 53713 1581 53726 1921
rect 54482 1921 54554 1965
rect 53654 1537 53726 1581
rect 54482 1581 54495 1921
rect 54541 1581 54554 1921
rect 54482 1537 54554 1581
rect 53654 1465 54554 1537
rect 1152 754 3072 826
rect 1152 710 1224 754
rect 1152 370 1165 710
rect 1211 370 1224 710
rect 1836 710 1908 754
rect 1152 326 1224 370
rect 1836 370 1849 710
rect 1895 370 1908 710
rect 2520 710 2592 754
rect 1836 326 1908 370
rect 2520 370 2533 710
rect 2579 370 2592 710
rect 3000 710 3072 754
rect 2520 326 2592 370
rect 3000 370 3013 710
rect 3059 370 3072 710
rect 3000 326 3072 370
rect 1152 254 3072 326
rect 10624 754 12544 826
rect 10624 710 10696 754
rect 10624 370 10637 710
rect 10683 370 10696 710
rect 11308 710 11380 754
rect 10624 326 10696 370
rect 11308 370 11321 710
rect 11367 370 11380 710
rect 11992 710 12064 754
rect 11308 326 11380 370
rect 11992 370 12005 710
rect 12051 370 12064 710
rect 12472 710 12544 754
rect 11992 326 12064 370
rect 12472 370 12485 710
rect 12531 370 12544 710
rect 12472 326 12544 370
rect 10624 254 12544 326
rect 20096 755 22016 827
rect 20096 711 20168 755
rect 20096 371 20109 711
rect 20155 371 20168 711
rect 20780 711 20852 755
rect 20096 327 20168 371
rect 20780 371 20793 711
rect 20839 371 20852 711
rect 21464 711 21536 755
rect 20780 327 20852 371
rect 21464 371 21477 711
rect 21523 371 21536 711
rect 21944 711 22016 755
rect 21464 327 21536 371
rect 21944 371 21957 711
rect 22003 371 22016 711
rect 21944 327 22016 371
rect 20096 255 22016 327
rect 29568 755 31488 827
rect 29568 711 29640 755
rect 29568 371 29581 711
rect 29627 371 29640 711
rect 30252 711 30324 755
rect 29568 327 29640 371
rect 30252 371 30265 711
rect 30311 371 30324 711
rect 30936 711 31008 755
rect 30252 327 30324 371
rect 30936 371 30949 711
rect 30995 371 31008 711
rect 31416 711 31488 755
rect 30936 327 31008 371
rect 31416 371 31429 711
rect 31475 371 31488 711
rect 31416 327 31488 371
rect 29568 255 31488 327
rect 39040 755 40960 827
rect 39040 711 39112 755
rect 39040 371 39053 711
rect 39099 371 39112 711
rect 39724 711 39796 755
rect 39040 327 39112 371
rect 39724 371 39737 711
rect 39783 371 39796 711
rect 40408 711 40480 755
rect 39724 327 39796 371
rect 40408 371 40421 711
rect 40467 371 40480 711
rect 40888 711 40960 755
rect 40408 327 40480 371
rect 40888 371 40901 711
rect 40947 371 40960 711
rect 40888 327 40960 371
rect 39040 255 40960 327
rect 48512 755 50432 827
rect 48512 711 48584 755
rect 48512 371 48525 711
rect 48571 371 48584 711
rect 49196 711 49268 755
rect 48512 327 48584 371
rect 49196 371 49209 711
rect 49255 371 49268 711
rect 49880 711 49952 755
rect 49196 327 49268 371
rect 49880 371 49893 711
rect 49939 371 49952 711
rect 50360 711 50432 755
rect 49880 327 49952 371
rect 50360 371 50373 711
rect 50419 371 50432 711
rect 50360 327 50432 371
rect 48512 255 50432 327
<< nsubdiff >>
rect 6294 9739 7194 9811
rect 6294 9695 6366 9739
rect 6294 9055 6307 9695
rect 6353 9055 6366 9695
rect 7122 9695 7194 9739
rect 6294 9011 6366 9055
rect 7122 9055 7135 9695
rect 7181 9055 7194 9695
rect 7122 9011 7194 9055
rect 6294 8939 7194 9011
rect 15766 9739 16666 9811
rect 15766 9695 15838 9739
rect 15766 9055 15779 9695
rect 15825 9055 15838 9695
rect 16594 9695 16666 9739
rect 15766 9011 15838 9055
rect 16594 9055 16607 9695
rect 16653 9055 16666 9695
rect 16594 9011 16666 9055
rect 15766 8939 16666 9011
rect 25238 9740 26138 9812
rect 25238 9696 25310 9740
rect 25238 9056 25251 9696
rect 25297 9056 25310 9696
rect 26066 9696 26138 9740
rect 25238 9012 25310 9056
rect 26066 9056 26079 9696
rect 26125 9056 26138 9696
rect 26066 9012 26138 9056
rect 25238 8940 26138 9012
rect 34710 9740 35610 9812
rect 34710 9696 34782 9740
rect 34710 9056 34723 9696
rect 34769 9056 34782 9696
rect 35538 9696 35610 9740
rect 34710 9012 34782 9056
rect 35538 9056 35551 9696
rect 35597 9056 35610 9696
rect 35538 9012 35610 9056
rect 34710 8940 35610 9012
rect 44182 9740 45082 9812
rect 44182 9696 44254 9740
rect 44182 9056 44195 9696
rect 44241 9056 44254 9696
rect 45010 9696 45082 9740
rect 44182 9012 44254 9056
rect 45010 9056 45023 9696
rect 45069 9056 45082 9696
rect 45010 9012 45082 9056
rect 44182 8940 45082 9012
rect 53654 9740 54554 9812
rect 53654 9696 53726 9740
rect 53654 9056 53667 9696
rect 53713 9056 53726 9696
rect 54482 9696 54554 9740
rect 53654 9012 53726 9056
rect 54482 9056 54495 9696
rect 54541 9056 54554 9696
rect 54482 9012 54554 9056
rect 53654 8940 54554 9012
rect 6294 7534 7194 7606
rect 6294 7490 6366 7534
rect 6294 6850 6307 7490
rect 6353 6850 6366 7490
rect 7122 7490 7194 7534
rect 6294 6806 6366 6850
rect 7122 6850 7135 7490
rect 7181 6850 7194 7490
rect 7122 6806 7194 6850
rect 6294 6734 7194 6806
rect 7780 7534 8680 7606
rect 7780 7490 7852 7534
rect 7780 6850 7793 7490
rect 7839 6850 7852 7490
rect 8608 7490 8680 7534
rect 7780 6806 7852 6850
rect 8608 6850 8621 7490
rect 8667 6850 8680 7490
rect 8608 6806 8680 6850
rect 7780 6734 8680 6806
rect 15766 7534 16666 7606
rect 15766 7490 15838 7534
rect 15766 6850 15779 7490
rect 15825 6850 15838 7490
rect 16594 7490 16666 7534
rect 15766 6806 15838 6850
rect 16594 6850 16607 7490
rect 16653 6850 16666 7490
rect 16594 6806 16666 6850
rect 15766 6734 16666 6806
rect 17252 7534 18152 7606
rect 17252 7490 17324 7534
rect 17252 6850 17265 7490
rect 17311 6850 17324 7490
rect 18080 7490 18152 7534
rect 17252 6806 17324 6850
rect 18080 6850 18093 7490
rect 18139 6850 18152 7490
rect 18080 6806 18152 6850
rect 17252 6734 18152 6806
rect 25238 7535 26138 7607
rect 25238 7491 25310 7535
rect 25238 6851 25251 7491
rect 25297 6851 25310 7491
rect 26066 7491 26138 7535
rect 25238 6807 25310 6851
rect 26066 6851 26079 7491
rect 26125 6851 26138 7491
rect 26066 6807 26138 6851
rect 25238 6735 26138 6807
rect 26724 7535 27624 7607
rect 26724 7491 26796 7535
rect 26724 6851 26737 7491
rect 26783 6851 26796 7491
rect 27552 7491 27624 7535
rect 26724 6807 26796 6851
rect 27552 6851 27565 7491
rect 27611 6851 27624 7491
rect 27552 6807 27624 6851
rect 26724 6735 27624 6807
rect 34710 7535 35610 7607
rect 34710 7491 34782 7535
rect 34710 6851 34723 7491
rect 34769 6851 34782 7491
rect 35538 7491 35610 7535
rect 34710 6807 34782 6851
rect 35538 6851 35551 7491
rect 35597 6851 35610 7491
rect 35538 6807 35610 6851
rect 34710 6735 35610 6807
rect 36196 7535 37096 7607
rect 36196 7491 36268 7535
rect 36196 6851 36209 7491
rect 36255 6851 36268 7491
rect 37024 7491 37096 7535
rect 36196 6807 36268 6851
rect 37024 6851 37037 7491
rect 37083 6851 37096 7491
rect 37024 6807 37096 6851
rect 36196 6735 37096 6807
rect 44182 7535 45082 7607
rect 44182 7491 44254 7535
rect 44182 6851 44195 7491
rect 44241 6851 44254 7491
rect 45010 7491 45082 7535
rect 44182 6807 44254 6851
rect 45010 6851 45023 7491
rect 45069 6851 45082 7491
rect 45010 6807 45082 6851
rect 44182 6735 45082 6807
rect 45668 7535 46568 7607
rect 45668 7491 45740 7535
rect 45668 6851 45681 7491
rect 45727 6851 45740 7491
rect 46496 7491 46568 7535
rect 45668 6807 45740 6851
rect 46496 6851 46509 7491
rect 46555 6851 46568 7491
rect 46496 6807 46568 6851
rect 45668 6735 46568 6807
rect 53654 7535 54554 7607
rect 53654 7491 53726 7535
rect 53654 6851 53667 7491
rect 53713 6851 53726 7491
rect 54482 7491 54554 7535
rect 53654 6807 53726 6851
rect 54482 6851 54495 7491
rect 54541 6851 54554 7491
rect 54482 6807 54554 6851
rect 53654 6735 54554 6807
rect 55140 7535 56040 7607
rect 55140 7491 55212 7535
rect 55140 6851 55153 7491
rect 55199 6851 55212 7491
rect 55968 7491 56040 7535
rect 55140 6807 55212 6851
rect 55968 6851 55981 7491
rect 56027 6851 56040 7491
rect 55968 6807 56040 6851
rect 55140 6735 56040 6807
rect 6294 5329 7194 5401
rect 6294 5285 6366 5329
rect 6294 4645 6307 5285
rect 6353 4645 6366 5285
rect 7122 5285 7194 5329
rect 6294 4601 6366 4645
rect 7122 4645 7135 5285
rect 7181 4645 7194 5285
rect 7122 4601 7194 4645
rect 6294 4529 7194 4601
rect 7780 5330 8680 5402
rect 7780 5286 7852 5330
rect 7780 4646 7793 5286
rect 7839 4646 7852 5286
rect 8608 5286 8680 5330
rect 7780 4602 7852 4646
rect 8608 4646 8621 5286
rect 8667 4646 8680 5286
rect 8608 4602 8680 4646
rect 7780 4530 8680 4602
rect 15766 5329 16666 5401
rect 15766 5285 15838 5329
rect 15766 4645 15779 5285
rect 15825 4645 15838 5285
rect 16594 5285 16666 5329
rect 15766 4601 15838 4645
rect 16594 4645 16607 5285
rect 16653 4645 16666 5285
rect 16594 4601 16666 4645
rect 15766 4529 16666 4601
rect 17252 5330 18152 5402
rect 17252 5286 17324 5330
rect 17252 4646 17265 5286
rect 17311 4646 17324 5286
rect 18080 5286 18152 5330
rect 17252 4602 17324 4646
rect 18080 4646 18093 5286
rect 18139 4646 18152 5286
rect 18080 4602 18152 4646
rect 17252 4530 18152 4602
rect 25238 5330 26138 5402
rect 25238 5286 25310 5330
rect 25238 4646 25251 5286
rect 25297 4646 25310 5286
rect 26066 5286 26138 5330
rect 25238 4602 25310 4646
rect 26066 4646 26079 5286
rect 26125 4646 26138 5286
rect 26066 4602 26138 4646
rect 25238 4530 26138 4602
rect 26724 5331 27624 5403
rect 26724 5287 26796 5331
rect 26724 4647 26737 5287
rect 26783 4647 26796 5287
rect 27552 5287 27624 5331
rect 26724 4603 26796 4647
rect 27552 4647 27565 5287
rect 27611 4647 27624 5287
rect 27552 4603 27624 4647
rect 26724 4531 27624 4603
rect 34710 5330 35610 5402
rect 34710 5286 34782 5330
rect 34710 4646 34723 5286
rect 34769 4646 34782 5286
rect 35538 5286 35610 5330
rect 34710 4602 34782 4646
rect 35538 4646 35551 5286
rect 35597 4646 35610 5286
rect 35538 4602 35610 4646
rect 34710 4530 35610 4602
rect 36196 5331 37096 5403
rect 36196 5287 36268 5331
rect 36196 4647 36209 5287
rect 36255 4647 36268 5287
rect 37024 5287 37096 5331
rect 36196 4603 36268 4647
rect 37024 4647 37037 5287
rect 37083 4647 37096 5287
rect 37024 4603 37096 4647
rect 36196 4531 37096 4603
rect 44182 5330 45082 5402
rect 44182 5286 44254 5330
rect 44182 4646 44195 5286
rect 44241 4646 44254 5286
rect 45010 5286 45082 5330
rect 44182 4602 44254 4646
rect 45010 4646 45023 5286
rect 45069 4646 45082 5286
rect 45010 4602 45082 4646
rect 44182 4530 45082 4602
rect 45668 5331 46568 5403
rect 45668 5287 45740 5331
rect 45668 4647 45681 5287
rect 45727 4647 45740 5287
rect 46496 5287 46568 5331
rect 45668 4603 45740 4647
rect 46496 4647 46509 5287
rect 46555 4647 46568 5287
rect 46496 4603 46568 4647
rect 45668 4531 46568 4603
rect 53654 5330 54554 5402
rect 53654 5286 53726 5330
rect 53654 4646 53667 5286
rect 53713 4646 53726 5286
rect 54482 5286 54554 5330
rect 53654 4602 53726 4646
rect 54482 4646 54495 5286
rect 54541 4646 54554 5286
rect 54482 4602 54554 4646
rect 53654 4530 54554 4602
rect 55140 5331 56040 5403
rect 55140 5287 55212 5331
rect 55140 4647 55153 5287
rect 55199 4647 55212 5287
rect 55968 5287 56040 5331
rect 55140 4603 55212 4647
rect 55968 4647 55981 5287
rect 56027 4647 56040 5287
rect 55968 4603 56040 4647
rect 55140 4531 56040 4603
rect 1152 4214 1704 4286
rect 1152 4170 1224 4214
rect 1152 3430 1165 4170
rect 1211 3430 1224 4170
rect 1632 4170 1704 4214
rect 1152 3386 1224 3430
rect 1632 3430 1645 4170
rect 1691 3430 1704 4170
rect 1632 3386 1704 3430
rect 1152 3314 1704 3386
rect 2040 4214 3072 4286
rect 2040 4170 2112 4214
rect 2040 3430 2053 4170
rect 2099 3430 2112 4170
rect 2520 4170 2592 4214
rect 2040 3386 2112 3430
rect 2520 3430 2533 4170
rect 2579 3430 2592 4170
rect 3000 4170 3072 4214
rect 2520 3386 2592 3430
rect 3000 3430 3013 4170
rect 3059 3430 3072 4170
rect 10624 4214 11176 4286
rect 10624 4170 10696 4214
rect 3000 3386 3072 3430
rect 2040 3314 3072 3386
rect 10624 3430 10637 4170
rect 10683 3430 10696 4170
rect 11104 4170 11176 4214
rect 10624 3386 10696 3430
rect 11104 3430 11117 4170
rect 11163 3430 11176 4170
rect 11104 3386 11176 3430
rect 10624 3314 11176 3386
rect 11512 4214 12544 4286
rect 11512 4170 11584 4214
rect 11512 3430 11525 4170
rect 11571 3430 11584 4170
rect 11992 4170 12064 4214
rect 11512 3386 11584 3430
rect 11992 3430 12005 4170
rect 12051 3430 12064 4170
rect 12472 4170 12544 4214
rect 11992 3386 12064 3430
rect 12472 3430 12485 4170
rect 12531 3430 12544 4170
rect 20096 4215 20648 4287
rect 20096 4171 20168 4215
rect 12472 3386 12544 3430
rect 11512 3314 12544 3386
rect 20096 3431 20109 4171
rect 20155 3431 20168 4171
rect 20576 4171 20648 4215
rect 20096 3387 20168 3431
rect 20576 3431 20589 4171
rect 20635 3431 20648 4171
rect 20576 3387 20648 3431
rect 20096 3315 20648 3387
rect 20984 4215 22016 4287
rect 20984 4171 21056 4215
rect 20984 3431 20997 4171
rect 21043 3431 21056 4171
rect 21464 4171 21536 4215
rect 20984 3387 21056 3431
rect 21464 3431 21477 4171
rect 21523 3431 21536 4171
rect 21944 4171 22016 4215
rect 21464 3387 21536 3431
rect 21944 3431 21957 4171
rect 22003 3431 22016 4171
rect 29568 4215 30120 4287
rect 29568 4171 29640 4215
rect 21944 3387 22016 3431
rect 20984 3315 22016 3387
rect 29568 3431 29581 4171
rect 29627 3431 29640 4171
rect 30048 4171 30120 4215
rect 29568 3387 29640 3431
rect 30048 3431 30061 4171
rect 30107 3431 30120 4171
rect 30048 3387 30120 3431
rect 29568 3315 30120 3387
rect 30456 4215 31488 4287
rect 30456 4171 30528 4215
rect 30456 3431 30469 4171
rect 30515 3431 30528 4171
rect 30936 4171 31008 4215
rect 30456 3387 30528 3431
rect 30936 3431 30949 4171
rect 30995 3431 31008 4171
rect 31416 4171 31488 4215
rect 30936 3387 31008 3431
rect 31416 3431 31429 4171
rect 31475 3431 31488 4171
rect 39040 4215 39592 4287
rect 39040 4171 39112 4215
rect 31416 3387 31488 3431
rect 30456 3315 31488 3387
rect 39040 3431 39053 4171
rect 39099 3431 39112 4171
rect 39520 4171 39592 4215
rect 39040 3387 39112 3431
rect 39520 3431 39533 4171
rect 39579 3431 39592 4171
rect 39520 3387 39592 3431
rect 39040 3315 39592 3387
rect 39928 4215 40960 4287
rect 39928 4171 40000 4215
rect 39928 3431 39941 4171
rect 39987 3431 40000 4171
rect 40408 4171 40480 4215
rect 39928 3387 40000 3431
rect 40408 3431 40421 4171
rect 40467 3431 40480 4171
rect 40888 4171 40960 4215
rect 40408 3387 40480 3431
rect 40888 3431 40901 4171
rect 40947 3431 40960 4171
rect 48512 4215 49064 4287
rect 48512 4171 48584 4215
rect 40888 3387 40960 3431
rect 39928 3315 40960 3387
rect 48512 3431 48525 4171
rect 48571 3431 48584 4171
rect 48992 4171 49064 4215
rect 48512 3387 48584 3431
rect 48992 3431 49005 4171
rect 49051 3431 49064 4171
rect 48992 3387 49064 3431
rect 48512 3315 49064 3387
rect 49400 4215 50432 4287
rect 49400 4171 49472 4215
rect 49400 3431 49413 4171
rect 49459 3431 49472 4171
rect 49880 4171 49952 4215
rect 49400 3387 49472 3431
rect 49880 3431 49893 4171
rect 49939 3431 49952 4171
rect 50360 4171 50432 4215
rect 49880 3387 49952 3431
rect 50360 3431 50373 4171
rect 50419 3431 50432 4171
rect 50360 3387 50432 3431
rect 49400 3315 50432 3387
rect 6294 3124 7194 3196
rect 258 2794 810 2866
rect 258 2750 330 2794
rect 258 2010 271 2750
rect 317 2010 330 2750
rect 738 2750 810 2794
rect 258 1966 330 2010
rect 738 2010 751 2750
rect 797 2010 810 2750
rect 3380 3038 5300 3110
rect 3380 2994 3452 3038
rect 3380 2254 3393 2994
rect 3439 2254 3452 2994
rect 4064 2994 4136 3038
rect 3380 2210 3452 2254
rect 4064 2254 4077 2994
rect 4123 2254 4136 2994
rect 4748 2994 4820 3038
rect 4064 2210 4136 2254
rect 4748 2254 4761 2994
rect 4807 2254 4820 2994
rect 5228 2994 5300 3038
rect 4748 2210 4820 2254
rect 5228 2254 5241 2994
rect 5287 2254 5300 2994
rect 6294 3080 6366 3124
rect 6294 2440 6307 3080
rect 6353 2440 6366 3080
rect 7122 3080 7194 3124
rect 6294 2396 6366 2440
rect 7122 2440 7135 3080
rect 7181 2440 7194 3080
rect 15766 3124 16666 3196
rect 7122 2396 7194 2440
rect 6294 2324 7194 2396
rect 9730 2794 10282 2866
rect 9730 2750 9802 2794
rect 5228 2210 5300 2254
rect 3380 2138 5300 2210
rect 738 1966 810 2010
rect 258 1894 810 1966
rect 1152 1874 1704 1946
rect 1152 1830 1224 1874
rect 1152 1090 1165 1830
rect 1211 1090 1224 1830
rect 1632 1830 1704 1874
rect 1152 1046 1224 1090
rect 1632 1090 1645 1830
rect 1691 1090 1704 1830
rect 1632 1046 1704 1090
rect 1152 974 1704 1046
rect 2040 1874 3072 1946
rect 2040 1830 2112 1874
rect 2040 1090 2053 1830
rect 2099 1090 2112 1830
rect 2520 1830 2592 1874
rect 2040 1046 2112 1090
rect 2520 1090 2533 1830
rect 2579 1090 2592 1830
rect 3000 1830 3072 1874
rect 2520 1046 2592 1090
rect 3000 1090 3013 1830
rect 3059 1090 3072 1830
rect 9730 2010 9743 2750
rect 9789 2010 9802 2750
rect 10210 2750 10282 2794
rect 9730 1966 9802 2010
rect 10210 2010 10223 2750
rect 10269 2010 10282 2750
rect 12852 3038 14772 3110
rect 12852 2994 12924 3038
rect 12852 2254 12865 2994
rect 12911 2254 12924 2994
rect 13536 2994 13608 3038
rect 12852 2210 12924 2254
rect 13536 2254 13549 2994
rect 13595 2254 13608 2994
rect 14220 2994 14292 3038
rect 13536 2210 13608 2254
rect 14220 2254 14233 2994
rect 14279 2254 14292 2994
rect 14700 2994 14772 3038
rect 14220 2210 14292 2254
rect 14700 2254 14713 2994
rect 14759 2254 14772 2994
rect 15766 3080 15838 3124
rect 15766 2440 15779 3080
rect 15825 2440 15838 3080
rect 16594 3080 16666 3124
rect 15766 2396 15838 2440
rect 16594 2440 16607 3080
rect 16653 2440 16666 3080
rect 25238 3125 26138 3197
rect 16594 2396 16666 2440
rect 15766 2324 16666 2396
rect 19202 2795 19754 2867
rect 19202 2751 19274 2795
rect 14700 2210 14772 2254
rect 12852 2138 14772 2210
rect 10210 1966 10282 2010
rect 9730 1894 10282 1966
rect 10624 1874 11176 1946
rect 10624 1830 10696 1874
rect 3000 1046 3072 1090
rect 2040 974 3072 1046
rect 10624 1090 10637 1830
rect 10683 1090 10696 1830
rect 11104 1830 11176 1874
rect 10624 1046 10696 1090
rect 11104 1090 11117 1830
rect 11163 1090 11176 1830
rect 11104 1046 11176 1090
rect 10624 974 11176 1046
rect 11512 1874 12544 1946
rect 11512 1830 11584 1874
rect 11512 1090 11525 1830
rect 11571 1090 11584 1830
rect 11992 1830 12064 1874
rect 11512 1046 11584 1090
rect 11992 1090 12005 1830
rect 12051 1090 12064 1830
rect 12472 1830 12544 1874
rect 11992 1046 12064 1090
rect 12472 1090 12485 1830
rect 12531 1090 12544 1830
rect 19202 2011 19215 2751
rect 19261 2011 19274 2751
rect 19682 2751 19754 2795
rect 19202 1967 19274 2011
rect 19682 2011 19695 2751
rect 19741 2011 19754 2751
rect 22324 3039 24244 3111
rect 22324 2995 22396 3039
rect 22324 2255 22337 2995
rect 22383 2255 22396 2995
rect 23008 2995 23080 3039
rect 22324 2211 22396 2255
rect 23008 2255 23021 2995
rect 23067 2255 23080 2995
rect 23692 2995 23764 3039
rect 23008 2211 23080 2255
rect 23692 2255 23705 2995
rect 23751 2255 23764 2995
rect 24172 2995 24244 3039
rect 23692 2211 23764 2255
rect 24172 2255 24185 2995
rect 24231 2255 24244 2995
rect 25238 3081 25310 3125
rect 25238 2441 25251 3081
rect 25297 2441 25310 3081
rect 26066 3081 26138 3125
rect 25238 2397 25310 2441
rect 26066 2441 26079 3081
rect 26125 2441 26138 3081
rect 34710 3125 35610 3197
rect 26066 2397 26138 2441
rect 25238 2325 26138 2397
rect 28674 2795 29226 2867
rect 28674 2751 28746 2795
rect 24172 2211 24244 2255
rect 22324 2139 24244 2211
rect 19682 1967 19754 2011
rect 19202 1895 19754 1967
rect 20096 1875 20648 1947
rect 20096 1831 20168 1875
rect 12472 1046 12544 1090
rect 11512 974 12544 1046
rect 20096 1091 20109 1831
rect 20155 1091 20168 1831
rect 20576 1831 20648 1875
rect 20096 1047 20168 1091
rect 20576 1091 20589 1831
rect 20635 1091 20648 1831
rect 20576 1047 20648 1091
rect 20096 975 20648 1047
rect 20984 1875 22016 1947
rect 20984 1831 21056 1875
rect 20984 1091 20997 1831
rect 21043 1091 21056 1831
rect 21464 1831 21536 1875
rect 20984 1047 21056 1091
rect 21464 1091 21477 1831
rect 21523 1091 21536 1831
rect 21944 1831 22016 1875
rect 21464 1047 21536 1091
rect 21944 1091 21957 1831
rect 22003 1091 22016 1831
rect 28674 2011 28687 2751
rect 28733 2011 28746 2751
rect 29154 2751 29226 2795
rect 28674 1967 28746 2011
rect 29154 2011 29167 2751
rect 29213 2011 29226 2751
rect 31796 3039 33716 3111
rect 31796 2995 31868 3039
rect 31796 2255 31809 2995
rect 31855 2255 31868 2995
rect 32480 2995 32552 3039
rect 31796 2211 31868 2255
rect 32480 2255 32493 2995
rect 32539 2255 32552 2995
rect 33164 2995 33236 3039
rect 32480 2211 32552 2255
rect 33164 2255 33177 2995
rect 33223 2255 33236 2995
rect 33644 2995 33716 3039
rect 33164 2211 33236 2255
rect 33644 2255 33657 2995
rect 33703 2255 33716 2995
rect 34710 3081 34782 3125
rect 34710 2441 34723 3081
rect 34769 2441 34782 3081
rect 35538 3081 35610 3125
rect 34710 2397 34782 2441
rect 35538 2441 35551 3081
rect 35597 2441 35610 3081
rect 44182 3125 45082 3197
rect 35538 2397 35610 2441
rect 34710 2325 35610 2397
rect 38146 2795 38698 2867
rect 38146 2751 38218 2795
rect 33644 2211 33716 2255
rect 31796 2139 33716 2211
rect 29154 1967 29226 2011
rect 28674 1895 29226 1967
rect 29568 1875 30120 1947
rect 29568 1831 29640 1875
rect 21944 1047 22016 1091
rect 20984 975 22016 1047
rect 29568 1091 29581 1831
rect 29627 1091 29640 1831
rect 30048 1831 30120 1875
rect 29568 1047 29640 1091
rect 30048 1091 30061 1831
rect 30107 1091 30120 1831
rect 30048 1047 30120 1091
rect 29568 975 30120 1047
rect 30456 1875 31488 1947
rect 30456 1831 30528 1875
rect 30456 1091 30469 1831
rect 30515 1091 30528 1831
rect 30936 1831 31008 1875
rect 30456 1047 30528 1091
rect 30936 1091 30949 1831
rect 30995 1091 31008 1831
rect 31416 1831 31488 1875
rect 30936 1047 31008 1091
rect 31416 1091 31429 1831
rect 31475 1091 31488 1831
rect 38146 2011 38159 2751
rect 38205 2011 38218 2751
rect 38626 2751 38698 2795
rect 38146 1967 38218 2011
rect 38626 2011 38639 2751
rect 38685 2011 38698 2751
rect 41268 3039 43188 3111
rect 41268 2995 41340 3039
rect 41268 2255 41281 2995
rect 41327 2255 41340 2995
rect 41952 2995 42024 3039
rect 41268 2211 41340 2255
rect 41952 2255 41965 2995
rect 42011 2255 42024 2995
rect 42636 2995 42708 3039
rect 41952 2211 42024 2255
rect 42636 2255 42649 2995
rect 42695 2255 42708 2995
rect 43116 2995 43188 3039
rect 42636 2211 42708 2255
rect 43116 2255 43129 2995
rect 43175 2255 43188 2995
rect 44182 3081 44254 3125
rect 44182 2441 44195 3081
rect 44241 2441 44254 3081
rect 45010 3081 45082 3125
rect 44182 2397 44254 2441
rect 45010 2441 45023 3081
rect 45069 2441 45082 3081
rect 53654 3125 54554 3197
rect 45010 2397 45082 2441
rect 44182 2325 45082 2397
rect 47618 2795 48170 2867
rect 47618 2751 47690 2795
rect 43116 2211 43188 2255
rect 41268 2139 43188 2211
rect 38626 1967 38698 2011
rect 38146 1895 38698 1967
rect 39040 1875 39592 1947
rect 39040 1831 39112 1875
rect 31416 1047 31488 1091
rect 30456 975 31488 1047
rect 39040 1091 39053 1831
rect 39099 1091 39112 1831
rect 39520 1831 39592 1875
rect 39040 1047 39112 1091
rect 39520 1091 39533 1831
rect 39579 1091 39592 1831
rect 39520 1047 39592 1091
rect 39040 975 39592 1047
rect 39928 1875 40960 1947
rect 39928 1831 40000 1875
rect 39928 1091 39941 1831
rect 39987 1091 40000 1831
rect 40408 1831 40480 1875
rect 39928 1047 40000 1091
rect 40408 1091 40421 1831
rect 40467 1091 40480 1831
rect 40888 1831 40960 1875
rect 40408 1047 40480 1091
rect 40888 1091 40901 1831
rect 40947 1091 40960 1831
rect 47618 2011 47631 2751
rect 47677 2011 47690 2751
rect 48098 2751 48170 2795
rect 47618 1967 47690 2011
rect 48098 2011 48111 2751
rect 48157 2011 48170 2751
rect 50740 3039 52660 3111
rect 50740 2995 50812 3039
rect 50740 2255 50753 2995
rect 50799 2255 50812 2995
rect 51424 2995 51496 3039
rect 50740 2211 50812 2255
rect 51424 2255 51437 2995
rect 51483 2255 51496 2995
rect 52108 2995 52180 3039
rect 51424 2211 51496 2255
rect 52108 2255 52121 2995
rect 52167 2255 52180 2995
rect 52588 2995 52660 3039
rect 52108 2211 52180 2255
rect 52588 2255 52601 2995
rect 52647 2255 52660 2995
rect 53654 3081 53726 3125
rect 53654 2441 53667 3081
rect 53713 2441 53726 3081
rect 54482 3081 54554 3125
rect 53654 2397 53726 2441
rect 54482 2441 54495 3081
rect 54541 2441 54554 3081
rect 54482 2397 54554 2441
rect 53654 2325 54554 2397
rect 52588 2211 52660 2255
rect 50740 2139 52660 2211
rect 48098 1967 48170 2011
rect 47618 1895 48170 1967
rect 48512 1875 49064 1947
rect 48512 1831 48584 1875
rect 40888 1047 40960 1091
rect 39928 975 40960 1047
rect 48512 1091 48525 1831
rect 48571 1091 48584 1831
rect 48992 1831 49064 1875
rect 48512 1047 48584 1091
rect 48992 1091 49005 1831
rect 49051 1091 49064 1831
rect 48992 1047 49064 1091
rect 48512 975 49064 1047
rect 49400 1875 50432 1947
rect 49400 1831 49472 1875
rect 49400 1091 49413 1831
rect 49459 1091 49472 1831
rect 49880 1831 49952 1875
rect 49400 1047 49472 1091
rect 49880 1091 49893 1831
rect 49939 1091 49952 1831
rect 50360 1831 50432 1875
rect 49880 1047 49952 1091
rect 50360 1091 50373 1831
rect 50419 1091 50432 1831
rect 50360 1047 50432 1091
rect 49400 975 50432 1047
<< psubdiffcont >>
rect 6307 8195 6353 8535
rect 7135 8195 7181 8535
rect 15779 8195 15825 8535
rect 16607 8195 16653 8535
rect 25251 8196 25297 8536
rect 26079 8196 26125 8536
rect 34723 8196 34769 8536
rect 35551 8196 35597 8536
rect 44195 8196 44241 8536
rect 45023 8196 45069 8536
rect 53667 8196 53713 8536
rect 54495 8196 54541 8536
rect 6307 5990 6353 6330
rect 7135 5990 7181 6330
rect 7793 5990 7839 6330
rect 8621 5990 8667 6330
rect 15779 5990 15825 6330
rect 16607 5990 16653 6330
rect 17265 5990 17311 6330
rect 18093 5990 18139 6330
rect 25251 5991 25297 6331
rect 26079 5991 26125 6331
rect 26737 5991 26783 6331
rect 27565 5991 27611 6331
rect 34723 5991 34769 6331
rect 35551 5991 35597 6331
rect 36209 5991 36255 6331
rect 37037 5991 37083 6331
rect 44195 5991 44241 6331
rect 45023 5991 45069 6331
rect 45681 5991 45727 6331
rect 46509 5991 46555 6331
rect 53667 5991 53713 6331
rect 54495 5991 54541 6331
rect 55153 5991 55199 6331
rect 55981 5991 56027 6331
rect 6307 3785 6353 4125
rect 7135 3785 7181 4125
rect 7793 3786 7839 4126
rect 8621 3786 8667 4126
rect 15779 3785 15825 4125
rect 16607 3785 16653 4125
rect 17265 3786 17311 4126
rect 18093 3786 18139 4126
rect 25251 3786 25297 4126
rect 26079 3786 26125 4126
rect 26737 3787 26783 4127
rect 27565 3787 27611 4127
rect 34723 3786 34769 4126
rect 35551 3786 35597 4126
rect 36209 3787 36255 4127
rect 37037 3787 37083 4127
rect 44195 3786 44241 4126
rect 45023 3786 45069 4126
rect 45681 3787 45727 4127
rect 46509 3787 46555 4127
rect 53667 3786 53713 4126
rect 54495 3786 54541 4126
rect 55153 3787 55199 4127
rect 55981 3787 56027 4127
rect 1165 2710 1211 3050
rect 1849 2710 1895 3050
rect 2533 2710 2579 3050
rect 3013 2710 3059 3050
rect 271 1290 317 1630
rect 751 1290 797 1630
rect 3393 1534 3439 1874
rect 3873 1534 3919 1874
rect 4077 1534 4123 1874
rect 4557 1534 4603 1874
rect 4761 1534 4807 1874
rect 5241 1534 5287 1874
rect 6307 1580 6353 1920
rect 7135 1580 7181 1920
rect 10637 2710 10683 3050
rect 11321 2710 11367 3050
rect 12005 2710 12051 3050
rect 12485 2710 12531 3050
rect 9743 1290 9789 1630
rect 10223 1290 10269 1630
rect 12865 1534 12911 1874
rect 13345 1534 13391 1874
rect 13549 1534 13595 1874
rect 14029 1534 14075 1874
rect 14233 1534 14279 1874
rect 14713 1534 14759 1874
rect 15779 1580 15825 1920
rect 16607 1580 16653 1920
rect 20109 2711 20155 3051
rect 20793 2711 20839 3051
rect 21477 2711 21523 3051
rect 21957 2711 22003 3051
rect 19215 1291 19261 1631
rect 19695 1291 19741 1631
rect 22337 1535 22383 1875
rect 22817 1535 22863 1875
rect 23021 1535 23067 1875
rect 23501 1535 23547 1875
rect 23705 1535 23751 1875
rect 24185 1535 24231 1875
rect 25251 1581 25297 1921
rect 26079 1581 26125 1921
rect 29581 2711 29627 3051
rect 30265 2711 30311 3051
rect 30949 2711 30995 3051
rect 31429 2711 31475 3051
rect 28687 1291 28733 1631
rect 29167 1291 29213 1631
rect 31809 1535 31855 1875
rect 32289 1535 32335 1875
rect 32493 1535 32539 1875
rect 32973 1535 33019 1875
rect 33177 1535 33223 1875
rect 33657 1535 33703 1875
rect 34723 1581 34769 1921
rect 35551 1581 35597 1921
rect 39053 2711 39099 3051
rect 39737 2711 39783 3051
rect 40421 2711 40467 3051
rect 40901 2711 40947 3051
rect 38159 1291 38205 1631
rect 38639 1291 38685 1631
rect 41281 1535 41327 1875
rect 41761 1535 41807 1875
rect 41965 1535 42011 1875
rect 42445 1535 42491 1875
rect 42649 1535 42695 1875
rect 43129 1535 43175 1875
rect 44195 1581 44241 1921
rect 45023 1581 45069 1921
rect 48525 2711 48571 3051
rect 49209 2711 49255 3051
rect 49893 2711 49939 3051
rect 50373 2711 50419 3051
rect 47631 1291 47677 1631
rect 48111 1291 48157 1631
rect 50753 1535 50799 1875
rect 51233 1535 51279 1875
rect 51437 1535 51483 1875
rect 51917 1535 51963 1875
rect 52121 1535 52167 1875
rect 52601 1535 52647 1875
rect 53667 1581 53713 1921
rect 54495 1581 54541 1921
rect 1165 370 1211 710
rect 1849 370 1895 710
rect 2533 370 2579 710
rect 3013 370 3059 710
rect 10637 370 10683 710
rect 11321 370 11367 710
rect 12005 370 12051 710
rect 12485 370 12531 710
rect 20109 371 20155 711
rect 20793 371 20839 711
rect 21477 371 21523 711
rect 21957 371 22003 711
rect 29581 371 29627 711
rect 30265 371 30311 711
rect 30949 371 30995 711
rect 31429 371 31475 711
rect 39053 371 39099 711
rect 39737 371 39783 711
rect 40421 371 40467 711
rect 40901 371 40947 711
rect 48525 371 48571 711
rect 49209 371 49255 711
rect 49893 371 49939 711
rect 50373 371 50419 711
<< nsubdiffcont >>
rect 6307 9055 6353 9695
rect 7135 9055 7181 9695
rect 15779 9055 15825 9695
rect 16607 9055 16653 9695
rect 25251 9056 25297 9696
rect 26079 9056 26125 9696
rect 34723 9056 34769 9696
rect 35551 9056 35597 9696
rect 44195 9056 44241 9696
rect 45023 9056 45069 9696
rect 53667 9056 53713 9696
rect 54495 9056 54541 9696
rect 6307 6850 6353 7490
rect 7135 6850 7181 7490
rect 7793 6850 7839 7490
rect 8621 6850 8667 7490
rect 15779 6850 15825 7490
rect 16607 6850 16653 7490
rect 17265 6850 17311 7490
rect 18093 6850 18139 7490
rect 25251 6851 25297 7491
rect 26079 6851 26125 7491
rect 26737 6851 26783 7491
rect 27565 6851 27611 7491
rect 34723 6851 34769 7491
rect 35551 6851 35597 7491
rect 36209 6851 36255 7491
rect 37037 6851 37083 7491
rect 44195 6851 44241 7491
rect 45023 6851 45069 7491
rect 45681 6851 45727 7491
rect 46509 6851 46555 7491
rect 53667 6851 53713 7491
rect 54495 6851 54541 7491
rect 55153 6851 55199 7491
rect 55981 6851 56027 7491
rect 6307 4645 6353 5285
rect 7135 4645 7181 5285
rect 7793 4646 7839 5286
rect 8621 4646 8667 5286
rect 15779 4645 15825 5285
rect 16607 4645 16653 5285
rect 17265 4646 17311 5286
rect 18093 4646 18139 5286
rect 25251 4646 25297 5286
rect 26079 4646 26125 5286
rect 26737 4647 26783 5287
rect 27565 4647 27611 5287
rect 34723 4646 34769 5286
rect 35551 4646 35597 5286
rect 36209 4647 36255 5287
rect 37037 4647 37083 5287
rect 44195 4646 44241 5286
rect 45023 4646 45069 5286
rect 45681 4647 45727 5287
rect 46509 4647 46555 5287
rect 53667 4646 53713 5286
rect 54495 4646 54541 5286
rect 55153 4647 55199 5287
rect 55981 4647 56027 5287
rect 1165 3430 1211 4170
rect 1645 3430 1691 4170
rect 2053 3430 2099 4170
rect 2533 3430 2579 4170
rect 3013 3430 3059 4170
rect 10637 3430 10683 4170
rect 11117 3430 11163 4170
rect 11525 3430 11571 4170
rect 12005 3430 12051 4170
rect 12485 3430 12531 4170
rect 20109 3431 20155 4171
rect 20589 3431 20635 4171
rect 20997 3431 21043 4171
rect 21477 3431 21523 4171
rect 21957 3431 22003 4171
rect 29581 3431 29627 4171
rect 30061 3431 30107 4171
rect 30469 3431 30515 4171
rect 30949 3431 30995 4171
rect 31429 3431 31475 4171
rect 39053 3431 39099 4171
rect 39533 3431 39579 4171
rect 39941 3431 39987 4171
rect 40421 3431 40467 4171
rect 40901 3431 40947 4171
rect 48525 3431 48571 4171
rect 49005 3431 49051 4171
rect 49413 3431 49459 4171
rect 49893 3431 49939 4171
rect 50373 3431 50419 4171
rect 271 2010 317 2750
rect 751 2010 797 2750
rect 3393 2254 3439 2994
rect 4077 2254 4123 2994
rect 4761 2254 4807 2994
rect 5241 2254 5287 2994
rect 6307 2440 6353 3080
rect 7135 2440 7181 3080
rect 1165 1090 1211 1830
rect 1645 1090 1691 1830
rect 2053 1090 2099 1830
rect 2533 1090 2579 1830
rect 3013 1090 3059 1830
rect 9743 2010 9789 2750
rect 10223 2010 10269 2750
rect 12865 2254 12911 2994
rect 13549 2254 13595 2994
rect 14233 2254 14279 2994
rect 14713 2254 14759 2994
rect 15779 2440 15825 3080
rect 16607 2440 16653 3080
rect 10637 1090 10683 1830
rect 11117 1090 11163 1830
rect 11525 1090 11571 1830
rect 12005 1090 12051 1830
rect 12485 1090 12531 1830
rect 19215 2011 19261 2751
rect 19695 2011 19741 2751
rect 22337 2255 22383 2995
rect 23021 2255 23067 2995
rect 23705 2255 23751 2995
rect 24185 2255 24231 2995
rect 25251 2441 25297 3081
rect 26079 2441 26125 3081
rect 20109 1091 20155 1831
rect 20589 1091 20635 1831
rect 20997 1091 21043 1831
rect 21477 1091 21523 1831
rect 21957 1091 22003 1831
rect 28687 2011 28733 2751
rect 29167 2011 29213 2751
rect 31809 2255 31855 2995
rect 32493 2255 32539 2995
rect 33177 2255 33223 2995
rect 33657 2255 33703 2995
rect 34723 2441 34769 3081
rect 35551 2441 35597 3081
rect 29581 1091 29627 1831
rect 30061 1091 30107 1831
rect 30469 1091 30515 1831
rect 30949 1091 30995 1831
rect 31429 1091 31475 1831
rect 38159 2011 38205 2751
rect 38639 2011 38685 2751
rect 41281 2255 41327 2995
rect 41965 2255 42011 2995
rect 42649 2255 42695 2995
rect 43129 2255 43175 2995
rect 44195 2441 44241 3081
rect 45023 2441 45069 3081
rect 39053 1091 39099 1831
rect 39533 1091 39579 1831
rect 39941 1091 39987 1831
rect 40421 1091 40467 1831
rect 40901 1091 40947 1831
rect 47631 2011 47677 2751
rect 48111 2011 48157 2751
rect 50753 2255 50799 2995
rect 51437 2255 51483 2995
rect 52121 2255 52167 2995
rect 52601 2255 52647 2995
rect 53667 2441 53713 3081
rect 54495 2441 54541 3081
rect 48525 1091 48571 1831
rect 49005 1091 49051 1831
rect 49413 1091 49459 1831
rect 49893 1091 49939 1831
rect 50373 1091 50419 1831
<< polysilicon >>
rect 6520 9704 6600 9717
rect 6520 9658 6533 9704
rect 6587 9658 6600 9704
rect 6520 9625 6600 9658
rect 6704 9704 6784 9717
rect 6704 9658 6717 9704
rect 6771 9658 6784 9704
rect 6704 9625 6784 9658
rect 6888 9704 6968 9717
rect 6888 9658 6901 9704
rect 6955 9658 6968 9704
rect 6888 9625 6968 9658
rect 6520 9092 6600 9125
rect 6520 9046 6533 9092
rect 6587 9046 6600 9092
rect 6520 9033 6600 9046
rect 6704 9092 6784 9125
rect 6704 9046 6717 9092
rect 6771 9046 6784 9092
rect 6704 9033 6784 9046
rect 6888 9092 6968 9125
rect 6888 9046 6901 9092
rect 6955 9046 6968 9092
rect 6888 9033 6968 9046
rect 15992 9704 16072 9717
rect 15992 9658 16005 9704
rect 16059 9658 16072 9704
rect 15992 9625 16072 9658
rect 16176 9704 16256 9717
rect 16176 9658 16189 9704
rect 16243 9658 16256 9704
rect 16176 9625 16256 9658
rect 16360 9704 16440 9717
rect 16360 9658 16373 9704
rect 16427 9658 16440 9704
rect 16360 9625 16440 9658
rect 15992 9092 16072 9125
rect 15992 9046 16005 9092
rect 16059 9046 16072 9092
rect 15992 9033 16072 9046
rect 16176 9092 16256 9125
rect 16176 9046 16189 9092
rect 16243 9046 16256 9092
rect 16176 9033 16256 9046
rect 16360 9092 16440 9125
rect 16360 9046 16373 9092
rect 16427 9046 16440 9092
rect 16360 9033 16440 9046
rect 25464 9705 25544 9718
rect 25464 9659 25477 9705
rect 25531 9659 25544 9705
rect 25464 9626 25544 9659
rect 25648 9705 25728 9718
rect 25648 9659 25661 9705
rect 25715 9659 25728 9705
rect 25648 9626 25728 9659
rect 25832 9705 25912 9718
rect 25832 9659 25845 9705
rect 25899 9659 25912 9705
rect 25832 9626 25912 9659
rect 25464 9093 25544 9126
rect 25464 9047 25477 9093
rect 25531 9047 25544 9093
rect 25464 9034 25544 9047
rect 25648 9093 25728 9126
rect 25648 9047 25661 9093
rect 25715 9047 25728 9093
rect 25648 9034 25728 9047
rect 25832 9093 25912 9126
rect 25832 9047 25845 9093
rect 25899 9047 25912 9093
rect 25832 9034 25912 9047
rect 34936 9705 35016 9718
rect 34936 9659 34949 9705
rect 35003 9659 35016 9705
rect 34936 9626 35016 9659
rect 35120 9705 35200 9718
rect 35120 9659 35133 9705
rect 35187 9659 35200 9705
rect 35120 9626 35200 9659
rect 35304 9705 35384 9718
rect 35304 9659 35317 9705
rect 35371 9659 35384 9705
rect 35304 9626 35384 9659
rect 34936 9093 35016 9126
rect 34936 9047 34949 9093
rect 35003 9047 35016 9093
rect 34936 9034 35016 9047
rect 35120 9093 35200 9126
rect 35120 9047 35133 9093
rect 35187 9047 35200 9093
rect 35120 9034 35200 9047
rect 35304 9093 35384 9126
rect 35304 9047 35317 9093
rect 35371 9047 35384 9093
rect 35304 9034 35384 9047
rect 44408 9705 44488 9718
rect 44408 9659 44421 9705
rect 44475 9659 44488 9705
rect 44408 9626 44488 9659
rect 44592 9705 44672 9718
rect 44592 9659 44605 9705
rect 44659 9659 44672 9705
rect 44592 9626 44672 9659
rect 44776 9705 44856 9718
rect 44776 9659 44789 9705
rect 44843 9659 44856 9705
rect 44776 9626 44856 9659
rect 44408 9093 44488 9126
rect 44408 9047 44421 9093
rect 44475 9047 44488 9093
rect 44408 9034 44488 9047
rect 44592 9093 44672 9126
rect 44592 9047 44605 9093
rect 44659 9047 44672 9093
rect 44592 9034 44672 9047
rect 44776 9093 44856 9126
rect 44776 9047 44789 9093
rect 44843 9047 44856 9093
rect 44776 9034 44856 9047
rect 53880 9705 53960 9718
rect 53880 9659 53893 9705
rect 53947 9659 53960 9705
rect 53880 9626 53960 9659
rect 54064 9705 54144 9718
rect 54064 9659 54077 9705
rect 54131 9659 54144 9705
rect 54064 9626 54144 9659
rect 54248 9705 54328 9718
rect 54248 9659 54261 9705
rect 54315 9659 54328 9705
rect 54248 9626 54328 9659
rect 53880 9093 53960 9126
rect 53880 9047 53893 9093
rect 53947 9047 53960 9093
rect 53880 9034 53960 9047
rect 54064 9093 54144 9126
rect 54064 9047 54077 9093
rect 54131 9047 54144 9093
rect 54064 9034 54144 9047
rect 54248 9093 54328 9126
rect 54248 9047 54261 9093
rect 54315 9047 54328 9093
rect 54248 9034 54328 9047
rect 6520 8544 6600 8557
rect 6520 8498 6533 8544
rect 6587 8498 6600 8544
rect 6520 8465 6600 8498
rect 6704 8544 6784 8557
rect 6704 8498 6717 8544
rect 6771 8498 6784 8544
rect 6704 8465 6784 8498
rect 6888 8544 6968 8557
rect 6888 8498 6901 8544
rect 6955 8498 6968 8544
rect 6888 8465 6968 8498
rect 6520 8232 6600 8265
rect 6520 8186 6533 8232
rect 6587 8186 6600 8232
rect 6520 8173 6600 8186
rect 6704 8232 6784 8265
rect 6704 8186 6717 8232
rect 6771 8186 6784 8232
rect 6704 8173 6784 8186
rect 6888 8232 6968 8265
rect 6888 8186 6901 8232
rect 6955 8186 6968 8232
rect 6888 8173 6968 8186
rect 15992 8544 16072 8557
rect 15992 8498 16005 8544
rect 16059 8498 16072 8544
rect 15992 8465 16072 8498
rect 16176 8544 16256 8557
rect 16176 8498 16189 8544
rect 16243 8498 16256 8544
rect 16176 8465 16256 8498
rect 16360 8544 16440 8557
rect 16360 8498 16373 8544
rect 16427 8498 16440 8544
rect 16360 8465 16440 8498
rect 15992 8232 16072 8265
rect 15992 8186 16005 8232
rect 16059 8186 16072 8232
rect 15992 8173 16072 8186
rect 16176 8232 16256 8265
rect 16176 8186 16189 8232
rect 16243 8186 16256 8232
rect 16176 8173 16256 8186
rect 16360 8232 16440 8265
rect 16360 8186 16373 8232
rect 16427 8186 16440 8232
rect 16360 8173 16440 8186
rect 25464 8545 25544 8558
rect 25464 8499 25477 8545
rect 25531 8499 25544 8545
rect 25464 8466 25544 8499
rect 25648 8545 25728 8558
rect 25648 8499 25661 8545
rect 25715 8499 25728 8545
rect 25648 8466 25728 8499
rect 25832 8545 25912 8558
rect 25832 8499 25845 8545
rect 25899 8499 25912 8545
rect 25832 8466 25912 8499
rect 25464 8233 25544 8266
rect 25464 8187 25477 8233
rect 25531 8187 25544 8233
rect 25464 8174 25544 8187
rect 25648 8233 25728 8266
rect 25648 8187 25661 8233
rect 25715 8187 25728 8233
rect 25648 8174 25728 8187
rect 25832 8233 25912 8266
rect 25832 8187 25845 8233
rect 25899 8187 25912 8233
rect 25832 8174 25912 8187
rect 34936 8545 35016 8558
rect 34936 8499 34949 8545
rect 35003 8499 35016 8545
rect 34936 8466 35016 8499
rect 35120 8545 35200 8558
rect 35120 8499 35133 8545
rect 35187 8499 35200 8545
rect 35120 8466 35200 8499
rect 35304 8545 35384 8558
rect 35304 8499 35317 8545
rect 35371 8499 35384 8545
rect 35304 8466 35384 8499
rect 34936 8233 35016 8266
rect 34936 8187 34949 8233
rect 35003 8187 35016 8233
rect 34936 8174 35016 8187
rect 35120 8233 35200 8266
rect 35120 8187 35133 8233
rect 35187 8187 35200 8233
rect 35120 8174 35200 8187
rect 35304 8233 35384 8266
rect 35304 8187 35317 8233
rect 35371 8187 35384 8233
rect 35304 8174 35384 8187
rect 44408 8545 44488 8558
rect 44408 8499 44421 8545
rect 44475 8499 44488 8545
rect 44408 8466 44488 8499
rect 44592 8545 44672 8558
rect 44592 8499 44605 8545
rect 44659 8499 44672 8545
rect 44592 8466 44672 8499
rect 44776 8545 44856 8558
rect 44776 8499 44789 8545
rect 44843 8499 44856 8545
rect 44776 8466 44856 8499
rect 44408 8233 44488 8266
rect 44408 8187 44421 8233
rect 44475 8187 44488 8233
rect 44408 8174 44488 8187
rect 44592 8233 44672 8266
rect 44592 8187 44605 8233
rect 44659 8187 44672 8233
rect 44592 8174 44672 8187
rect 44776 8233 44856 8266
rect 44776 8187 44789 8233
rect 44843 8187 44856 8233
rect 44776 8174 44856 8187
rect 53880 8545 53960 8558
rect 53880 8499 53893 8545
rect 53947 8499 53960 8545
rect 53880 8466 53960 8499
rect 54064 8545 54144 8558
rect 54064 8499 54077 8545
rect 54131 8499 54144 8545
rect 54064 8466 54144 8499
rect 54248 8545 54328 8558
rect 54248 8499 54261 8545
rect 54315 8499 54328 8545
rect 54248 8466 54328 8499
rect 53880 8233 53960 8266
rect 53880 8187 53893 8233
rect 53947 8187 53960 8233
rect 53880 8174 53960 8187
rect 54064 8233 54144 8266
rect 54064 8187 54077 8233
rect 54131 8187 54144 8233
rect 54064 8174 54144 8187
rect 54248 8233 54328 8266
rect 54248 8187 54261 8233
rect 54315 8187 54328 8233
rect 54248 8174 54328 8187
rect 6520 7499 6600 7512
rect 6520 7453 6533 7499
rect 6587 7453 6600 7499
rect 6520 7420 6600 7453
rect 6704 7499 6784 7512
rect 6704 7453 6717 7499
rect 6771 7453 6784 7499
rect 6704 7420 6784 7453
rect 6888 7499 6968 7512
rect 6888 7453 6901 7499
rect 6955 7453 6968 7499
rect 6888 7420 6968 7453
rect 6520 6887 6600 6920
rect 6520 6841 6533 6887
rect 6587 6841 6600 6887
rect 6520 6828 6600 6841
rect 6704 6887 6784 6920
rect 6704 6841 6717 6887
rect 6771 6841 6784 6887
rect 6704 6828 6784 6841
rect 6888 6887 6968 6920
rect 6888 6841 6901 6887
rect 6955 6841 6968 6887
rect 6888 6828 6968 6841
rect 8006 7499 8086 7512
rect 8006 7453 8019 7499
rect 8073 7453 8086 7499
rect 8006 7420 8086 7453
rect 8190 7499 8270 7512
rect 8190 7453 8203 7499
rect 8257 7453 8270 7499
rect 8190 7420 8270 7453
rect 8374 7499 8454 7512
rect 8374 7453 8387 7499
rect 8441 7453 8454 7499
rect 8374 7420 8454 7453
rect 8006 6887 8086 6920
rect 8006 6841 8019 6887
rect 8073 6841 8086 6887
rect 8006 6828 8086 6841
rect 8190 6887 8270 6920
rect 8190 6841 8203 6887
rect 8257 6841 8270 6887
rect 8190 6828 8270 6841
rect 8374 6887 8454 6920
rect 8374 6841 8387 6887
rect 8441 6841 8454 6887
rect 8374 6828 8454 6841
rect 15992 7499 16072 7512
rect 15992 7453 16005 7499
rect 16059 7453 16072 7499
rect 15992 7420 16072 7453
rect 16176 7499 16256 7512
rect 16176 7453 16189 7499
rect 16243 7453 16256 7499
rect 16176 7420 16256 7453
rect 16360 7499 16440 7512
rect 16360 7453 16373 7499
rect 16427 7453 16440 7499
rect 16360 7420 16440 7453
rect 15992 6887 16072 6920
rect 15992 6841 16005 6887
rect 16059 6841 16072 6887
rect 15992 6828 16072 6841
rect 16176 6887 16256 6920
rect 16176 6841 16189 6887
rect 16243 6841 16256 6887
rect 16176 6828 16256 6841
rect 16360 6887 16440 6920
rect 16360 6841 16373 6887
rect 16427 6841 16440 6887
rect 16360 6828 16440 6841
rect 17478 7499 17558 7512
rect 17478 7453 17491 7499
rect 17545 7453 17558 7499
rect 17478 7420 17558 7453
rect 17662 7499 17742 7512
rect 17662 7453 17675 7499
rect 17729 7453 17742 7499
rect 17662 7420 17742 7453
rect 17846 7499 17926 7512
rect 17846 7453 17859 7499
rect 17913 7453 17926 7499
rect 17846 7420 17926 7453
rect 17478 6887 17558 6920
rect 17478 6841 17491 6887
rect 17545 6841 17558 6887
rect 17478 6828 17558 6841
rect 17662 6887 17742 6920
rect 17662 6841 17675 6887
rect 17729 6841 17742 6887
rect 17662 6828 17742 6841
rect 17846 6887 17926 6920
rect 17846 6841 17859 6887
rect 17913 6841 17926 6887
rect 17846 6828 17926 6841
rect 25464 7500 25544 7513
rect 25464 7454 25477 7500
rect 25531 7454 25544 7500
rect 25464 7421 25544 7454
rect 25648 7500 25728 7513
rect 25648 7454 25661 7500
rect 25715 7454 25728 7500
rect 25648 7421 25728 7454
rect 25832 7500 25912 7513
rect 25832 7454 25845 7500
rect 25899 7454 25912 7500
rect 25832 7421 25912 7454
rect 25464 6888 25544 6921
rect 25464 6842 25477 6888
rect 25531 6842 25544 6888
rect 25464 6829 25544 6842
rect 25648 6888 25728 6921
rect 25648 6842 25661 6888
rect 25715 6842 25728 6888
rect 25648 6829 25728 6842
rect 25832 6888 25912 6921
rect 25832 6842 25845 6888
rect 25899 6842 25912 6888
rect 25832 6829 25912 6842
rect 26950 7500 27030 7513
rect 26950 7454 26963 7500
rect 27017 7454 27030 7500
rect 26950 7421 27030 7454
rect 27134 7500 27214 7513
rect 27134 7454 27147 7500
rect 27201 7454 27214 7500
rect 27134 7421 27214 7454
rect 27318 7500 27398 7513
rect 27318 7454 27331 7500
rect 27385 7454 27398 7500
rect 27318 7421 27398 7454
rect 26950 6888 27030 6921
rect 26950 6842 26963 6888
rect 27017 6842 27030 6888
rect 26950 6829 27030 6842
rect 27134 6888 27214 6921
rect 27134 6842 27147 6888
rect 27201 6842 27214 6888
rect 27134 6829 27214 6842
rect 27318 6888 27398 6921
rect 27318 6842 27331 6888
rect 27385 6842 27398 6888
rect 27318 6829 27398 6842
rect 34936 7500 35016 7513
rect 34936 7454 34949 7500
rect 35003 7454 35016 7500
rect 34936 7421 35016 7454
rect 35120 7500 35200 7513
rect 35120 7454 35133 7500
rect 35187 7454 35200 7500
rect 35120 7421 35200 7454
rect 35304 7500 35384 7513
rect 35304 7454 35317 7500
rect 35371 7454 35384 7500
rect 35304 7421 35384 7454
rect 34936 6888 35016 6921
rect 34936 6842 34949 6888
rect 35003 6842 35016 6888
rect 34936 6829 35016 6842
rect 35120 6888 35200 6921
rect 35120 6842 35133 6888
rect 35187 6842 35200 6888
rect 35120 6829 35200 6842
rect 35304 6888 35384 6921
rect 35304 6842 35317 6888
rect 35371 6842 35384 6888
rect 35304 6829 35384 6842
rect 36422 7500 36502 7513
rect 36422 7454 36435 7500
rect 36489 7454 36502 7500
rect 36422 7421 36502 7454
rect 36606 7500 36686 7513
rect 36606 7454 36619 7500
rect 36673 7454 36686 7500
rect 36606 7421 36686 7454
rect 36790 7500 36870 7513
rect 36790 7454 36803 7500
rect 36857 7454 36870 7500
rect 36790 7421 36870 7454
rect 36422 6888 36502 6921
rect 36422 6842 36435 6888
rect 36489 6842 36502 6888
rect 36422 6829 36502 6842
rect 36606 6888 36686 6921
rect 36606 6842 36619 6888
rect 36673 6842 36686 6888
rect 36606 6829 36686 6842
rect 36790 6888 36870 6921
rect 36790 6842 36803 6888
rect 36857 6842 36870 6888
rect 36790 6829 36870 6842
rect 44408 7500 44488 7513
rect 44408 7454 44421 7500
rect 44475 7454 44488 7500
rect 44408 7421 44488 7454
rect 44592 7500 44672 7513
rect 44592 7454 44605 7500
rect 44659 7454 44672 7500
rect 44592 7421 44672 7454
rect 44776 7500 44856 7513
rect 44776 7454 44789 7500
rect 44843 7454 44856 7500
rect 44776 7421 44856 7454
rect 44408 6888 44488 6921
rect 44408 6842 44421 6888
rect 44475 6842 44488 6888
rect 44408 6829 44488 6842
rect 44592 6888 44672 6921
rect 44592 6842 44605 6888
rect 44659 6842 44672 6888
rect 44592 6829 44672 6842
rect 44776 6888 44856 6921
rect 44776 6842 44789 6888
rect 44843 6842 44856 6888
rect 44776 6829 44856 6842
rect 45894 7500 45974 7513
rect 45894 7454 45907 7500
rect 45961 7454 45974 7500
rect 45894 7421 45974 7454
rect 46078 7500 46158 7513
rect 46078 7454 46091 7500
rect 46145 7454 46158 7500
rect 46078 7421 46158 7454
rect 46262 7500 46342 7513
rect 46262 7454 46275 7500
rect 46329 7454 46342 7500
rect 46262 7421 46342 7454
rect 45894 6888 45974 6921
rect 45894 6842 45907 6888
rect 45961 6842 45974 6888
rect 45894 6829 45974 6842
rect 46078 6888 46158 6921
rect 46078 6842 46091 6888
rect 46145 6842 46158 6888
rect 46078 6829 46158 6842
rect 46262 6888 46342 6921
rect 46262 6842 46275 6888
rect 46329 6842 46342 6888
rect 46262 6829 46342 6842
rect 53880 7500 53960 7513
rect 53880 7454 53893 7500
rect 53947 7454 53960 7500
rect 53880 7421 53960 7454
rect 54064 7500 54144 7513
rect 54064 7454 54077 7500
rect 54131 7454 54144 7500
rect 54064 7421 54144 7454
rect 54248 7500 54328 7513
rect 54248 7454 54261 7500
rect 54315 7454 54328 7500
rect 54248 7421 54328 7454
rect 53880 6888 53960 6921
rect 53880 6842 53893 6888
rect 53947 6842 53960 6888
rect 53880 6829 53960 6842
rect 54064 6888 54144 6921
rect 54064 6842 54077 6888
rect 54131 6842 54144 6888
rect 54064 6829 54144 6842
rect 54248 6888 54328 6921
rect 54248 6842 54261 6888
rect 54315 6842 54328 6888
rect 54248 6829 54328 6842
rect 55366 7500 55446 7513
rect 55366 7454 55379 7500
rect 55433 7454 55446 7500
rect 55366 7421 55446 7454
rect 55550 7500 55630 7513
rect 55550 7454 55563 7500
rect 55617 7454 55630 7500
rect 55550 7421 55630 7454
rect 55734 7500 55814 7513
rect 55734 7454 55747 7500
rect 55801 7454 55814 7500
rect 55734 7421 55814 7454
rect 55366 6888 55446 6921
rect 55366 6842 55379 6888
rect 55433 6842 55446 6888
rect 55366 6829 55446 6842
rect 55550 6888 55630 6921
rect 55550 6842 55563 6888
rect 55617 6842 55630 6888
rect 55550 6829 55630 6842
rect 55734 6888 55814 6921
rect 55734 6842 55747 6888
rect 55801 6842 55814 6888
rect 55734 6829 55814 6842
rect 6520 6339 6600 6352
rect 6520 6293 6533 6339
rect 6587 6293 6600 6339
rect 6520 6260 6600 6293
rect 6704 6339 6784 6352
rect 6704 6293 6717 6339
rect 6771 6293 6784 6339
rect 6704 6260 6784 6293
rect 6888 6339 6968 6352
rect 6888 6293 6901 6339
rect 6955 6293 6968 6339
rect 6888 6260 6968 6293
rect 6520 6027 6600 6060
rect 6520 5981 6533 6027
rect 6587 5981 6600 6027
rect 6520 5968 6600 5981
rect 6704 6027 6784 6060
rect 6704 5981 6717 6027
rect 6771 5981 6784 6027
rect 6704 5968 6784 5981
rect 6888 6027 6968 6060
rect 6888 5981 6901 6027
rect 6955 5981 6968 6027
rect 6888 5968 6968 5981
rect 8006 6339 8086 6352
rect 8006 6293 8019 6339
rect 8073 6293 8086 6339
rect 8006 6260 8086 6293
rect 8190 6339 8270 6352
rect 8190 6293 8203 6339
rect 8257 6293 8270 6339
rect 8190 6260 8270 6293
rect 8374 6339 8454 6352
rect 8374 6293 8387 6339
rect 8441 6293 8454 6339
rect 8374 6260 8454 6293
rect 8006 6027 8086 6060
rect 8006 5981 8019 6027
rect 8073 5981 8086 6027
rect 8006 5968 8086 5981
rect 8190 6027 8270 6060
rect 8190 5981 8203 6027
rect 8257 5981 8270 6027
rect 8190 5968 8270 5981
rect 8374 6027 8454 6060
rect 8374 5981 8387 6027
rect 8441 5981 8454 6027
rect 8374 5968 8454 5981
rect 15992 6339 16072 6352
rect 15992 6293 16005 6339
rect 16059 6293 16072 6339
rect 15992 6260 16072 6293
rect 16176 6339 16256 6352
rect 16176 6293 16189 6339
rect 16243 6293 16256 6339
rect 16176 6260 16256 6293
rect 16360 6339 16440 6352
rect 16360 6293 16373 6339
rect 16427 6293 16440 6339
rect 16360 6260 16440 6293
rect 15992 6027 16072 6060
rect 15992 5981 16005 6027
rect 16059 5981 16072 6027
rect 15992 5968 16072 5981
rect 16176 6027 16256 6060
rect 16176 5981 16189 6027
rect 16243 5981 16256 6027
rect 16176 5968 16256 5981
rect 16360 6027 16440 6060
rect 16360 5981 16373 6027
rect 16427 5981 16440 6027
rect 16360 5968 16440 5981
rect 17478 6339 17558 6352
rect 17478 6293 17491 6339
rect 17545 6293 17558 6339
rect 17478 6260 17558 6293
rect 17662 6339 17742 6352
rect 17662 6293 17675 6339
rect 17729 6293 17742 6339
rect 17662 6260 17742 6293
rect 17846 6339 17926 6352
rect 17846 6293 17859 6339
rect 17913 6293 17926 6339
rect 17846 6260 17926 6293
rect 17478 6027 17558 6060
rect 17478 5981 17491 6027
rect 17545 5981 17558 6027
rect 17478 5968 17558 5981
rect 17662 6027 17742 6060
rect 17662 5981 17675 6027
rect 17729 5981 17742 6027
rect 17662 5968 17742 5981
rect 17846 6027 17926 6060
rect 17846 5981 17859 6027
rect 17913 5981 17926 6027
rect 17846 5968 17926 5981
rect 25464 6340 25544 6353
rect 25464 6294 25477 6340
rect 25531 6294 25544 6340
rect 25464 6261 25544 6294
rect 25648 6340 25728 6353
rect 25648 6294 25661 6340
rect 25715 6294 25728 6340
rect 25648 6261 25728 6294
rect 25832 6340 25912 6353
rect 25832 6294 25845 6340
rect 25899 6294 25912 6340
rect 25832 6261 25912 6294
rect 25464 6028 25544 6061
rect 25464 5982 25477 6028
rect 25531 5982 25544 6028
rect 25464 5969 25544 5982
rect 25648 6028 25728 6061
rect 25648 5982 25661 6028
rect 25715 5982 25728 6028
rect 25648 5969 25728 5982
rect 25832 6028 25912 6061
rect 25832 5982 25845 6028
rect 25899 5982 25912 6028
rect 25832 5969 25912 5982
rect 26950 6340 27030 6353
rect 26950 6294 26963 6340
rect 27017 6294 27030 6340
rect 26950 6261 27030 6294
rect 27134 6340 27214 6353
rect 27134 6294 27147 6340
rect 27201 6294 27214 6340
rect 27134 6261 27214 6294
rect 27318 6340 27398 6353
rect 27318 6294 27331 6340
rect 27385 6294 27398 6340
rect 27318 6261 27398 6294
rect 26950 6028 27030 6061
rect 26950 5982 26963 6028
rect 27017 5982 27030 6028
rect 26950 5969 27030 5982
rect 27134 6028 27214 6061
rect 27134 5982 27147 6028
rect 27201 5982 27214 6028
rect 27134 5969 27214 5982
rect 27318 6028 27398 6061
rect 27318 5982 27331 6028
rect 27385 5982 27398 6028
rect 27318 5969 27398 5982
rect 34936 6340 35016 6353
rect 34936 6294 34949 6340
rect 35003 6294 35016 6340
rect 34936 6261 35016 6294
rect 35120 6340 35200 6353
rect 35120 6294 35133 6340
rect 35187 6294 35200 6340
rect 35120 6261 35200 6294
rect 35304 6340 35384 6353
rect 35304 6294 35317 6340
rect 35371 6294 35384 6340
rect 35304 6261 35384 6294
rect 34936 6028 35016 6061
rect 34936 5982 34949 6028
rect 35003 5982 35016 6028
rect 34936 5969 35016 5982
rect 35120 6028 35200 6061
rect 35120 5982 35133 6028
rect 35187 5982 35200 6028
rect 35120 5969 35200 5982
rect 35304 6028 35384 6061
rect 35304 5982 35317 6028
rect 35371 5982 35384 6028
rect 35304 5969 35384 5982
rect 36422 6340 36502 6353
rect 36422 6294 36435 6340
rect 36489 6294 36502 6340
rect 36422 6261 36502 6294
rect 36606 6340 36686 6353
rect 36606 6294 36619 6340
rect 36673 6294 36686 6340
rect 36606 6261 36686 6294
rect 36790 6340 36870 6353
rect 36790 6294 36803 6340
rect 36857 6294 36870 6340
rect 36790 6261 36870 6294
rect 36422 6028 36502 6061
rect 36422 5982 36435 6028
rect 36489 5982 36502 6028
rect 36422 5969 36502 5982
rect 36606 6028 36686 6061
rect 36606 5982 36619 6028
rect 36673 5982 36686 6028
rect 36606 5969 36686 5982
rect 36790 6028 36870 6061
rect 36790 5982 36803 6028
rect 36857 5982 36870 6028
rect 36790 5969 36870 5982
rect 44408 6340 44488 6353
rect 44408 6294 44421 6340
rect 44475 6294 44488 6340
rect 44408 6261 44488 6294
rect 44592 6340 44672 6353
rect 44592 6294 44605 6340
rect 44659 6294 44672 6340
rect 44592 6261 44672 6294
rect 44776 6340 44856 6353
rect 44776 6294 44789 6340
rect 44843 6294 44856 6340
rect 44776 6261 44856 6294
rect 44408 6028 44488 6061
rect 44408 5982 44421 6028
rect 44475 5982 44488 6028
rect 44408 5969 44488 5982
rect 44592 6028 44672 6061
rect 44592 5982 44605 6028
rect 44659 5982 44672 6028
rect 44592 5969 44672 5982
rect 44776 6028 44856 6061
rect 44776 5982 44789 6028
rect 44843 5982 44856 6028
rect 44776 5969 44856 5982
rect 45894 6340 45974 6353
rect 45894 6294 45907 6340
rect 45961 6294 45974 6340
rect 45894 6261 45974 6294
rect 46078 6340 46158 6353
rect 46078 6294 46091 6340
rect 46145 6294 46158 6340
rect 46078 6261 46158 6294
rect 46262 6340 46342 6353
rect 46262 6294 46275 6340
rect 46329 6294 46342 6340
rect 46262 6261 46342 6294
rect 45894 6028 45974 6061
rect 45894 5982 45907 6028
rect 45961 5982 45974 6028
rect 45894 5969 45974 5982
rect 46078 6028 46158 6061
rect 46078 5982 46091 6028
rect 46145 5982 46158 6028
rect 46078 5969 46158 5982
rect 46262 6028 46342 6061
rect 46262 5982 46275 6028
rect 46329 5982 46342 6028
rect 46262 5969 46342 5982
rect 53880 6340 53960 6353
rect 53880 6294 53893 6340
rect 53947 6294 53960 6340
rect 53880 6261 53960 6294
rect 54064 6340 54144 6353
rect 54064 6294 54077 6340
rect 54131 6294 54144 6340
rect 54064 6261 54144 6294
rect 54248 6340 54328 6353
rect 54248 6294 54261 6340
rect 54315 6294 54328 6340
rect 54248 6261 54328 6294
rect 53880 6028 53960 6061
rect 53880 5982 53893 6028
rect 53947 5982 53960 6028
rect 53880 5969 53960 5982
rect 54064 6028 54144 6061
rect 54064 5982 54077 6028
rect 54131 5982 54144 6028
rect 54064 5969 54144 5982
rect 54248 6028 54328 6061
rect 54248 5982 54261 6028
rect 54315 5982 54328 6028
rect 54248 5969 54328 5982
rect 55366 6340 55446 6353
rect 55366 6294 55379 6340
rect 55433 6294 55446 6340
rect 55366 6261 55446 6294
rect 55550 6340 55630 6353
rect 55550 6294 55563 6340
rect 55617 6294 55630 6340
rect 55550 6261 55630 6294
rect 55734 6340 55814 6353
rect 55734 6294 55747 6340
rect 55801 6294 55814 6340
rect 55734 6261 55814 6294
rect 55366 6028 55446 6061
rect 55366 5982 55379 6028
rect 55433 5982 55446 6028
rect 55366 5969 55446 5982
rect 55550 6028 55630 6061
rect 55550 5982 55563 6028
rect 55617 5982 55630 6028
rect 55550 5969 55630 5982
rect 55734 6028 55814 6061
rect 55734 5982 55747 6028
rect 55801 5982 55814 6028
rect 55734 5969 55814 5982
rect 6520 5294 6600 5307
rect 6520 5248 6533 5294
rect 6587 5248 6600 5294
rect 6520 5215 6600 5248
rect 6704 5294 6784 5307
rect 6704 5248 6717 5294
rect 6771 5248 6784 5294
rect 6704 5215 6784 5248
rect 6888 5294 6968 5307
rect 6888 5248 6901 5294
rect 6955 5248 6968 5294
rect 6888 5215 6968 5248
rect 6520 4682 6600 4715
rect 6520 4636 6533 4682
rect 6587 4636 6600 4682
rect 6520 4623 6600 4636
rect 6704 4682 6784 4715
rect 6704 4636 6717 4682
rect 6771 4636 6784 4682
rect 6704 4623 6784 4636
rect 6888 4682 6968 4715
rect 6888 4636 6901 4682
rect 6955 4636 6968 4682
rect 6888 4623 6968 4636
rect 8006 5295 8086 5308
rect 8006 5249 8019 5295
rect 8073 5249 8086 5295
rect 8006 5216 8086 5249
rect 8190 5295 8270 5308
rect 8190 5249 8203 5295
rect 8257 5249 8270 5295
rect 8190 5216 8270 5249
rect 8374 5295 8454 5308
rect 8374 5249 8387 5295
rect 8441 5249 8454 5295
rect 8374 5216 8454 5249
rect 8006 4683 8086 4716
rect 8006 4637 8019 4683
rect 8073 4637 8086 4683
rect 8006 4624 8086 4637
rect 8190 4683 8270 4716
rect 8190 4637 8203 4683
rect 8257 4637 8270 4683
rect 8190 4624 8270 4637
rect 8374 4683 8454 4716
rect 8374 4637 8387 4683
rect 8441 4637 8454 4683
rect 8374 4624 8454 4637
rect 15992 5294 16072 5307
rect 15992 5248 16005 5294
rect 16059 5248 16072 5294
rect 15992 5215 16072 5248
rect 16176 5294 16256 5307
rect 16176 5248 16189 5294
rect 16243 5248 16256 5294
rect 16176 5215 16256 5248
rect 16360 5294 16440 5307
rect 16360 5248 16373 5294
rect 16427 5248 16440 5294
rect 16360 5215 16440 5248
rect 15992 4682 16072 4715
rect 15992 4636 16005 4682
rect 16059 4636 16072 4682
rect 15992 4623 16072 4636
rect 16176 4682 16256 4715
rect 16176 4636 16189 4682
rect 16243 4636 16256 4682
rect 16176 4623 16256 4636
rect 16360 4682 16440 4715
rect 16360 4636 16373 4682
rect 16427 4636 16440 4682
rect 16360 4623 16440 4636
rect 17478 5295 17558 5308
rect 17478 5249 17491 5295
rect 17545 5249 17558 5295
rect 17478 5216 17558 5249
rect 17662 5295 17742 5308
rect 17662 5249 17675 5295
rect 17729 5249 17742 5295
rect 17662 5216 17742 5249
rect 17846 5295 17926 5308
rect 17846 5249 17859 5295
rect 17913 5249 17926 5295
rect 17846 5216 17926 5249
rect 17478 4683 17558 4716
rect 17478 4637 17491 4683
rect 17545 4637 17558 4683
rect 17478 4624 17558 4637
rect 17662 4683 17742 4716
rect 17662 4637 17675 4683
rect 17729 4637 17742 4683
rect 17662 4624 17742 4637
rect 17846 4683 17926 4716
rect 17846 4637 17859 4683
rect 17913 4637 17926 4683
rect 17846 4624 17926 4637
rect 25464 5295 25544 5308
rect 25464 5249 25477 5295
rect 25531 5249 25544 5295
rect 25464 5216 25544 5249
rect 25648 5295 25728 5308
rect 25648 5249 25661 5295
rect 25715 5249 25728 5295
rect 25648 5216 25728 5249
rect 25832 5295 25912 5308
rect 25832 5249 25845 5295
rect 25899 5249 25912 5295
rect 25832 5216 25912 5249
rect 25464 4683 25544 4716
rect 25464 4637 25477 4683
rect 25531 4637 25544 4683
rect 25464 4624 25544 4637
rect 25648 4683 25728 4716
rect 25648 4637 25661 4683
rect 25715 4637 25728 4683
rect 25648 4624 25728 4637
rect 25832 4683 25912 4716
rect 25832 4637 25845 4683
rect 25899 4637 25912 4683
rect 25832 4624 25912 4637
rect 26950 5296 27030 5309
rect 26950 5250 26963 5296
rect 27017 5250 27030 5296
rect 26950 5217 27030 5250
rect 27134 5296 27214 5309
rect 27134 5250 27147 5296
rect 27201 5250 27214 5296
rect 27134 5217 27214 5250
rect 27318 5296 27398 5309
rect 27318 5250 27331 5296
rect 27385 5250 27398 5296
rect 27318 5217 27398 5250
rect 26950 4684 27030 4717
rect 26950 4638 26963 4684
rect 27017 4638 27030 4684
rect 26950 4625 27030 4638
rect 27134 4684 27214 4717
rect 27134 4638 27147 4684
rect 27201 4638 27214 4684
rect 27134 4625 27214 4638
rect 27318 4684 27398 4717
rect 27318 4638 27331 4684
rect 27385 4638 27398 4684
rect 27318 4625 27398 4638
rect 34936 5295 35016 5308
rect 34936 5249 34949 5295
rect 35003 5249 35016 5295
rect 34936 5216 35016 5249
rect 35120 5295 35200 5308
rect 35120 5249 35133 5295
rect 35187 5249 35200 5295
rect 35120 5216 35200 5249
rect 35304 5295 35384 5308
rect 35304 5249 35317 5295
rect 35371 5249 35384 5295
rect 35304 5216 35384 5249
rect 34936 4683 35016 4716
rect 34936 4637 34949 4683
rect 35003 4637 35016 4683
rect 34936 4624 35016 4637
rect 35120 4683 35200 4716
rect 35120 4637 35133 4683
rect 35187 4637 35200 4683
rect 35120 4624 35200 4637
rect 35304 4683 35384 4716
rect 35304 4637 35317 4683
rect 35371 4637 35384 4683
rect 35304 4624 35384 4637
rect 36422 5296 36502 5309
rect 36422 5250 36435 5296
rect 36489 5250 36502 5296
rect 36422 5217 36502 5250
rect 36606 5296 36686 5309
rect 36606 5250 36619 5296
rect 36673 5250 36686 5296
rect 36606 5217 36686 5250
rect 36790 5296 36870 5309
rect 36790 5250 36803 5296
rect 36857 5250 36870 5296
rect 36790 5217 36870 5250
rect 36422 4684 36502 4717
rect 36422 4638 36435 4684
rect 36489 4638 36502 4684
rect 36422 4625 36502 4638
rect 36606 4684 36686 4717
rect 36606 4638 36619 4684
rect 36673 4638 36686 4684
rect 36606 4625 36686 4638
rect 36790 4684 36870 4717
rect 36790 4638 36803 4684
rect 36857 4638 36870 4684
rect 36790 4625 36870 4638
rect 44408 5295 44488 5308
rect 44408 5249 44421 5295
rect 44475 5249 44488 5295
rect 44408 5216 44488 5249
rect 44592 5295 44672 5308
rect 44592 5249 44605 5295
rect 44659 5249 44672 5295
rect 44592 5216 44672 5249
rect 44776 5295 44856 5308
rect 44776 5249 44789 5295
rect 44843 5249 44856 5295
rect 44776 5216 44856 5249
rect 44408 4683 44488 4716
rect 44408 4637 44421 4683
rect 44475 4637 44488 4683
rect 44408 4624 44488 4637
rect 44592 4683 44672 4716
rect 44592 4637 44605 4683
rect 44659 4637 44672 4683
rect 44592 4624 44672 4637
rect 44776 4683 44856 4716
rect 44776 4637 44789 4683
rect 44843 4637 44856 4683
rect 44776 4624 44856 4637
rect 45894 5296 45974 5309
rect 45894 5250 45907 5296
rect 45961 5250 45974 5296
rect 45894 5217 45974 5250
rect 46078 5296 46158 5309
rect 46078 5250 46091 5296
rect 46145 5250 46158 5296
rect 46078 5217 46158 5250
rect 46262 5296 46342 5309
rect 46262 5250 46275 5296
rect 46329 5250 46342 5296
rect 46262 5217 46342 5250
rect 45894 4684 45974 4717
rect 45894 4638 45907 4684
rect 45961 4638 45974 4684
rect 45894 4625 45974 4638
rect 46078 4684 46158 4717
rect 46078 4638 46091 4684
rect 46145 4638 46158 4684
rect 46078 4625 46158 4638
rect 46262 4684 46342 4717
rect 46262 4638 46275 4684
rect 46329 4638 46342 4684
rect 46262 4625 46342 4638
rect 53880 5295 53960 5308
rect 53880 5249 53893 5295
rect 53947 5249 53960 5295
rect 53880 5216 53960 5249
rect 54064 5295 54144 5308
rect 54064 5249 54077 5295
rect 54131 5249 54144 5295
rect 54064 5216 54144 5249
rect 54248 5295 54328 5308
rect 54248 5249 54261 5295
rect 54315 5249 54328 5295
rect 54248 5216 54328 5249
rect 53880 4683 53960 4716
rect 53880 4637 53893 4683
rect 53947 4637 53960 4683
rect 53880 4624 53960 4637
rect 54064 4683 54144 4716
rect 54064 4637 54077 4683
rect 54131 4637 54144 4683
rect 54064 4624 54144 4637
rect 54248 4683 54328 4716
rect 54248 4637 54261 4683
rect 54315 4637 54328 4683
rect 54248 4624 54328 4637
rect 55366 5296 55446 5309
rect 55366 5250 55379 5296
rect 55433 5250 55446 5296
rect 55366 5217 55446 5250
rect 55550 5296 55630 5309
rect 55550 5250 55563 5296
rect 55617 5250 55630 5296
rect 55550 5217 55630 5250
rect 55734 5296 55814 5309
rect 55734 5250 55747 5296
rect 55801 5250 55814 5296
rect 55734 5217 55814 5250
rect 55366 4684 55446 4717
rect 55366 4638 55379 4684
rect 55433 4638 55446 4684
rect 55366 4625 55446 4638
rect 55550 4684 55630 4717
rect 55550 4638 55563 4684
rect 55617 4638 55630 4684
rect 55550 4625 55630 4638
rect 55734 4684 55814 4717
rect 55734 4638 55747 4684
rect 55801 4638 55814 4684
rect 55734 4625 55814 4638
rect 1378 4179 1478 4192
rect 1378 4133 1391 4179
rect 1465 4133 1478 4179
rect 1378 4100 1478 4133
rect 1378 3467 1478 3500
rect 1378 3421 1391 3467
rect 1465 3421 1478 3467
rect 1378 3408 1478 3421
rect 2266 4179 2366 4192
rect 2266 4133 2279 4179
rect 2353 4133 2366 4179
rect 2266 4100 2366 4133
rect 2266 3467 2366 3500
rect 2266 3421 2279 3467
rect 2353 3421 2366 3467
rect 2266 3408 2366 3421
rect 2746 4179 2846 4192
rect 2746 4133 2759 4179
rect 2833 4133 2846 4179
rect 2746 4100 2846 4133
rect 2746 3467 2846 3500
rect 2746 3421 2759 3467
rect 2833 3421 2846 3467
rect 2746 3408 2846 3421
rect 6520 4134 6600 4147
rect 6520 4088 6533 4134
rect 6587 4088 6600 4134
rect 6520 4055 6600 4088
rect 6704 4134 6784 4147
rect 6704 4088 6717 4134
rect 6771 4088 6784 4134
rect 6704 4055 6784 4088
rect 6888 4134 6968 4147
rect 6888 4088 6901 4134
rect 6955 4088 6968 4134
rect 6888 4055 6968 4088
rect 6520 3822 6600 3855
rect 6520 3776 6533 3822
rect 6587 3776 6600 3822
rect 6520 3763 6600 3776
rect 6704 3822 6784 3855
rect 6704 3776 6717 3822
rect 6771 3776 6784 3822
rect 6704 3763 6784 3776
rect 6888 3822 6968 3855
rect 6888 3776 6901 3822
rect 6955 3776 6968 3822
rect 6888 3763 6968 3776
rect 8006 4135 8086 4148
rect 8006 4089 8019 4135
rect 8073 4089 8086 4135
rect 8006 4056 8086 4089
rect 8190 4135 8270 4148
rect 8190 4089 8203 4135
rect 8257 4089 8270 4135
rect 8190 4056 8270 4089
rect 8374 4135 8454 4148
rect 8374 4089 8387 4135
rect 8441 4089 8454 4135
rect 8374 4056 8454 4089
rect 8006 3823 8086 3856
rect 8006 3777 8019 3823
rect 8073 3777 8086 3823
rect 8006 3764 8086 3777
rect 8190 3823 8270 3856
rect 8190 3777 8203 3823
rect 8257 3777 8270 3823
rect 8190 3764 8270 3777
rect 8374 3823 8454 3856
rect 8374 3777 8387 3823
rect 8441 3777 8454 3823
rect 8374 3764 8454 3777
rect 10850 4179 10950 4192
rect 10850 4133 10863 4179
rect 10937 4133 10950 4179
rect 10850 4100 10950 4133
rect 10850 3467 10950 3500
rect 10850 3421 10863 3467
rect 10937 3421 10950 3467
rect 10850 3408 10950 3421
rect 11738 4179 11838 4192
rect 11738 4133 11751 4179
rect 11825 4133 11838 4179
rect 11738 4100 11838 4133
rect 11738 3467 11838 3500
rect 11738 3421 11751 3467
rect 11825 3421 11838 3467
rect 11738 3408 11838 3421
rect 12218 4179 12318 4192
rect 12218 4133 12231 4179
rect 12305 4133 12318 4179
rect 12218 4100 12318 4133
rect 12218 3467 12318 3500
rect 12218 3421 12231 3467
rect 12305 3421 12318 3467
rect 12218 3408 12318 3421
rect 15992 4134 16072 4147
rect 15992 4088 16005 4134
rect 16059 4088 16072 4134
rect 15992 4055 16072 4088
rect 16176 4134 16256 4147
rect 16176 4088 16189 4134
rect 16243 4088 16256 4134
rect 16176 4055 16256 4088
rect 16360 4134 16440 4147
rect 16360 4088 16373 4134
rect 16427 4088 16440 4134
rect 16360 4055 16440 4088
rect 15992 3822 16072 3855
rect 15992 3776 16005 3822
rect 16059 3776 16072 3822
rect 15992 3763 16072 3776
rect 16176 3822 16256 3855
rect 16176 3776 16189 3822
rect 16243 3776 16256 3822
rect 16176 3763 16256 3776
rect 16360 3822 16440 3855
rect 16360 3776 16373 3822
rect 16427 3776 16440 3822
rect 16360 3763 16440 3776
rect 17478 4135 17558 4148
rect 17478 4089 17491 4135
rect 17545 4089 17558 4135
rect 17478 4056 17558 4089
rect 17662 4135 17742 4148
rect 17662 4089 17675 4135
rect 17729 4089 17742 4135
rect 17662 4056 17742 4089
rect 17846 4135 17926 4148
rect 17846 4089 17859 4135
rect 17913 4089 17926 4135
rect 17846 4056 17926 4089
rect 17478 3823 17558 3856
rect 17478 3777 17491 3823
rect 17545 3777 17558 3823
rect 17478 3764 17558 3777
rect 17662 3823 17742 3856
rect 17662 3777 17675 3823
rect 17729 3777 17742 3823
rect 17662 3764 17742 3777
rect 17846 3823 17926 3856
rect 17846 3777 17859 3823
rect 17913 3777 17926 3823
rect 17846 3764 17926 3777
rect 20322 4180 20422 4193
rect 20322 4134 20335 4180
rect 20409 4134 20422 4180
rect 20322 4101 20422 4134
rect 20322 3468 20422 3501
rect 20322 3422 20335 3468
rect 20409 3422 20422 3468
rect 20322 3409 20422 3422
rect 21210 4180 21310 4193
rect 21210 4134 21223 4180
rect 21297 4134 21310 4180
rect 21210 4101 21310 4134
rect 21210 3468 21310 3501
rect 21210 3422 21223 3468
rect 21297 3422 21310 3468
rect 21210 3409 21310 3422
rect 21690 4180 21790 4193
rect 21690 4134 21703 4180
rect 21777 4134 21790 4180
rect 21690 4101 21790 4134
rect 21690 3468 21790 3501
rect 21690 3422 21703 3468
rect 21777 3422 21790 3468
rect 21690 3409 21790 3422
rect 25464 4135 25544 4148
rect 25464 4089 25477 4135
rect 25531 4089 25544 4135
rect 25464 4056 25544 4089
rect 25648 4135 25728 4148
rect 25648 4089 25661 4135
rect 25715 4089 25728 4135
rect 25648 4056 25728 4089
rect 25832 4135 25912 4148
rect 25832 4089 25845 4135
rect 25899 4089 25912 4135
rect 25832 4056 25912 4089
rect 25464 3823 25544 3856
rect 25464 3777 25477 3823
rect 25531 3777 25544 3823
rect 25464 3764 25544 3777
rect 25648 3823 25728 3856
rect 25648 3777 25661 3823
rect 25715 3777 25728 3823
rect 25648 3764 25728 3777
rect 25832 3823 25912 3856
rect 25832 3777 25845 3823
rect 25899 3777 25912 3823
rect 25832 3764 25912 3777
rect 26950 4136 27030 4149
rect 26950 4090 26963 4136
rect 27017 4090 27030 4136
rect 26950 4057 27030 4090
rect 27134 4136 27214 4149
rect 27134 4090 27147 4136
rect 27201 4090 27214 4136
rect 27134 4057 27214 4090
rect 27318 4136 27398 4149
rect 27318 4090 27331 4136
rect 27385 4090 27398 4136
rect 27318 4057 27398 4090
rect 26950 3824 27030 3857
rect 26950 3778 26963 3824
rect 27017 3778 27030 3824
rect 26950 3765 27030 3778
rect 27134 3824 27214 3857
rect 27134 3778 27147 3824
rect 27201 3778 27214 3824
rect 27134 3765 27214 3778
rect 27318 3824 27398 3857
rect 27318 3778 27331 3824
rect 27385 3778 27398 3824
rect 27318 3765 27398 3778
rect 29794 4180 29894 4193
rect 29794 4134 29807 4180
rect 29881 4134 29894 4180
rect 29794 4101 29894 4134
rect 29794 3468 29894 3501
rect 29794 3422 29807 3468
rect 29881 3422 29894 3468
rect 29794 3409 29894 3422
rect 30682 4180 30782 4193
rect 30682 4134 30695 4180
rect 30769 4134 30782 4180
rect 30682 4101 30782 4134
rect 30682 3468 30782 3501
rect 30682 3422 30695 3468
rect 30769 3422 30782 3468
rect 30682 3409 30782 3422
rect 31162 4180 31262 4193
rect 31162 4134 31175 4180
rect 31249 4134 31262 4180
rect 31162 4101 31262 4134
rect 31162 3468 31262 3501
rect 31162 3422 31175 3468
rect 31249 3422 31262 3468
rect 31162 3409 31262 3422
rect 34936 4135 35016 4148
rect 34936 4089 34949 4135
rect 35003 4089 35016 4135
rect 34936 4056 35016 4089
rect 35120 4135 35200 4148
rect 35120 4089 35133 4135
rect 35187 4089 35200 4135
rect 35120 4056 35200 4089
rect 35304 4135 35384 4148
rect 35304 4089 35317 4135
rect 35371 4089 35384 4135
rect 35304 4056 35384 4089
rect 34936 3823 35016 3856
rect 34936 3777 34949 3823
rect 35003 3777 35016 3823
rect 34936 3764 35016 3777
rect 35120 3823 35200 3856
rect 35120 3777 35133 3823
rect 35187 3777 35200 3823
rect 35120 3764 35200 3777
rect 35304 3823 35384 3856
rect 35304 3777 35317 3823
rect 35371 3777 35384 3823
rect 35304 3764 35384 3777
rect 36422 4136 36502 4149
rect 36422 4090 36435 4136
rect 36489 4090 36502 4136
rect 36422 4057 36502 4090
rect 36606 4136 36686 4149
rect 36606 4090 36619 4136
rect 36673 4090 36686 4136
rect 36606 4057 36686 4090
rect 36790 4136 36870 4149
rect 36790 4090 36803 4136
rect 36857 4090 36870 4136
rect 36790 4057 36870 4090
rect 36422 3824 36502 3857
rect 36422 3778 36435 3824
rect 36489 3778 36502 3824
rect 36422 3765 36502 3778
rect 36606 3824 36686 3857
rect 36606 3778 36619 3824
rect 36673 3778 36686 3824
rect 36606 3765 36686 3778
rect 36790 3824 36870 3857
rect 36790 3778 36803 3824
rect 36857 3778 36870 3824
rect 36790 3765 36870 3778
rect 39266 4180 39366 4193
rect 39266 4134 39279 4180
rect 39353 4134 39366 4180
rect 39266 4101 39366 4134
rect 39266 3468 39366 3501
rect 39266 3422 39279 3468
rect 39353 3422 39366 3468
rect 39266 3409 39366 3422
rect 40154 4180 40254 4193
rect 40154 4134 40167 4180
rect 40241 4134 40254 4180
rect 40154 4101 40254 4134
rect 40154 3468 40254 3501
rect 40154 3422 40167 3468
rect 40241 3422 40254 3468
rect 40154 3409 40254 3422
rect 40634 4180 40734 4193
rect 40634 4134 40647 4180
rect 40721 4134 40734 4180
rect 40634 4101 40734 4134
rect 40634 3468 40734 3501
rect 40634 3422 40647 3468
rect 40721 3422 40734 3468
rect 40634 3409 40734 3422
rect 44408 4135 44488 4148
rect 44408 4089 44421 4135
rect 44475 4089 44488 4135
rect 44408 4056 44488 4089
rect 44592 4135 44672 4148
rect 44592 4089 44605 4135
rect 44659 4089 44672 4135
rect 44592 4056 44672 4089
rect 44776 4135 44856 4148
rect 44776 4089 44789 4135
rect 44843 4089 44856 4135
rect 44776 4056 44856 4089
rect 44408 3823 44488 3856
rect 44408 3777 44421 3823
rect 44475 3777 44488 3823
rect 44408 3764 44488 3777
rect 44592 3823 44672 3856
rect 44592 3777 44605 3823
rect 44659 3777 44672 3823
rect 44592 3764 44672 3777
rect 44776 3823 44856 3856
rect 44776 3777 44789 3823
rect 44843 3777 44856 3823
rect 44776 3764 44856 3777
rect 45894 4136 45974 4149
rect 45894 4090 45907 4136
rect 45961 4090 45974 4136
rect 45894 4057 45974 4090
rect 46078 4136 46158 4149
rect 46078 4090 46091 4136
rect 46145 4090 46158 4136
rect 46078 4057 46158 4090
rect 46262 4136 46342 4149
rect 46262 4090 46275 4136
rect 46329 4090 46342 4136
rect 46262 4057 46342 4090
rect 45894 3824 45974 3857
rect 45894 3778 45907 3824
rect 45961 3778 45974 3824
rect 45894 3765 45974 3778
rect 46078 3824 46158 3857
rect 46078 3778 46091 3824
rect 46145 3778 46158 3824
rect 46078 3765 46158 3778
rect 46262 3824 46342 3857
rect 46262 3778 46275 3824
rect 46329 3778 46342 3824
rect 46262 3765 46342 3778
rect 48738 4180 48838 4193
rect 48738 4134 48751 4180
rect 48825 4134 48838 4180
rect 48738 4101 48838 4134
rect 48738 3468 48838 3501
rect 48738 3422 48751 3468
rect 48825 3422 48838 3468
rect 48738 3409 48838 3422
rect 49626 4180 49726 4193
rect 49626 4134 49639 4180
rect 49713 4134 49726 4180
rect 49626 4101 49726 4134
rect 49626 3468 49726 3501
rect 49626 3422 49639 3468
rect 49713 3422 49726 3468
rect 49626 3409 49726 3422
rect 50106 4180 50206 4193
rect 50106 4134 50119 4180
rect 50193 4134 50206 4180
rect 50106 4101 50206 4134
rect 50106 3468 50206 3501
rect 50106 3422 50119 3468
rect 50193 3422 50206 3468
rect 50106 3409 50206 3422
rect 53880 4135 53960 4148
rect 53880 4089 53893 4135
rect 53947 4089 53960 4135
rect 53880 4056 53960 4089
rect 54064 4135 54144 4148
rect 54064 4089 54077 4135
rect 54131 4089 54144 4135
rect 54064 4056 54144 4089
rect 54248 4135 54328 4148
rect 54248 4089 54261 4135
rect 54315 4089 54328 4135
rect 54248 4056 54328 4089
rect 53880 3823 53960 3856
rect 53880 3777 53893 3823
rect 53947 3777 53960 3823
rect 53880 3764 53960 3777
rect 54064 3823 54144 3856
rect 54064 3777 54077 3823
rect 54131 3777 54144 3823
rect 54064 3764 54144 3777
rect 54248 3823 54328 3856
rect 54248 3777 54261 3823
rect 54315 3777 54328 3823
rect 54248 3764 54328 3777
rect 55366 4136 55446 4149
rect 55366 4090 55379 4136
rect 55433 4090 55446 4136
rect 55366 4057 55446 4090
rect 55550 4136 55630 4149
rect 55550 4090 55563 4136
rect 55617 4090 55630 4136
rect 55550 4057 55630 4090
rect 55734 4136 55814 4149
rect 55734 4090 55747 4136
rect 55801 4090 55814 4136
rect 55734 4057 55814 4090
rect 55366 3824 55446 3857
rect 55366 3778 55379 3824
rect 55433 3778 55446 3824
rect 55366 3765 55446 3778
rect 55550 3824 55630 3857
rect 55550 3778 55563 3824
rect 55617 3778 55630 3824
rect 55550 3765 55630 3778
rect 55734 3824 55814 3857
rect 55734 3778 55747 3824
rect 55801 3778 55814 3824
rect 55734 3765 55814 3778
rect 484 2759 584 2772
rect 484 2713 497 2759
rect 571 2713 584 2759
rect 484 2680 584 2713
rect 484 2047 584 2080
rect 484 2001 497 2047
rect 571 2001 584 2047
rect 484 1988 584 2001
rect 1378 3059 1478 3072
rect 1378 3013 1391 3059
rect 1465 3013 1478 3059
rect 1378 2980 1478 3013
rect 1582 3059 1682 3072
rect 1582 3013 1595 3059
rect 1669 3013 1682 3059
rect 1582 2980 1682 3013
rect 1378 2747 1478 2780
rect 1378 2701 1391 2747
rect 1465 2701 1478 2747
rect 1378 2688 1478 2701
rect 1582 2747 1682 2780
rect 1582 2701 1595 2747
rect 1669 2701 1682 2747
rect 1582 2688 1682 2701
rect 2062 3059 2162 3072
rect 2062 3013 2075 3059
rect 2149 3013 2162 3059
rect 2062 2980 2162 3013
rect 2266 3059 2366 3072
rect 2266 3013 2279 3059
rect 2353 3013 2366 3059
rect 2266 2980 2366 3013
rect 2062 2747 2162 2780
rect 2062 2701 2075 2747
rect 2149 2701 2162 2747
rect 2062 2688 2162 2701
rect 2266 2747 2366 2780
rect 2266 2701 2279 2747
rect 2353 2701 2366 2747
rect 2266 2688 2366 2701
rect 2746 3059 2846 3072
rect 2746 3013 2759 3059
rect 2833 3013 2846 3059
rect 2746 2980 2846 3013
rect 2746 2747 2846 2780
rect 2746 2701 2759 2747
rect 2833 2701 2846 2747
rect 2746 2688 2846 2701
rect 3606 3003 3706 3016
rect 3606 2957 3619 3003
rect 3693 2957 3706 3003
rect 3606 2924 3706 2957
rect 3810 3003 3910 3016
rect 3810 2957 3823 3003
rect 3897 2957 3910 3003
rect 3810 2924 3910 2957
rect 3606 2291 3706 2324
rect 3606 2245 3619 2291
rect 3693 2245 3706 2291
rect 3606 2232 3706 2245
rect 3810 2291 3910 2324
rect 3810 2245 3823 2291
rect 3897 2245 3910 2291
rect 3810 2232 3910 2245
rect 4290 3003 4390 3016
rect 4290 2957 4303 3003
rect 4377 2957 4390 3003
rect 4290 2924 4390 2957
rect 4494 3003 4594 3016
rect 4494 2957 4507 3003
rect 4581 2957 4594 3003
rect 4494 2924 4594 2957
rect 4290 2291 4390 2324
rect 4290 2245 4303 2291
rect 4377 2245 4390 2291
rect 4290 2232 4390 2245
rect 4494 2291 4594 2324
rect 4494 2245 4507 2291
rect 4581 2245 4594 2291
rect 4494 2232 4594 2245
rect 4974 3003 5074 3016
rect 4974 2957 4987 3003
rect 5061 2957 5074 3003
rect 4974 2924 5074 2957
rect 4974 2291 5074 2324
rect 4974 2245 4987 2291
rect 5061 2245 5074 2291
rect 4974 2232 5074 2245
rect 6520 3089 6600 3102
rect 6520 3043 6533 3089
rect 6587 3043 6600 3089
rect 6520 3010 6600 3043
rect 6704 3089 6784 3102
rect 6704 3043 6717 3089
rect 6771 3043 6784 3089
rect 6704 3010 6784 3043
rect 6888 3089 6968 3102
rect 6888 3043 6901 3089
rect 6955 3043 6968 3089
rect 6888 3010 6968 3043
rect 6520 2477 6600 2510
rect 6520 2431 6533 2477
rect 6587 2431 6600 2477
rect 6520 2418 6600 2431
rect 6704 2477 6784 2510
rect 6704 2431 6717 2477
rect 6771 2431 6784 2477
rect 6704 2418 6784 2431
rect 6888 2477 6968 2510
rect 6888 2431 6901 2477
rect 6955 2431 6968 2477
rect 6888 2418 6968 2431
rect 484 1639 584 1652
rect 484 1593 497 1639
rect 571 1593 584 1639
rect 484 1560 584 1593
rect 484 1327 584 1360
rect 484 1281 497 1327
rect 571 1281 584 1327
rect 484 1268 584 1281
rect 1378 1839 1478 1852
rect 1378 1793 1391 1839
rect 1465 1793 1478 1839
rect 1378 1760 1478 1793
rect 1378 1127 1478 1160
rect 1378 1081 1391 1127
rect 1465 1081 1478 1127
rect 1378 1068 1478 1081
rect 2266 1839 2366 1852
rect 2266 1793 2279 1839
rect 2353 1793 2366 1839
rect 2266 1760 2366 1793
rect 2266 1127 2366 1160
rect 2266 1081 2279 1127
rect 2353 1081 2366 1127
rect 2266 1068 2366 1081
rect 2746 1839 2846 1852
rect 2746 1793 2759 1839
rect 2833 1793 2846 1839
rect 2746 1760 2846 1793
rect 2746 1127 2846 1160
rect 2746 1081 2759 1127
rect 2833 1081 2846 1127
rect 2746 1068 2846 1081
rect 3606 1883 3706 1896
rect 3606 1837 3619 1883
rect 3693 1837 3706 1883
rect 3606 1804 3706 1837
rect 3606 1571 3706 1604
rect 3606 1525 3619 1571
rect 3693 1525 3706 1571
rect 3606 1512 3706 1525
rect 4290 1883 4390 1896
rect 4290 1837 4303 1883
rect 4377 1837 4390 1883
rect 4290 1804 4390 1837
rect 4290 1571 4390 1604
rect 4290 1525 4303 1571
rect 4377 1525 4390 1571
rect 4290 1512 4390 1525
rect 4974 1883 5074 1896
rect 4974 1837 4987 1883
rect 5061 1837 5074 1883
rect 4974 1804 5074 1837
rect 4974 1571 5074 1604
rect 4974 1525 4987 1571
rect 5061 1525 5074 1571
rect 4974 1512 5074 1525
rect 6520 1929 6600 1942
rect 6520 1883 6533 1929
rect 6587 1883 6600 1929
rect 6520 1850 6600 1883
rect 6704 1929 6784 1942
rect 6704 1883 6717 1929
rect 6771 1883 6784 1929
rect 6704 1850 6784 1883
rect 6888 1929 6968 1942
rect 6888 1883 6901 1929
rect 6955 1883 6968 1929
rect 6888 1850 6968 1883
rect 6520 1617 6600 1650
rect 6520 1571 6533 1617
rect 6587 1571 6600 1617
rect 6520 1558 6600 1571
rect 6704 1617 6784 1650
rect 6704 1571 6717 1617
rect 6771 1571 6784 1617
rect 6704 1558 6784 1571
rect 6888 1617 6968 1650
rect 6888 1571 6901 1617
rect 6955 1571 6968 1617
rect 6888 1558 6968 1571
rect 9956 2759 10056 2772
rect 9956 2713 9969 2759
rect 10043 2713 10056 2759
rect 9956 2680 10056 2713
rect 9956 2047 10056 2080
rect 9956 2001 9969 2047
rect 10043 2001 10056 2047
rect 9956 1988 10056 2001
rect 10850 3059 10950 3072
rect 10850 3013 10863 3059
rect 10937 3013 10950 3059
rect 10850 2980 10950 3013
rect 11054 3059 11154 3072
rect 11054 3013 11067 3059
rect 11141 3013 11154 3059
rect 11054 2980 11154 3013
rect 10850 2747 10950 2780
rect 10850 2701 10863 2747
rect 10937 2701 10950 2747
rect 10850 2688 10950 2701
rect 11054 2747 11154 2780
rect 11054 2701 11067 2747
rect 11141 2701 11154 2747
rect 11054 2688 11154 2701
rect 11534 3059 11634 3072
rect 11534 3013 11547 3059
rect 11621 3013 11634 3059
rect 11534 2980 11634 3013
rect 11738 3059 11838 3072
rect 11738 3013 11751 3059
rect 11825 3013 11838 3059
rect 11738 2980 11838 3013
rect 11534 2747 11634 2780
rect 11534 2701 11547 2747
rect 11621 2701 11634 2747
rect 11534 2688 11634 2701
rect 11738 2747 11838 2780
rect 11738 2701 11751 2747
rect 11825 2701 11838 2747
rect 11738 2688 11838 2701
rect 12218 3059 12318 3072
rect 12218 3013 12231 3059
rect 12305 3013 12318 3059
rect 12218 2980 12318 3013
rect 12218 2747 12318 2780
rect 12218 2701 12231 2747
rect 12305 2701 12318 2747
rect 12218 2688 12318 2701
rect 13078 3003 13178 3016
rect 13078 2957 13091 3003
rect 13165 2957 13178 3003
rect 13078 2924 13178 2957
rect 13282 3003 13382 3016
rect 13282 2957 13295 3003
rect 13369 2957 13382 3003
rect 13282 2924 13382 2957
rect 13078 2291 13178 2324
rect 13078 2245 13091 2291
rect 13165 2245 13178 2291
rect 13078 2232 13178 2245
rect 13282 2291 13382 2324
rect 13282 2245 13295 2291
rect 13369 2245 13382 2291
rect 13282 2232 13382 2245
rect 13762 3003 13862 3016
rect 13762 2957 13775 3003
rect 13849 2957 13862 3003
rect 13762 2924 13862 2957
rect 13966 3003 14066 3016
rect 13966 2957 13979 3003
rect 14053 2957 14066 3003
rect 13966 2924 14066 2957
rect 13762 2291 13862 2324
rect 13762 2245 13775 2291
rect 13849 2245 13862 2291
rect 13762 2232 13862 2245
rect 13966 2291 14066 2324
rect 13966 2245 13979 2291
rect 14053 2245 14066 2291
rect 13966 2232 14066 2245
rect 14446 3003 14546 3016
rect 14446 2957 14459 3003
rect 14533 2957 14546 3003
rect 14446 2924 14546 2957
rect 14446 2291 14546 2324
rect 14446 2245 14459 2291
rect 14533 2245 14546 2291
rect 14446 2232 14546 2245
rect 15992 3089 16072 3102
rect 15992 3043 16005 3089
rect 16059 3043 16072 3089
rect 15992 3010 16072 3043
rect 16176 3089 16256 3102
rect 16176 3043 16189 3089
rect 16243 3043 16256 3089
rect 16176 3010 16256 3043
rect 16360 3089 16440 3102
rect 16360 3043 16373 3089
rect 16427 3043 16440 3089
rect 16360 3010 16440 3043
rect 15992 2477 16072 2510
rect 15992 2431 16005 2477
rect 16059 2431 16072 2477
rect 15992 2418 16072 2431
rect 16176 2477 16256 2510
rect 16176 2431 16189 2477
rect 16243 2431 16256 2477
rect 16176 2418 16256 2431
rect 16360 2477 16440 2510
rect 16360 2431 16373 2477
rect 16427 2431 16440 2477
rect 16360 2418 16440 2431
rect 9956 1639 10056 1652
rect 9956 1593 9969 1639
rect 10043 1593 10056 1639
rect 9956 1560 10056 1593
rect 9956 1327 10056 1360
rect 9956 1281 9969 1327
rect 10043 1281 10056 1327
rect 9956 1268 10056 1281
rect 10850 1839 10950 1852
rect 10850 1793 10863 1839
rect 10937 1793 10950 1839
rect 10850 1760 10950 1793
rect 10850 1127 10950 1160
rect 10850 1081 10863 1127
rect 10937 1081 10950 1127
rect 10850 1068 10950 1081
rect 11738 1839 11838 1852
rect 11738 1793 11751 1839
rect 11825 1793 11838 1839
rect 11738 1760 11838 1793
rect 11738 1127 11838 1160
rect 11738 1081 11751 1127
rect 11825 1081 11838 1127
rect 11738 1068 11838 1081
rect 12218 1839 12318 1852
rect 12218 1793 12231 1839
rect 12305 1793 12318 1839
rect 12218 1760 12318 1793
rect 12218 1127 12318 1160
rect 12218 1081 12231 1127
rect 12305 1081 12318 1127
rect 12218 1068 12318 1081
rect 13078 1883 13178 1896
rect 13078 1837 13091 1883
rect 13165 1837 13178 1883
rect 13078 1804 13178 1837
rect 13078 1571 13178 1604
rect 13078 1525 13091 1571
rect 13165 1525 13178 1571
rect 13078 1512 13178 1525
rect 13762 1883 13862 1896
rect 13762 1837 13775 1883
rect 13849 1837 13862 1883
rect 13762 1804 13862 1837
rect 13762 1571 13862 1604
rect 13762 1525 13775 1571
rect 13849 1525 13862 1571
rect 13762 1512 13862 1525
rect 14446 1883 14546 1896
rect 14446 1837 14459 1883
rect 14533 1837 14546 1883
rect 14446 1804 14546 1837
rect 14446 1571 14546 1604
rect 14446 1525 14459 1571
rect 14533 1525 14546 1571
rect 14446 1512 14546 1525
rect 15992 1929 16072 1942
rect 15992 1883 16005 1929
rect 16059 1883 16072 1929
rect 15992 1850 16072 1883
rect 16176 1929 16256 1942
rect 16176 1883 16189 1929
rect 16243 1883 16256 1929
rect 16176 1850 16256 1883
rect 16360 1929 16440 1942
rect 16360 1883 16373 1929
rect 16427 1883 16440 1929
rect 16360 1850 16440 1883
rect 15992 1617 16072 1650
rect 15992 1571 16005 1617
rect 16059 1571 16072 1617
rect 15992 1558 16072 1571
rect 16176 1617 16256 1650
rect 16176 1571 16189 1617
rect 16243 1571 16256 1617
rect 16176 1558 16256 1571
rect 16360 1617 16440 1650
rect 16360 1571 16373 1617
rect 16427 1571 16440 1617
rect 16360 1558 16440 1571
rect 19428 2760 19528 2773
rect 19428 2714 19441 2760
rect 19515 2714 19528 2760
rect 19428 2681 19528 2714
rect 19428 2048 19528 2081
rect 19428 2002 19441 2048
rect 19515 2002 19528 2048
rect 19428 1989 19528 2002
rect 20322 3060 20422 3073
rect 20322 3014 20335 3060
rect 20409 3014 20422 3060
rect 20322 2981 20422 3014
rect 20526 3060 20626 3073
rect 20526 3014 20539 3060
rect 20613 3014 20626 3060
rect 20526 2981 20626 3014
rect 20322 2748 20422 2781
rect 20322 2702 20335 2748
rect 20409 2702 20422 2748
rect 20322 2689 20422 2702
rect 20526 2748 20626 2781
rect 20526 2702 20539 2748
rect 20613 2702 20626 2748
rect 20526 2689 20626 2702
rect 21006 3060 21106 3073
rect 21006 3014 21019 3060
rect 21093 3014 21106 3060
rect 21006 2981 21106 3014
rect 21210 3060 21310 3073
rect 21210 3014 21223 3060
rect 21297 3014 21310 3060
rect 21210 2981 21310 3014
rect 21006 2748 21106 2781
rect 21006 2702 21019 2748
rect 21093 2702 21106 2748
rect 21006 2689 21106 2702
rect 21210 2748 21310 2781
rect 21210 2702 21223 2748
rect 21297 2702 21310 2748
rect 21210 2689 21310 2702
rect 21690 3060 21790 3073
rect 21690 3014 21703 3060
rect 21777 3014 21790 3060
rect 21690 2981 21790 3014
rect 21690 2748 21790 2781
rect 21690 2702 21703 2748
rect 21777 2702 21790 2748
rect 21690 2689 21790 2702
rect 22550 3004 22650 3017
rect 22550 2958 22563 3004
rect 22637 2958 22650 3004
rect 22550 2925 22650 2958
rect 22754 3004 22854 3017
rect 22754 2958 22767 3004
rect 22841 2958 22854 3004
rect 22754 2925 22854 2958
rect 22550 2292 22650 2325
rect 22550 2246 22563 2292
rect 22637 2246 22650 2292
rect 22550 2233 22650 2246
rect 22754 2292 22854 2325
rect 22754 2246 22767 2292
rect 22841 2246 22854 2292
rect 22754 2233 22854 2246
rect 23234 3004 23334 3017
rect 23234 2958 23247 3004
rect 23321 2958 23334 3004
rect 23234 2925 23334 2958
rect 23438 3004 23538 3017
rect 23438 2958 23451 3004
rect 23525 2958 23538 3004
rect 23438 2925 23538 2958
rect 23234 2292 23334 2325
rect 23234 2246 23247 2292
rect 23321 2246 23334 2292
rect 23234 2233 23334 2246
rect 23438 2292 23538 2325
rect 23438 2246 23451 2292
rect 23525 2246 23538 2292
rect 23438 2233 23538 2246
rect 23918 3004 24018 3017
rect 23918 2958 23931 3004
rect 24005 2958 24018 3004
rect 23918 2925 24018 2958
rect 23918 2292 24018 2325
rect 23918 2246 23931 2292
rect 24005 2246 24018 2292
rect 23918 2233 24018 2246
rect 25464 3090 25544 3103
rect 25464 3044 25477 3090
rect 25531 3044 25544 3090
rect 25464 3011 25544 3044
rect 25648 3090 25728 3103
rect 25648 3044 25661 3090
rect 25715 3044 25728 3090
rect 25648 3011 25728 3044
rect 25832 3090 25912 3103
rect 25832 3044 25845 3090
rect 25899 3044 25912 3090
rect 25832 3011 25912 3044
rect 25464 2478 25544 2511
rect 25464 2432 25477 2478
rect 25531 2432 25544 2478
rect 25464 2419 25544 2432
rect 25648 2478 25728 2511
rect 25648 2432 25661 2478
rect 25715 2432 25728 2478
rect 25648 2419 25728 2432
rect 25832 2478 25912 2511
rect 25832 2432 25845 2478
rect 25899 2432 25912 2478
rect 25832 2419 25912 2432
rect 19428 1640 19528 1653
rect 19428 1594 19441 1640
rect 19515 1594 19528 1640
rect 19428 1561 19528 1594
rect 19428 1328 19528 1361
rect 19428 1282 19441 1328
rect 19515 1282 19528 1328
rect 19428 1269 19528 1282
rect 20322 1840 20422 1853
rect 20322 1794 20335 1840
rect 20409 1794 20422 1840
rect 20322 1761 20422 1794
rect 20322 1128 20422 1161
rect 20322 1082 20335 1128
rect 20409 1082 20422 1128
rect 20322 1069 20422 1082
rect 21210 1840 21310 1853
rect 21210 1794 21223 1840
rect 21297 1794 21310 1840
rect 21210 1761 21310 1794
rect 21210 1128 21310 1161
rect 21210 1082 21223 1128
rect 21297 1082 21310 1128
rect 21210 1069 21310 1082
rect 21690 1840 21790 1853
rect 21690 1794 21703 1840
rect 21777 1794 21790 1840
rect 21690 1761 21790 1794
rect 21690 1128 21790 1161
rect 21690 1082 21703 1128
rect 21777 1082 21790 1128
rect 21690 1069 21790 1082
rect 22550 1884 22650 1897
rect 22550 1838 22563 1884
rect 22637 1838 22650 1884
rect 22550 1805 22650 1838
rect 22550 1572 22650 1605
rect 22550 1526 22563 1572
rect 22637 1526 22650 1572
rect 22550 1513 22650 1526
rect 23234 1884 23334 1897
rect 23234 1838 23247 1884
rect 23321 1838 23334 1884
rect 23234 1805 23334 1838
rect 23234 1572 23334 1605
rect 23234 1526 23247 1572
rect 23321 1526 23334 1572
rect 23234 1513 23334 1526
rect 23918 1884 24018 1897
rect 23918 1838 23931 1884
rect 24005 1838 24018 1884
rect 23918 1805 24018 1838
rect 23918 1572 24018 1605
rect 23918 1526 23931 1572
rect 24005 1526 24018 1572
rect 23918 1513 24018 1526
rect 25464 1930 25544 1943
rect 25464 1884 25477 1930
rect 25531 1884 25544 1930
rect 25464 1851 25544 1884
rect 25648 1930 25728 1943
rect 25648 1884 25661 1930
rect 25715 1884 25728 1930
rect 25648 1851 25728 1884
rect 25832 1930 25912 1943
rect 25832 1884 25845 1930
rect 25899 1884 25912 1930
rect 25832 1851 25912 1884
rect 25464 1618 25544 1651
rect 25464 1572 25477 1618
rect 25531 1572 25544 1618
rect 25464 1559 25544 1572
rect 25648 1618 25728 1651
rect 25648 1572 25661 1618
rect 25715 1572 25728 1618
rect 25648 1559 25728 1572
rect 25832 1618 25912 1651
rect 25832 1572 25845 1618
rect 25899 1572 25912 1618
rect 25832 1559 25912 1572
rect 28900 2760 29000 2773
rect 28900 2714 28913 2760
rect 28987 2714 29000 2760
rect 28900 2681 29000 2714
rect 28900 2048 29000 2081
rect 28900 2002 28913 2048
rect 28987 2002 29000 2048
rect 28900 1989 29000 2002
rect 29794 3060 29894 3073
rect 29794 3014 29807 3060
rect 29881 3014 29894 3060
rect 29794 2981 29894 3014
rect 29998 3060 30098 3073
rect 29998 3014 30011 3060
rect 30085 3014 30098 3060
rect 29998 2981 30098 3014
rect 29794 2748 29894 2781
rect 29794 2702 29807 2748
rect 29881 2702 29894 2748
rect 29794 2689 29894 2702
rect 29998 2748 30098 2781
rect 29998 2702 30011 2748
rect 30085 2702 30098 2748
rect 29998 2689 30098 2702
rect 30478 3060 30578 3073
rect 30478 3014 30491 3060
rect 30565 3014 30578 3060
rect 30478 2981 30578 3014
rect 30682 3060 30782 3073
rect 30682 3014 30695 3060
rect 30769 3014 30782 3060
rect 30682 2981 30782 3014
rect 30478 2748 30578 2781
rect 30478 2702 30491 2748
rect 30565 2702 30578 2748
rect 30478 2689 30578 2702
rect 30682 2748 30782 2781
rect 30682 2702 30695 2748
rect 30769 2702 30782 2748
rect 30682 2689 30782 2702
rect 31162 3060 31262 3073
rect 31162 3014 31175 3060
rect 31249 3014 31262 3060
rect 31162 2981 31262 3014
rect 31162 2748 31262 2781
rect 31162 2702 31175 2748
rect 31249 2702 31262 2748
rect 31162 2689 31262 2702
rect 32022 3004 32122 3017
rect 32022 2958 32035 3004
rect 32109 2958 32122 3004
rect 32022 2925 32122 2958
rect 32226 3004 32326 3017
rect 32226 2958 32239 3004
rect 32313 2958 32326 3004
rect 32226 2925 32326 2958
rect 32022 2292 32122 2325
rect 32022 2246 32035 2292
rect 32109 2246 32122 2292
rect 32022 2233 32122 2246
rect 32226 2292 32326 2325
rect 32226 2246 32239 2292
rect 32313 2246 32326 2292
rect 32226 2233 32326 2246
rect 32706 3004 32806 3017
rect 32706 2958 32719 3004
rect 32793 2958 32806 3004
rect 32706 2925 32806 2958
rect 32910 3004 33010 3017
rect 32910 2958 32923 3004
rect 32997 2958 33010 3004
rect 32910 2925 33010 2958
rect 32706 2292 32806 2325
rect 32706 2246 32719 2292
rect 32793 2246 32806 2292
rect 32706 2233 32806 2246
rect 32910 2292 33010 2325
rect 32910 2246 32923 2292
rect 32997 2246 33010 2292
rect 32910 2233 33010 2246
rect 33390 3004 33490 3017
rect 33390 2958 33403 3004
rect 33477 2958 33490 3004
rect 33390 2925 33490 2958
rect 33390 2292 33490 2325
rect 33390 2246 33403 2292
rect 33477 2246 33490 2292
rect 33390 2233 33490 2246
rect 34936 3090 35016 3103
rect 34936 3044 34949 3090
rect 35003 3044 35016 3090
rect 34936 3011 35016 3044
rect 35120 3090 35200 3103
rect 35120 3044 35133 3090
rect 35187 3044 35200 3090
rect 35120 3011 35200 3044
rect 35304 3090 35384 3103
rect 35304 3044 35317 3090
rect 35371 3044 35384 3090
rect 35304 3011 35384 3044
rect 34936 2478 35016 2511
rect 34936 2432 34949 2478
rect 35003 2432 35016 2478
rect 34936 2419 35016 2432
rect 35120 2478 35200 2511
rect 35120 2432 35133 2478
rect 35187 2432 35200 2478
rect 35120 2419 35200 2432
rect 35304 2478 35384 2511
rect 35304 2432 35317 2478
rect 35371 2432 35384 2478
rect 35304 2419 35384 2432
rect 28900 1640 29000 1653
rect 28900 1594 28913 1640
rect 28987 1594 29000 1640
rect 28900 1561 29000 1594
rect 28900 1328 29000 1361
rect 28900 1282 28913 1328
rect 28987 1282 29000 1328
rect 28900 1269 29000 1282
rect 29794 1840 29894 1853
rect 29794 1794 29807 1840
rect 29881 1794 29894 1840
rect 29794 1761 29894 1794
rect 29794 1128 29894 1161
rect 29794 1082 29807 1128
rect 29881 1082 29894 1128
rect 29794 1069 29894 1082
rect 30682 1840 30782 1853
rect 30682 1794 30695 1840
rect 30769 1794 30782 1840
rect 30682 1761 30782 1794
rect 30682 1128 30782 1161
rect 30682 1082 30695 1128
rect 30769 1082 30782 1128
rect 30682 1069 30782 1082
rect 31162 1840 31262 1853
rect 31162 1794 31175 1840
rect 31249 1794 31262 1840
rect 31162 1761 31262 1794
rect 31162 1128 31262 1161
rect 31162 1082 31175 1128
rect 31249 1082 31262 1128
rect 31162 1069 31262 1082
rect 32022 1884 32122 1897
rect 32022 1838 32035 1884
rect 32109 1838 32122 1884
rect 32022 1805 32122 1838
rect 32022 1572 32122 1605
rect 32022 1526 32035 1572
rect 32109 1526 32122 1572
rect 32022 1513 32122 1526
rect 32706 1884 32806 1897
rect 32706 1838 32719 1884
rect 32793 1838 32806 1884
rect 32706 1805 32806 1838
rect 32706 1572 32806 1605
rect 32706 1526 32719 1572
rect 32793 1526 32806 1572
rect 32706 1513 32806 1526
rect 33390 1884 33490 1897
rect 33390 1838 33403 1884
rect 33477 1838 33490 1884
rect 33390 1805 33490 1838
rect 33390 1572 33490 1605
rect 33390 1526 33403 1572
rect 33477 1526 33490 1572
rect 33390 1513 33490 1526
rect 34936 1930 35016 1943
rect 34936 1884 34949 1930
rect 35003 1884 35016 1930
rect 34936 1851 35016 1884
rect 35120 1930 35200 1943
rect 35120 1884 35133 1930
rect 35187 1884 35200 1930
rect 35120 1851 35200 1884
rect 35304 1930 35384 1943
rect 35304 1884 35317 1930
rect 35371 1884 35384 1930
rect 35304 1851 35384 1884
rect 34936 1618 35016 1651
rect 34936 1572 34949 1618
rect 35003 1572 35016 1618
rect 34936 1559 35016 1572
rect 35120 1618 35200 1651
rect 35120 1572 35133 1618
rect 35187 1572 35200 1618
rect 35120 1559 35200 1572
rect 35304 1618 35384 1651
rect 35304 1572 35317 1618
rect 35371 1572 35384 1618
rect 35304 1559 35384 1572
rect 38372 2760 38472 2773
rect 38372 2714 38385 2760
rect 38459 2714 38472 2760
rect 38372 2681 38472 2714
rect 38372 2048 38472 2081
rect 38372 2002 38385 2048
rect 38459 2002 38472 2048
rect 38372 1989 38472 2002
rect 39266 3060 39366 3073
rect 39266 3014 39279 3060
rect 39353 3014 39366 3060
rect 39266 2981 39366 3014
rect 39470 3060 39570 3073
rect 39470 3014 39483 3060
rect 39557 3014 39570 3060
rect 39470 2981 39570 3014
rect 39266 2748 39366 2781
rect 39266 2702 39279 2748
rect 39353 2702 39366 2748
rect 39266 2689 39366 2702
rect 39470 2748 39570 2781
rect 39470 2702 39483 2748
rect 39557 2702 39570 2748
rect 39470 2689 39570 2702
rect 39950 3060 40050 3073
rect 39950 3014 39963 3060
rect 40037 3014 40050 3060
rect 39950 2981 40050 3014
rect 40154 3060 40254 3073
rect 40154 3014 40167 3060
rect 40241 3014 40254 3060
rect 40154 2981 40254 3014
rect 39950 2748 40050 2781
rect 39950 2702 39963 2748
rect 40037 2702 40050 2748
rect 39950 2689 40050 2702
rect 40154 2748 40254 2781
rect 40154 2702 40167 2748
rect 40241 2702 40254 2748
rect 40154 2689 40254 2702
rect 40634 3060 40734 3073
rect 40634 3014 40647 3060
rect 40721 3014 40734 3060
rect 40634 2981 40734 3014
rect 40634 2748 40734 2781
rect 40634 2702 40647 2748
rect 40721 2702 40734 2748
rect 40634 2689 40734 2702
rect 41494 3004 41594 3017
rect 41494 2958 41507 3004
rect 41581 2958 41594 3004
rect 41494 2925 41594 2958
rect 41698 3004 41798 3017
rect 41698 2958 41711 3004
rect 41785 2958 41798 3004
rect 41698 2925 41798 2958
rect 41494 2292 41594 2325
rect 41494 2246 41507 2292
rect 41581 2246 41594 2292
rect 41494 2233 41594 2246
rect 41698 2292 41798 2325
rect 41698 2246 41711 2292
rect 41785 2246 41798 2292
rect 41698 2233 41798 2246
rect 42178 3004 42278 3017
rect 42178 2958 42191 3004
rect 42265 2958 42278 3004
rect 42178 2925 42278 2958
rect 42382 3004 42482 3017
rect 42382 2958 42395 3004
rect 42469 2958 42482 3004
rect 42382 2925 42482 2958
rect 42178 2292 42278 2325
rect 42178 2246 42191 2292
rect 42265 2246 42278 2292
rect 42178 2233 42278 2246
rect 42382 2292 42482 2325
rect 42382 2246 42395 2292
rect 42469 2246 42482 2292
rect 42382 2233 42482 2246
rect 42862 3004 42962 3017
rect 42862 2958 42875 3004
rect 42949 2958 42962 3004
rect 42862 2925 42962 2958
rect 42862 2292 42962 2325
rect 42862 2246 42875 2292
rect 42949 2246 42962 2292
rect 42862 2233 42962 2246
rect 44408 3090 44488 3103
rect 44408 3044 44421 3090
rect 44475 3044 44488 3090
rect 44408 3011 44488 3044
rect 44592 3090 44672 3103
rect 44592 3044 44605 3090
rect 44659 3044 44672 3090
rect 44592 3011 44672 3044
rect 44776 3090 44856 3103
rect 44776 3044 44789 3090
rect 44843 3044 44856 3090
rect 44776 3011 44856 3044
rect 44408 2478 44488 2511
rect 44408 2432 44421 2478
rect 44475 2432 44488 2478
rect 44408 2419 44488 2432
rect 44592 2478 44672 2511
rect 44592 2432 44605 2478
rect 44659 2432 44672 2478
rect 44592 2419 44672 2432
rect 44776 2478 44856 2511
rect 44776 2432 44789 2478
rect 44843 2432 44856 2478
rect 44776 2419 44856 2432
rect 38372 1640 38472 1653
rect 38372 1594 38385 1640
rect 38459 1594 38472 1640
rect 38372 1561 38472 1594
rect 38372 1328 38472 1361
rect 38372 1282 38385 1328
rect 38459 1282 38472 1328
rect 38372 1269 38472 1282
rect 39266 1840 39366 1853
rect 39266 1794 39279 1840
rect 39353 1794 39366 1840
rect 39266 1761 39366 1794
rect 39266 1128 39366 1161
rect 39266 1082 39279 1128
rect 39353 1082 39366 1128
rect 39266 1069 39366 1082
rect 40154 1840 40254 1853
rect 40154 1794 40167 1840
rect 40241 1794 40254 1840
rect 40154 1761 40254 1794
rect 40154 1128 40254 1161
rect 40154 1082 40167 1128
rect 40241 1082 40254 1128
rect 40154 1069 40254 1082
rect 40634 1840 40734 1853
rect 40634 1794 40647 1840
rect 40721 1794 40734 1840
rect 40634 1761 40734 1794
rect 40634 1128 40734 1161
rect 40634 1082 40647 1128
rect 40721 1082 40734 1128
rect 40634 1069 40734 1082
rect 41494 1884 41594 1897
rect 41494 1838 41507 1884
rect 41581 1838 41594 1884
rect 41494 1805 41594 1838
rect 41494 1572 41594 1605
rect 41494 1526 41507 1572
rect 41581 1526 41594 1572
rect 41494 1513 41594 1526
rect 42178 1884 42278 1897
rect 42178 1838 42191 1884
rect 42265 1838 42278 1884
rect 42178 1805 42278 1838
rect 42178 1572 42278 1605
rect 42178 1526 42191 1572
rect 42265 1526 42278 1572
rect 42178 1513 42278 1526
rect 42862 1884 42962 1897
rect 42862 1838 42875 1884
rect 42949 1838 42962 1884
rect 42862 1805 42962 1838
rect 42862 1572 42962 1605
rect 42862 1526 42875 1572
rect 42949 1526 42962 1572
rect 42862 1513 42962 1526
rect 44408 1930 44488 1943
rect 44408 1884 44421 1930
rect 44475 1884 44488 1930
rect 44408 1851 44488 1884
rect 44592 1930 44672 1943
rect 44592 1884 44605 1930
rect 44659 1884 44672 1930
rect 44592 1851 44672 1884
rect 44776 1930 44856 1943
rect 44776 1884 44789 1930
rect 44843 1884 44856 1930
rect 44776 1851 44856 1884
rect 44408 1618 44488 1651
rect 44408 1572 44421 1618
rect 44475 1572 44488 1618
rect 44408 1559 44488 1572
rect 44592 1618 44672 1651
rect 44592 1572 44605 1618
rect 44659 1572 44672 1618
rect 44592 1559 44672 1572
rect 44776 1618 44856 1651
rect 44776 1572 44789 1618
rect 44843 1572 44856 1618
rect 44776 1559 44856 1572
rect 47844 2760 47944 2773
rect 47844 2714 47857 2760
rect 47931 2714 47944 2760
rect 47844 2681 47944 2714
rect 47844 2048 47944 2081
rect 47844 2002 47857 2048
rect 47931 2002 47944 2048
rect 47844 1989 47944 2002
rect 48738 3060 48838 3073
rect 48738 3014 48751 3060
rect 48825 3014 48838 3060
rect 48738 2981 48838 3014
rect 48942 3060 49042 3073
rect 48942 3014 48955 3060
rect 49029 3014 49042 3060
rect 48942 2981 49042 3014
rect 48738 2748 48838 2781
rect 48738 2702 48751 2748
rect 48825 2702 48838 2748
rect 48738 2689 48838 2702
rect 48942 2748 49042 2781
rect 48942 2702 48955 2748
rect 49029 2702 49042 2748
rect 48942 2689 49042 2702
rect 49422 3060 49522 3073
rect 49422 3014 49435 3060
rect 49509 3014 49522 3060
rect 49422 2981 49522 3014
rect 49626 3060 49726 3073
rect 49626 3014 49639 3060
rect 49713 3014 49726 3060
rect 49626 2981 49726 3014
rect 49422 2748 49522 2781
rect 49422 2702 49435 2748
rect 49509 2702 49522 2748
rect 49422 2689 49522 2702
rect 49626 2748 49726 2781
rect 49626 2702 49639 2748
rect 49713 2702 49726 2748
rect 49626 2689 49726 2702
rect 50106 3060 50206 3073
rect 50106 3014 50119 3060
rect 50193 3014 50206 3060
rect 50106 2981 50206 3014
rect 50106 2748 50206 2781
rect 50106 2702 50119 2748
rect 50193 2702 50206 2748
rect 50106 2689 50206 2702
rect 50966 3004 51066 3017
rect 50966 2958 50979 3004
rect 51053 2958 51066 3004
rect 50966 2925 51066 2958
rect 51170 3004 51270 3017
rect 51170 2958 51183 3004
rect 51257 2958 51270 3004
rect 51170 2925 51270 2958
rect 50966 2292 51066 2325
rect 50966 2246 50979 2292
rect 51053 2246 51066 2292
rect 50966 2233 51066 2246
rect 51170 2292 51270 2325
rect 51170 2246 51183 2292
rect 51257 2246 51270 2292
rect 51170 2233 51270 2246
rect 51650 3004 51750 3017
rect 51650 2958 51663 3004
rect 51737 2958 51750 3004
rect 51650 2925 51750 2958
rect 51854 3004 51954 3017
rect 51854 2958 51867 3004
rect 51941 2958 51954 3004
rect 51854 2925 51954 2958
rect 51650 2292 51750 2325
rect 51650 2246 51663 2292
rect 51737 2246 51750 2292
rect 51650 2233 51750 2246
rect 51854 2292 51954 2325
rect 51854 2246 51867 2292
rect 51941 2246 51954 2292
rect 51854 2233 51954 2246
rect 52334 3004 52434 3017
rect 52334 2958 52347 3004
rect 52421 2958 52434 3004
rect 52334 2925 52434 2958
rect 52334 2292 52434 2325
rect 52334 2246 52347 2292
rect 52421 2246 52434 2292
rect 52334 2233 52434 2246
rect 53880 3090 53960 3103
rect 53880 3044 53893 3090
rect 53947 3044 53960 3090
rect 53880 3011 53960 3044
rect 54064 3090 54144 3103
rect 54064 3044 54077 3090
rect 54131 3044 54144 3090
rect 54064 3011 54144 3044
rect 54248 3090 54328 3103
rect 54248 3044 54261 3090
rect 54315 3044 54328 3090
rect 54248 3011 54328 3044
rect 53880 2478 53960 2511
rect 53880 2432 53893 2478
rect 53947 2432 53960 2478
rect 53880 2419 53960 2432
rect 54064 2478 54144 2511
rect 54064 2432 54077 2478
rect 54131 2432 54144 2478
rect 54064 2419 54144 2432
rect 54248 2478 54328 2511
rect 54248 2432 54261 2478
rect 54315 2432 54328 2478
rect 54248 2419 54328 2432
rect 47844 1640 47944 1653
rect 47844 1594 47857 1640
rect 47931 1594 47944 1640
rect 47844 1561 47944 1594
rect 47844 1328 47944 1361
rect 47844 1282 47857 1328
rect 47931 1282 47944 1328
rect 47844 1269 47944 1282
rect 48738 1840 48838 1853
rect 48738 1794 48751 1840
rect 48825 1794 48838 1840
rect 48738 1761 48838 1794
rect 48738 1128 48838 1161
rect 48738 1082 48751 1128
rect 48825 1082 48838 1128
rect 48738 1069 48838 1082
rect 49626 1840 49726 1853
rect 49626 1794 49639 1840
rect 49713 1794 49726 1840
rect 49626 1761 49726 1794
rect 49626 1128 49726 1161
rect 49626 1082 49639 1128
rect 49713 1082 49726 1128
rect 49626 1069 49726 1082
rect 50106 1840 50206 1853
rect 50106 1794 50119 1840
rect 50193 1794 50206 1840
rect 50106 1761 50206 1794
rect 50106 1128 50206 1161
rect 50106 1082 50119 1128
rect 50193 1082 50206 1128
rect 50106 1069 50206 1082
rect 50966 1884 51066 1897
rect 50966 1838 50979 1884
rect 51053 1838 51066 1884
rect 50966 1805 51066 1838
rect 50966 1572 51066 1605
rect 50966 1526 50979 1572
rect 51053 1526 51066 1572
rect 50966 1513 51066 1526
rect 51650 1884 51750 1897
rect 51650 1838 51663 1884
rect 51737 1838 51750 1884
rect 51650 1805 51750 1838
rect 51650 1572 51750 1605
rect 51650 1526 51663 1572
rect 51737 1526 51750 1572
rect 51650 1513 51750 1526
rect 52334 1884 52434 1897
rect 52334 1838 52347 1884
rect 52421 1838 52434 1884
rect 52334 1805 52434 1838
rect 52334 1572 52434 1605
rect 52334 1526 52347 1572
rect 52421 1526 52434 1572
rect 52334 1513 52434 1526
rect 53880 1930 53960 1943
rect 53880 1884 53893 1930
rect 53947 1884 53960 1930
rect 53880 1851 53960 1884
rect 54064 1930 54144 1943
rect 54064 1884 54077 1930
rect 54131 1884 54144 1930
rect 54064 1851 54144 1884
rect 54248 1930 54328 1943
rect 54248 1884 54261 1930
rect 54315 1884 54328 1930
rect 54248 1851 54328 1884
rect 53880 1618 53960 1651
rect 53880 1572 53893 1618
rect 53947 1572 53960 1618
rect 53880 1559 53960 1572
rect 54064 1618 54144 1651
rect 54064 1572 54077 1618
rect 54131 1572 54144 1618
rect 54064 1559 54144 1572
rect 54248 1618 54328 1651
rect 54248 1572 54261 1618
rect 54315 1572 54328 1618
rect 54248 1559 54328 1572
rect 1378 719 1478 732
rect 1378 673 1391 719
rect 1465 673 1478 719
rect 1378 640 1478 673
rect 1582 719 1682 732
rect 1582 673 1595 719
rect 1669 673 1682 719
rect 1582 640 1682 673
rect 1378 407 1478 440
rect 1378 361 1391 407
rect 1465 361 1478 407
rect 1378 348 1478 361
rect 1582 407 1682 440
rect 1582 361 1595 407
rect 1669 361 1682 407
rect 1582 348 1682 361
rect 2062 719 2162 732
rect 2062 673 2075 719
rect 2149 673 2162 719
rect 2062 640 2162 673
rect 2266 719 2366 732
rect 2266 673 2279 719
rect 2353 673 2366 719
rect 2266 640 2366 673
rect 2062 407 2162 440
rect 2062 361 2075 407
rect 2149 361 2162 407
rect 2062 348 2162 361
rect 2266 407 2366 440
rect 2266 361 2279 407
rect 2353 361 2366 407
rect 2266 348 2366 361
rect 2746 719 2846 732
rect 2746 673 2759 719
rect 2833 673 2846 719
rect 2746 640 2846 673
rect 2746 407 2846 440
rect 2746 361 2759 407
rect 2833 361 2846 407
rect 2746 348 2846 361
rect 10850 719 10950 732
rect 10850 673 10863 719
rect 10937 673 10950 719
rect 10850 640 10950 673
rect 11054 719 11154 732
rect 11054 673 11067 719
rect 11141 673 11154 719
rect 11054 640 11154 673
rect 10850 407 10950 440
rect 10850 361 10863 407
rect 10937 361 10950 407
rect 10850 348 10950 361
rect 11054 407 11154 440
rect 11054 361 11067 407
rect 11141 361 11154 407
rect 11054 348 11154 361
rect 11534 719 11634 732
rect 11534 673 11547 719
rect 11621 673 11634 719
rect 11534 640 11634 673
rect 11738 719 11838 732
rect 11738 673 11751 719
rect 11825 673 11838 719
rect 11738 640 11838 673
rect 11534 407 11634 440
rect 11534 361 11547 407
rect 11621 361 11634 407
rect 11534 348 11634 361
rect 11738 407 11838 440
rect 11738 361 11751 407
rect 11825 361 11838 407
rect 11738 348 11838 361
rect 12218 719 12318 732
rect 12218 673 12231 719
rect 12305 673 12318 719
rect 12218 640 12318 673
rect 12218 407 12318 440
rect 12218 361 12231 407
rect 12305 361 12318 407
rect 12218 348 12318 361
rect 20322 720 20422 733
rect 20322 674 20335 720
rect 20409 674 20422 720
rect 20322 641 20422 674
rect 20526 720 20626 733
rect 20526 674 20539 720
rect 20613 674 20626 720
rect 20526 641 20626 674
rect 20322 408 20422 441
rect 20322 362 20335 408
rect 20409 362 20422 408
rect 20322 349 20422 362
rect 20526 408 20626 441
rect 20526 362 20539 408
rect 20613 362 20626 408
rect 20526 349 20626 362
rect 21006 720 21106 733
rect 21006 674 21019 720
rect 21093 674 21106 720
rect 21006 641 21106 674
rect 21210 720 21310 733
rect 21210 674 21223 720
rect 21297 674 21310 720
rect 21210 641 21310 674
rect 21006 408 21106 441
rect 21006 362 21019 408
rect 21093 362 21106 408
rect 21006 349 21106 362
rect 21210 408 21310 441
rect 21210 362 21223 408
rect 21297 362 21310 408
rect 21210 349 21310 362
rect 21690 720 21790 733
rect 21690 674 21703 720
rect 21777 674 21790 720
rect 21690 641 21790 674
rect 21690 408 21790 441
rect 21690 362 21703 408
rect 21777 362 21790 408
rect 21690 349 21790 362
rect 29794 720 29894 733
rect 29794 674 29807 720
rect 29881 674 29894 720
rect 29794 641 29894 674
rect 29998 720 30098 733
rect 29998 674 30011 720
rect 30085 674 30098 720
rect 29998 641 30098 674
rect 29794 408 29894 441
rect 29794 362 29807 408
rect 29881 362 29894 408
rect 29794 349 29894 362
rect 29998 408 30098 441
rect 29998 362 30011 408
rect 30085 362 30098 408
rect 29998 349 30098 362
rect 30478 720 30578 733
rect 30478 674 30491 720
rect 30565 674 30578 720
rect 30478 641 30578 674
rect 30682 720 30782 733
rect 30682 674 30695 720
rect 30769 674 30782 720
rect 30682 641 30782 674
rect 30478 408 30578 441
rect 30478 362 30491 408
rect 30565 362 30578 408
rect 30478 349 30578 362
rect 30682 408 30782 441
rect 30682 362 30695 408
rect 30769 362 30782 408
rect 30682 349 30782 362
rect 31162 720 31262 733
rect 31162 674 31175 720
rect 31249 674 31262 720
rect 31162 641 31262 674
rect 31162 408 31262 441
rect 31162 362 31175 408
rect 31249 362 31262 408
rect 31162 349 31262 362
rect 39266 720 39366 733
rect 39266 674 39279 720
rect 39353 674 39366 720
rect 39266 641 39366 674
rect 39470 720 39570 733
rect 39470 674 39483 720
rect 39557 674 39570 720
rect 39470 641 39570 674
rect 39266 408 39366 441
rect 39266 362 39279 408
rect 39353 362 39366 408
rect 39266 349 39366 362
rect 39470 408 39570 441
rect 39470 362 39483 408
rect 39557 362 39570 408
rect 39470 349 39570 362
rect 39950 720 40050 733
rect 39950 674 39963 720
rect 40037 674 40050 720
rect 39950 641 40050 674
rect 40154 720 40254 733
rect 40154 674 40167 720
rect 40241 674 40254 720
rect 40154 641 40254 674
rect 39950 408 40050 441
rect 39950 362 39963 408
rect 40037 362 40050 408
rect 39950 349 40050 362
rect 40154 408 40254 441
rect 40154 362 40167 408
rect 40241 362 40254 408
rect 40154 349 40254 362
rect 40634 720 40734 733
rect 40634 674 40647 720
rect 40721 674 40734 720
rect 40634 641 40734 674
rect 40634 408 40734 441
rect 40634 362 40647 408
rect 40721 362 40734 408
rect 40634 349 40734 362
rect 48738 720 48838 733
rect 48738 674 48751 720
rect 48825 674 48838 720
rect 48738 641 48838 674
rect 48942 720 49042 733
rect 48942 674 48955 720
rect 49029 674 49042 720
rect 48942 641 49042 674
rect 48738 408 48838 441
rect 48738 362 48751 408
rect 48825 362 48838 408
rect 48738 349 48838 362
rect 48942 408 49042 441
rect 48942 362 48955 408
rect 49029 362 49042 408
rect 48942 349 49042 362
rect 49422 720 49522 733
rect 49422 674 49435 720
rect 49509 674 49522 720
rect 49422 641 49522 674
rect 49626 720 49726 733
rect 49626 674 49639 720
rect 49713 674 49726 720
rect 49626 641 49726 674
rect 49422 408 49522 441
rect 49422 362 49435 408
rect 49509 362 49522 408
rect 49422 349 49522 362
rect 49626 408 49726 441
rect 49626 362 49639 408
rect 49713 362 49726 408
rect 49626 349 49726 362
rect 50106 720 50206 733
rect 50106 674 50119 720
rect 50193 674 50206 720
rect 50106 641 50206 674
rect 50106 408 50206 441
rect 50106 362 50119 408
rect 50193 362 50206 408
rect 50106 349 50206 362
<< polycontact >>
rect 6533 9658 6587 9704
rect 6717 9658 6771 9704
rect 6901 9658 6955 9704
rect 6533 9046 6587 9092
rect 6717 9046 6771 9092
rect 6901 9046 6955 9092
rect 16005 9658 16059 9704
rect 16189 9658 16243 9704
rect 16373 9658 16427 9704
rect 16005 9046 16059 9092
rect 16189 9046 16243 9092
rect 16373 9046 16427 9092
rect 25477 9659 25531 9705
rect 25661 9659 25715 9705
rect 25845 9659 25899 9705
rect 25477 9047 25531 9093
rect 25661 9047 25715 9093
rect 25845 9047 25899 9093
rect 34949 9659 35003 9705
rect 35133 9659 35187 9705
rect 35317 9659 35371 9705
rect 34949 9047 35003 9093
rect 35133 9047 35187 9093
rect 35317 9047 35371 9093
rect 44421 9659 44475 9705
rect 44605 9659 44659 9705
rect 44789 9659 44843 9705
rect 44421 9047 44475 9093
rect 44605 9047 44659 9093
rect 44789 9047 44843 9093
rect 53893 9659 53947 9705
rect 54077 9659 54131 9705
rect 54261 9659 54315 9705
rect 53893 9047 53947 9093
rect 54077 9047 54131 9093
rect 54261 9047 54315 9093
rect 6533 8498 6587 8544
rect 6717 8498 6771 8544
rect 6901 8498 6955 8544
rect 6533 8186 6587 8232
rect 6717 8186 6771 8232
rect 6901 8186 6955 8232
rect 16005 8498 16059 8544
rect 16189 8498 16243 8544
rect 16373 8498 16427 8544
rect 16005 8186 16059 8232
rect 16189 8186 16243 8232
rect 16373 8186 16427 8232
rect 25477 8499 25531 8545
rect 25661 8499 25715 8545
rect 25845 8499 25899 8545
rect 25477 8187 25531 8233
rect 25661 8187 25715 8233
rect 25845 8187 25899 8233
rect 34949 8499 35003 8545
rect 35133 8499 35187 8545
rect 35317 8499 35371 8545
rect 34949 8187 35003 8233
rect 35133 8187 35187 8233
rect 35317 8187 35371 8233
rect 44421 8499 44475 8545
rect 44605 8499 44659 8545
rect 44789 8499 44843 8545
rect 44421 8187 44475 8233
rect 44605 8187 44659 8233
rect 44789 8187 44843 8233
rect 53893 8499 53947 8545
rect 54077 8499 54131 8545
rect 54261 8499 54315 8545
rect 53893 8187 53947 8233
rect 54077 8187 54131 8233
rect 54261 8187 54315 8233
rect 6533 7453 6587 7499
rect 6717 7453 6771 7499
rect 6901 7453 6955 7499
rect 6533 6841 6587 6887
rect 6717 6841 6771 6887
rect 6901 6841 6955 6887
rect 8019 7453 8073 7499
rect 8203 7453 8257 7499
rect 8387 7453 8441 7499
rect 8019 6841 8073 6887
rect 8203 6841 8257 6887
rect 8387 6841 8441 6887
rect 16005 7453 16059 7499
rect 16189 7453 16243 7499
rect 16373 7453 16427 7499
rect 16005 6841 16059 6887
rect 16189 6841 16243 6887
rect 16373 6841 16427 6887
rect 17491 7453 17545 7499
rect 17675 7453 17729 7499
rect 17859 7453 17913 7499
rect 17491 6841 17545 6887
rect 17675 6841 17729 6887
rect 17859 6841 17913 6887
rect 25477 7454 25531 7500
rect 25661 7454 25715 7500
rect 25845 7454 25899 7500
rect 25477 6842 25531 6888
rect 25661 6842 25715 6888
rect 25845 6842 25899 6888
rect 26963 7454 27017 7500
rect 27147 7454 27201 7500
rect 27331 7454 27385 7500
rect 26963 6842 27017 6888
rect 27147 6842 27201 6888
rect 27331 6842 27385 6888
rect 34949 7454 35003 7500
rect 35133 7454 35187 7500
rect 35317 7454 35371 7500
rect 34949 6842 35003 6888
rect 35133 6842 35187 6888
rect 35317 6842 35371 6888
rect 36435 7454 36489 7500
rect 36619 7454 36673 7500
rect 36803 7454 36857 7500
rect 36435 6842 36489 6888
rect 36619 6842 36673 6888
rect 36803 6842 36857 6888
rect 44421 7454 44475 7500
rect 44605 7454 44659 7500
rect 44789 7454 44843 7500
rect 44421 6842 44475 6888
rect 44605 6842 44659 6888
rect 44789 6842 44843 6888
rect 45907 7454 45961 7500
rect 46091 7454 46145 7500
rect 46275 7454 46329 7500
rect 45907 6842 45961 6888
rect 46091 6842 46145 6888
rect 46275 6842 46329 6888
rect 53893 7454 53947 7500
rect 54077 7454 54131 7500
rect 54261 7454 54315 7500
rect 53893 6842 53947 6888
rect 54077 6842 54131 6888
rect 54261 6842 54315 6888
rect 55379 7454 55433 7500
rect 55563 7454 55617 7500
rect 55747 7454 55801 7500
rect 55379 6842 55433 6888
rect 55563 6842 55617 6888
rect 55747 6842 55801 6888
rect 6533 6293 6587 6339
rect 6717 6293 6771 6339
rect 6901 6293 6955 6339
rect 6533 5981 6587 6027
rect 6717 5981 6771 6027
rect 6901 5981 6955 6027
rect 8019 6293 8073 6339
rect 8203 6293 8257 6339
rect 8387 6293 8441 6339
rect 8019 5981 8073 6027
rect 8203 5981 8257 6027
rect 8387 5981 8441 6027
rect 16005 6293 16059 6339
rect 16189 6293 16243 6339
rect 16373 6293 16427 6339
rect 16005 5981 16059 6027
rect 16189 5981 16243 6027
rect 16373 5981 16427 6027
rect 17491 6293 17545 6339
rect 17675 6293 17729 6339
rect 17859 6293 17913 6339
rect 17491 5981 17545 6027
rect 17675 5981 17729 6027
rect 17859 5981 17913 6027
rect 25477 6294 25531 6340
rect 25661 6294 25715 6340
rect 25845 6294 25899 6340
rect 25477 5982 25531 6028
rect 25661 5982 25715 6028
rect 25845 5982 25899 6028
rect 26963 6294 27017 6340
rect 27147 6294 27201 6340
rect 27331 6294 27385 6340
rect 26963 5982 27017 6028
rect 27147 5982 27201 6028
rect 27331 5982 27385 6028
rect 34949 6294 35003 6340
rect 35133 6294 35187 6340
rect 35317 6294 35371 6340
rect 34949 5982 35003 6028
rect 35133 5982 35187 6028
rect 35317 5982 35371 6028
rect 36435 6294 36489 6340
rect 36619 6294 36673 6340
rect 36803 6294 36857 6340
rect 36435 5982 36489 6028
rect 36619 5982 36673 6028
rect 36803 5982 36857 6028
rect 44421 6294 44475 6340
rect 44605 6294 44659 6340
rect 44789 6294 44843 6340
rect 44421 5982 44475 6028
rect 44605 5982 44659 6028
rect 44789 5982 44843 6028
rect 45907 6294 45961 6340
rect 46091 6294 46145 6340
rect 46275 6294 46329 6340
rect 45907 5982 45961 6028
rect 46091 5982 46145 6028
rect 46275 5982 46329 6028
rect 53893 6294 53947 6340
rect 54077 6294 54131 6340
rect 54261 6294 54315 6340
rect 53893 5982 53947 6028
rect 54077 5982 54131 6028
rect 54261 5982 54315 6028
rect 55379 6294 55433 6340
rect 55563 6294 55617 6340
rect 55747 6294 55801 6340
rect 55379 5982 55433 6028
rect 55563 5982 55617 6028
rect 55747 5982 55801 6028
rect 6533 5248 6587 5294
rect 6717 5248 6771 5294
rect 6901 5248 6955 5294
rect 6533 4636 6587 4682
rect 6717 4636 6771 4682
rect 6901 4636 6955 4682
rect 8019 5249 8073 5295
rect 8203 5249 8257 5295
rect 8387 5249 8441 5295
rect 8019 4637 8073 4683
rect 8203 4637 8257 4683
rect 8387 4637 8441 4683
rect 16005 5248 16059 5294
rect 16189 5248 16243 5294
rect 16373 5248 16427 5294
rect 16005 4636 16059 4682
rect 16189 4636 16243 4682
rect 16373 4636 16427 4682
rect 17491 5249 17545 5295
rect 17675 5249 17729 5295
rect 17859 5249 17913 5295
rect 17491 4637 17545 4683
rect 17675 4637 17729 4683
rect 17859 4637 17913 4683
rect 25477 5249 25531 5295
rect 25661 5249 25715 5295
rect 25845 5249 25899 5295
rect 25477 4637 25531 4683
rect 25661 4637 25715 4683
rect 25845 4637 25899 4683
rect 26963 5250 27017 5296
rect 27147 5250 27201 5296
rect 27331 5250 27385 5296
rect 26963 4638 27017 4684
rect 27147 4638 27201 4684
rect 27331 4638 27385 4684
rect 34949 5249 35003 5295
rect 35133 5249 35187 5295
rect 35317 5249 35371 5295
rect 34949 4637 35003 4683
rect 35133 4637 35187 4683
rect 35317 4637 35371 4683
rect 36435 5250 36489 5296
rect 36619 5250 36673 5296
rect 36803 5250 36857 5296
rect 36435 4638 36489 4684
rect 36619 4638 36673 4684
rect 36803 4638 36857 4684
rect 44421 5249 44475 5295
rect 44605 5249 44659 5295
rect 44789 5249 44843 5295
rect 44421 4637 44475 4683
rect 44605 4637 44659 4683
rect 44789 4637 44843 4683
rect 45907 5250 45961 5296
rect 46091 5250 46145 5296
rect 46275 5250 46329 5296
rect 45907 4638 45961 4684
rect 46091 4638 46145 4684
rect 46275 4638 46329 4684
rect 53893 5249 53947 5295
rect 54077 5249 54131 5295
rect 54261 5249 54315 5295
rect 53893 4637 53947 4683
rect 54077 4637 54131 4683
rect 54261 4637 54315 4683
rect 55379 5250 55433 5296
rect 55563 5250 55617 5296
rect 55747 5250 55801 5296
rect 55379 4638 55433 4684
rect 55563 4638 55617 4684
rect 55747 4638 55801 4684
rect 1391 4133 1465 4179
rect 1391 3421 1465 3467
rect 2279 4133 2353 4179
rect 2279 3421 2353 3467
rect 2759 4133 2833 4179
rect 2759 3421 2833 3467
rect 6533 4088 6587 4134
rect 6717 4088 6771 4134
rect 6901 4088 6955 4134
rect 6533 3776 6587 3822
rect 6717 3776 6771 3822
rect 6901 3776 6955 3822
rect 8019 4089 8073 4135
rect 8203 4089 8257 4135
rect 8387 4089 8441 4135
rect 8019 3777 8073 3823
rect 8203 3777 8257 3823
rect 8387 3777 8441 3823
rect 10863 4133 10937 4179
rect 10863 3421 10937 3467
rect 11751 4133 11825 4179
rect 11751 3421 11825 3467
rect 12231 4133 12305 4179
rect 12231 3421 12305 3467
rect 16005 4088 16059 4134
rect 16189 4088 16243 4134
rect 16373 4088 16427 4134
rect 16005 3776 16059 3822
rect 16189 3776 16243 3822
rect 16373 3776 16427 3822
rect 17491 4089 17545 4135
rect 17675 4089 17729 4135
rect 17859 4089 17913 4135
rect 17491 3777 17545 3823
rect 17675 3777 17729 3823
rect 17859 3777 17913 3823
rect 20335 4134 20409 4180
rect 20335 3422 20409 3468
rect 21223 4134 21297 4180
rect 21223 3422 21297 3468
rect 21703 4134 21777 4180
rect 21703 3422 21777 3468
rect 25477 4089 25531 4135
rect 25661 4089 25715 4135
rect 25845 4089 25899 4135
rect 25477 3777 25531 3823
rect 25661 3777 25715 3823
rect 25845 3777 25899 3823
rect 26963 4090 27017 4136
rect 27147 4090 27201 4136
rect 27331 4090 27385 4136
rect 26963 3778 27017 3824
rect 27147 3778 27201 3824
rect 27331 3778 27385 3824
rect 29807 4134 29881 4180
rect 29807 3422 29881 3468
rect 30695 4134 30769 4180
rect 30695 3422 30769 3468
rect 31175 4134 31249 4180
rect 31175 3422 31249 3468
rect 34949 4089 35003 4135
rect 35133 4089 35187 4135
rect 35317 4089 35371 4135
rect 34949 3777 35003 3823
rect 35133 3777 35187 3823
rect 35317 3777 35371 3823
rect 36435 4090 36489 4136
rect 36619 4090 36673 4136
rect 36803 4090 36857 4136
rect 36435 3778 36489 3824
rect 36619 3778 36673 3824
rect 36803 3778 36857 3824
rect 39279 4134 39353 4180
rect 39279 3422 39353 3468
rect 40167 4134 40241 4180
rect 40167 3422 40241 3468
rect 40647 4134 40721 4180
rect 40647 3422 40721 3468
rect 44421 4089 44475 4135
rect 44605 4089 44659 4135
rect 44789 4089 44843 4135
rect 44421 3777 44475 3823
rect 44605 3777 44659 3823
rect 44789 3777 44843 3823
rect 45907 4090 45961 4136
rect 46091 4090 46145 4136
rect 46275 4090 46329 4136
rect 45907 3778 45961 3824
rect 46091 3778 46145 3824
rect 46275 3778 46329 3824
rect 48751 4134 48825 4180
rect 48751 3422 48825 3468
rect 49639 4134 49713 4180
rect 49639 3422 49713 3468
rect 50119 4134 50193 4180
rect 50119 3422 50193 3468
rect 53893 4089 53947 4135
rect 54077 4089 54131 4135
rect 54261 4089 54315 4135
rect 53893 3777 53947 3823
rect 54077 3777 54131 3823
rect 54261 3777 54315 3823
rect 55379 4090 55433 4136
rect 55563 4090 55617 4136
rect 55747 4090 55801 4136
rect 55379 3778 55433 3824
rect 55563 3778 55617 3824
rect 55747 3778 55801 3824
rect 497 2713 571 2759
rect 497 2001 571 2047
rect 1391 3013 1465 3059
rect 1595 3013 1669 3059
rect 1391 2701 1465 2747
rect 1595 2701 1669 2747
rect 2075 3013 2149 3059
rect 2279 3013 2353 3059
rect 2075 2701 2149 2747
rect 2279 2701 2353 2747
rect 2759 3013 2833 3059
rect 2759 2701 2833 2747
rect 3619 2957 3693 3003
rect 3823 2957 3897 3003
rect 3619 2245 3693 2291
rect 3823 2245 3897 2291
rect 4303 2957 4377 3003
rect 4507 2957 4581 3003
rect 4303 2245 4377 2291
rect 4507 2245 4581 2291
rect 4987 2957 5061 3003
rect 4987 2245 5061 2291
rect 6533 3043 6587 3089
rect 6717 3043 6771 3089
rect 6901 3043 6955 3089
rect 6533 2431 6587 2477
rect 6717 2431 6771 2477
rect 6901 2431 6955 2477
rect 497 1593 571 1639
rect 497 1281 571 1327
rect 1391 1793 1465 1839
rect 1391 1081 1465 1127
rect 2279 1793 2353 1839
rect 2279 1081 2353 1127
rect 2759 1793 2833 1839
rect 2759 1081 2833 1127
rect 3619 1837 3693 1883
rect 3619 1525 3693 1571
rect 4303 1837 4377 1883
rect 4303 1525 4377 1571
rect 4987 1837 5061 1883
rect 4987 1525 5061 1571
rect 6533 1883 6587 1929
rect 6717 1883 6771 1929
rect 6901 1883 6955 1929
rect 6533 1571 6587 1617
rect 6717 1571 6771 1617
rect 6901 1571 6955 1617
rect 9969 2713 10043 2759
rect 9969 2001 10043 2047
rect 10863 3013 10937 3059
rect 11067 3013 11141 3059
rect 10863 2701 10937 2747
rect 11067 2701 11141 2747
rect 11547 3013 11621 3059
rect 11751 3013 11825 3059
rect 11547 2701 11621 2747
rect 11751 2701 11825 2747
rect 12231 3013 12305 3059
rect 12231 2701 12305 2747
rect 13091 2957 13165 3003
rect 13295 2957 13369 3003
rect 13091 2245 13165 2291
rect 13295 2245 13369 2291
rect 13775 2957 13849 3003
rect 13979 2957 14053 3003
rect 13775 2245 13849 2291
rect 13979 2245 14053 2291
rect 14459 2957 14533 3003
rect 14459 2245 14533 2291
rect 16005 3043 16059 3089
rect 16189 3043 16243 3089
rect 16373 3043 16427 3089
rect 16005 2431 16059 2477
rect 16189 2431 16243 2477
rect 16373 2431 16427 2477
rect 9969 1593 10043 1639
rect 9969 1281 10043 1327
rect 10863 1793 10937 1839
rect 10863 1081 10937 1127
rect 11751 1793 11825 1839
rect 11751 1081 11825 1127
rect 12231 1793 12305 1839
rect 12231 1081 12305 1127
rect 13091 1837 13165 1883
rect 13091 1525 13165 1571
rect 13775 1837 13849 1883
rect 13775 1525 13849 1571
rect 14459 1837 14533 1883
rect 14459 1525 14533 1571
rect 16005 1883 16059 1929
rect 16189 1883 16243 1929
rect 16373 1883 16427 1929
rect 16005 1571 16059 1617
rect 16189 1571 16243 1617
rect 16373 1571 16427 1617
rect 19441 2714 19515 2760
rect 19441 2002 19515 2048
rect 20335 3014 20409 3060
rect 20539 3014 20613 3060
rect 20335 2702 20409 2748
rect 20539 2702 20613 2748
rect 21019 3014 21093 3060
rect 21223 3014 21297 3060
rect 21019 2702 21093 2748
rect 21223 2702 21297 2748
rect 21703 3014 21777 3060
rect 21703 2702 21777 2748
rect 22563 2958 22637 3004
rect 22767 2958 22841 3004
rect 22563 2246 22637 2292
rect 22767 2246 22841 2292
rect 23247 2958 23321 3004
rect 23451 2958 23525 3004
rect 23247 2246 23321 2292
rect 23451 2246 23525 2292
rect 23931 2958 24005 3004
rect 23931 2246 24005 2292
rect 25477 3044 25531 3090
rect 25661 3044 25715 3090
rect 25845 3044 25899 3090
rect 25477 2432 25531 2478
rect 25661 2432 25715 2478
rect 25845 2432 25899 2478
rect 19441 1594 19515 1640
rect 19441 1282 19515 1328
rect 20335 1794 20409 1840
rect 20335 1082 20409 1128
rect 21223 1794 21297 1840
rect 21223 1082 21297 1128
rect 21703 1794 21777 1840
rect 21703 1082 21777 1128
rect 22563 1838 22637 1884
rect 22563 1526 22637 1572
rect 23247 1838 23321 1884
rect 23247 1526 23321 1572
rect 23931 1838 24005 1884
rect 23931 1526 24005 1572
rect 25477 1884 25531 1930
rect 25661 1884 25715 1930
rect 25845 1884 25899 1930
rect 25477 1572 25531 1618
rect 25661 1572 25715 1618
rect 25845 1572 25899 1618
rect 28913 2714 28987 2760
rect 28913 2002 28987 2048
rect 29807 3014 29881 3060
rect 30011 3014 30085 3060
rect 29807 2702 29881 2748
rect 30011 2702 30085 2748
rect 30491 3014 30565 3060
rect 30695 3014 30769 3060
rect 30491 2702 30565 2748
rect 30695 2702 30769 2748
rect 31175 3014 31249 3060
rect 31175 2702 31249 2748
rect 32035 2958 32109 3004
rect 32239 2958 32313 3004
rect 32035 2246 32109 2292
rect 32239 2246 32313 2292
rect 32719 2958 32793 3004
rect 32923 2958 32997 3004
rect 32719 2246 32793 2292
rect 32923 2246 32997 2292
rect 33403 2958 33477 3004
rect 33403 2246 33477 2292
rect 34949 3044 35003 3090
rect 35133 3044 35187 3090
rect 35317 3044 35371 3090
rect 34949 2432 35003 2478
rect 35133 2432 35187 2478
rect 35317 2432 35371 2478
rect 28913 1594 28987 1640
rect 28913 1282 28987 1328
rect 29807 1794 29881 1840
rect 29807 1082 29881 1128
rect 30695 1794 30769 1840
rect 30695 1082 30769 1128
rect 31175 1794 31249 1840
rect 31175 1082 31249 1128
rect 32035 1838 32109 1884
rect 32035 1526 32109 1572
rect 32719 1838 32793 1884
rect 32719 1526 32793 1572
rect 33403 1838 33477 1884
rect 33403 1526 33477 1572
rect 34949 1884 35003 1930
rect 35133 1884 35187 1930
rect 35317 1884 35371 1930
rect 34949 1572 35003 1618
rect 35133 1572 35187 1618
rect 35317 1572 35371 1618
rect 38385 2714 38459 2760
rect 38385 2002 38459 2048
rect 39279 3014 39353 3060
rect 39483 3014 39557 3060
rect 39279 2702 39353 2748
rect 39483 2702 39557 2748
rect 39963 3014 40037 3060
rect 40167 3014 40241 3060
rect 39963 2702 40037 2748
rect 40167 2702 40241 2748
rect 40647 3014 40721 3060
rect 40647 2702 40721 2748
rect 41507 2958 41581 3004
rect 41711 2958 41785 3004
rect 41507 2246 41581 2292
rect 41711 2246 41785 2292
rect 42191 2958 42265 3004
rect 42395 2958 42469 3004
rect 42191 2246 42265 2292
rect 42395 2246 42469 2292
rect 42875 2958 42949 3004
rect 42875 2246 42949 2292
rect 44421 3044 44475 3090
rect 44605 3044 44659 3090
rect 44789 3044 44843 3090
rect 44421 2432 44475 2478
rect 44605 2432 44659 2478
rect 44789 2432 44843 2478
rect 38385 1594 38459 1640
rect 38385 1282 38459 1328
rect 39279 1794 39353 1840
rect 39279 1082 39353 1128
rect 40167 1794 40241 1840
rect 40167 1082 40241 1128
rect 40647 1794 40721 1840
rect 40647 1082 40721 1128
rect 41507 1838 41581 1884
rect 41507 1526 41581 1572
rect 42191 1838 42265 1884
rect 42191 1526 42265 1572
rect 42875 1838 42949 1884
rect 42875 1526 42949 1572
rect 44421 1884 44475 1930
rect 44605 1884 44659 1930
rect 44789 1884 44843 1930
rect 44421 1572 44475 1618
rect 44605 1572 44659 1618
rect 44789 1572 44843 1618
rect 47857 2714 47931 2760
rect 47857 2002 47931 2048
rect 48751 3014 48825 3060
rect 48955 3014 49029 3060
rect 48751 2702 48825 2748
rect 48955 2702 49029 2748
rect 49435 3014 49509 3060
rect 49639 3014 49713 3060
rect 49435 2702 49509 2748
rect 49639 2702 49713 2748
rect 50119 3014 50193 3060
rect 50119 2702 50193 2748
rect 50979 2958 51053 3004
rect 51183 2958 51257 3004
rect 50979 2246 51053 2292
rect 51183 2246 51257 2292
rect 51663 2958 51737 3004
rect 51867 2958 51941 3004
rect 51663 2246 51737 2292
rect 51867 2246 51941 2292
rect 52347 2958 52421 3004
rect 52347 2246 52421 2292
rect 53893 3044 53947 3090
rect 54077 3044 54131 3090
rect 54261 3044 54315 3090
rect 53893 2432 53947 2478
rect 54077 2432 54131 2478
rect 54261 2432 54315 2478
rect 47857 1594 47931 1640
rect 47857 1282 47931 1328
rect 48751 1794 48825 1840
rect 48751 1082 48825 1128
rect 49639 1794 49713 1840
rect 49639 1082 49713 1128
rect 50119 1794 50193 1840
rect 50119 1082 50193 1128
rect 50979 1838 51053 1884
rect 50979 1526 51053 1572
rect 51663 1838 51737 1884
rect 51663 1526 51737 1572
rect 52347 1838 52421 1884
rect 52347 1526 52421 1572
rect 53893 1884 53947 1930
rect 54077 1884 54131 1930
rect 54261 1884 54315 1930
rect 53893 1572 53947 1618
rect 54077 1572 54131 1618
rect 54261 1572 54315 1618
rect 1391 673 1465 719
rect 1595 673 1669 719
rect 1391 361 1465 407
rect 1595 361 1669 407
rect 2075 673 2149 719
rect 2279 673 2353 719
rect 2075 361 2149 407
rect 2279 361 2353 407
rect 2759 673 2833 719
rect 2759 361 2833 407
rect 10863 673 10937 719
rect 11067 673 11141 719
rect 10863 361 10937 407
rect 11067 361 11141 407
rect 11547 673 11621 719
rect 11751 673 11825 719
rect 11547 361 11621 407
rect 11751 361 11825 407
rect 12231 673 12305 719
rect 12231 361 12305 407
rect 20335 674 20409 720
rect 20539 674 20613 720
rect 20335 362 20409 408
rect 20539 362 20613 408
rect 21019 674 21093 720
rect 21223 674 21297 720
rect 21019 362 21093 408
rect 21223 362 21297 408
rect 21703 674 21777 720
rect 21703 362 21777 408
rect 29807 674 29881 720
rect 30011 674 30085 720
rect 29807 362 29881 408
rect 30011 362 30085 408
rect 30491 674 30565 720
rect 30695 674 30769 720
rect 30491 362 30565 408
rect 30695 362 30769 408
rect 31175 674 31249 720
rect 31175 362 31249 408
rect 39279 674 39353 720
rect 39483 674 39557 720
rect 39279 362 39353 408
rect 39483 362 39557 408
rect 39963 674 40037 720
rect 40167 674 40241 720
rect 39963 362 40037 408
rect 40167 362 40241 408
rect 40647 674 40721 720
rect 40647 362 40721 408
rect 48751 674 48825 720
rect 48955 674 49029 720
rect 48751 362 48825 408
rect 48955 362 49029 408
rect 49435 674 49509 720
rect 49639 674 49713 720
rect 49435 362 49509 408
rect 49639 362 49713 408
rect 50119 674 50193 720
rect 50119 362 50193 408
<< metal1 >>
rect 6127 9960 7674 10016
rect 5630 8939 5718 8951
rect 6127 8939 6183 9960
rect 6796 9908 6882 9912
rect 6796 9852 6808 9908
rect 6864 9852 6882 9908
rect 6796 9840 6882 9852
rect 6307 9695 6353 9706
rect 6522 9704 6598 9737
rect 6522 9658 6533 9704
rect 6587 9658 6598 9704
rect 6706 9704 6782 9737
rect 6706 9658 6717 9704
rect 6771 9658 6782 9704
rect 6890 9704 6966 9737
rect 6890 9658 6901 9704
rect 6955 9658 6966 9704
rect 7135 9695 7181 9706
rect 6445 9612 6491 9623
rect 6428 9585 6445 9587
rect 6629 9612 6675 9623
rect 6491 9585 6508 9587
rect 6353 9465 6440 9585
rect 6496 9465 6508 9585
rect 6428 9463 6445 9465
rect 6353 9165 6445 9285
rect 6491 9463 6508 9465
rect 6612 9285 6629 9287
rect 6813 9612 6859 9623
rect 6796 9585 6813 9587
rect 6997 9612 7043 9623
rect 6859 9585 6876 9587
rect 6796 9465 6808 9585
rect 6864 9465 6876 9585
rect 6796 9463 6813 9465
rect 6675 9285 6692 9287
rect 6612 9165 6624 9285
rect 6680 9165 6692 9285
rect 6612 9163 6629 9165
rect 6445 9127 6491 9138
rect 6675 9163 6692 9165
rect 6629 9127 6675 9138
rect 6859 9463 6876 9465
rect 6980 9285 6997 9287
rect 7118 9585 7135 9587
rect 7181 9585 7198 9587
rect 7118 9464 7130 9585
rect 7186 9464 7198 9585
rect 7118 9462 7135 9464
rect 7043 9285 7060 9287
rect 6980 9165 6992 9285
rect 7048 9165 7060 9285
rect 6980 9163 6997 9165
rect 6813 9127 6859 9138
rect 7043 9163 7060 9165
rect 6997 9127 7043 9138
rect 6522 9089 6533 9092
rect 6587 9089 6598 9092
rect 6706 9089 6717 9092
rect 6771 9089 6782 9092
rect 6890 9089 6901 9092
rect 6955 9089 6966 9092
rect 6307 9044 6353 9055
rect 6520 9033 6532 9089
rect 6588 9033 6600 9089
rect 6520 9019 6600 9033
rect 6704 9033 6716 9089
rect 6772 9033 6784 9089
rect 6704 9019 6784 9033
rect 6888 9033 6900 9089
rect 6956 9033 6968 9089
rect 7181 9462 7198 9464
rect 7135 9044 7181 9055
rect 6888 9019 6968 9033
rect 6520 8939 6600 8941
rect 5630 8883 5644 8939
rect 5700 8883 6532 8939
rect 6588 8883 6600 8939
rect 5630 8871 5718 8883
rect 6520 8881 6600 8883
rect 5848 8823 5918 8835
rect 6704 8823 6784 8825
rect 5848 8767 5860 8823
rect 5916 8767 6716 8823
rect 6772 8767 6784 8823
rect 5848 8755 5918 8767
rect 6704 8765 6784 8767
rect 7033 8823 7113 8825
rect 7300 8823 7370 8835
rect 7033 8767 7045 8823
rect 7101 8767 7302 8823
rect 7358 8767 7370 8823
rect 7033 8765 7113 8767
rect 7300 8757 7370 8767
rect 6888 8707 6968 8709
rect 6132 8651 6900 8707
rect 6956 8651 6968 8707
rect 6132 7920 6188 8651
rect 6888 8649 6968 8651
rect 6520 8557 6600 8571
rect 6307 8535 6353 8546
rect 6520 8501 6532 8557
rect 6588 8501 6600 8557
rect 6704 8557 6784 8571
rect 6704 8501 6716 8557
rect 6772 8501 6784 8557
rect 6888 8557 6968 8571
rect 6888 8501 6900 8557
rect 6956 8501 6968 8557
rect 7135 8535 7181 8546
rect 6522 8498 6533 8501
rect 6587 8498 6598 8501
rect 6706 8498 6717 8501
rect 6771 8498 6782 8501
rect 6890 8498 6901 8501
rect 6955 8498 6966 8501
rect 6445 8452 6491 8463
rect 6353 8278 6445 8452
rect 6445 8267 6491 8278
rect 6629 8452 6675 8463
rect 6629 8267 6675 8278
rect 6813 8452 6859 8463
rect 6997 8452 7043 8463
rect 6980 8425 6997 8427
rect 7043 8425 7060 8427
rect 6980 8305 6992 8425
rect 7048 8305 7060 8425
rect 6980 8303 6997 8305
rect 6813 8267 6859 8278
rect 7043 8303 7060 8305
rect 6997 8267 7043 8278
rect 6307 8050 6353 8195
rect 6522 8186 6533 8232
rect 6587 8186 6598 8232
rect 6522 8153 6598 8186
rect 6706 8186 6717 8232
rect 6771 8186 6782 8232
rect 6706 8153 6782 8186
rect 6890 8186 6901 8232
rect 6955 8186 6966 8232
rect 6890 8153 6966 8186
rect 7135 8050 7181 8195
rect 6295 8038 6375 8050
rect 6295 7982 6307 8038
rect 6363 7982 6375 8038
rect 6295 7970 6375 7982
rect 7113 8038 7193 8050
rect 7113 7982 7125 8038
rect 7181 7982 7193 8038
rect 7113 7970 7193 7982
rect 7466 7920 7546 7930
rect 6132 7864 7478 7920
rect 7534 7864 7546 7920
rect 7466 7862 7546 7864
rect 7300 7811 7370 7813
rect 6132 7810 7370 7811
rect 6132 7756 7302 7810
rect 7358 7756 7370 7810
rect 6132 7755 7370 7756
rect 6132 6734 6188 7755
rect 7300 7747 7370 7755
rect 6796 7703 6882 7707
rect 6796 7647 6808 7703
rect 6864 7647 6882 7703
rect 6796 7635 6882 7647
rect 6307 7490 6353 7501
rect 6522 7499 6598 7532
rect 6522 7453 6533 7499
rect 6587 7453 6598 7499
rect 6706 7499 6782 7532
rect 6706 7453 6717 7499
rect 6771 7453 6782 7499
rect 6890 7499 6966 7532
rect 6890 7453 6901 7499
rect 6955 7453 6966 7499
rect 7135 7490 7181 7501
rect 6445 7407 6491 7418
rect 6428 7380 6445 7382
rect 6629 7407 6675 7418
rect 6491 7380 6508 7382
rect 6353 7260 6440 7380
rect 6496 7260 6508 7380
rect 6428 7258 6445 7260
rect 6353 6960 6445 7080
rect 6491 7258 6508 7260
rect 6612 7080 6629 7082
rect 6813 7407 6859 7418
rect 6796 7380 6813 7382
rect 6997 7407 7043 7418
rect 6859 7380 6876 7382
rect 6796 7260 6808 7380
rect 6864 7260 6876 7380
rect 6796 7258 6813 7260
rect 6675 7080 6692 7082
rect 6612 6960 6624 7080
rect 6680 6960 6692 7080
rect 6612 6958 6629 6960
rect 6445 6922 6491 6933
rect 6675 6958 6692 6960
rect 6629 6922 6675 6933
rect 6859 7258 6876 7260
rect 6980 7080 6997 7082
rect 7118 7380 7135 7382
rect 7181 7380 7198 7382
rect 7118 7259 7130 7380
rect 7186 7259 7198 7380
rect 7118 7257 7135 7259
rect 7043 7080 7060 7082
rect 6980 6960 6992 7080
rect 7048 6960 7060 7080
rect 6980 6958 6997 6960
rect 6813 6922 6859 6933
rect 7043 6958 7060 6960
rect 6997 6922 7043 6933
rect 6522 6884 6533 6887
rect 6587 6884 6598 6887
rect 6706 6884 6717 6887
rect 6771 6884 6782 6887
rect 6890 6884 6901 6887
rect 6955 6884 6966 6887
rect 6307 6839 6353 6850
rect 6520 6828 6532 6884
rect 6588 6828 6600 6884
rect 6520 6814 6600 6828
rect 6704 6828 6716 6884
rect 6772 6828 6784 6884
rect 6704 6814 6784 6828
rect 6888 6828 6900 6884
rect 6956 6828 6968 6884
rect 7181 7257 7198 7259
rect 7135 6839 7181 6850
rect 6888 6814 6968 6828
rect 6520 6734 6600 6736
rect 6132 6678 6532 6734
rect 6588 6678 6600 6734
rect 7618 6734 7674 9960
rect 15599 9960 17146 10016
rect 15102 8939 15190 8951
rect 15599 8939 15655 9960
rect 16268 9908 16354 9912
rect 16268 9852 16280 9908
rect 16336 9852 16354 9908
rect 16268 9840 16354 9852
rect 15779 9695 15825 9706
rect 15994 9704 16070 9737
rect 15994 9658 16005 9704
rect 16059 9658 16070 9704
rect 16178 9704 16254 9737
rect 16178 9658 16189 9704
rect 16243 9658 16254 9704
rect 16362 9704 16438 9737
rect 16362 9658 16373 9704
rect 16427 9658 16438 9704
rect 16607 9695 16653 9706
rect 15917 9612 15963 9623
rect 15900 9585 15917 9587
rect 16101 9612 16147 9623
rect 15963 9585 15980 9587
rect 15825 9465 15912 9585
rect 15968 9465 15980 9585
rect 15900 9463 15917 9465
rect 15825 9165 15917 9285
rect 15963 9463 15980 9465
rect 16084 9285 16101 9287
rect 16285 9612 16331 9623
rect 16268 9585 16285 9587
rect 16469 9612 16515 9623
rect 16331 9585 16348 9587
rect 16268 9465 16280 9585
rect 16336 9465 16348 9585
rect 16268 9463 16285 9465
rect 16147 9285 16164 9287
rect 16084 9165 16096 9285
rect 16152 9165 16164 9285
rect 16084 9163 16101 9165
rect 15917 9127 15963 9138
rect 16147 9163 16164 9165
rect 16101 9127 16147 9138
rect 16331 9463 16348 9465
rect 16452 9285 16469 9287
rect 16590 9585 16607 9587
rect 16653 9585 16670 9587
rect 16590 9464 16602 9585
rect 16658 9464 16670 9585
rect 16590 9462 16607 9464
rect 16515 9285 16532 9287
rect 16452 9165 16464 9285
rect 16520 9165 16532 9285
rect 16452 9163 16469 9165
rect 16285 9127 16331 9138
rect 16515 9163 16532 9165
rect 16469 9127 16515 9138
rect 15994 9089 16005 9092
rect 16059 9089 16070 9092
rect 16178 9089 16189 9092
rect 16243 9089 16254 9092
rect 16362 9089 16373 9092
rect 16427 9089 16438 9092
rect 15779 9044 15825 9055
rect 15992 9033 16004 9089
rect 16060 9033 16072 9089
rect 15992 9019 16072 9033
rect 16176 9033 16188 9089
rect 16244 9033 16256 9089
rect 16176 9019 16256 9033
rect 16360 9033 16372 9089
rect 16428 9033 16440 9089
rect 16653 9462 16670 9464
rect 16607 9044 16653 9055
rect 16360 9019 16440 9033
rect 15992 8939 16072 8941
rect 15102 8883 15116 8939
rect 15172 8883 16004 8939
rect 16060 8883 16072 8939
rect 15102 8871 15190 8883
rect 15992 8881 16072 8883
rect 15320 8823 15390 8835
rect 16176 8823 16256 8825
rect 15320 8767 15332 8823
rect 15388 8767 16188 8823
rect 16244 8767 16256 8823
rect 15320 8755 15390 8767
rect 16176 8765 16256 8767
rect 16505 8823 16585 8825
rect 16772 8823 16842 8835
rect 16505 8767 16517 8823
rect 16573 8767 16774 8823
rect 16830 8767 16842 8823
rect 16505 8765 16585 8767
rect 16772 8757 16842 8767
rect 16360 8707 16440 8709
rect 15604 8651 16372 8707
rect 16428 8651 16440 8707
rect 15604 7920 15660 8651
rect 16360 8649 16440 8651
rect 15992 8557 16072 8571
rect 15779 8535 15825 8546
rect 15992 8501 16004 8557
rect 16060 8501 16072 8557
rect 16176 8557 16256 8571
rect 16176 8501 16188 8557
rect 16244 8501 16256 8557
rect 16360 8557 16440 8571
rect 16360 8501 16372 8557
rect 16428 8501 16440 8557
rect 16607 8535 16653 8546
rect 15994 8498 16005 8501
rect 16059 8498 16070 8501
rect 16178 8498 16189 8501
rect 16243 8498 16254 8501
rect 16362 8498 16373 8501
rect 16427 8498 16438 8501
rect 15917 8452 15963 8463
rect 15825 8278 15917 8452
rect 15917 8267 15963 8278
rect 16101 8452 16147 8463
rect 16101 8267 16147 8278
rect 16285 8452 16331 8463
rect 16469 8452 16515 8463
rect 16452 8425 16469 8427
rect 16515 8425 16532 8427
rect 16452 8305 16464 8425
rect 16520 8305 16532 8425
rect 16452 8303 16469 8305
rect 16285 8267 16331 8278
rect 16515 8303 16532 8305
rect 16469 8267 16515 8278
rect 15779 8050 15825 8195
rect 15994 8186 16005 8232
rect 16059 8186 16070 8232
rect 15994 8153 16070 8186
rect 16178 8186 16189 8232
rect 16243 8186 16254 8232
rect 16178 8153 16254 8186
rect 16362 8186 16373 8232
rect 16427 8186 16438 8232
rect 16362 8153 16438 8186
rect 16607 8050 16653 8195
rect 15767 8038 15847 8050
rect 15767 7982 15779 8038
rect 15835 7982 15847 8038
rect 15767 7970 15847 7982
rect 16585 8038 16665 8050
rect 16585 7982 16597 8038
rect 16653 7982 16665 8038
rect 16585 7970 16665 7982
rect 16938 7920 17018 7930
rect 15604 7864 16950 7920
rect 17006 7864 17018 7920
rect 16938 7862 17018 7864
rect 16772 7811 16842 7813
rect 15604 7810 16842 7811
rect 15604 7756 16774 7810
rect 16830 7756 16842 7810
rect 15604 7755 16842 7756
rect 8282 7703 8368 7707
rect 8282 7647 8294 7703
rect 8350 7647 8368 7703
rect 8282 7635 8368 7647
rect 7793 7490 7839 7501
rect 8008 7499 8084 7532
rect 8008 7453 8019 7499
rect 8073 7453 8084 7499
rect 8192 7499 8268 7532
rect 8192 7453 8203 7499
rect 8257 7453 8268 7499
rect 8376 7499 8452 7532
rect 8376 7453 8387 7499
rect 8441 7453 8452 7499
rect 8621 7490 8667 7501
rect 7931 7407 7977 7418
rect 7914 7380 7931 7382
rect 8115 7407 8161 7418
rect 7977 7380 7994 7382
rect 7839 7260 7926 7380
rect 7982 7260 7994 7380
rect 7914 7258 7931 7260
rect 7839 6960 7931 7080
rect 7977 7258 7994 7260
rect 8098 7080 8115 7082
rect 8299 7407 8345 7418
rect 8282 7380 8299 7382
rect 8483 7407 8529 7418
rect 8345 7380 8362 7382
rect 8282 7260 8294 7380
rect 8350 7260 8362 7380
rect 8282 7258 8299 7260
rect 8161 7080 8178 7082
rect 8098 6960 8110 7080
rect 8166 6960 8178 7080
rect 8098 6958 8115 6960
rect 7931 6922 7977 6933
rect 8161 6958 8178 6960
rect 8115 6922 8161 6933
rect 8345 7258 8362 7260
rect 8466 7080 8483 7082
rect 8604 7380 8621 7382
rect 8667 7380 8684 7382
rect 8604 7259 8616 7380
rect 8672 7259 8684 7380
rect 8604 7257 8621 7259
rect 8529 7080 8546 7082
rect 8466 6960 8478 7080
rect 8534 6960 8546 7080
rect 8466 6958 8483 6960
rect 8299 6922 8345 6933
rect 8529 6958 8546 6960
rect 8483 6922 8529 6933
rect 8008 6884 8019 6887
rect 8073 6884 8084 6887
rect 8192 6884 8203 6887
rect 8257 6884 8268 6887
rect 8376 6884 8387 6887
rect 8441 6884 8452 6887
rect 7793 6839 7839 6850
rect 8006 6828 8018 6884
rect 8074 6828 8086 6884
rect 8006 6814 8086 6828
rect 8190 6828 8202 6884
rect 8258 6828 8270 6884
rect 8190 6814 8270 6828
rect 8374 6828 8386 6884
rect 8442 6828 8454 6884
rect 8667 7257 8684 7259
rect 8621 6839 8667 6850
rect 8374 6814 8454 6828
rect 8006 6734 8086 6736
rect 7618 6678 8018 6734
rect 8074 6678 8086 6734
rect 15604 6734 15660 7755
rect 16772 7747 16842 7755
rect 16268 7703 16354 7707
rect 16268 7647 16280 7703
rect 16336 7647 16354 7703
rect 16268 7635 16354 7647
rect 15779 7490 15825 7501
rect 15994 7499 16070 7532
rect 15994 7453 16005 7499
rect 16059 7453 16070 7499
rect 16178 7499 16254 7532
rect 16178 7453 16189 7499
rect 16243 7453 16254 7499
rect 16362 7499 16438 7532
rect 16362 7453 16373 7499
rect 16427 7453 16438 7499
rect 16607 7490 16653 7501
rect 15917 7407 15963 7418
rect 15900 7380 15917 7382
rect 16101 7407 16147 7418
rect 15963 7380 15980 7382
rect 15825 7260 15912 7380
rect 15968 7260 15980 7380
rect 15900 7258 15917 7260
rect 15825 6960 15917 7080
rect 15963 7258 15980 7260
rect 16084 7080 16101 7082
rect 16285 7407 16331 7418
rect 16268 7380 16285 7382
rect 16469 7407 16515 7418
rect 16331 7380 16348 7382
rect 16268 7260 16280 7380
rect 16336 7260 16348 7380
rect 16268 7258 16285 7260
rect 16147 7080 16164 7082
rect 16084 6960 16096 7080
rect 16152 6960 16164 7080
rect 16084 6958 16101 6960
rect 15917 6922 15963 6933
rect 16147 6958 16164 6960
rect 16101 6922 16147 6933
rect 16331 7258 16348 7260
rect 16452 7080 16469 7082
rect 16590 7380 16607 7382
rect 16653 7380 16670 7382
rect 16590 7259 16602 7380
rect 16658 7259 16670 7380
rect 16590 7257 16607 7259
rect 16515 7080 16532 7082
rect 16452 6960 16464 7080
rect 16520 6960 16532 7080
rect 16452 6958 16469 6960
rect 16285 6922 16331 6933
rect 16515 6958 16532 6960
rect 16469 6922 16515 6933
rect 15994 6884 16005 6887
rect 16059 6884 16070 6887
rect 16178 6884 16189 6887
rect 16243 6884 16254 6887
rect 16362 6884 16373 6887
rect 16427 6884 16438 6887
rect 15779 6839 15825 6850
rect 15992 6828 16004 6884
rect 16060 6828 16072 6884
rect 15992 6814 16072 6828
rect 16176 6828 16188 6884
rect 16244 6828 16256 6884
rect 16176 6814 16256 6828
rect 16360 6828 16372 6884
rect 16428 6828 16440 6884
rect 16653 7257 16670 7259
rect 16607 6839 16653 6850
rect 16360 6814 16440 6828
rect 15992 6734 16072 6736
rect 15604 6678 16004 6734
rect 16060 6678 16072 6734
rect 17090 6734 17146 9960
rect 25071 9961 26618 10017
rect 24574 8940 24662 8952
rect 25071 8940 25127 9961
rect 25740 9909 25826 9913
rect 25740 9853 25752 9909
rect 25808 9853 25826 9909
rect 25740 9841 25826 9853
rect 25251 9696 25297 9707
rect 25466 9705 25542 9738
rect 25466 9659 25477 9705
rect 25531 9659 25542 9705
rect 25650 9705 25726 9738
rect 25650 9659 25661 9705
rect 25715 9659 25726 9705
rect 25834 9705 25910 9738
rect 25834 9659 25845 9705
rect 25899 9659 25910 9705
rect 26079 9696 26125 9707
rect 25389 9613 25435 9624
rect 25372 9586 25389 9588
rect 25573 9613 25619 9624
rect 25435 9586 25452 9588
rect 25297 9466 25384 9586
rect 25440 9466 25452 9586
rect 25372 9464 25389 9466
rect 25297 9166 25389 9286
rect 25435 9464 25452 9466
rect 25556 9286 25573 9288
rect 25757 9613 25803 9624
rect 25740 9586 25757 9588
rect 25941 9613 25987 9624
rect 25803 9586 25820 9588
rect 25740 9466 25752 9586
rect 25808 9466 25820 9586
rect 25740 9464 25757 9466
rect 25619 9286 25636 9288
rect 25556 9166 25568 9286
rect 25624 9166 25636 9286
rect 25556 9164 25573 9166
rect 25389 9128 25435 9139
rect 25619 9164 25636 9166
rect 25573 9128 25619 9139
rect 25803 9464 25820 9466
rect 25924 9286 25941 9288
rect 26062 9586 26079 9588
rect 26125 9586 26142 9588
rect 26062 9465 26074 9586
rect 26130 9465 26142 9586
rect 26062 9463 26079 9465
rect 25987 9286 26004 9288
rect 25924 9166 25936 9286
rect 25992 9166 26004 9286
rect 25924 9164 25941 9166
rect 25757 9128 25803 9139
rect 25987 9164 26004 9166
rect 25941 9128 25987 9139
rect 25466 9090 25477 9093
rect 25531 9090 25542 9093
rect 25650 9090 25661 9093
rect 25715 9090 25726 9093
rect 25834 9090 25845 9093
rect 25899 9090 25910 9093
rect 25251 9045 25297 9056
rect 25464 9034 25476 9090
rect 25532 9034 25544 9090
rect 25464 9020 25544 9034
rect 25648 9034 25660 9090
rect 25716 9034 25728 9090
rect 25648 9020 25728 9034
rect 25832 9034 25844 9090
rect 25900 9034 25912 9090
rect 26125 9463 26142 9465
rect 26079 9045 26125 9056
rect 25832 9020 25912 9034
rect 25464 8940 25544 8942
rect 24574 8884 24588 8940
rect 24644 8884 25476 8940
rect 25532 8884 25544 8940
rect 24574 8872 24662 8884
rect 25464 8882 25544 8884
rect 24792 8824 24862 8836
rect 25648 8824 25728 8826
rect 24792 8768 24804 8824
rect 24860 8768 25660 8824
rect 25716 8768 25728 8824
rect 24792 8756 24862 8768
rect 25648 8766 25728 8768
rect 25977 8824 26057 8826
rect 26244 8824 26314 8836
rect 25977 8768 25989 8824
rect 26045 8768 26246 8824
rect 26302 8768 26314 8824
rect 25977 8766 26057 8768
rect 26244 8758 26314 8768
rect 25832 8708 25912 8710
rect 25076 8652 25844 8708
rect 25900 8652 25912 8708
rect 25076 7921 25132 8652
rect 25832 8650 25912 8652
rect 25464 8558 25544 8572
rect 25251 8536 25297 8547
rect 25464 8502 25476 8558
rect 25532 8502 25544 8558
rect 25648 8558 25728 8572
rect 25648 8502 25660 8558
rect 25716 8502 25728 8558
rect 25832 8558 25912 8572
rect 25832 8502 25844 8558
rect 25900 8502 25912 8558
rect 26079 8536 26125 8547
rect 25466 8499 25477 8502
rect 25531 8499 25542 8502
rect 25650 8499 25661 8502
rect 25715 8499 25726 8502
rect 25834 8499 25845 8502
rect 25899 8499 25910 8502
rect 25389 8453 25435 8464
rect 25297 8279 25389 8453
rect 25389 8268 25435 8279
rect 25573 8453 25619 8464
rect 25573 8268 25619 8279
rect 25757 8453 25803 8464
rect 25941 8453 25987 8464
rect 25924 8426 25941 8428
rect 25987 8426 26004 8428
rect 25924 8306 25936 8426
rect 25992 8306 26004 8426
rect 25924 8304 25941 8306
rect 25757 8268 25803 8279
rect 25987 8304 26004 8306
rect 25941 8268 25987 8279
rect 25251 8051 25297 8196
rect 25466 8187 25477 8233
rect 25531 8187 25542 8233
rect 25466 8154 25542 8187
rect 25650 8187 25661 8233
rect 25715 8187 25726 8233
rect 25650 8154 25726 8187
rect 25834 8187 25845 8233
rect 25899 8187 25910 8233
rect 25834 8154 25910 8187
rect 26079 8051 26125 8196
rect 25239 8039 25319 8051
rect 25239 7983 25251 8039
rect 25307 7983 25319 8039
rect 25239 7971 25319 7983
rect 26057 8039 26137 8051
rect 26057 7983 26069 8039
rect 26125 7983 26137 8039
rect 26057 7971 26137 7983
rect 26410 7921 26490 7931
rect 25076 7865 26422 7921
rect 26478 7865 26490 7921
rect 26410 7863 26490 7865
rect 26244 7812 26314 7814
rect 25076 7811 26314 7812
rect 25076 7757 26246 7811
rect 26302 7757 26314 7811
rect 25076 7756 26314 7757
rect 17754 7703 17840 7707
rect 17754 7647 17766 7703
rect 17822 7647 17840 7703
rect 17754 7635 17840 7647
rect 17265 7490 17311 7501
rect 17480 7499 17556 7532
rect 17480 7453 17491 7499
rect 17545 7453 17556 7499
rect 17664 7499 17740 7532
rect 17664 7453 17675 7499
rect 17729 7453 17740 7499
rect 17848 7499 17924 7532
rect 17848 7453 17859 7499
rect 17913 7453 17924 7499
rect 18093 7490 18139 7501
rect 17403 7407 17449 7418
rect 17386 7380 17403 7382
rect 17587 7407 17633 7418
rect 17449 7380 17466 7382
rect 17311 7260 17398 7380
rect 17454 7260 17466 7380
rect 17386 7258 17403 7260
rect 17311 6960 17403 7080
rect 17449 7258 17466 7260
rect 17570 7080 17587 7082
rect 17771 7407 17817 7418
rect 17754 7380 17771 7382
rect 17955 7407 18001 7418
rect 17817 7380 17834 7382
rect 17754 7260 17766 7380
rect 17822 7260 17834 7380
rect 17754 7258 17771 7260
rect 17633 7080 17650 7082
rect 17570 6960 17582 7080
rect 17638 6960 17650 7080
rect 17570 6958 17587 6960
rect 17403 6922 17449 6933
rect 17633 6958 17650 6960
rect 17587 6922 17633 6933
rect 17817 7258 17834 7260
rect 17938 7080 17955 7082
rect 18076 7380 18093 7382
rect 18139 7380 18156 7382
rect 18076 7259 18088 7380
rect 18144 7259 18156 7380
rect 18076 7257 18093 7259
rect 18001 7080 18018 7082
rect 17938 6960 17950 7080
rect 18006 6960 18018 7080
rect 17938 6958 17955 6960
rect 17771 6922 17817 6933
rect 18001 6958 18018 6960
rect 17955 6922 18001 6933
rect 17480 6884 17491 6887
rect 17545 6884 17556 6887
rect 17664 6884 17675 6887
rect 17729 6884 17740 6887
rect 17848 6884 17859 6887
rect 17913 6884 17924 6887
rect 17265 6839 17311 6850
rect 17478 6828 17490 6884
rect 17546 6828 17558 6884
rect 17478 6814 17558 6828
rect 17662 6828 17674 6884
rect 17730 6828 17742 6884
rect 17662 6814 17742 6828
rect 17846 6828 17858 6884
rect 17914 6828 17926 6884
rect 18139 7257 18156 7259
rect 18093 6839 18139 6850
rect 17846 6814 17926 6828
rect 17478 6734 17558 6736
rect 17090 6678 17490 6734
rect 17546 6678 17558 6734
rect 25076 6735 25132 7756
rect 26244 7748 26314 7756
rect 25740 7704 25826 7708
rect 25740 7648 25752 7704
rect 25808 7648 25826 7704
rect 25740 7636 25826 7648
rect 25251 7491 25297 7502
rect 25466 7500 25542 7533
rect 25466 7454 25477 7500
rect 25531 7454 25542 7500
rect 25650 7500 25726 7533
rect 25650 7454 25661 7500
rect 25715 7454 25726 7500
rect 25834 7500 25910 7533
rect 25834 7454 25845 7500
rect 25899 7454 25910 7500
rect 26079 7491 26125 7502
rect 25389 7408 25435 7419
rect 25372 7381 25389 7383
rect 25573 7408 25619 7419
rect 25435 7381 25452 7383
rect 25297 7261 25384 7381
rect 25440 7261 25452 7381
rect 25372 7259 25389 7261
rect 25297 6961 25389 7081
rect 25435 7259 25452 7261
rect 25556 7081 25573 7083
rect 25757 7408 25803 7419
rect 25740 7381 25757 7383
rect 25941 7408 25987 7419
rect 25803 7381 25820 7383
rect 25740 7261 25752 7381
rect 25808 7261 25820 7381
rect 25740 7259 25757 7261
rect 25619 7081 25636 7083
rect 25556 6961 25568 7081
rect 25624 6961 25636 7081
rect 25556 6959 25573 6961
rect 25389 6923 25435 6934
rect 25619 6959 25636 6961
rect 25573 6923 25619 6934
rect 25803 7259 25820 7261
rect 25924 7081 25941 7083
rect 26062 7381 26079 7383
rect 26125 7381 26142 7383
rect 26062 7260 26074 7381
rect 26130 7260 26142 7381
rect 26062 7258 26079 7260
rect 25987 7081 26004 7083
rect 25924 6961 25936 7081
rect 25992 6961 26004 7081
rect 25924 6959 25941 6961
rect 25757 6923 25803 6934
rect 25987 6959 26004 6961
rect 25941 6923 25987 6934
rect 25466 6885 25477 6888
rect 25531 6885 25542 6888
rect 25650 6885 25661 6888
rect 25715 6885 25726 6888
rect 25834 6885 25845 6888
rect 25899 6885 25910 6888
rect 25251 6840 25297 6851
rect 25464 6829 25476 6885
rect 25532 6829 25544 6885
rect 25464 6815 25544 6829
rect 25648 6829 25660 6885
rect 25716 6829 25728 6885
rect 25648 6815 25728 6829
rect 25832 6829 25844 6885
rect 25900 6829 25912 6885
rect 26125 7258 26142 7260
rect 26079 6840 26125 6851
rect 25832 6815 25912 6829
rect 25464 6735 25544 6737
rect 25076 6679 25476 6735
rect 25532 6679 25544 6735
rect 26562 6735 26618 9961
rect 34543 9961 36090 10017
rect 34046 8940 34134 8952
rect 34543 8940 34599 9961
rect 35212 9909 35298 9913
rect 35212 9853 35224 9909
rect 35280 9853 35298 9909
rect 35212 9841 35298 9853
rect 34723 9696 34769 9707
rect 34938 9705 35014 9738
rect 34938 9659 34949 9705
rect 35003 9659 35014 9705
rect 35122 9705 35198 9738
rect 35122 9659 35133 9705
rect 35187 9659 35198 9705
rect 35306 9705 35382 9738
rect 35306 9659 35317 9705
rect 35371 9659 35382 9705
rect 35551 9696 35597 9707
rect 34861 9613 34907 9624
rect 34844 9586 34861 9588
rect 35045 9613 35091 9624
rect 34907 9586 34924 9588
rect 34769 9466 34856 9586
rect 34912 9466 34924 9586
rect 34844 9464 34861 9466
rect 34769 9166 34861 9286
rect 34907 9464 34924 9466
rect 35028 9286 35045 9288
rect 35229 9613 35275 9624
rect 35212 9586 35229 9588
rect 35413 9613 35459 9624
rect 35275 9586 35292 9588
rect 35212 9466 35224 9586
rect 35280 9466 35292 9586
rect 35212 9464 35229 9466
rect 35091 9286 35108 9288
rect 35028 9166 35040 9286
rect 35096 9166 35108 9286
rect 35028 9164 35045 9166
rect 34861 9128 34907 9139
rect 35091 9164 35108 9166
rect 35045 9128 35091 9139
rect 35275 9464 35292 9466
rect 35396 9286 35413 9288
rect 35534 9586 35551 9588
rect 35597 9586 35614 9588
rect 35534 9465 35546 9586
rect 35602 9465 35614 9586
rect 35534 9463 35551 9465
rect 35459 9286 35476 9288
rect 35396 9166 35408 9286
rect 35464 9166 35476 9286
rect 35396 9164 35413 9166
rect 35229 9128 35275 9139
rect 35459 9164 35476 9166
rect 35413 9128 35459 9139
rect 34938 9090 34949 9093
rect 35003 9090 35014 9093
rect 35122 9090 35133 9093
rect 35187 9090 35198 9093
rect 35306 9090 35317 9093
rect 35371 9090 35382 9093
rect 34723 9045 34769 9056
rect 34936 9034 34948 9090
rect 35004 9034 35016 9090
rect 34936 9020 35016 9034
rect 35120 9034 35132 9090
rect 35188 9034 35200 9090
rect 35120 9020 35200 9034
rect 35304 9034 35316 9090
rect 35372 9034 35384 9090
rect 35597 9463 35614 9465
rect 35551 9045 35597 9056
rect 35304 9020 35384 9034
rect 34936 8940 35016 8942
rect 34046 8884 34060 8940
rect 34116 8884 34948 8940
rect 35004 8884 35016 8940
rect 34046 8872 34134 8884
rect 34936 8882 35016 8884
rect 34264 8824 34334 8836
rect 35120 8824 35200 8826
rect 34264 8768 34276 8824
rect 34332 8768 35132 8824
rect 35188 8768 35200 8824
rect 34264 8756 34334 8768
rect 35120 8766 35200 8768
rect 35449 8824 35529 8826
rect 35716 8824 35786 8836
rect 35449 8768 35461 8824
rect 35517 8768 35718 8824
rect 35774 8768 35786 8824
rect 35449 8766 35529 8768
rect 35716 8758 35786 8768
rect 35304 8708 35384 8710
rect 34548 8652 35316 8708
rect 35372 8652 35384 8708
rect 34548 7921 34604 8652
rect 35304 8650 35384 8652
rect 34936 8558 35016 8572
rect 34723 8536 34769 8547
rect 34936 8502 34948 8558
rect 35004 8502 35016 8558
rect 35120 8558 35200 8572
rect 35120 8502 35132 8558
rect 35188 8502 35200 8558
rect 35304 8558 35384 8572
rect 35304 8502 35316 8558
rect 35372 8502 35384 8558
rect 35551 8536 35597 8547
rect 34938 8499 34949 8502
rect 35003 8499 35014 8502
rect 35122 8499 35133 8502
rect 35187 8499 35198 8502
rect 35306 8499 35317 8502
rect 35371 8499 35382 8502
rect 34861 8453 34907 8464
rect 34769 8279 34861 8453
rect 34861 8268 34907 8279
rect 35045 8453 35091 8464
rect 35045 8268 35091 8279
rect 35229 8453 35275 8464
rect 35413 8453 35459 8464
rect 35396 8426 35413 8428
rect 35459 8426 35476 8428
rect 35396 8306 35408 8426
rect 35464 8306 35476 8426
rect 35396 8304 35413 8306
rect 35229 8268 35275 8279
rect 35459 8304 35476 8306
rect 35413 8268 35459 8279
rect 34723 8051 34769 8196
rect 34938 8187 34949 8233
rect 35003 8187 35014 8233
rect 34938 8154 35014 8187
rect 35122 8187 35133 8233
rect 35187 8187 35198 8233
rect 35122 8154 35198 8187
rect 35306 8187 35317 8233
rect 35371 8187 35382 8233
rect 35306 8154 35382 8187
rect 35551 8051 35597 8196
rect 34711 8039 34791 8051
rect 34711 7983 34723 8039
rect 34779 7983 34791 8039
rect 34711 7971 34791 7983
rect 35529 8039 35609 8051
rect 35529 7983 35541 8039
rect 35597 7983 35609 8039
rect 35529 7971 35609 7983
rect 35882 7921 35962 7931
rect 34548 7865 35894 7921
rect 35950 7865 35962 7921
rect 35882 7863 35962 7865
rect 35716 7812 35786 7814
rect 34548 7811 35786 7812
rect 34548 7757 35718 7811
rect 35774 7757 35786 7811
rect 34548 7756 35786 7757
rect 27226 7704 27312 7708
rect 27226 7648 27238 7704
rect 27294 7648 27312 7704
rect 27226 7636 27312 7648
rect 26737 7491 26783 7502
rect 26952 7500 27028 7533
rect 26952 7454 26963 7500
rect 27017 7454 27028 7500
rect 27136 7500 27212 7533
rect 27136 7454 27147 7500
rect 27201 7454 27212 7500
rect 27320 7500 27396 7533
rect 27320 7454 27331 7500
rect 27385 7454 27396 7500
rect 27565 7491 27611 7502
rect 26875 7408 26921 7419
rect 26858 7381 26875 7383
rect 27059 7408 27105 7419
rect 26921 7381 26938 7383
rect 26783 7261 26870 7381
rect 26926 7261 26938 7381
rect 26858 7259 26875 7261
rect 26783 6961 26875 7081
rect 26921 7259 26938 7261
rect 27042 7081 27059 7083
rect 27243 7408 27289 7419
rect 27226 7381 27243 7383
rect 27427 7408 27473 7419
rect 27289 7381 27306 7383
rect 27226 7261 27238 7381
rect 27294 7261 27306 7381
rect 27226 7259 27243 7261
rect 27105 7081 27122 7083
rect 27042 6961 27054 7081
rect 27110 6961 27122 7081
rect 27042 6959 27059 6961
rect 26875 6923 26921 6934
rect 27105 6959 27122 6961
rect 27059 6923 27105 6934
rect 27289 7259 27306 7261
rect 27410 7081 27427 7083
rect 27548 7381 27565 7383
rect 27611 7381 27628 7383
rect 27548 7260 27560 7381
rect 27616 7260 27628 7381
rect 27548 7258 27565 7260
rect 27473 7081 27490 7083
rect 27410 6961 27422 7081
rect 27478 6961 27490 7081
rect 27410 6959 27427 6961
rect 27243 6923 27289 6934
rect 27473 6959 27490 6961
rect 27427 6923 27473 6934
rect 26952 6885 26963 6888
rect 27017 6885 27028 6888
rect 27136 6885 27147 6888
rect 27201 6885 27212 6888
rect 27320 6885 27331 6888
rect 27385 6885 27396 6888
rect 26737 6840 26783 6851
rect 26950 6829 26962 6885
rect 27018 6829 27030 6885
rect 26950 6815 27030 6829
rect 27134 6829 27146 6885
rect 27202 6829 27214 6885
rect 27134 6815 27214 6829
rect 27318 6829 27330 6885
rect 27386 6829 27398 6885
rect 27611 7258 27628 7260
rect 27565 6840 27611 6851
rect 27318 6815 27398 6829
rect 26950 6735 27030 6737
rect 26562 6679 26962 6735
rect 27018 6679 27030 6735
rect 34548 6735 34604 7756
rect 35716 7748 35786 7756
rect 35212 7704 35298 7708
rect 35212 7648 35224 7704
rect 35280 7648 35298 7704
rect 35212 7636 35298 7648
rect 34723 7491 34769 7502
rect 34938 7500 35014 7533
rect 34938 7454 34949 7500
rect 35003 7454 35014 7500
rect 35122 7500 35198 7533
rect 35122 7454 35133 7500
rect 35187 7454 35198 7500
rect 35306 7500 35382 7533
rect 35306 7454 35317 7500
rect 35371 7454 35382 7500
rect 35551 7491 35597 7502
rect 34861 7408 34907 7419
rect 34844 7381 34861 7383
rect 35045 7408 35091 7419
rect 34907 7381 34924 7383
rect 34769 7261 34856 7381
rect 34912 7261 34924 7381
rect 34844 7259 34861 7261
rect 34769 6961 34861 7081
rect 34907 7259 34924 7261
rect 35028 7081 35045 7083
rect 35229 7408 35275 7419
rect 35212 7381 35229 7383
rect 35413 7408 35459 7419
rect 35275 7381 35292 7383
rect 35212 7261 35224 7381
rect 35280 7261 35292 7381
rect 35212 7259 35229 7261
rect 35091 7081 35108 7083
rect 35028 6961 35040 7081
rect 35096 6961 35108 7081
rect 35028 6959 35045 6961
rect 34861 6923 34907 6934
rect 35091 6959 35108 6961
rect 35045 6923 35091 6934
rect 35275 7259 35292 7261
rect 35396 7081 35413 7083
rect 35534 7381 35551 7383
rect 35597 7381 35614 7383
rect 35534 7260 35546 7381
rect 35602 7260 35614 7381
rect 35534 7258 35551 7260
rect 35459 7081 35476 7083
rect 35396 6961 35408 7081
rect 35464 6961 35476 7081
rect 35396 6959 35413 6961
rect 35229 6923 35275 6934
rect 35459 6959 35476 6961
rect 35413 6923 35459 6934
rect 34938 6885 34949 6888
rect 35003 6885 35014 6888
rect 35122 6885 35133 6888
rect 35187 6885 35198 6888
rect 35306 6885 35317 6888
rect 35371 6885 35382 6888
rect 34723 6840 34769 6851
rect 34936 6829 34948 6885
rect 35004 6829 35016 6885
rect 34936 6815 35016 6829
rect 35120 6829 35132 6885
rect 35188 6829 35200 6885
rect 35120 6815 35200 6829
rect 35304 6829 35316 6885
rect 35372 6829 35384 6885
rect 35597 7258 35614 7260
rect 35551 6840 35597 6851
rect 35304 6815 35384 6829
rect 34936 6735 35016 6737
rect 34548 6679 34948 6735
rect 35004 6679 35016 6735
rect 36034 6735 36090 9961
rect 44015 9961 45562 10017
rect 43518 8940 43606 8952
rect 44015 8940 44071 9961
rect 44684 9909 44770 9913
rect 44684 9853 44696 9909
rect 44752 9853 44770 9909
rect 44684 9841 44770 9853
rect 44195 9696 44241 9707
rect 44410 9705 44486 9738
rect 44410 9659 44421 9705
rect 44475 9659 44486 9705
rect 44594 9705 44670 9738
rect 44594 9659 44605 9705
rect 44659 9659 44670 9705
rect 44778 9705 44854 9738
rect 44778 9659 44789 9705
rect 44843 9659 44854 9705
rect 45023 9696 45069 9707
rect 44333 9613 44379 9624
rect 44316 9586 44333 9588
rect 44517 9613 44563 9624
rect 44379 9586 44396 9588
rect 44241 9466 44328 9586
rect 44384 9466 44396 9586
rect 44316 9464 44333 9466
rect 44241 9166 44333 9286
rect 44379 9464 44396 9466
rect 44500 9286 44517 9288
rect 44701 9613 44747 9624
rect 44684 9586 44701 9588
rect 44885 9613 44931 9624
rect 44747 9586 44764 9588
rect 44684 9466 44696 9586
rect 44752 9466 44764 9586
rect 44684 9464 44701 9466
rect 44563 9286 44580 9288
rect 44500 9166 44512 9286
rect 44568 9166 44580 9286
rect 44500 9164 44517 9166
rect 44333 9128 44379 9139
rect 44563 9164 44580 9166
rect 44517 9128 44563 9139
rect 44747 9464 44764 9466
rect 44868 9286 44885 9288
rect 45006 9586 45023 9588
rect 45069 9586 45086 9588
rect 45006 9465 45018 9586
rect 45074 9465 45086 9586
rect 45006 9463 45023 9465
rect 44931 9286 44948 9288
rect 44868 9166 44880 9286
rect 44936 9166 44948 9286
rect 44868 9164 44885 9166
rect 44701 9128 44747 9139
rect 44931 9164 44948 9166
rect 44885 9128 44931 9139
rect 44410 9090 44421 9093
rect 44475 9090 44486 9093
rect 44594 9090 44605 9093
rect 44659 9090 44670 9093
rect 44778 9090 44789 9093
rect 44843 9090 44854 9093
rect 44195 9045 44241 9056
rect 44408 9034 44420 9090
rect 44476 9034 44488 9090
rect 44408 9020 44488 9034
rect 44592 9034 44604 9090
rect 44660 9034 44672 9090
rect 44592 9020 44672 9034
rect 44776 9034 44788 9090
rect 44844 9034 44856 9090
rect 45069 9463 45086 9465
rect 45023 9045 45069 9056
rect 44776 9020 44856 9034
rect 44408 8940 44488 8942
rect 43518 8884 43532 8940
rect 43588 8884 44420 8940
rect 44476 8884 44488 8940
rect 43518 8872 43606 8884
rect 44408 8882 44488 8884
rect 43736 8824 43806 8836
rect 44592 8824 44672 8826
rect 43736 8768 43748 8824
rect 43804 8768 44604 8824
rect 44660 8768 44672 8824
rect 43736 8756 43806 8768
rect 44592 8766 44672 8768
rect 44921 8824 45001 8826
rect 45188 8824 45258 8836
rect 44921 8768 44933 8824
rect 44989 8768 45190 8824
rect 45246 8768 45258 8824
rect 44921 8766 45001 8768
rect 45188 8758 45258 8768
rect 44776 8708 44856 8710
rect 44020 8652 44788 8708
rect 44844 8652 44856 8708
rect 44020 7921 44076 8652
rect 44776 8650 44856 8652
rect 44408 8558 44488 8572
rect 44195 8536 44241 8547
rect 44408 8502 44420 8558
rect 44476 8502 44488 8558
rect 44592 8558 44672 8572
rect 44592 8502 44604 8558
rect 44660 8502 44672 8558
rect 44776 8558 44856 8572
rect 44776 8502 44788 8558
rect 44844 8502 44856 8558
rect 45023 8536 45069 8547
rect 44410 8499 44421 8502
rect 44475 8499 44486 8502
rect 44594 8499 44605 8502
rect 44659 8499 44670 8502
rect 44778 8499 44789 8502
rect 44843 8499 44854 8502
rect 44333 8453 44379 8464
rect 44241 8279 44333 8453
rect 44333 8268 44379 8279
rect 44517 8453 44563 8464
rect 44517 8268 44563 8279
rect 44701 8453 44747 8464
rect 44885 8453 44931 8464
rect 44868 8426 44885 8428
rect 44931 8426 44948 8428
rect 44868 8306 44880 8426
rect 44936 8306 44948 8426
rect 44868 8304 44885 8306
rect 44701 8268 44747 8279
rect 44931 8304 44948 8306
rect 44885 8268 44931 8279
rect 44195 8051 44241 8196
rect 44410 8187 44421 8233
rect 44475 8187 44486 8233
rect 44410 8154 44486 8187
rect 44594 8187 44605 8233
rect 44659 8187 44670 8233
rect 44594 8154 44670 8187
rect 44778 8187 44789 8233
rect 44843 8187 44854 8233
rect 44778 8154 44854 8187
rect 45023 8051 45069 8196
rect 44183 8039 44263 8051
rect 44183 7983 44195 8039
rect 44251 7983 44263 8039
rect 44183 7971 44263 7983
rect 45001 8039 45081 8051
rect 45001 7983 45013 8039
rect 45069 7983 45081 8039
rect 45001 7971 45081 7983
rect 45354 7921 45434 7931
rect 44020 7865 45366 7921
rect 45422 7865 45434 7921
rect 45354 7863 45434 7865
rect 45188 7812 45258 7814
rect 44020 7811 45258 7812
rect 44020 7757 45190 7811
rect 45246 7757 45258 7811
rect 44020 7756 45258 7757
rect 36698 7704 36784 7708
rect 36698 7648 36710 7704
rect 36766 7648 36784 7704
rect 36698 7636 36784 7648
rect 36209 7491 36255 7502
rect 36424 7500 36500 7533
rect 36424 7454 36435 7500
rect 36489 7454 36500 7500
rect 36608 7500 36684 7533
rect 36608 7454 36619 7500
rect 36673 7454 36684 7500
rect 36792 7500 36868 7533
rect 36792 7454 36803 7500
rect 36857 7454 36868 7500
rect 37037 7491 37083 7502
rect 36347 7408 36393 7419
rect 36330 7381 36347 7383
rect 36531 7408 36577 7419
rect 36393 7381 36410 7383
rect 36255 7261 36342 7381
rect 36398 7261 36410 7381
rect 36330 7259 36347 7261
rect 36255 6961 36347 7081
rect 36393 7259 36410 7261
rect 36514 7081 36531 7083
rect 36715 7408 36761 7419
rect 36698 7381 36715 7383
rect 36899 7408 36945 7419
rect 36761 7381 36778 7383
rect 36698 7261 36710 7381
rect 36766 7261 36778 7381
rect 36698 7259 36715 7261
rect 36577 7081 36594 7083
rect 36514 6961 36526 7081
rect 36582 6961 36594 7081
rect 36514 6959 36531 6961
rect 36347 6923 36393 6934
rect 36577 6959 36594 6961
rect 36531 6923 36577 6934
rect 36761 7259 36778 7261
rect 36882 7081 36899 7083
rect 37020 7381 37037 7383
rect 37083 7381 37100 7383
rect 37020 7260 37032 7381
rect 37088 7260 37100 7381
rect 37020 7258 37037 7260
rect 36945 7081 36962 7083
rect 36882 6961 36894 7081
rect 36950 6961 36962 7081
rect 36882 6959 36899 6961
rect 36715 6923 36761 6934
rect 36945 6959 36962 6961
rect 36899 6923 36945 6934
rect 36424 6885 36435 6888
rect 36489 6885 36500 6888
rect 36608 6885 36619 6888
rect 36673 6885 36684 6888
rect 36792 6885 36803 6888
rect 36857 6885 36868 6888
rect 36209 6840 36255 6851
rect 36422 6829 36434 6885
rect 36490 6829 36502 6885
rect 36422 6815 36502 6829
rect 36606 6829 36618 6885
rect 36674 6829 36686 6885
rect 36606 6815 36686 6829
rect 36790 6829 36802 6885
rect 36858 6829 36870 6885
rect 37083 7258 37100 7260
rect 37037 6840 37083 6851
rect 36790 6815 36870 6829
rect 36422 6735 36502 6737
rect 36034 6679 36434 6735
rect 36490 6679 36502 6735
rect 44020 6735 44076 7756
rect 45188 7748 45258 7756
rect 44684 7704 44770 7708
rect 44684 7648 44696 7704
rect 44752 7648 44770 7704
rect 44684 7636 44770 7648
rect 44195 7491 44241 7502
rect 44410 7500 44486 7533
rect 44410 7454 44421 7500
rect 44475 7454 44486 7500
rect 44594 7500 44670 7533
rect 44594 7454 44605 7500
rect 44659 7454 44670 7500
rect 44778 7500 44854 7533
rect 44778 7454 44789 7500
rect 44843 7454 44854 7500
rect 45023 7491 45069 7502
rect 44333 7408 44379 7419
rect 44316 7381 44333 7383
rect 44517 7408 44563 7419
rect 44379 7381 44396 7383
rect 44241 7261 44328 7381
rect 44384 7261 44396 7381
rect 44316 7259 44333 7261
rect 44241 6961 44333 7081
rect 44379 7259 44396 7261
rect 44500 7081 44517 7083
rect 44701 7408 44747 7419
rect 44684 7381 44701 7383
rect 44885 7408 44931 7419
rect 44747 7381 44764 7383
rect 44684 7261 44696 7381
rect 44752 7261 44764 7381
rect 44684 7259 44701 7261
rect 44563 7081 44580 7083
rect 44500 6961 44512 7081
rect 44568 6961 44580 7081
rect 44500 6959 44517 6961
rect 44333 6923 44379 6934
rect 44563 6959 44580 6961
rect 44517 6923 44563 6934
rect 44747 7259 44764 7261
rect 44868 7081 44885 7083
rect 45006 7381 45023 7383
rect 45069 7381 45086 7383
rect 45006 7260 45018 7381
rect 45074 7260 45086 7381
rect 45006 7258 45023 7260
rect 44931 7081 44948 7083
rect 44868 6961 44880 7081
rect 44936 6961 44948 7081
rect 44868 6959 44885 6961
rect 44701 6923 44747 6934
rect 44931 6959 44948 6961
rect 44885 6923 44931 6934
rect 44410 6885 44421 6888
rect 44475 6885 44486 6888
rect 44594 6885 44605 6888
rect 44659 6885 44670 6888
rect 44778 6885 44789 6888
rect 44843 6885 44854 6888
rect 44195 6840 44241 6851
rect 44408 6829 44420 6885
rect 44476 6829 44488 6885
rect 44408 6815 44488 6829
rect 44592 6829 44604 6885
rect 44660 6829 44672 6885
rect 44592 6815 44672 6829
rect 44776 6829 44788 6885
rect 44844 6829 44856 6885
rect 45069 7258 45086 7260
rect 45023 6840 45069 6851
rect 44776 6815 44856 6829
rect 44408 6735 44488 6737
rect 44020 6679 44420 6735
rect 44476 6679 44488 6735
rect 45506 6735 45562 9961
rect 53487 9961 55034 10017
rect 52990 8940 53078 8952
rect 53487 8940 53543 9961
rect 54156 9909 54242 9913
rect 54156 9853 54168 9909
rect 54224 9853 54242 9909
rect 54156 9841 54242 9853
rect 53667 9696 53713 9707
rect 53882 9705 53958 9738
rect 53882 9659 53893 9705
rect 53947 9659 53958 9705
rect 54066 9705 54142 9738
rect 54066 9659 54077 9705
rect 54131 9659 54142 9705
rect 54250 9705 54326 9738
rect 54250 9659 54261 9705
rect 54315 9659 54326 9705
rect 54495 9696 54541 9707
rect 53805 9613 53851 9624
rect 53788 9586 53805 9588
rect 53989 9613 54035 9624
rect 53851 9586 53868 9588
rect 53713 9466 53800 9586
rect 53856 9466 53868 9586
rect 53788 9464 53805 9466
rect 53713 9166 53805 9286
rect 53851 9464 53868 9466
rect 53972 9286 53989 9288
rect 54173 9613 54219 9624
rect 54156 9586 54173 9588
rect 54357 9613 54403 9624
rect 54219 9586 54236 9588
rect 54156 9466 54168 9586
rect 54224 9466 54236 9586
rect 54156 9464 54173 9466
rect 54035 9286 54052 9288
rect 53972 9166 53984 9286
rect 54040 9166 54052 9286
rect 53972 9164 53989 9166
rect 53805 9128 53851 9139
rect 54035 9164 54052 9166
rect 53989 9128 54035 9139
rect 54219 9464 54236 9466
rect 54340 9286 54357 9288
rect 54478 9586 54495 9588
rect 54541 9586 54558 9588
rect 54478 9465 54490 9586
rect 54546 9465 54558 9586
rect 54478 9463 54495 9465
rect 54403 9286 54420 9288
rect 54340 9166 54352 9286
rect 54408 9166 54420 9286
rect 54340 9164 54357 9166
rect 54173 9128 54219 9139
rect 54403 9164 54420 9166
rect 54357 9128 54403 9139
rect 53882 9090 53893 9093
rect 53947 9090 53958 9093
rect 54066 9090 54077 9093
rect 54131 9090 54142 9093
rect 54250 9090 54261 9093
rect 54315 9090 54326 9093
rect 53667 9045 53713 9056
rect 53880 9034 53892 9090
rect 53948 9034 53960 9090
rect 53880 9020 53960 9034
rect 54064 9034 54076 9090
rect 54132 9034 54144 9090
rect 54064 9020 54144 9034
rect 54248 9034 54260 9090
rect 54316 9034 54328 9090
rect 54541 9463 54558 9465
rect 54495 9045 54541 9056
rect 54248 9020 54328 9034
rect 53880 8940 53960 8942
rect 52990 8884 53004 8940
rect 53060 8884 53892 8940
rect 53948 8884 53960 8940
rect 52990 8872 53078 8884
rect 53880 8882 53960 8884
rect 53208 8824 53278 8836
rect 54064 8824 54144 8826
rect 53208 8768 53220 8824
rect 53276 8768 54076 8824
rect 54132 8768 54144 8824
rect 53208 8756 53278 8768
rect 54064 8766 54144 8768
rect 54393 8824 54473 8826
rect 54660 8824 54730 8836
rect 54393 8768 54405 8824
rect 54461 8768 54662 8824
rect 54718 8768 54730 8824
rect 54393 8766 54473 8768
rect 54660 8758 54730 8768
rect 54248 8708 54328 8710
rect 53492 8652 54260 8708
rect 54316 8652 54328 8708
rect 53492 7921 53548 8652
rect 54248 8650 54328 8652
rect 53880 8558 53960 8572
rect 53667 8536 53713 8547
rect 53880 8502 53892 8558
rect 53948 8502 53960 8558
rect 54064 8558 54144 8572
rect 54064 8502 54076 8558
rect 54132 8502 54144 8558
rect 54248 8558 54328 8572
rect 54248 8502 54260 8558
rect 54316 8502 54328 8558
rect 54495 8536 54541 8547
rect 53882 8499 53893 8502
rect 53947 8499 53958 8502
rect 54066 8499 54077 8502
rect 54131 8499 54142 8502
rect 54250 8499 54261 8502
rect 54315 8499 54326 8502
rect 53805 8453 53851 8464
rect 53713 8279 53805 8453
rect 53805 8268 53851 8279
rect 53989 8453 54035 8464
rect 53989 8268 54035 8279
rect 54173 8453 54219 8464
rect 54357 8453 54403 8464
rect 54340 8426 54357 8428
rect 54403 8426 54420 8428
rect 54340 8306 54352 8426
rect 54408 8306 54420 8426
rect 54340 8304 54357 8306
rect 54173 8268 54219 8279
rect 54403 8304 54420 8306
rect 54357 8268 54403 8279
rect 53667 8051 53713 8196
rect 53882 8187 53893 8233
rect 53947 8187 53958 8233
rect 53882 8154 53958 8187
rect 54066 8187 54077 8233
rect 54131 8187 54142 8233
rect 54066 8154 54142 8187
rect 54250 8187 54261 8233
rect 54315 8187 54326 8233
rect 54250 8154 54326 8187
rect 54495 8051 54541 8196
rect 53655 8039 53735 8051
rect 53655 7983 53667 8039
rect 53723 7983 53735 8039
rect 53655 7971 53735 7983
rect 54473 8039 54553 8051
rect 54473 7983 54485 8039
rect 54541 7983 54553 8039
rect 54473 7971 54553 7983
rect 54826 7921 54906 7931
rect 53492 7865 54838 7921
rect 54894 7865 54906 7921
rect 54826 7863 54906 7865
rect 54660 7812 54730 7814
rect 53492 7811 54730 7812
rect 53492 7757 54662 7811
rect 54718 7757 54730 7811
rect 53492 7756 54730 7757
rect 46170 7704 46256 7708
rect 46170 7648 46182 7704
rect 46238 7648 46256 7704
rect 46170 7636 46256 7648
rect 45681 7491 45727 7502
rect 45896 7500 45972 7533
rect 45896 7454 45907 7500
rect 45961 7454 45972 7500
rect 46080 7500 46156 7533
rect 46080 7454 46091 7500
rect 46145 7454 46156 7500
rect 46264 7500 46340 7533
rect 46264 7454 46275 7500
rect 46329 7454 46340 7500
rect 46509 7491 46555 7502
rect 45819 7408 45865 7419
rect 45802 7381 45819 7383
rect 46003 7408 46049 7419
rect 45865 7381 45882 7383
rect 45727 7261 45814 7381
rect 45870 7261 45882 7381
rect 45802 7259 45819 7261
rect 45727 6961 45819 7081
rect 45865 7259 45882 7261
rect 45986 7081 46003 7083
rect 46187 7408 46233 7419
rect 46170 7381 46187 7383
rect 46371 7408 46417 7419
rect 46233 7381 46250 7383
rect 46170 7261 46182 7381
rect 46238 7261 46250 7381
rect 46170 7259 46187 7261
rect 46049 7081 46066 7083
rect 45986 6961 45998 7081
rect 46054 6961 46066 7081
rect 45986 6959 46003 6961
rect 45819 6923 45865 6934
rect 46049 6959 46066 6961
rect 46003 6923 46049 6934
rect 46233 7259 46250 7261
rect 46354 7081 46371 7083
rect 46492 7381 46509 7383
rect 46555 7381 46572 7383
rect 46492 7260 46504 7381
rect 46560 7260 46572 7381
rect 46492 7258 46509 7260
rect 46417 7081 46434 7083
rect 46354 6961 46366 7081
rect 46422 6961 46434 7081
rect 46354 6959 46371 6961
rect 46187 6923 46233 6934
rect 46417 6959 46434 6961
rect 46371 6923 46417 6934
rect 45896 6885 45907 6888
rect 45961 6885 45972 6888
rect 46080 6885 46091 6888
rect 46145 6885 46156 6888
rect 46264 6885 46275 6888
rect 46329 6885 46340 6888
rect 45681 6840 45727 6851
rect 45894 6829 45906 6885
rect 45962 6829 45974 6885
rect 45894 6815 45974 6829
rect 46078 6829 46090 6885
rect 46146 6829 46158 6885
rect 46078 6815 46158 6829
rect 46262 6829 46274 6885
rect 46330 6829 46342 6885
rect 46555 7258 46572 7260
rect 46509 6840 46555 6851
rect 46262 6815 46342 6829
rect 45894 6735 45974 6737
rect 45506 6679 45906 6735
rect 45962 6679 45974 6735
rect 53492 6735 53548 7756
rect 54660 7748 54730 7756
rect 54156 7704 54242 7708
rect 54156 7648 54168 7704
rect 54224 7648 54242 7704
rect 54156 7636 54242 7648
rect 53667 7491 53713 7502
rect 53882 7500 53958 7533
rect 53882 7454 53893 7500
rect 53947 7454 53958 7500
rect 54066 7500 54142 7533
rect 54066 7454 54077 7500
rect 54131 7454 54142 7500
rect 54250 7500 54326 7533
rect 54250 7454 54261 7500
rect 54315 7454 54326 7500
rect 54495 7491 54541 7502
rect 53805 7408 53851 7419
rect 53788 7381 53805 7383
rect 53989 7408 54035 7419
rect 53851 7381 53868 7383
rect 53713 7261 53800 7381
rect 53856 7261 53868 7381
rect 53788 7259 53805 7261
rect 53713 6961 53805 7081
rect 53851 7259 53868 7261
rect 53972 7081 53989 7083
rect 54173 7408 54219 7419
rect 54156 7381 54173 7383
rect 54357 7408 54403 7419
rect 54219 7381 54236 7383
rect 54156 7261 54168 7381
rect 54224 7261 54236 7381
rect 54156 7259 54173 7261
rect 54035 7081 54052 7083
rect 53972 6961 53984 7081
rect 54040 6961 54052 7081
rect 53972 6959 53989 6961
rect 53805 6923 53851 6934
rect 54035 6959 54052 6961
rect 53989 6923 54035 6934
rect 54219 7259 54236 7261
rect 54340 7081 54357 7083
rect 54478 7381 54495 7383
rect 54541 7381 54558 7383
rect 54478 7260 54490 7381
rect 54546 7260 54558 7381
rect 54478 7258 54495 7260
rect 54403 7081 54420 7083
rect 54340 6961 54352 7081
rect 54408 6961 54420 7081
rect 54340 6959 54357 6961
rect 54173 6923 54219 6934
rect 54403 6959 54420 6961
rect 54357 6923 54403 6934
rect 53882 6885 53893 6888
rect 53947 6885 53958 6888
rect 54066 6885 54077 6888
rect 54131 6885 54142 6888
rect 54250 6885 54261 6888
rect 54315 6885 54326 6888
rect 53667 6840 53713 6851
rect 53880 6829 53892 6885
rect 53948 6829 53960 6885
rect 53880 6815 53960 6829
rect 54064 6829 54076 6885
rect 54132 6829 54144 6885
rect 54064 6815 54144 6829
rect 54248 6829 54260 6885
rect 54316 6829 54328 6885
rect 54541 7258 54558 7260
rect 54495 6840 54541 6851
rect 54248 6815 54328 6829
rect 53880 6735 53960 6737
rect 53492 6679 53892 6735
rect 53948 6679 53960 6735
rect 54978 6735 55034 9961
rect 55642 7704 55728 7708
rect 55642 7648 55654 7704
rect 55710 7648 55728 7704
rect 55642 7636 55728 7648
rect 55153 7491 55199 7502
rect 55368 7500 55444 7533
rect 55368 7454 55379 7500
rect 55433 7454 55444 7500
rect 55552 7500 55628 7533
rect 55552 7454 55563 7500
rect 55617 7454 55628 7500
rect 55736 7500 55812 7533
rect 55736 7454 55747 7500
rect 55801 7454 55812 7500
rect 55981 7491 56027 7502
rect 55291 7408 55337 7419
rect 55274 7381 55291 7383
rect 55475 7408 55521 7419
rect 55337 7381 55354 7383
rect 55199 7261 55286 7381
rect 55342 7261 55354 7381
rect 55274 7259 55291 7261
rect 55199 6961 55291 7081
rect 55337 7259 55354 7261
rect 55458 7081 55475 7083
rect 55659 7408 55705 7419
rect 55642 7381 55659 7383
rect 55843 7408 55889 7419
rect 55705 7381 55722 7383
rect 55642 7261 55654 7381
rect 55710 7261 55722 7381
rect 55642 7259 55659 7261
rect 55521 7081 55538 7083
rect 55458 6961 55470 7081
rect 55526 6961 55538 7081
rect 55458 6959 55475 6961
rect 55291 6923 55337 6934
rect 55521 6959 55538 6961
rect 55475 6923 55521 6934
rect 55705 7259 55722 7261
rect 55826 7081 55843 7083
rect 55964 7381 55981 7383
rect 56027 7381 56044 7383
rect 55964 7260 55976 7381
rect 56032 7260 56044 7381
rect 55964 7258 55981 7260
rect 55889 7081 55906 7083
rect 55826 6961 55838 7081
rect 55894 6961 55906 7081
rect 55826 6959 55843 6961
rect 55659 6923 55705 6934
rect 55889 6959 55906 6961
rect 55843 6923 55889 6934
rect 55368 6885 55379 6888
rect 55433 6885 55444 6888
rect 55552 6885 55563 6888
rect 55617 6885 55628 6888
rect 55736 6885 55747 6888
rect 55801 6885 55812 6888
rect 55153 6840 55199 6851
rect 55366 6829 55378 6885
rect 55434 6829 55446 6885
rect 55366 6815 55446 6829
rect 55550 6829 55562 6885
rect 55618 6829 55630 6885
rect 55550 6815 55630 6829
rect 55734 6829 55746 6885
rect 55802 6829 55814 6885
rect 56027 7258 56044 7260
rect 55981 6840 56027 6851
rect 55734 6815 55814 6829
rect 55366 6735 55446 6737
rect 54978 6679 55378 6735
rect 55434 6679 55446 6735
rect 6520 6676 6600 6678
rect 8006 6676 8086 6678
rect 15992 6676 16072 6678
rect 17478 6676 17558 6678
rect 25464 6677 25544 6679
rect 26950 6677 27030 6679
rect 34936 6677 35016 6679
rect 36422 6677 36502 6679
rect 44408 6677 44488 6679
rect 45894 6677 45974 6679
rect 53880 6677 53960 6679
rect 55366 6677 55446 6679
rect 5712 6618 5782 6632
rect 6704 6618 6784 6620
rect 5712 6562 5724 6618
rect 5780 6562 6716 6618
rect 6772 6562 6784 6618
rect 5712 6550 5782 6562
rect 6704 6560 6784 6562
rect 7033 6618 7113 6620
rect 7476 6618 7536 6628
rect 8190 6618 8270 6620
rect 7033 6562 7045 6618
rect 7101 6562 7478 6618
rect 7534 6562 8202 6618
rect 8258 6562 8270 6618
rect 7033 6560 7113 6562
rect 7476 6550 7536 6562
rect 8190 6560 8270 6562
rect 8519 6618 8599 6620
rect 8786 6618 8856 6630
rect 8519 6562 8531 6618
rect 8587 6562 8788 6618
rect 8844 6562 8856 6618
rect 8519 6560 8599 6562
rect 8786 6552 8856 6562
rect 15184 6618 15254 6632
rect 16176 6618 16256 6620
rect 15184 6562 15196 6618
rect 15252 6562 16188 6618
rect 16244 6562 16256 6618
rect 15184 6550 15254 6562
rect 16176 6560 16256 6562
rect 16505 6618 16585 6620
rect 16948 6618 17008 6628
rect 17662 6618 17742 6620
rect 16505 6562 16517 6618
rect 16573 6562 16950 6618
rect 17006 6562 17674 6618
rect 17730 6562 17742 6618
rect 16505 6560 16585 6562
rect 16948 6550 17008 6562
rect 17662 6560 17742 6562
rect 17991 6618 18071 6620
rect 18258 6618 18328 6630
rect 17991 6562 18003 6618
rect 18059 6562 18260 6618
rect 18316 6562 18328 6618
rect 17991 6560 18071 6562
rect 18258 6552 18328 6562
rect 24656 6619 24726 6633
rect 25648 6619 25728 6621
rect 24656 6563 24668 6619
rect 24724 6563 25660 6619
rect 25716 6563 25728 6619
rect 24656 6551 24726 6563
rect 25648 6561 25728 6563
rect 25977 6619 26057 6621
rect 26420 6619 26480 6629
rect 27134 6619 27214 6621
rect 25977 6563 25989 6619
rect 26045 6563 26422 6619
rect 26478 6563 27146 6619
rect 27202 6563 27214 6619
rect 25977 6561 26057 6563
rect 26420 6551 26480 6563
rect 27134 6561 27214 6563
rect 27463 6619 27543 6621
rect 27730 6619 27800 6631
rect 27463 6563 27475 6619
rect 27531 6563 27732 6619
rect 27788 6563 27800 6619
rect 27463 6561 27543 6563
rect 27730 6553 27800 6563
rect 34128 6619 34198 6633
rect 35120 6619 35200 6621
rect 34128 6563 34140 6619
rect 34196 6563 35132 6619
rect 35188 6563 35200 6619
rect 34128 6551 34198 6563
rect 35120 6561 35200 6563
rect 35449 6619 35529 6621
rect 35892 6619 35952 6629
rect 36606 6619 36686 6621
rect 35449 6563 35461 6619
rect 35517 6563 35894 6619
rect 35950 6563 36618 6619
rect 36674 6563 36686 6619
rect 35449 6561 35529 6563
rect 35892 6551 35952 6563
rect 36606 6561 36686 6563
rect 36935 6619 37015 6621
rect 37202 6619 37272 6631
rect 36935 6563 36947 6619
rect 37003 6563 37204 6619
rect 37260 6563 37272 6619
rect 36935 6561 37015 6563
rect 37202 6553 37272 6563
rect 43600 6619 43670 6633
rect 44592 6619 44672 6621
rect 43600 6563 43612 6619
rect 43668 6563 44604 6619
rect 44660 6563 44672 6619
rect 43600 6551 43670 6563
rect 44592 6561 44672 6563
rect 44921 6619 45001 6621
rect 45364 6619 45424 6629
rect 46078 6619 46158 6621
rect 44921 6563 44933 6619
rect 44989 6563 45366 6619
rect 45422 6563 46090 6619
rect 46146 6563 46158 6619
rect 44921 6561 45001 6563
rect 45364 6551 45424 6563
rect 46078 6561 46158 6563
rect 46407 6619 46487 6621
rect 46674 6619 46744 6631
rect 46407 6563 46419 6619
rect 46475 6563 46676 6619
rect 46732 6563 46744 6619
rect 46407 6561 46487 6563
rect 46674 6553 46744 6563
rect 53072 6619 53142 6633
rect 54064 6619 54144 6621
rect 53072 6563 53084 6619
rect 53140 6563 54076 6619
rect 54132 6563 54144 6619
rect 53072 6551 53142 6563
rect 54064 6561 54144 6563
rect 54393 6619 54473 6621
rect 54836 6619 54896 6629
rect 55550 6619 55630 6621
rect 54393 6563 54405 6619
rect 54461 6563 54838 6619
rect 54894 6563 55562 6619
rect 55618 6563 55630 6619
rect 54393 6561 54473 6563
rect 54836 6551 54896 6563
rect 55550 6561 55630 6563
rect 55879 6619 55959 6621
rect 56146 6619 56216 6631
rect 55879 6563 55891 6619
rect 55947 6563 56148 6619
rect 56204 6563 56216 6619
rect 55879 6561 55959 6563
rect 56146 6553 56216 6563
rect 6888 6502 6968 6504
rect 8374 6502 8454 6504
rect 16360 6502 16440 6504
rect 17846 6502 17926 6504
rect 25832 6503 25912 6505
rect 27318 6503 27398 6505
rect 35304 6503 35384 6505
rect 36790 6503 36870 6505
rect 44776 6503 44856 6505
rect 46262 6503 46342 6505
rect 54248 6503 54328 6505
rect 55734 6503 55814 6505
rect 5996 6446 6900 6502
rect 6956 6446 6968 6502
rect 5430 5716 5512 5728
rect 5996 5716 6052 6446
rect 6888 6444 6968 6446
rect 7618 6446 8386 6502
rect 8442 6446 8454 6502
rect 6520 6352 6600 6366
rect 6307 6330 6353 6341
rect 6520 6296 6532 6352
rect 6588 6296 6600 6352
rect 6704 6352 6784 6366
rect 6704 6296 6716 6352
rect 6772 6296 6784 6352
rect 6888 6352 6968 6366
rect 6888 6296 6900 6352
rect 6956 6296 6968 6352
rect 7135 6330 7181 6341
rect 6522 6293 6533 6296
rect 6587 6293 6598 6296
rect 6706 6293 6717 6296
rect 6771 6293 6782 6296
rect 6890 6293 6901 6296
rect 6955 6293 6966 6296
rect 6445 6247 6491 6258
rect 6353 6073 6445 6247
rect 6445 6062 6491 6073
rect 6629 6247 6675 6258
rect 6629 6062 6675 6073
rect 6813 6247 6859 6258
rect 6997 6247 7043 6258
rect 6980 6220 6997 6222
rect 7043 6220 7060 6222
rect 6980 6100 6992 6220
rect 7048 6100 7060 6220
rect 6980 6098 6997 6100
rect 6813 6062 6859 6073
rect 7043 6098 7060 6100
rect 6997 6062 7043 6073
rect 6307 5845 6353 5990
rect 6522 5981 6533 6027
rect 6587 5981 6598 6027
rect 6522 5948 6598 5981
rect 6706 5981 6717 6027
rect 6771 5981 6782 6027
rect 6706 5948 6782 5981
rect 6890 5981 6901 6027
rect 6955 5981 6966 6027
rect 6890 5948 6966 5981
rect 7135 5845 7181 5990
rect 6295 5833 6375 5845
rect 6295 5777 6307 5833
rect 6363 5777 6375 5833
rect 6295 5765 6375 5777
rect 7113 5833 7191 5845
rect 7113 5777 7125 5833
rect 7181 5777 7191 5833
rect 7113 5765 7191 5777
rect 5430 5660 5444 5716
rect 5500 5660 6052 5716
rect 7618 5716 7674 6446
rect 8374 6444 8454 6446
rect 15468 6446 16372 6502
rect 16428 6446 16440 6502
rect 8006 6352 8086 6366
rect 7793 6330 7839 6341
rect 8006 6296 8018 6352
rect 8074 6296 8086 6352
rect 8190 6352 8270 6366
rect 8190 6296 8202 6352
rect 8258 6296 8270 6352
rect 8374 6352 8454 6366
rect 8374 6296 8386 6352
rect 8442 6296 8454 6352
rect 8621 6330 8667 6341
rect 8008 6293 8019 6296
rect 8073 6293 8084 6296
rect 8192 6293 8203 6296
rect 8257 6293 8268 6296
rect 8376 6293 8387 6296
rect 8441 6293 8452 6296
rect 7931 6247 7977 6258
rect 7839 6073 7931 6247
rect 7931 6062 7977 6073
rect 8115 6247 8161 6258
rect 8115 6062 8161 6073
rect 8299 6247 8345 6258
rect 8483 6247 8529 6258
rect 8466 6220 8483 6222
rect 8529 6220 8546 6222
rect 8466 6100 8478 6220
rect 8534 6100 8546 6220
rect 8466 6098 8483 6100
rect 8299 6062 8345 6073
rect 8529 6098 8546 6100
rect 8483 6062 8529 6073
rect 7793 5845 7839 5990
rect 8008 5981 8019 6027
rect 8073 5981 8084 6027
rect 8008 5948 8084 5981
rect 8192 5981 8203 6027
rect 8257 5981 8268 6027
rect 8192 5948 8268 5981
rect 8376 5981 8387 6027
rect 8441 5981 8452 6027
rect 8376 5948 8452 5981
rect 8621 5845 8667 5990
rect 7781 5833 7861 5845
rect 7781 5777 7793 5833
rect 7849 5777 7861 5833
rect 7781 5765 7861 5777
rect 8599 5833 8677 5845
rect 8599 5777 8611 5833
rect 8667 5777 8677 5833
rect 8599 5765 8677 5777
rect 8952 5716 9032 5726
rect 7618 5660 8964 5716
rect 9020 5660 9032 5716
rect 5430 5648 5512 5660
rect 230 4310 5324 4510
rect 5996 4413 6052 5660
rect 8952 5658 9032 5660
rect 14902 5716 14984 5728
rect 15468 5716 15524 6446
rect 16360 6444 16440 6446
rect 17090 6446 17858 6502
rect 17914 6446 17926 6502
rect 15992 6352 16072 6366
rect 15779 6330 15825 6341
rect 15992 6296 16004 6352
rect 16060 6296 16072 6352
rect 16176 6352 16256 6366
rect 16176 6296 16188 6352
rect 16244 6296 16256 6352
rect 16360 6352 16440 6366
rect 16360 6296 16372 6352
rect 16428 6296 16440 6352
rect 16607 6330 16653 6341
rect 15994 6293 16005 6296
rect 16059 6293 16070 6296
rect 16178 6293 16189 6296
rect 16243 6293 16254 6296
rect 16362 6293 16373 6296
rect 16427 6293 16438 6296
rect 15917 6247 15963 6258
rect 15825 6073 15917 6247
rect 15917 6062 15963 6073
rect 16101 6247 16147 6258
rect 16101 6062 16147 6073
rect 16285 6247 16331 6258
rect 16469 6247 16515 6258
rect 16452 6220 16469 6222
rect 16515 6220 16532 6222
rect 16452 6100 16464 6220
rect 16520 6100 16532 6220
rect 16452 6098 16469 6100
rect 16285 6062 16331 6073
rect 16515 6098 16532 6100
rect 16469 6062 16515 6073
rect 15779 5845 15825 5990
rect 15994 5981 16005 6027
rect 16059 5981 16070 6027
rect 15994 5948 16070 5981
rect 16178 5981 16189 6027
rect 16243 5981 16254 6027
rect 16178 5948 16254 5981
rect 16362 5981 16373 6027
rect 16427 5981 16438 6027
rect 16362 5948 16438 5981
rect 16607 5845 16653 5990
rect 15767 5833 15847 5845
rect 15767 5777 15779 5833
rect 15835 5777 15847 5833
rect 15767 5765 15847 5777
rect 16585 5833 16663 5845
rect 16585 5777 16597 5833
rect 16653 5777 16663 5833
rect 16585 5765 16663 5777
rect 14902 5660 14916 5716
rect 14972 5660 15524 5716
rect 17090 5716 17146 6446
rect 17846 6444 17926 6446
rect 24940 6447 25844 6503
rect 25900 6447 25912 6503
rect 17478 6352 17558 6366
rect 17265 6330 17311 6341
rect 17478 6296 17490 6352
rect 17546 6296 17558 6352
rect 17662 6352 17742 6366
rect 17662 6296 17674 6352
rect 17730 6296 17742 6352
rect 17846 6352 17926 6366
rect 17846 6296 17858 6352
rect 17914 6296 17926 6352
rect 18093 6330 18139 6341
rect 17480 6293 17491 6296
rect 17545 6293 17556 6296
rect 17664 6293 17675 6296
rect 17729 6293 17740 6296
rect 17848 6293 17859 6296
rect 17913 6293 17924 6296
rect 17403 6247 17449 6258
rect 17311 6073 17403 6247
rect 17403 6062 17449 6073
rect 17587 6247 17633 6258
rect 17587 6062 17633 6073
rect 17771 6247 17817 6258
rect 17955 6247 18001 6258
rect 17938 6220 17955 6222
rect 18001 6220 18018 6222
rect 17938 6100 17950 6220
rect 18006 6100 18018 6220
rect 17938 6098 17955 6100
rect 17771 6062 17817 6073
rect 18001 6098 18018 6100
rect 17955 6062 18001 6073
rect 17265 5845 17311 5990
rect 17480 5981 17491 6027
rect 17545 5981 17556 6027
rect 17480 5948 17556 5981
rect 17664 5981 17675 6027
rect 17729 5981 17740 6027
rect 17664 5948 17740 5981
rect 17848 5981 17859 6027
rect 17913 5981 17924 6027
rect 17848 5948 17924 5981
rect 18093 5845 18139 5990
rect 17253 5833 17333 5845
rect 17253 5777 17265 5833
rect 17321 5777 17333 5833
rect 17253 5765 17333 5777
rect 18071 5833 18149 5845
rect 18071 5777 18083 5833
rect 18139 5777 18149 5833
rect 18071 5765 18149 5777
rect 18424 5716 18504 5726
rect 17090 5660 18436 5716
rect 18492 5660 18504 5716
rect 14902 5648 14984 5660
rect 7476 5605 7546 5607
rect 8776 5606 8856 5608
rect 6132 5549 7478 5605
rect 7534 5549 7546 5605
rect 6132 4529 6188 5549
rect 7476 5537 7546 5549
rect 7618 5550 8788 5606
rect 8844 5550 8856 5606
rect 6796 5498 6882 5502
rect 6796 5442 6808 5498
rect 6864 5442 6882 5498
rect 6796 5430 6882 5442
rect 6307 5285 6353 5296
rect 6522 5294 6598 5327
rect 6522 5248 6533 5294
rect 6587 5248 6598 5294
rect 6706 5294 6782 5327
rect 6706 5248 6717 5294
rect 6771 5248 6782 5294
rect 6890 5294 6966 5327
rect 6890 5248 6901 5294
rect 6955 5248 6966 5294
rect 7135 5285 7181 5296
rect 6445 5202 6491 5213
rect 6428 5175 6445 5177
rect 6629 5202 6675 5213
rect 6491 5175 6508 5177
rect 6353 5055 6440 5175
rect 6496 5055 6508 5175
rect 6428 5053 6445 5055
rect 6353 4755 6445 4875
rect 6491 5053 6508 5055
rect 6612 4875 6629 4877
rect 6813 5202 6859 5213
rect 6796 5175 6813 5177
rect 6997 5202 7043 5213
rect 6859 5175 6876 5177
rect 6796 5055 6808 5175
rect 6864 5055 6876 5175
rect 6796 5053 6813 5055
rect 6675 4875 6692 4877
rect 6612 4755 6624 4875
rect 6680 4755 6692 4875
rect 6612 4753 6629 4755
rect 6445 4717 6491 4728
rect 6675 4753 6692 4755
rect 6629 4717 6675 4728
rect 6859 5053 6876 5055
rect 6980 4875 6997 4877
rect 7118 5175 7135 5177
rect 7181 5175 7198 5177
rect 7118 5054 7130 5175
rect 7186 5054 7198 5175
rect 7118 5052 7135 5054
rect 7043 4875 7060 4877
rect 6980 4755 6992 4875
rect 7048 4755 7060 4875
rect 6980 4753 6997 4755
rect 6813 4717 6859 4728
rect 7043 4753 7060 4755
rect 6997 4717 7043 4728
rect 6522 4679 6533 4682
rect 6587 4679 6598 4682
rect 6706 4679 6717 4682
rect 6771 4679 6782 4682
rect 6890 4679 6901 4682
rect 6955 4679 6966 4682
rect 6307 4634 6353 4645
rect 6520 4623 6532 4679
rect 6588 4623 6600 4679
rect 6520 4609 6600 4623
rect 6704 4623 6716 4679
rect 6772 4623 6784 4679
rect 6704 4609 6784 4623
rect 6888 4623 6900 4679
rect 6956 4623 6968 4679
rect 7181 5052 7198 5054
rect 7135 4634 7181 4645
rect 6888 4609 6968 4623
rect 6520 4529 6600 4531
rect 6132 4473 6532 4529
rect 6588 4473 6600 4529
rect 7618 4530 7674 5550
rect 8776 5538 8856 5550
rect 8282 5499 8368 5503
rect 8282 5443 8294 5499
rect 8350 5443 8368 5499
rect 8282 5431 8368 5443
rect 7793 5286 7839 5297
rect 8008 5295 8084 5328
rect 8008 5249 8019 5295
rect 8073 5249 8084 5295
rect 8192 5295 8268 5328
rect 8192 5249 8203 5295
rect 8257 5249 8268 5295
rect 8376 5295 8452 5328
rect 8376 5249 8387 5295
rect 8441 5249 8452 5295
rect 8621 5286 8667 5297
rect 7931 5203 7977 5214
rect 7914 5176 7931 5178
rect 8115 5203 8161 5214
rect 7977 5176 7994 5178
rect 7839 5056 7926 5176
rect 7982 5056 7994 5176
rect 7914 5054 7931 5056
rect 7839 4756 7931 4876
rect 7977 5054 7994 5056
rect 8098 4876 8115 4878
rect 8299 5203 8345 5214
rect 8282 5176 8299 5178
rect 8483 5203 8529 5214
rect 8345 5176 8362 5178
rect 8282 5056 8294 5176
rect 8350 5056 8362 5176
rect 8282 5054 8299 5056
rect 8161 4876 8178 4878
rect 8098 4756 8110 4876
rect 8166 4756 8178 4876
rect 8098 4754 8115 4756
rect 7931 4718 7977 4729
rect 8161 4754 8178 4756
rect 8115 4718 8161 4729
rect 8345 5054 8362 5056
rect 8466 4876 8483 4878
rect 8604 5176 8621 5178
rect 8667 5176 8684 5178
rect 8604 5055 8616 5176
rect 8672 5055 8684 5176
rect 8604 5053 8621 5055
rect 8529 4876 8546 4878
rect 8466 4756 8478 4876
rect 8534 4756 8546 4876
rect 8466 4754 8483 4756
rect 8299 4718 8345 4729
rect 8529 4754 8546 4756
rect 8483 4718 8529 4729
rect 8008 4680 8019 4683
rect 8073 4680 8084 4683
rect 8192 4680 8203 4683
rect 8257 4680 8268 4683
rect 8376 4680 8387 4683
rect 8441 4680 8452 4683
rect 7793 4635 7839 4646
rect 8006 4624 8018 4680
rect 8074 4624 8086 4680
rect 8006 4610 8086 4624
rect 8190 4624 8202 4680
rect 8258 4624 8270 4680
rect 8190 4610 8270 4624
rect 8374 4624 8386 4680
rect 8442 4624 8454 4680
rect 8667 5053 8684 5055
rect 8621 4635 8667 4646
rect 8374 4610 8454 4624
rect 8006 4530 8086 4532
rect 7618 4474 8018 4530
rect 8074 4474 8086 4530
rect 6520 4471 6600 4473
rect 8006 4472 8086 4474
rect 6704 4413 6784 4415
rect 5996 4357 6716 4413
rect 6772 4357 6784 4413
rect 6704 4355 6784 4357
rect 7033 4413 7113 4415
rect 7300 4414 7370 4425
rect 8190 4414 8270 4416
rect 7300 4413 8202 4414
rect 7033 4357 7045 4413
rect 7101 4357 7302 4413
rect 7358 4358 8202 4413
rect 8258 4358 8270 4414
rect 7358 4357 7618 4358
rect 7033 4355 7113 4357
rect 7300 4347 7370 4357
rect 8190 4356 8270 4358
rect 8519 4414 8599 4416
rect 8962 4414 9032 4424
rect 8519 4358 8531 4414
rect 8587 4358 8964 4414
rect 9020 4358 9032 4414
rect 8519 4356 8599 4358
rect 8962 4346 9032 4358
rect 230 2890 834 4310
rect 1165 4170 1211 4181
rect 1380 4179 1476 4210
rect 1380 4133 1391 4179
rect 1465 4133 1476 4179
rect 1645 4170 2099 4310
rect 1303 4087 1349 4098
rect 1286 3803 1303 3813
rect 1507 4087 1645 4098
rect 1349 3803 1366 3813
rect 1286 3563 1298 3803
rect 1354 3563 1366 3803
rect 1286 3553 1303 3563
rect 1349 3553 1366 3563
rect 1303 3502 1349 3513
rect 1553 3513 1645 4087
rect 1507 3502 1645 3513
rect 1165 3419 1211 3430
rect 1380 3421 1391 3467
rect 1465 3421 1476 3467
rect 940 3346 1020 3356
rect 940 3290 952 3346
rect 1008 3290 1020 3346
rect 940 3280 1020 3290
rect 1380 3346 1476 3421
rect 1691 3502 2053 4170
rect 1645 3419 1691 3430
rect 2268 4179 2364 4210
rect 2268 4133 2279 4179
rect 2353 4133 2364 4179
rect 2533 4170 2579 4310
rect 2099 4087 2237 4098
rect 2099 3513 2191 4087
rect 2395 4087 2441 4098
rect 2378 3803 2395 3813
rect 2441 3803 2458 3813
rect 2378 3563 2390 3803
rect 2446 3563 2458 3803
rect 2378 3553 2395 3563
rect 2099 3502 2237 3513
rect 2441 3553 2458 3563
rect 2395 3502 2441 3513
rect 2053 3419 2099 3430
rect 2268 3421 2279 3467
rect 2353 3421 2364 3467
rect 1380 3290 1400 3346
rect 1456 3290 1476 3346
rect 1380 3072 1476 3290
rect 2268 3202 2364 3421
rect 2748 4179 2844 4210
rect 2748 4133 2759 4179
rect 2833 4133 2844 4179
rect 3013 4170 3059 4310
rect 2579 4087 2717 4098
rect 2579 3513 2671 4087
rect 2875 4087 2921 4098
rect 2858 3803 2875 3813
rect 2921 3803 2938 3813
rect 2858 3563 2870 3803
rect 2926 3563 2938 3803
rect 2858 3553 2875 3563
rect 2579 3502 2717 3513
rect 2921 3553 2938 3563
rect 2875 3502 2921 3513
rect 2533 3419 2579 3430
rect 2748 3421 2759 3467
rect 2833 3421 2844 3467
rect 2748 3280 2844 3421
rect 3013 3419 3059 3430
rect 3356 3510 4824 4310
rect 5124 3510 5324 4310
rect 9706 4310 14796 4510
rect 15468 4413 15524 5660
rect 18424 5658 18504 5660
rect 24374 5717 24456 5729
rect 24940 5717 24996 6447
rect 25832 6445 25912 6447
rect 26562 6447 27330 6503
rect 27386 6447 27398 6503
rect 25464 6353 25544 6367
rect 25251 6331 25297 6342
rect 25464 6297 25476 6353
rect 25532 6297 25544 6353
rect 25648 6353 25728 6367
rect 25648 6297 25660 6353
rect 25716 6297 25728 6353
rect 25832 6353 25912 6367
rect 25832 6297 25844 6353
rect 25900 6297 25912 6353
rect 26079 6331 26125 6342
rect 25466 6294 25477 6297
rect 25531 6294 25542 6297
rect 25650 6294 25661 6297
rect 25715 6294 25726 6297
rect 25834 6294 25845 6297
rect 25899 6294 25910 6297
rect 25389 6248 25435 6259
rect 25297 6074 25389 6248
rect 25389 6063 25435 6074
rect 25573 6248 25619 6259
rect 25573 6063 25619 6074
rect 25757 6248 25803 6259
rect 25941 6248 25987 6259
rect 25924 6221 25941 6223
rect 25987 6221 26004 6223
rect 25924 6101 25936 6221
rect 25992 6101 26004 6221
rect 25924 6099 25941 6101
rect 25757 6063 25803 6074
rect 25987 6099 26004 6101
rect 25941 6063 25987 6074
rect 25251 5846 25297 5991
rect 25466 5982 25477 6028
rect 25531 5982 25542 6028
rect 25466 5949 25542 5982
rect 25650 5982 25661 6028
rect 25715 5982 25726 6028
rect 25650 5949 25726 5982
rect 25834 5982 25845 6028
rect 25899 5982 25910 6028
rect 25834 5949 25910 5982
rect 26079 5846 26125 5991
rect 25239 5834 25319 5846
rect 25239 5778 25251 5834
rect 25307 5778 25319 5834
rect 25239 5766 25319 5778
rect 26057 5834 26135 5846
rect 26057 5778 26069 5834
rect 26125 5778 26135 5834
rect 26057 5766 26135 5778
rect 24374 5661 24388 5717
rect 24444 5661 24996 5717
rect 26562 5717 26618 6447
rect 27318 6445 27398 6447
rect 34412 6447 35316 6503
rect 35372 6447 35384 6503
rect 26950 6353 27030 6367
rect 26737 6331 26783 6342
rect 26950 6297 26962 6353
rect 27018 6297 27030 6353
rect 27134 6353 27214 6367
rect 27134 6297 27146 6353
rect 27202 6297 27214 6353
rect 27318 6353 27398 6367
rect 27318 6297 27330 6353
rect 27386 6297 27398 6353
rect 27565 6331 27611 6342
rect 26952 6294 26963 6297
rect 27017 6294 27028 6297
rect 27136 6294 27147 6297
rect 27201 6294 27212 6297
rect 27320 6294 27331 6297
rect 27385 6294 27396 6297
rect 26875 6248 26921 6259
rect 26783 6074 26875 6248
rect 26875 6063 26921 6074
rect 27059 6248 27105 6259
rect 27059 6063 27105 6074
rect 27243 6248 27289 6259
rect 27427 6248 27473 6259
rect 27410 6221 27427 6223
rect 27473 6221 27490 6223
rect 27410 6101 27422 6221
rect 27478 6101 27490 6221
rect 27410 6099 27427 6101
rect 27243 6063 27289 6074
rect 27473 6099 27490 6101
rect 27427 6063 27473 6074
rect 26737 5846 26783 5991
rect 26952 5982 26963 6028
rect 27017 5982 27028 6028
rect 26952 5949 27028 5982
rect 27136 5982 27147 6028
rect 27201 5982 27212 6028
rect 27136 5949 27212 5982
rect 27320 5982 27331 6028
rect 27385 5982 27396 6028
rect 27320 5949 27396 5982
rect 27565 5846 27611 5991
rect 26725 5834 26805 5846
rect 26725 5778 26737 5834
rect 26793 5778 26805 5834
rect 26725 5766 26805 5778
rect 27543 5834 27621 5846
rect 27543 5778 27555 5834
rect 27611 5778 27621 5834
rect 27543 5766 27621 5778
rect 27896 5717 27976 5727
rect 26562 5661 27908 5717
rect 27964 5661 27976 5717
rect 24374 5649 24456 5661
rect 16948 5605 17018 5607
rect 18248 5606 18328 5608
rect 15604 5549 16950 5605
rect 17006 5549 17018 5605
rect 15604 4529 15660 5549
rect 16948 5537 17018 5549
rect 17090 5550 18260 5606
rect 18316 5550 18328 5606
rect 16268 5498 16354 5502
rect 16268 5442 16280 5498
rect 16336 5442 16354 5498
rect 16268 5430 16354 5442
rect 15779 5285 15825 5296
rect 15994 5294 16070 5327
rect 15994 5248 16005 5294
rect 16059 5248 16070 5294
rect 16178 5294 16254 5327
rect 16178 5248 16189 5294
rect 16243 5248 16254 5294
rect 16362 5294 16438 5327
rect 16362 5248 16373 5294
rect 16427 5248 16438 5294
rect 16607 5285 16653 5296
rect 15917 5202 15963 5213
rect 15900 5175 15917 5177
rect 16101 5202 16147 5213
rect 15963 5175 15980 5177
rect 15825 5055 15912 5175
rect 15968 5055 15980 5175
rect 15900 5053 15917 5055
rect 15825 4755 15917 4875
rect 15963 5053 15980 5055
rect 16084 4875 16101 4877
rect 16285 5202 16331 5213
rect 16268 5175 16285 5177
rect 16469 5202 16515 5213
rect 16331 5175 16348 5177
rect 16268 5055 16280 5175
rect 16336 5055 16348 5175
rect 16268 5053 16285 5055
rect 16147 4875 16164 4877
rect 16084 4755 16096 4875
rect 16152 4755 16164 4875
rect 16084 4753 16101 4755
rect 15917 4717 15963 4728
rect 16147 4753 16164 4755
rect 16101 4717 16147 4728
rect 16331 5053 16348 5055
rect 16452 4875 16469 4877
rect 16590 5175 16607 5177
rect 16653 5175 16670 5177
rect 16590 5054 16602 5175
rect 16658 5054 16670 5175
rect 16590 5052 16607 5054
rect 16515 4875 16532 4877
rect 16452 4755 16464 4875
rect 16520 4755 16532 4875
rect 16452 4753 16469 4755
rect 16285 4717 16331 4728
rect 16515 4753 16532 4755
rect 16469 4717 16515 4728
rect 15994 4679 16005 4682
rect 16059 4679 16070 4682
rect 16178 4679 16189 4682
rect 16243 4679 16254 4682
rect 16362 4679 16373 4682
rect 16427 4679 16438 4682
rect 15779 4634 15825 4645
rect 15992 4623 16004 4679
rect 16060 4623 16072 4679
rect 15992 4609 16072 4623
rect 16176 4623 16188 4679
rect 16244 4623 16256 4679
rect 16176 4609 16256 4623
rect 16360 4623 16372 4679
rect 16428 4623 16440 4679
rect 16653 5052 16670 5054
rect 16607 4634 16653 4645
rect 16360 4609 16440 4623
rect 15992 4529 16072 4531
rect 15604 4473 16004 4529
rect 16060 4473 16072 4529
rect 17090 4530 17146 5550
rect 18248 5538 18328 5550
rect 17754 5499 17840 5503
rect 17754 5443 17766 5499
rect 17822 5443 17840 5499
rect 17754 5431 17840 5443
rect 17265 5286 17311 5297
rect 17480 5295 17556 5328
rect 17480 5249 17491 5295
rect 17545 5249 17556 5295
rect 17664 5295 17740 5328
rect 17664 5249 17675 5295
rect 17729 5249 17740 5295
rect 17848 5295 17924 5328
rect 17848 5249 17859 5295
rect 17913 5249 17924 5295
rect 18093 5286 18139 5297
rect 17403 5203 17449 5214
rect 17386 5176 17403 5178
rect 17587 5203 17633 5214
rect 17449 5176 17466 5178
rect 17311 5056 17398 5176
rect 17454 5056 17466 5176
rect 17386 5054 17403 5056
rect 17311 4756 17403 4876
rect 17449 5054 17466 5056
rect 17570 4876 17587 4878
rect 17771 5203 17817 5214
rect 17754 5176 17771 5178
rect 17955 5203 18001 5214
rect 17817 5176 17834 5178
rect 17754 5056 17766 5176
rect 17822 5056 17834 5176
rect 17754 5054 17771 5056
rect 17633 4876 17650 4878
rect 17570 4756 17582 4876
rect 17638 4756 17650 4876
rect 17570 4754 17587 4756
rect 17403 4718 17449 4729
rect 17633 4754 17650 4756
rect 17587 4718 17633 4729
rect 17817 5054 17834 5056
rect 17938 4876 17955 4878
rect 18076 5176 18093 5178
rect 18139 5176 18156 5178
rect 18076 5055 18088 5176
rect 18144 5055 18156 5176
rect 18076 5053 18093 5055
rect 18001 4876 18018 4878
rect 17938 4756 17950 4876
rect 18006 4756 18018 4876
rect 17938 4754 17955 4756
rect 17771 4718 17817 4729
rect 18001 4754 18018 4756
rect 17955 4718 18001 4729
rect 17480 4680 17491 4683
rect 17545 4680 17556 4683
rect 17664 4680 17675 4683
rect 17729 4680 17740 4683
rect 17848 4680 17859 4683
rect 17913 4680 17924 4683
rect 17265 4635 17311 4646
rect 17478 4624 17490 4680
rect 17546 4624 17558 4680
rect 17478 4610 17558 4624
rect 17662 4624 17674 4680
rect 17730 4624 17742 4680
rect 17662 4610 17742 4624
rect 17846 4624 17858 4680
rect 17914 4624 17926 4680
rect 18139 5053 18156 5055
rect 18093 4635 18139 4646
rect 17846 4610 17926 4624
rect 17478 4530 17558 4532
rect 17090 4474 17490 4530
rect 17546 4474 17558 4530
rect 15992 4471 16072 4473
rect 17478 4472 17558 4474
rect 16176 4413 16256 4415
rect 15468 4357 16188 4413
rect 16244 4357 16256 4413
rect 16176 4355 16256 4357
rect 16505 4413 16585 4415
rect 16772 4414 16842 4425
rect 17662 4414 17742 4416
rect 16772 4413 17674 4414
rect 16505 4357 16517 4413
rect 16573 4357 16774 4413
rect 16830 4358 17674 4413
rect 17730 4358 17742 4414
rect 16830 4357 17090 4358
rect 16505 4355 16585 4357
rect 16772 4347 16842 4357
rect 17662 4356 17742 4358
rect 17991 4414 18071 4416
rect 18434 4414 18504 4424
rect 17991 4358 18003 4414
rect 18059 4358 18436 4414
rect 18492 4358 18504 4414
rect 17991 4356 18071 4358
rect 18434 4346 18504 4358
rect 5848 4297 5918 4309
rect 6888 4297 6968 4299
rect 8374 4298 8454 4300
rect 5848 4241 5860 4297
rect 5916 4241 6900 4297
rect 6956 4241 6968 4297
rect 5848 4229 5918 4241
rect 2200 3190 2364 3202
rect 2680 3268 2844 3280
rect 2680 3212 2692 3268
rect 2748 3212 2844 3268
rect 2680 3200 2844 3212
rect 2200 3134 2212 3190
rect 2268 3134 2364 3190
rect 2200 3122 2364 3134
rect 2268 3072 2364 3122
rect 1165 3050 1211 3061
rect 271 2750 317 2890
rect 486 2759 582 2790
rect 486 2713 497 2759
rect 571 2713 582 2759
rect 751 2750 797 2890
rect 317 2667 455 2678
rect 317 2093 409 2667
rect 613 2667 659 2678
rect 596 2383 613 2393
rect 659 2383 676 2393
rect 596 2143 608 2383
rect 664 2143 676 2383
rect 596 2133 613 2143
rect 317 2082 455 2093
rect 659 2133 676 2143
rect 613 2082 659 2093
rect 271 1999 317 2010
rect 486 2001 497 2047
rect 571 2001 582 2047
rect 486 1860 582 2001
rect 1380 3059 1680 3072
rect 1380 3013 1391 3059
rect 1465 3026 1595 3059
rect 1465 3013 1476 3026
rect 1584 3013 1595 3026
rect 1669 3013 1680 3059
rect 1849 3050 1895 3061
rect 1211 2967 1349 2978
rect 1211 2793 1303 2967
rect 1507 2967 1553 2978
rect 1490 2908 1507 2918
rect 1711 2967 1849 2978
rect 1553 2908 1570 2918
rect 1490 2852 1502 2908
rect 1558 2852 1570 2908
rect 1490 2842 1507 2852
rect 1211 2782 1349 2793
rect 1553 2842 1570 2852
rect 1507 2782 1553 2793
rect 1757 2793 1849 2967
rect 1711 2782 1849 2793
rect 1165 2570 1211 2710
rect 1380 2701 1391 2747
rect 1465 2701 1476 2747
rect 1380 2670 1476 2701
rect 1584 2701 1595 2747
rect 1669 2701 1680 2747
rect 1584 2670 1680 2701
rect 2064 3059 2364 3072
rect 2064 3013 2075 3059
rect 2149 3026 2279 3059
rect 2149 3013 2160 3026
rect 2268 3013 2279 3026
rect 2353 3013 2364 3059
rect 2533 3050 2579 3061
rect 1987 2967 2033 2978
rect 1970 2908 1987 2918
rect 2191 2967 2237 2978
rect 2033 2908 2050 2918
rect 1970 2852 1982 2908
rect 2038 2852 2050 2908
rect 1970 2842 1987 2852
rect 2033 2842 2050 2852
rect 2174 2908 2191 2918
rect 2395 2967 2441 2978
rect 2237 2908 2254 2918
rect 2174 2852 2186 2908
rect 2242 2852 2254 2908
rect 2174 2842 2191 2852
rect 1987 2782 2033 2793
rect 2237 2842 2254 2852
rect 2378 2908 2395 2918
rect 2441 2908 2458 2918
rect 2378 2852 2390 2908
rect 2446 2852 2458 2908
rect 2378 2842 2395 2852
rect 2191 2782 2237 2793
rect 2441 2842 2458 2852
rect 2395 2782 2441 2793
rect 1849 2570 1895 2710
rect 2064 2701 2075 2747
rect 2149 2701 2160 2747
rect 2064 2670 2160 2701
rect 2268 2701 2279 2747
rect 2353 2701 2364 2747
rect 2268 2670 2364 2701
rect 2748 3059 2844 3200
rect 3356 3314 5324 3510
rect 6132 3510 6188 4241
rect 6888 4239 6968 4241
rect 7618 4242 8386 4298
rect 8442 4242 8454 4298
rect 6520 4147 6600 4161
rect 6307 4125 6353 4136
rect 6520 4091 6532 4147
rect 6588 4091 6600 4147
rect 6704 4147 6784 4161
rect 6704 4091 6716 4147
rect 6772 4091 6784 4147
rect 6888 4147 6968 4161
rect 6888 4091 6900 4147
rect 6956 4091 6968 4147
rect 7135 4125 7181 4136
rect 6522 4088 6533 4091
rect 6587 4088 6598 4091
rect 6706 4088 6717 4091
rect 6771 4088 6782 4091
rect 6890 4088 6901 4091
rect 6955 4088 6966 4091
rect 6445 4042 6491 4053
rect 6353 3868 6445 4042
rect 6445 3857 6491 3868
rect 6629 4042 6675 4053
rect 6629 3857 6675 3868
rect 6813 4042 6859 4053
rect 6997 4042 7043 4053
rect 6980 4015 6997 4017
rect 7043 4015 7060 4017
rect 6980 3895 6992 4015
rect 7048 3895 7060 4015
rect 6980 3893 6997 3895
rect 6813 3857 6859 3868
rect 7043 3893 7060 3895
rect 6997 3857 7043 3868
rect 6307 3640 6353 3785
rect 6522 3776 6533 3822
rect 6587 3776 6598 3822
rect 6522 3743 6598 3776
rect 6706 3776 6717 3822
rect 6771 3776 6782 3822
rect 6706 3743 6782 3776
rect 6890 3776 6901 3822
rect 6955 3776 6966 3822
rect 6890 3743 6966 3776
rect 7135 3640 7181 3785
rect 6295 3628 6375 3640
rect 6295 3572 6307 3628
rect 6363 3572 6375 3628
rect 6295 3560 6375 3572
rect 7113 3628 7191 3640
rect 7113 3572 7125 3628
rect 7181 3572 7191 3628
rect 7113 3560 7191 3572
rect 7466 3510 7546 3520
rect 6132 3454 7478 3510
rect 7534 3454 7546 3510
rect 7466 3452 7546 3454
rect 7300 3401 7370 3403
rect 3356 3174 3456 3314
rect 5224 3174 5324 3314
rect 3356 3134 5324 3174
rect 6132 3400 7370 3401
rect 6132 3346 7302 3400
rect 7358 3346 7370 3400
rect 6132 3345 7370 3346
rect 2748 3013 2759 3059
rect 2833 3013 2844 3059
rect 3013 3050 3059 3061
rect 2579 2967 2717 2978
rect 2579 2793 2671 2967
rect 2875 2967 2921 2978
rect 2858 2908 2875 2918
rect 2921 2908 2938 2918
rect 2858 2852 2870 2908
rect 2926 2852 2938 2908
rect 2858 2842 2875 2852
rect 2579 2782 2717 2793
rect 2921 2842 2938 2852
rect 2875 2782 2921 2793
rect 2533 2570 2579 2710
rect 2748 2701 2759 2747
rect 2833 2701 2844 2747
rect 2748 2670 2844 2701
rect 3013 2570 3059 2710
rect 3393 2994 3439 3134
rect 1128 2540 3096 2570
rect 1128 2507 2396 2540
rect 1128 2431 1166 2507
rect 1246 2431 2396 2507
rect 1128 2400 2396 2431
rect 2996 2400 3096 2540
rect 1128 2370 3096 2400
rect 3608 3003 3704 3034
rect 3608 2957 3619 3003
rect 3693 2957 3704 3003
rect 3812 3003 3908 3034
rect 3812 2957 3823 3003
rect 3897 2957 3908 3003
rect 4077 2994 4123 3134
rect 3439 2911 3577 2922
rect 3735 2911 3781 2922
rect 3939 2911 4077 2922
rect 3439 2337 3531 2911
rect 3718 2671 3730 2911
rect 3786 2671 3798 2911
rect 3439 2326 3577 2337
rect 3735 2326 3781 2337
rect 3985 2337 4077 2911
rect 3939 2326 4077 2337
rect 3393 2243 3439 2254
rect 3608 2245 3619 2291
rect 3693 2271 3704 2291
rect 3812 2271 3823 2291
rect 3693 2245 3823 2271
rect 3897 2245 3908 2291
rect 3608 2218 3908 2245
rect 4292 3003 4388 3034
rect 4292 2957 4303 3003
rect 4377 2957 4388 3003
rect 4496 3003 4592 3034
rect 4496 2957 4507 3003
rect 4581 2957 4592 3003
rect 4761 2994 4807 3134
rect 4215 2911 4261 2922
rect 4419 2911 4465 2922
rect 4623 2911 4669 2922
rect 4402 2671 4414 2911
rect 4470 2671 4482 2911
rect 4198 2337 4210 2577
rect 4266 2337 4278 2577
rect 4606 2337 4618 2577
rect 4674 2337 4686 2577
rect 4215 2326 4261 2337
rect 4419 2326 4465 2337
rect 4623 2326 4669 2337
rect 4077 2243 4123 2254
rect 4292 2245 4303 2291
rect 4377 2271 4388 2291
rect 4496 2271 4507 2291
rect 4377 2245 4507 2271
rect 4581 2245 4592 2291
rect 4292 2218 4592 2245
rect 4976 3003 5072 3034
rect 4976 2957 4987 3003
rect 5061 2957 5072 3003
rect 5241 2994 5287 3134
rect 4807 2911 4945 2922
rect 4807 2337 4899 2911
rect 5103 2911 5149 2922
rect 5086 2627 5103 2637
rect 5149 2627 5166 2637
rect 5086 2387 5098 2627
rect 5154 2387 5166 2627
rect 5086 2377 5103 2387
rect 4807 2326 4945 2337
rect 5149 2377 5166 2387
rect 5103 2326 5149 2337
rect 4761 2243 4807 2254
rect 4976 2245 4987 2291
rect 5061 2245 5072 2291
rect 3608 2170 3704 2218
rect 751 1999 797 2010
rect 1128 2140 3096 2170
rect 1128 2000 2396 2140
rect 2996 2000 3096 2140
rect 1128 1970 3096 2000
rect 3608 2114 3628 2170
rect 3684 2114 3704 2170
rect 418 1848 582 1860
rect 418 1792 430 1848
rect 486 1792 582 1848
rect 418 1780 582 1792
rect 271 1630 317 1641
rect 486 1639 582 1780
rect 1165 1830 1211 1841
rect 486 1593 497 1639
rect 571 1593 582 1639
rect 751 1630 797 1641
rect 317 1547 455 1558
rect 317 1373 409 1547
rect 613 1547 659 1558
rect 596 1488 613 1498
rect 659 1488 676 1498
rect 596 1432 608 1488
rect 664 1432 676 1488
rect 596 1422 613 1432
rect 317 1362 455 1373
rect 659 1422 676 1432
rect 613 1362 659 1373
rect 271 1150 317 1290
rect 486 1281 497 1327
rect 571 1281 582 1327
rect 486 1250 582 1281
rect 751 1150 797 1290
rect 230 230 834 1150
rect 1380 1839 1476 1870
rect 1380 1793 1391 1839
rect 1465 1793 1476 1839
rect 1645 1830 2099 1970
rect 1303 1747 1349 1758
rect 1286 1463 1303 1473
rect 1507 1747 1645 1758
rect 1349 1463 1366 1473
rect 1286 1223 1298 1463
rect 1354 1223 1366 1463
rect 1286 1213 1303 1223
rect 1349 1213 1366 1223
rect 1303 1162 1349 1173
rect 1553 1173 1645 1747
rect 1507 1162 1645 1173
rect 1165 1079 1211 1090
rect 1380 1081 1391 1127
rect 1465 1081 1476 1127
rect 1380 1006 1476 1081
rect 1691 1162 2053 1830
rect 1645 1079 1691 1090
rect 2268 1839 2364 1870
rect 2268 1793 2279 1839
rect 2353 1793 2364 1839
rect 2533 1830 2579 1970
rect 2099 1747 2237 1758
rect 2099 1173 2191 1747
rect 2395 1747 2441 1758
rect 2378 1463 2395 1473
rect 2441 1463 2458 1473
rect 2378 1223 2390 1463
rect 2446 1223 2458 1463
rect 2378 1213 2395 1223
rect 2099 1162 2237 1173
rect 2441 1213 2458 1223
rect 2395 1162 2441 1173
rect 2053 1079 2099 1090
rect 2268 1081 2279 1127
rect 2353 1081 2364 1127
rect 1380 950 1400 1006
rect 1456 950 1476 1006
rect 1380 732 1476 950
rect 2268 862 2364 1081
rect 2748 1839 2844 1870
rect 2748 1793 2759 1839
rect 2833 1793 2844 1839
rect 3013 1830 3059 1970
rect 2579 1747 2717 1758
rect 2579 1173 2671 1747
rect 2875 1747 2921 1758
rect 2858 1463 2875 1473
rect 2921 1463 2938 1473
rect 2858 1223 2870 1463
rect 2926 1223 2938 1463
rect 2858 1213 2875 1223
rect 2579 1162 2717 1173
rect 2921 1213 2938 1223
rect 2875 1162 2921 1173
rect 2533 1079 2579 1090
rect 2748 1081 2759 1127
rect 2833 1081 2844 1127
rect 2748 940 2844 1081
rect 3393 1874 3439 1885
rect 3608 1883 3704 2114
rect 4292 2014 4388 2218
rect 4976 2104 5072 2245
rect 6132 2324 6188 3345
rect 7300 3337 7370 3345
rect 6796 3293 6882 3297
rect 6796 3237 6808 3293
rect 6864 3237 6882 3293
rect 6796 3225 6882 3237
rect 6307 3080 6353 3091
rect 6522 3089 6598 3122
rect 6522 3043 6533 3089
rect 6587 3043 6598 3089
rect 6706 3089 6782 3122
rect 6706 3043 6717 3089
rect 6771 3043 6782 3089
rect 6890 3089 6966 3122
rect 6890 3043 6901 3089
rect 6955 3043 6966 3089
rect 7135 3080 7181 3091
rect 6445 2997 6491 3008
rect 6428 2970 6445 2972
rect 6629 2997 6675 3008
rect 6491 2970 6508 2972
rect 6353 2850 6440 2970
rect 6496 2850 6508 2970
rect 6428 2848 6445 2850
rect 6353 2550 6445 2670
rect 6491 2848 6508 2850
rect 6612 2670 6629 2672
rect 6813 2997 6859 3008
rect 6796 2970 6813 2972
rect 6997 2997 7043 3008
rect 6859 2970 6876 2972
rect 6796 2850 6808 2970
rect 6864 2850 6876 2970
rect 6796 2848 6813 2850
rect 6675 2670 6692 2672
rect 6612 2550 6624 2670
rect 6680 2550 6692 2670
rect 6612 2548 6629 2550
rect 6445 2512 6491 2523
rect 6675 2548 6692 2550
rect 6629 2512 6675 2523
rect 6859 2848 6876 2850
rect 6980 2670 6997 2672
rect 7118 2970 7135 2972
rect 7181 2970 7198 2972
rect 7118 2849 7130 2970
rect 7186 2849 7198 2970
rect 7118 2847 7135 2849
rect 7043 2670 7060 2672
rect 6980 2550 6992 2670
rect 7048 2550 7060 2670
rect 6980 2548 6997 2550
rect 6813 2512 6859 2523
rect 7043 2548 7060 2550
rect 6997 2512 7043 2523
rect 6522 2474 6533 2477
rect 6587 2474 6598 2477
rect 6706 2474 6717 2477
rect 6771 2474 6782 2477
rect 6890 2474 6901 2477
rect 6955 2474 6966 2477
rect 6307 2429 6353 2440
rect 6520 2418 6532 2474
rect 6588 2418 6600 2474
rect 6520 2404 6600 2418
rect 6704 2418 6716 2474
rect 6772 2418 6784 2474
rect 6704 2404 6784 2418
rect 6888 2418 6900 2474
rect 6956 2418 6968 2474
rect 7181 2847 7198 2849
rect 7135 2429 7181 2440
rect 6888 2404 6968 2418
rect 6520 2324 6600 2326
rect 6132 2268 6532 2324
rect 6588 2268 6600 2324
rect 6520 2266 6600 2268
rect 5241 2243 5287 2254
rect 5712 2208 5782 2222
rect 6704 2208 6784 2210
rect 5712 2152 5724 2208
rect 5780 2152 6716 2208
rect 6772 2152 6784 2208
rect 5712 2140 5782 2152
rect 6704 2150 6784 2152
rect 7033 2208 7113 2210
rect 7476 2208 7536 2220
rect 7033 2152 7045 2208
rect 7101 2152 7478 2208
rect 7534 2152 7536 2208
rect 7033 2150 7113 2152
rect 7476 2140 7536 2152
rect 4908 2092 5072 2104
rect 4908 2036 4920 2092
rect 4976 2036 5072 2092
rect 4908 2024 5072 2036
rect 5478 2092 5556 2103
rect 6888 2092 6968 2094
rect 5478 2091 6900 2092
rect 5478 2037 5490 2091
rect 5544 2037 6900 2091
rect 5478 2036 6900 2037
rect 6956 2036 6968 2092
rect 5478 2025 5556 2036
rect 6888 2034 6968 2036
rect 4292 1958 4312 2014
rect 4368 1958 4388 2014
rect 3608 1837 3619 1883
rect 3693 1837 3704 1883
rect 3873 1874 4123 1885
rect 3531 1791 3577 1802
rect 3514 1732 3531 1742
rect 3735 1791 3873 1802
rect 3577 1732 3594 1742
rect 3514 1676 3526 1732
rect 3582 1676 3594 1732
rect 3514 1666 3531 1676
rect 3577 1666 3594 1676
rect 3531 1606 3577 1617
rect 3781 1617 3873 1791
rect 3735 1606 3873 1617
rect 3393 1394 3439 1534
rect 3608 1525 3619 1571
rect 3693 1525 3704 1571
rect 3608 1494 3704 1525
rect 3919 1534 4077 1874
rect 4292 1883 4388 1958
rect 4292 1837 4303 1883
rect 4377 1837 4388 1883
rect 4557 1874 4603 1885
rect 4123 1791 4261 1802
rect 4123 1617 4215 1791
rect 4419 1791 4465 1802
rect 4402 1732 4419 1742
rect 4465 1732 4482 1742
rect 4402 1676 4414 1732
rect 4470 1676 4482 1732
rect 4402 1666 4419 1676
rect 4123 1606 4261 1617
rect 4465 1666 4482 1676
rect 4419 1606 4465 1617
rect 3873 1523 4123 1534
rect 4292 1525 4303 1571
rect 4377 1525 4388 1571
rect 3919 1394 4077 1523
rect 4292 1494 4388 1525
rect 4557 1394 4603 1534
rect 4761 1874 4807 1885
rect 4976 1883 5072 2024
rect 6520 1942 6600 1956
rect 6307 1920 6353 1931
rect 4976 1837 4987 1883
rect 5061 1837 5072 1883
rect 5241 1874 5287 1885
rect 4807 1791 4945 1802
rect 4807 1617 4899 1791
rect 5103 1791 5149 1802
rect 5086 1732 5103 1742
rect 5149 1732 5166 1742
rect 5086 1676 5098 1732
rect 5154 1676 5166 1732
rect 5086 1666 5103 1676
rect 4807 1606 4945 1617
rect 5149 1666 5166 1676
rect 5103 1606 5149 1617
rect 4761 1394 4807 1534
rect 4976 1525 4987 1571
rect 5061 1525 5072 1571
rect 4976 1494 5072 1525
rect 5241 1394 5287 1534
rect 6520 1886 6532 1942
rect 6588 1886 6600 1942
rect 6704 1942 6784 1956
rect 6704 1886 6716 1942
rect 6772 1886 6784 1942
rect 6888 1942 6968 1956
rect 6888 1886 6900 1942
rect 6956 1886 6968 1942
rect 7135 1920 7181 1931
rect 6522 1883 6533 1886
rect 6587 1883 6598 1886
rect 6706 1883 6717 1886
rect 6771 1883 6782 1886
rect 6890 1883 6901 1886
rect 6955 1883 6966 1886
rect 6445 1837 6491 1848
rect 6353 1663 6445 1837
rect 6445 1652 6491 1663
rect 6629 1837 6675 1848
rect 6629 1652 6675 1663
rect 6813 1837 6859 1848
rect 6997 1837 7043 1848
rect 6980 1810 6997 1812
rect 7043 1810 7060 1812
rect 6980 1690 6992 1810
rect 7048 1690 7060 1810
rect 6980 1688 6997 1690
rect 6813 1652 6859 1663
rect 7043 1688 7060 1690
rect 6997 1652 7043 1663
rect 6307 1435 6353 1580
rect 6522 1571 6533 1617
rect 6587 1571 6598 1617
rect 6522 1538 6598 1571
rect 6706 1571 6717 1617
rect 6771 1571 6782 1617
rect 6706 1538 6782 1571
rect 6890 1571 6901 1617
rect 6955 1571 6966 1617
rect 6890 1538 6966 1571
rect 7135 1435 7181 1580
rect 6295 1423 6375 1435
rect 3013 1079 3059 1090
rect 3356 1354 5324 1394
rect 6295 1367 6307 1423
rect 6363 1367 6375 1423
rect 6295 1355 6375 1367
rect 7113 1423 7193 1435
rect 7113 1367 7125 1423
rect 7181 1367 7193 1423
rect 7113 1355 7193 1367
rect 3356 1214 3456 1354
rect 5224 1214 5324 1354
rect 5529 1305 5615 1317
rect 5722 1305 5782 1309
rect 7618 1305 7674 4242
rect 8374 4240 8454 4242
rect 8006 4148 8086 4162
rect 7793 4126 7839 4137
rect 8006 4092 8018 4148
rect 8074 4092 8086 4148
rect 8190 4148 8270 4162
rect 8190 4092 8202 4148
rect 8258 4092 8270 4148
rect 8374 4148 8454 4162
rect 8374 4092 8386 4148
rect 8442 4092 8454 4148
rect 8621 4126 8667 4137
rect 8008 4089 8019 4092
rect 8073 4089 8084 4092
rect 8192 4089 8203 4092
rect 8257 4089 8268 4092
rect 8376 4089 8387 4092
rect 8441 4089 8452 4092
rect 7931 4043 7977 4054
rect 7839 3869 7931 4043
rect 7931 3858 7977 3869
rect 8115 4043 8161 4054
rect 8115 3858 8161 3869
rect 8299 4043 8345 4054
rect 8483 4043 8529 4054
rect 8466 4016 8483 4018
rect 8529 4016 8546 4018
rect 8466 3896 8478 4016
rect 8534 3896 8546 4016
rect 8466 3894 8483 3896
rect 8299 3858 8345 3869
rect 8529 3894 8546 3896
rect 8483 3858 8529 3869
rect 7793 3641 7839 3786
rect 8008 3777 8019 3823
rect 8073 3777 8084 3823
rect 8008 3744 8084 3777
rect 8192 3777 8203 3823
rect 8257 3777 8268 3823
rect 8192 3744 8268 3777
rect 8376 3777 8387 3823
rect 8441 3777 8452 3823
rect 8376 3744 8452 3777
rect 8621 3641 8667 3786
rect 7781 3629 7861 3641
rect 7781 3573 7793 3629
rect 7849 3573 7861 3629
rect 7781 3561 7861 3573
rect 8599 3629 8677 3641
rect 8599 3573 8611 3629
rect 8667 3573 8677 3629
rect 8599 3561 8677 3573
rect 9706 3510 9906 4310
rect 10106 3510 10306 4310
rect 9706 2890 10306 3510
rect 10637 4170 10683 4181
rect 10852 4179 10948 4210
rect 10852 4133 10863 4179
rect 10937 4133 10948 4179
rect 11117 4170 11571 4310
rect 10775 4087 10821 4098
rect 10758 3803 10775 3813
rect 10979 4087 11117 4098
rect 10821 3803 10838 3813
rect 10758 3563 10770 3803
rect 10826 3563 10838 3803
rect 10758 3553 10775 3563
rect 10821 3553 10838 3563
rect 10775 3502 10821 3513
rect 11025 3513 11117 4087
rect 10979 3502 11117 3513
rect 10637 3419 10683 3430
rect 10852 3421 10863 3467
rect 10937 3421 10948 3467
rect 10852 3346 10948 3421
rect 11163 3502 11525 4170
rect 11117 3419 11163 3430
rect 11740 4179 11836 4210
rect 11740 4133 11751 4179
rect 11825 4133 11836 4179
rect 12005 4170 12051 4310
rect 11571 4087 11709 4098
rect 11571 3513 11663 4087
rect 11867 4087 11913 4098
rect 11850 3803 11867 3813
rect 11913 3803 11930 3813
rect 11850 3563 11862 3803
rect 11918 3563 11930 3803
rect 11850 3553 11867 3563
rect 11571 3502 11709 3513
rect 11913 3553 11930 3563
rect 11867 3502 11913 3513
rect 11525 3419 11571 3430
rect 11740 3421 11751 3467
rect 11825 3421 11836 3467
rect 10852 3290 10872 3346
rect 10928 3290 10948 3346
rect 10852 3072 10948 3290
rect 11740 3202 11836 3421
rect 12220 4179 12316 4210
rect 12220 4133 12231 4179
rect 12305 4133 12316 4179
rect 12485 4170 12531 4310
rect 12051 4087 12189 4098
rect 12051 3513 12143 4087
rect 12347 4087 12393 4098
rect 12330 3803 12347 3813
rect 12393 3803 12410 3813
rect 12330 3563 12342 3803
rect 12398 3563 12410 3803
rect 12330 3553 12347 3563
rect 12051 3502 12189 3513
rect 12393 3553 12410 3563
rect 12347 3502 12393 3513
rect 12005 3419 12051 3430
rect 12220 3421 12231 3467
rect 12305 3421 12316 3467
rect 12220 3280 12316 3421
rect 12485 3419 12531 3430
rect 12828 3510 14296 4310
rect 14596 3510 14796 4310
rect 19178 4311 24268 4511
rect 24940 4414 24996 5661
rect 27896 5659 27976 5661
rect 33846 5717 33928 5729
rect 34412 5717 34468 6447
rect 35304 6445 35384 6447
rect 36034 6447 36802 6503
rect 36858 6447 36870 6503
rect 34936 6353 35016 6367
rect 34723 6331 34769 6342
rect 34936 6297 34948 6353
rect 35004 6297 35016 6353
rect 35120 6353 35200 6367
rect 35120 6297 35132 6353
rect 35188 6297 35200 6353
rect 35304 6353 35384 6367
rect 35304 6297 35316 6353
rect 35372 6297 35384 6353
rect 35551 6331 35597 6342
rect 34938 6294 34949 6297
rect 35003 6294 35014 6297
rect 35122 6294 35133 6297
rect 35187 6294 35198 6297
rect 35306 6294 35317 6297
rect 35371 6294 35382 6297
rect 34861 6248 34907 6259
rect 34769 6074 34861 6248
rect 34861 6063 34907 6074
rect 35045 6248 35091 6259
rect 35045 6063 35091 6074
rect 35229 6248 35275 6259
rect 35413 6248 35459 6259
rect 35396 6221 35413 6223
rect 35459 6221 35476 6223
rect 35396 6101 35408 6221
rect 35464 6101 35476 6221
rect 35396 6099 35413 6101
rect 35229 6063 35275 6074
rect 35459 6099 35476 6101
rect 35413 6063 35459 6074
rect 34723 5846 34769 5991
rect 34938 5982 34949 6028
rect 35003 5982 35014 6028
rect 34938 5949 35014 5982
rect 35122 5982 35133 6028
rect 35187 5982 35198 6028
rect 35122 5949 35198 5982
rect 35306 5982 35317 6028
rect 35371 5982 35382 6028
rect 35306 5949 35382 5982
rect 35551 5846 35597 5991
rect 34711 5834 34791 5846
rect 34711 5778 34723 5834
rect 34779 5778 34791 5834
rect 34711 5766 34791 5778
rect 35529 5834 35607 5846
rect 35529 5778 35541 5834
rect 35597 5778 35607 5834
rect 35529 5766 35607 5778
rect 33846 5661 33860 5717
rect 33916 5661 34468 5717
rect 36034 5717 36090 6447
rect 36790 6445 36870 6447
rect 43884 6447 44788 6503
rect 44844 6447 44856 6503
rect 36422 6353 36502 6367
rect 36209 6331 36255 6342
rect 36422 6297 36434 6353
rect 36490 6297 36502 6353
rect 36606 6353 36686 6367
rect 36606 6297 36618 6353
rect 36674 6297 36686 6353
rect 36790 6353 36870 6367
rect 36790 6297 36802 6353
rect 36858 6297 36870 6353
rect 37037 6331 37083 6342
rect 36424 6294 36435 6297
rect 36489 6294 36500 6297
rect 36608 6294 36619 6297
rect 36673 6294 36684 6297
rect 36792 6294 36803 6297
rect 36857 6294 36868 6297
rect 36347 6248 36393 6259
rect 36255 6074 36347 6248
rect 36347 6063 36393 6074
rect 36531 6248 36577 6259
rect 36531 6063 36577 6074
rect 36715 6248 36761 6259
rect 36899 6248 36945 6259
rect 36882 6221 36899 6223
rect 36945 6221 36962 6223
rect 36882 6101 36894 6221
rect 36950 6101 36962 6221
rect 36882 6099 36899 6101
rect 36715 6063 36761 6074
rect 36945 6099 36962 6101
rect 36899 6063 36945 6074
rect 36209 5846 36255 5991
rect 36424 5982 36435 6028
rect 36489 5982 36500 6028
rect 36424 5949 36500 5982
rect 36608 5982 36619 6028
rect 36673 5982 36684 6028
rect 36608 5949 36684 5982
rect 36792 5982 36803 6028
rect 36857 5982 36868 6028
rect 36792 5949 36868 5982
rect 37037 5846 37083 5991
rect 36197 5834 36277 5846
rect 36197 5778 36209 5834
rect 36265 5778 36277 5834
rect 36197 5766 36277 5778
rect 37015 5834 37093 5846
rect 37015 5778 37027 5834
rect 37083 5778 37093 5834
rect 37015 5766 37093 5778
rect 37368 5717 37448 5727
rect 36034 5661 37380 5717
rect 37436 5661 37448 5717
rect 33846 5649 33928 5661
rect 26420 5606 26490 5608
rect 27720 5607 27800 5609
rect 25076 5550 26422 5606
rect 26478 5550 26490 5606
rect 25076 4530 25132 5550
rect 26420 5538 26490 5550
rect 26562 5551 27732 5607
rect 27788 5551 27800 5607
rect 25740 5499 25826 5503
rect 25740 5443 25752 5499
rect 25808 5443 25826 5499
rect 25740 5431 25826 5443
rect 25251 5286 25297 5297
rect 25466 5295 25542 5328
rect 25466 5249 25477 5295
rect 25531 5249 25542 5295
rect 25650 5295 25726 5328
rect 25650 5249 25661 5295
rect 25715 5249 25726 5295
rect 25834 5295 25910 5328
rect 25834 5249 25845 5295
rect 25899 5249 25910 5295
rect 26079 5286 26125 5297
rect 25389 5203 25435 5214
rect 25372 5176 25389 5178
rect 25573 5203 25619 5214
rect 25435 5176 25452 5178
rect 25297 5056 25384 5176
rect 25440 5056 25452 5176
rect 25372 5054 25389 5056
rect 25297 4756 25389 4876
rect 25435 5054 25452 5056
rect 25556 4876 25573 4878
rect 25757 5203 25803 5214
rect 25740 5176 25757 5178
rect 25941 5203 25987 5214
rect 25803 5176 25820 5178
rect 25740 5056 25752 5176
rect 25808 5056 25820 5176
rect 25740 5054 25757 5056
rect 25619 4876 25636 4878
rect 25556 4756 25568 4876
rect 25624 4756 25636 4876
rect 25556 4754 25573 4756
rect 25389 4718 25435 4729
rect 25619 4754 25636 4756
rect 25573 4718 25619 4729
rect 25803 5054 25820 5056
rect 25924 4876 25941 4878
rect 26062 5176 26079 5178
rect 26125 5176 26142 5178
rect 26062 5055 26074 5176
rect 26130 5055 26142 5176
rect 26062 5053 26079 5055
rect 25987 4876 26004 4878
rect 25924 4756 25936 4876
rect 25992 4756 26004 4876
rect 25924 4754 25941 4756
rect 25757 4718 25803 4729
rect 25987 4754 26004 4756
rect 25941 4718 25987 4729
rect 25466 4680 25477 4683
rect 25531 4680 25542 4683
rect 25650 4680 25661 4683
rect 25715 4680 25726 4683
rect 25834 4680 25845 4683
rect 25899 4680 25910 4683
rect 25251 4635 25297 4646
rect 25464 4624 25476 4680
rect 25532 4624 25544 4680
rect 25464 4610 25544 4624
rect 25648 4624 25660 4680
rect 25716 4624 25728 4680
rect 25648 4610 25728 4624
rect 25832 4624 25844 4680
rect 25900 4624 25912 4680
rect 26125 5053 26142 5055
rect 26079 4635 26125 4646
rect 25832 4610 25912 4624
rect 25464 4530 25544 4532
rect 25076 4474 25476 4530
rect 25532 4474 25544 4530
rect 26562 4531 26618 5551
rect 27720 5539 27800 5551
rect 27226 5500 27312 5504
rect 27226 5444 27238 5500
rect 27294 5444 27312 5500
rect 27226 5432 27312 5444
rect 26737 5287 26783 5298
rect 26952 5296 27028 5329
rect 26952 5250 26963 5296
rect 27017 5250 27028 5296
rect 27136 5296 27212 5329
rect 27136 5250 27147 5296
rect 27201 5250 27212 5296
rect 27320 5296 27396 5329
rect 27320 5250 27331 5296
rect 27385 5250 27396 5296
rect 27565 5287 27611 5298
rect 26875 5204 26921 5215
rect 26858 5177 26875 5179
rect 27059 5204 27105 5215
rect 26921 5177 26938 5179
rect 26783 5057 26870 5177
rect 26926 5057 26938 5177
rect 26858 5055 26875 5057
rect 26783 4757 26875 4877
rect 26921 5055 26938 5057
rect 27042 4877 27059 4879
rect 27243 5204 27289 5215
rect 27226 5177 27243 5179
rect 27427 5204 27473 5215
rect 27289 5177 27306 5179
rect 27226 5057 27238 5177
rect 27294 5057 27306 5177
rect 27226 5055 27243 5057
rect 27105 4877 27122 4879
rect 27042 4757 27054 4877
rect 27110 4757 27122 4877
rect 27042 4755 27059 4757
rect 26875 4719 26921 4730
rect 27105 4755 27122 4757
rect 27059 4719 27105 4730
rect 27289 5055 27306 5057
rect 27410 4877 27427 4879
rect 27548 5177 27565 5179
rect 27611 5177 27628 5179
rect 27548 5056 27560 5177
rect 27616 5056 27628 5177
rect 27548 5054 27565 5056
rect 27473 4877 27490 4879
rect 27410 4757 27422 4877
rect 27478 4757 27490 4877
rect 27410 4755 27427 4757
rect 27243 4719 27289 4730
rect 27473 4755 27490 4757
rect 27427 4719 27473 4730
rect 26952 4681 26963 4684
rect 27017 4681 27028 4684
rect 27136 4681 27147 4684
rect 27201 4681 27212 4684
rect 27320 4681 27331 4684
rect 27385 4681 27396 4684
rect 26737 4636 26783 4647
rect 26950 4625 26962 4681
rect 27018 4625 27030 4681
rect 26950 4611 27030 4625
rect 27134 4625 27146 4681
rect 27202 4625 27214 4681
rect 27134 4611 27214 4625
rect 27318 4625 27330 4681
rect 27386 4625 27398 4681
rect 27611 5054 27628 5056
rect 27565 4636 27611 4647
rect 27318 4611 27398 4625
rect 26950 4531 27030 4533
rect 26562 4475 26962 4531
rect 27018 4475 27030 4531
rect 25464 4472 25544 4474
rect 26950 4473 27030 4475
rect 25648 4414 25728 4416
rect 24940 4358 25660 4414
rect 25716 4358 25728 4414
rect 25648 4356 25728 4358
rect 25977 4414 26057 4416
rect 26244 4415 26314 4426
rect 27134 4415 27214 4417
rect 26244 4414 27146 4415
rect 25977 4358 25989 4414
rect 26045 4358 26246 4414
rect 26302 4359 27146 4414
rect 27202 4359 27214 4415
rect 26302 4358 26562 4359
rect 25977 4356 26057 4358
rect 26244 4348 26314 4358
rect 27134 4357 27214 4359
rect 27463 4415 27543 4417
rect 27906 4415 27976 4425
rect 27463 4359 27475 4415
rect 27531 4359 27908 4415
rect 27964 4359 27976 4415
rect 27463 4357 27543 4359
rect 27906 4347 27976 4359
rect 15320 4297 15390 4309
rect 16360 4297 16440 4299
rect 17846 4298 17926 4300
rect 15320 4241 15332 4297
rect 15388 4241 16372 4297
rect 16428 4241 16440 4297
rect 15320 4229 15390 4241
rect 11672 3190 11836 3202
rect 12152 3268 12316 3280
rect 12152 3212 12164 3268
rect 12220 3212 12316 3268
rect 12152 3200 12316 3212
rect 11672 3134 11684 3190
rect 11740 3134 11836 3190
rect 11672 3122 11836 3134
rect 11740 3072 11836 3122
rect 10637 3050 10683 3061
rect 9743 2750 9789 2890
rect 9958 2759 10054 2790
rect 9958 2713 9969 2759
rect 10043 2713 10054 2759
rect 10223 2750 10269 2890
rect 9789 2667 9927 2678
rect 9789 2093 9881 2667
rect 10085 2667 10131 2678
rect 10068 2383 10085 2393
rect 10131 2383 10148 2393
rect 10068 2143 10080 2383
rect 10136 2143 10148 2383
rect 10068 2133 10085 2143
rect 9789 2082 9927 2093
rect 10131 2133 10148 2143
rect 10085 2082 10131 2093
rect 9743 1999 9789 2010
rect 9958 2001 9969 2047
rect 10043 2001 10054 2047
rect 9958 1860 10054 2001
rect 10852 3059 11152 3072
rect 10852 3013 10863 3059
rect 10937 3026 11067 3059
rect 10937 3013 10948 3026
rect 11056 3013 11067 3026
rect 11141 3013 11152 3059
rect 11321 3050 11367 3061
rect 10683 2967 10821 2978
rect 10683 2793 10775 2967
rect 10979 2967 11025 2978
rect 10962 2908 10979 2918
rect 11183 2967 11321 2978
rect 11025 2908 11042 2918
rect 10962 2852 10974 2908
rect 11030 2852 11042 2908
rect 10962 2842 10979 2852
rect 10683 2782 10821 2793
rect 11025 2842 11042 2852
rect 10979 2782 11025 2793
rect 11229 2793 11321 2967
rect 11183 2782 11321 2793
rect 10637 2570 10683 2710
rect 10852 2701 10863 2747
rect 10937 2701 10948 2747
rect 10852 2670 10948 2701
rect 11056 2701 11067 2747
rect 11141 2701 11152 2747
rect 11056 2670 11152 2701
rect 11536 3059 11836 3072
rect 11536 3013 11547 3059
rect 11621 3026 11751 3059
rect 11621 3013 11632 3026
rect 11740 3013 11751 3026
rect 11825 3013 11836 3059
rect 12005 3050 12051 3061
rect 11459 2967 11505 2978
rect 11442 2908 11459 2918
rect 11663 2967 11709 2978
rect 11505 2908 11522 2918
rect 11442 2852 11454 2908
rect 11510 2852 11522 2908
rect 11442 2842 11459 2852
rect 11505 2842 11522 2852
rect 11646 2908 11663 2918
rect 11867 2967 11913 2978
rect 11709 2908 11726 2918
rect 11646 2852 11658 2908
rect 11714 2852 11726 2908
rect 11646 2842 11663 2852
rect 11459 2782 11505 2793
rect 11709 2842 11726 2852
rect 11850 2908 11867 2918
rect 11913 2908 11930 2918
rect 11850 2852 11862 2908
rect 11918 2852 11930 2908
rect 11850 2842 11867 2852
rect 11663 2782 11709 2793
rect 11913 2842 11930 2852
rect 11867 2782 11913 2793
rect 11321 2570 11367 2710
rect 11536 2701 11547 2747
rect 11621 2701 11632 2747
rect 11536 2670 11632 2701
rect 11740 2701 11751 2747
rect 11825 2701 11836 2747
rect 11740 2670 11836 2701
rect 12220 3059 12316 3200
rect 12828 3314 14796 3510
rect 15604 3510 15660 4241
rect 16360 4239 16440 4241
rect 17090 4242 17858 4298
rect 17914 4242 17926 4298
rect 15992 4147 16072 4161
rect 15779 4125 15825 4136
rect 15992 4091 16004 4147
rect 16060 4091 16072 4147
rect 16176 4147 16256 4161
rect 16176 4091 16188 4147
rect 16244 4091 16256 4147
rect 16360 4147 16440 4161
rect 16360 4091 16372 4147
rect 16428 4091 16440 4147
rect 16607 4125 16653 4136
rect 15994 4088 16005 4091
rect 16059 4088 16070 4091
rect 16178 4088 16189 4091
rect 16243 4088 16254 4091
rect 16362 4088 16373 4091
rect 16427 4088 16438 4091
rect 15917 4042 15963 4053
rect 15825 3868 15917 4042
rect 15917 3857 15963 3868
rect 16101 4042 16147 4053
rect 16101 3857 16147 3868
rect 16285 4042 16331 4053
rect 16469 4042 16515 4053
rect 16452 4015 16469 4017
rect 16515 4015 16532 4017
rect 16452 3895 16464 4015
rect 16520 3895 16532 4015
rect 16452 3893 16469 3895
rect 16285 3857 16331 3868
rect 16515 3893 16532 3895
rect 16469 3857 16515 3868
rect 15779 3640 15825 3785
rect 15994 3776 16005 3822
rect 16059 3776 16070 3822
rect 15994 3743 16070 3776
rect 16178 3776 16189 3822
rect 16243 3776 16254 3822
rect 16178 3743 16254 3776
rect 16362 3776 16373 3822
rect 16427 3776 16438 3822
rect 16362 3743 16438 3776
rect 16607 3640 16653 3785
rect 15767 3628 15847 3640
rect 15767 3572 15779 3628
rect 15835 3572 15847 3628
rect 15767 3560 15847 3572
rect 16585 3628 16663 3640
rect 16585 3572 16597 3628
rect 16653 3572 16663 3628
rect 16585 3560 16663 3572
rect 16938 3510 17018 3520
rect 15604 3454 16950 3510
rect 17006 3454 17018 3510
rect 16938 3452 17018 3454
rect 16772 3401 16842 3403
rect 12828 3174 12928 3314
rect 14696 3174 14796 3314
rect 12828 3134 14796 3174
rect 15604 3400 16842 3401
rect 15604 3346 16774 3400
rect 16830 3346 16842 3400
rect 15604 3345 16842 3346
rect 12220 3013 12231 3059
rect 12305 3013 12316 3059
rect 12485 3050 12531 3061
rect 12051 2967 12189 2978
rect 12051 2793 12143 2967
rect 12347 2967 12393 2978
rect 12330 2908 12347 2918
rect 12393 2908 12410 2918
rect 12330 2852 12342 2908
rect 12398 2852 12410 2908
rect 12330 2842 12347 2852
rect 12051 2782 12189 2793
rect 12393 2842 12410 2852
rect 12347 2782 12393 2793
rect 12005 2570 12051 2710
rect 12220 2701 12231 2747
rect 12305 2701 12316 2747
rect 12220 2670 12316 2701
rect 12485 2570 12531 2710
rect 12865 2994 12911 3134
rect 10600 2540 12568 2570
rect 10600 2400 11868 2540
rect 12468 2400 12568 2540
rect 10600 2370 12568 2400
rect 13080 3003 13176 3034
rect 13080 2957 13091 3003
rect 13165 2957 13176 3003
rect 13284 3003 13380 3034
rect 13284 2957 13295 3003
rect 13369 2957 13380 3003
rect 13549 2994 13595 3134
rect 12911 2911 13049 2922
rect 13207 2911 13253 2922
rect 13411 2911 13549 2922
rect 12911 2337 13003 2911
rect 13190 2671 13202 2911
rect 13258 2671 13270 2911
rect 12911 2326 13049 2337
rect 13207 2326 13253 2337
rect 13457 2337 13549 2911
rect 13411 2326 13549 2337
rect 12865 2243 12911 2254
rect 13080 2245 13091 2291
rect 13165 2271 13176 2291
rect 13284 2271 13295 2291
rect 13165 2245 13295 2271
rect 13369 2245 13380 2291
rect 13080 2218 13380 2245
rect 13764 3003 13860 3034
rect 13764 2957 13775 3003
rect 13849 2957 13860 3003
rect 13968 3003 14064 3034
rect 13968 2957 13979 3003
rect 14053 2957 14064 3003
rect 14233 2994 14279 3134
rect 13687 2911 13733 2922
rect 13891 2911 13937 2922
rect 14095 2911 14141 2922
rect 13874 2671 13886 2911
rect 13942 2671 13954 2911
rect 13670 2337 13682 2577
rect 13738 2337 13750 2577
rect 14078 2337 14090 2577
rect 14146 2337 14158 2577
rect 13687 2326 13733 2337
rect 13891 2326 13937 2337
rect 14095 2326 14141 2337
rect 13549 2243 13595 2254
rect 13764 2245 13775 2291
rect 13849 2271 13860 2291
rect 13968 2271 13979 2291
rect 13849 2245 13979 2271
rect 14053 2245 14064 2291
rect 13764 2218 14064 2245
rect 14448 3003 14544 3034
rect 14448 2957 14459 3003
rect 14533 2957 14544 3003
rect 14713 2994 14759 3134
rect 14279 2911 14417 2922
rect 14279 2337 14371 2911
rect 14575 2911 14621 2922
rect 14558 2627 14575 2637
rect 14621 2627 14638 2637
rect 14558 2387 14570 2627
rect 14626 2387 14638 2627
rect 14558 2377 14575 2387
rect 14279 2326 14417 2337
rect 14621 2377 14638 2387
rect 14575 2326 14621 2337
rect 14233 2243 14279 2254
rect 14448 2245 14459 2291
rect 14533 2245 14544 2291
rect 13080 2170 13176 2218
rect 10223 1999 10269 2010
rect 10600 2140 12568 2170
rect 10600 2000 11868 2140
rect 12468 2000 12568 2140
rect 10600 1970 12568 2000
rect 13080 2114 13100 2170
rect 13156 2114 13176 2170
rect 9890 1848 10054 1860
rect 9890 1792 9902 1848
rect 9958 1792 10054 1848
rect 9890 1780 10054 1792
rect 5529 1249 5541 1305
rect 5597 1249 5724 1305
rect 5780 1249 7674 1305
rect 9743 1630 9789 1641
rect 9958 1639 10054 1780
rect 10637 1830 10683 1841
rect 9958 1593 9969 1639
rect 10043 1593 10054 1639
rect 10223 1630 10269 1641
rect 9789 1547 9927 1558
rect 9789 1373 9881 1547
rect 10085 1547 10131 1558
rect 10068 1488 10085 1498
rect 10131 1488 10148 1498
rect 10068 1432 10080 1488
rect 10136 1432 10148 1488
rect 10068 1422 10085 1432
rect 9789 1362 9927 1373
rect 10131 1422 10148 1432
rect 10085 1362 10131 1373
rect 5529 1237 5615 1249
rect 5722 1237 5782 1249
rect 2200 850 2364 862
rect 2680 928 2844 940
rect 2680 872 2692 928
rect 2748 872 2844 928
rect 2680 860 2844 872
rect 2200 794 2212 850
rect 2268 794 2364 850
rect 2200 782 2364 794
rect 2268 732 2364 782
rect 1165 710 1211 721
rect 1380 719 1680 732
rect 1380 673 1391 719
rect 1465 686 1595 719
rect 1465 673 1476 686
rect 1584 673 1595 686
rect 1669 673 1680 719
rect 1849 710 1895 721
rect 1211 627 1349 638
rect 1211 453 1303 627
rect 1507 627 1553 638
rect 1490 568 1507 578
rect 1711 627 1849 638
rect 1553 568 1570 578
rect 1490 512 1502 568
rect 1558 512 1570 568
rect 1490 502 1507 512
rect 1211 442 1349 453
rect 1553 502 1570 512
rect 1507 442 1553 453
rect 1757 453 1849 627
rect 1711 442 1849 453
rect 1165 230 1211 370
rect 1380 361 1391 407
rect 1465 361 1476 407
rect 1380 330 1476 361
rect 1584 361 1595 407
rect 1669 361 1680 407
rect 1584 330 1680 361
rect 2064 719 2364 732
rect 2064 673 2075 719
rect 2149 686 2279 719
rect 2149 673 2160 686
rect 2268 673 2279 686
rect 2353 673 2364 719
rect 2533 710 2579 721
rect 1987 627 2033 638
rect 1970 568 1987 578
rect 2191 627 2237 638
rect 2033 568 2050 578
rect 1970 512 1982 568
rect 2038 512 2050 568
rect 1970 502 1987 512
rect 2033 502 2050 512
rect 2174 568 2191 578
rect 2395 627 2441 638
rect 2237 568 2254 578
rect 2174 512 2186 568
rect 2242 512 2254 568
rect 2174 502 2191 512
rect 1987 442 2033 453
rect 2237 502 2254 512
rect 2378 568 2395 578
rect 2441 568 2458 578
rect 2378 512 2390 568
rect 2446 512 2458 568
rect 2378 502 2395 512
rect 2191 442 2237 453
rect 2441 502 2458 512
rect 2395 442 2441 453
rect 1849 230 1895 370
rect 2064 361 2075 407
rect 2149 361 2160 407
rect 2064 330 2160 361
rect 2268 361 2279 407
rect 2353 361 2364 407
rect 2268 330 2364 361
rect 2748 719 2844 860
rect 3356 1030 5324 1214
rect 9743 1150 9789 1290
rect 9958 1281 9969 1327
rect 10043 1281 10054 1327
rect 9958 1250 10054 1281
rect 10223 1150 10269 1290
rect 2748 673 2759 719
rect 2833 673 2844 719
rect 3013 710 3059 721
rect 2579 627 2717 638
rect 2579 453 2671 627
rect 2875 627 2921 638
rect 2858 568 2875 578
rect 2921 568 2938 578
rect 2858 512 2870 568
rect 2926 512 2938 568
rect 2858 502 2875 512
rect 2579 442 2717 453
rect 2921 502 2938 512
rect 2875 442 2921 453
rect 2533 230 2579 370
rect 2748 361 2759 407
rect 2833 361 2844 407
rect 2748 330 2844 361
rect 3013 230 3059 370
rect 3356 230 4824 1030
rect 5124 430 5324 1030
rect 9706 430 10306 1150
rect 10852 1839 10948 1870
rect 10852 1793 10863 1839
rect 10937 1793 10948 1839
rect 11117 1830 11571 1970
rect 10775 1747 10821 1758
rect 10758 1463 10775 1473
rect 10979 1747 11117 1758
rect 10821 1463 10838 1473
rect 10758 1223 10770 1463
rect 10826 1223 10838 1463
rect 10758 1213 10775 1223
rect 10821 1213 10838 1223
rect 10775 1162 10821 1173
rect 11025 1173 11117 1747
rect 10979 1162 11117 1173
rect 10637 1079 10683 1090
rect 10852 1081 10863 1127
rect 10937 1081 10948 1127
rect 10852 1006 10948 1081
rect 11163 1162 11525 1830
rect 11117 1079 11163 1090
rect 11740 1839 11836 1870
rect 11740 1793 11751 1839
rect 11825 1793 11836 1839
rect 12005 1830 12051 1970
rect 11571 1747 11709 1758
rect 11571 1173 11663 1747
rect 11867 1747 11913 1758
rect 11850 1463 11867 1473
rect 11913 1463 11930 1473
rect 11850 1223 11862 1463
rect 11918 1223 11930 1463
rect 11850 1213 11867 1223
rect 11571 1162 11709 1173
rect 11913 1213 11930 1223
rect 11867 1162 11913 1173
rect 11525 1079 11571 1090
rect 11740 1081 11751 1127
rect 11825 1081 11836 1127
rect 10852 950 10872 1006
rect 10928 950 10948 1006
rect 10852 732 10948 950
rect 11740 862 11836 1081
rect 12220 1839 12316 1870
rect 12220 1793 12231 1839
rect 12305 1793 12316 1839
rect 12485 1830 12531 1970
rect 12051 1747 12189 1758
rect 12051 1173 12143 1747
rect 12347 1747 12393 1758
rect 12330 1463 12347 1473
rect 12393 1463 12410 1473
rect 12330 1223 12342 1463
rect 12398 1223 12410 1463
rect 12330 1213 12347 1223
rect 12051 1162 12189 1173
rect 12393 1213 12410 1223
rect 12347 1162 12393 1173
rect 12005 1079 12051 1090
rect 12220 1081 12231 1127
rect 12305 1081 12316 1127
rect 12220 940 12316 1081
rect 12865 1874 12911 1885
rect 13080 1883 13176 2114
rect 13764 2014 13860 2218
rect 14448 2104 14544 2245
rect 15604 2324 15660 3345
rect 16772 3337 16842 3345
rect 16268 3293 16354 3297
rect 16268 3237 16280 3293
rect 16336 3237 16354 3293
rect 16268 3225 16354 3237
rect 15779 3080 15825 3091
rect 15994 3089 16070 3122
rect 15994 3043 16005 3089
rect 16059 3043 16070 3089
rect 16178 3089 16254 3122
rect 16178 3043 16189 3089
rect 16243 3043 16254 3089
rect 16362 3089 16438 3122
rect 16362 3043 16373 3089
rect 16427 3043 16438 3089
rect 16607 3080 16653 3091
rect 15917 2997 15963 3008
rect 15900 2970 15917 2972
rect 16101 2997 16147 3008
rect 15963 2970 15980 2972
rect 15825 2850 15912 2970
rect 15968 2850 15980 2970
rect 15900 2848 15917 2850
rect 15825 2550 15917 2670
rect 15963 2848 15980 2850
rect 16084 2670 16101 2672
rect 16285 2997 16331 3008
rect 16268 2970 16285 2972
rect 16469 2997 16515 3008
rect 16331 2970 16348 2972
rect 16268 2850 16280 2970
rect 16336 2850 16348 2970
rect 16268 2848 16285 2850
rect 16147 2670 16164 2672
rect 16084 2550 16096 2670
rect 16152 2550 16164 2670
rect 16084 2548 16101 2550
rect 15917 2512 15963 2523
rect 16147 2548 16164 2550
rect 16101 2512 16147 2523
rect 16331 2848 16348 2850
rect 16452 2670 16469 2672
rect 16590 2970 16607 2972
rect 16653 2970 16670 2972
rect 16590 2849 16602 2970
rect 16658 2849 16670 2970
rect 16590 2847 16607 2849
rect 16515 2670 16532 2672
rect 16452 2550 16464 2670
rect 16520 2550 16532 2670
rect 16452 2548 16469 2550
rect 16285 2512 16331 2523
rect 16515 2548 16532 2550
rect 16469 2512 16515 2523
rect 15994 2474 16005 2477
rect 16059 2474 16070 2477
rect 16178 2474 16189 2477
rect 16243 2474 16254 2477
rect 16362 2474 16373 2477
rect 16427 2474 16438 2477
rect 15779 2429 15825 2440
rect 15992 2418 16004 2474
rect 16060 2418 16072 2474
rect 15992 2404 16072 2418
rect 16176 2418 16188 2474
rect 16244 2418 16256 2474
rect 16176 2404 16256 2418
rect 16360 2418 16372 2474
rect 16428 2418 16440 2474
rect 16653 2847 16670 2849
rect 16607 2429 16653 2440
rect 16360 2404 16440 2418
rect 15992 2324 16072 2326
rect 15604 2268 16004 2324
rect 16060 2268 16072 2324
rect 15992 2266 16072 2268
rect 14713 2243 14759 2254
rect 15184 2208 15254 2222
rect 16176 2208 16256 2210
rect 15184 2152 15196 2208
rect 15252 2152 16188 2208
rect 16244 2152 16256 2208
rect 15184 2140 15254 2152
rect 16176 2150 16256 2152
rect 16505 2208 16585 2210
rect 16948 2208 17008 2220
rect 16505 2152 16517 2208
rect 16573 2152 16950 2208
rect 17006 2152 17008 2208
rect 16505 2150 16585 2152
rect 16948 2140 17008 2152
rect 14380 2092 14544 2104
rect 14380 2036 14392 2092
rect 14448 2036 14544 2092
rect 14380 2024 14544 2036
rect 14950 2092 15028 2103
rect 16360 2092 16440 2094
rect 14950 2091 16372 2092
rect 14950 2037 14962 2091
rect 15016 2037 16372 2091
rect 14950 2036 16372 2037
rect 16428 2036 16440 2092
rect 14950 2025 15028 2036
rect 16360 2034 16440 2036
rect 13764 1958 13784 2014
rect 13840 1958 13860 2014
rect 13080 1837 13091 1883
rect 13165 1837 13176 1883
rect 13345 1874 13595 1885
rect 13003 1791 13049 1802
rect 12986 1732 13003 1742
rect 13207 1791 13345 1802
rect 13049 1732 13066 1742
rect 12986 1676 12998 1732
rect 13054 1676 13066 1732
rect 12986 1666 13003 1676
rect 13049 1666 13066 1676
rect 13003 1606 13049 1617
rect 13253 1617 13345 1791
rect 13207 1606 13345 1617
rect 12865 1394 12911 1534
rect 13080 1525 13091 1571
rect 13165 1525 13176 1571
rect 13080 1494 13176 1525
rect 13391 1534 13549 1874
rect 13764 1883 13860 1958
rect 13764 1837 13775 1883
rect 13849 1837 13860 1883
rect 14029 1874 14075 1885
rect 13595 1791 13733 1802
rect 13595 1617 13687 1791
rect 13891 1791 13937 1802
rect 13874 1732 13891 1742
rect 13937 1732 13954 1742
rect 13874 1676 13886 1732
rect 13942 1676 13954 1732
rect 13874 1666 13891 1676
rect 13595 1606 13733 1617
rect 13937 1666 13954 1676
rect 13891 1606 13937 1617
rect 13345 1523 13595 1534
rect 13764 1525 13775 1571
rect 13849 1525 13860 1571
rect 13391 1394 13549 1523
rect 13764 1494 13860 1525
rect 14029 1394 14075 1534
rect 14233 1874 14279 1885
rect 14448 1883 14544 2024
rect 15992 1942 16072 1956
rect 15779 1920 15825 1931
rect 14448 1837 14459 1883
rect 14533 1837 14544 1883
rect 14713 1874 14759 1885
rect 14279 1791 14417 1802
rect 14279 1617 14371 1791
rect 14575 1791 14621 1802
rect 14558 1732 14575 1742
rect 14621 1732 14638 1742
rect 14558 1676 14570 1732
rect 14626 1676 14638 1732
rect 14558 1666 14575 1676
rect 14279 1606 14417 1617
rect 14621 1666 14638 1676
rect 14575 1606 14621 1617
rect 14233 1394 14279 1534
rect 14448 1525 14459 1571
rect 14533 1525 14544 1571
rect 14448 1494 14544 1525
rect 14713 1394 14759 1534
rect 15992 1886 16004 1942
rect 16060 1886 16072 1942
rect 16176 1942 16256 1956
rect 16176 1886 16188 1942
rect 16244 1886 16256 1942
rect 16360 1942 16440 1956
rect 16360 1886 16372 1942
rect 16428 1886 16440 1942
rect 16607 1920 16653 1931
rect 15994 1883 16005 1886
rect 16059 1883 16070 1886
rect 16178 1883 16189 1886
rect 16243 1883 16254 1886
rect 16362 1883 16373 1886
rect 16427 1883 16438 1886
rect 15917 1837 15963 1848
rect 15825 1663 15917 1837
rect 15917 1652 15963 1663
rect 16101 1837 16147 1848
rect 16101 1652 16147 1663
rect 16285 1837 16331 1848
rect 16469 1837 16515 1848
rect 16452 1810 16469 1812
rect 16515 1810 16532 1812
rect 16452 1690 16464 1810
rect 16520 1690 16532 1810
rect 16452 1688 16469 1690
rect 16285 1652 16331 1663
rect 16515 1688 16532 1690
rect 16469 1652 16515 1663
rect 15779 1435 15825 1580
rect 15994 1571 16005 1617
rect 16059 1571 16070 1617
rect 15994 1538 16070 1571
rect 16178 1571 16189 1617
rect 16243 1571 16254 1617
rect 16178 1538 16254 1571
rect 16362 1571 16373 1617
rect 16427 1571 16438 1617
rect 16362 1538 16438 1571
rect 16607 1435 16653 1580
rect 15767 1423 15847 1435
rect 12485 1079 12531 1090
rect 12828 1354 14796 1394
rect 15767 1367 15779 1423
rect 15835 1367 15847 1423
rect 15767 1355 15847 1367
rect 16585 1423 16665 1435
rect 16585 1367 16597 1423
rect 16653 1367 16665 1423
rect 16585 1355 16665 1367
rect 12828 1214 12928 1354
rect 14696 1214 14796 1354
rect 15001 1305 15087 1317
rect 15194 1305 15254 1309
rect 17090 1305 17146 4242
rect 17846 4240 17926 4242
rect 17478 4148 17558 4162
rect 17265 4126 17311 4137
rect 17478 4092 17490 4148
rect 17546 4092 17558 4148
rect 17662 4148 17742 4162
rect 17662 4092 17674 4148
rect 17730 4092 17742 4148
rect 17846 4148 17926 4162
rect 17846 4092 17858 4148
rect 17914 4092 17926 4148
rect 18093 4126 18139 4137
rect 17480 4089 17491 4092
rect 17545 4089 17556 4092
rect 17664 4089 17675 4092
rect 17729 4089 17740 4092
rect 17848 4089 17859 4092
rect 17913 4089 17924 4092
rect 17403 4043 17449 4054
rect 17311 3869 17403 4043
rect 17403 3858 17449 3869
rect 17587 4043 17633 4054
rect 17587 3858 17633 3869
rect 17771 4043 17817 4054
rect 17955 4043 18001 4054
rect 17938 4016 17955 4018
rect 18001 4016 18018 4018
rect 17938 3896 17950 4016
rect 18006 3896 18018 4016
rect 17938 3894 17955 3896
rect 17771 3858 17817 3869
rect 18001 3894 18018 3896
rect 17955 3858 18001 3869
rect 17265 3641 17311 3786
rect 17480 3777 17491 3823
rect 17545 3777 17556 3823
rect 17480 3744 17556 3777
rect 17664 3777 17675 3823
rect 17729 3777 17740 3823
rect 17664 3744 17740 3777
rect 17848 3777 17859 3823
rect 17913 3777 17924 3823
rect 17848 3744 17924 3777
rect 18093 3641 18139 3786
rect 17253 3629 17333 3641
rect 17253 3573 17265 3629
rect 17321 3573 17333 3629
rect 17253 3561 17333 3573
rect 18071 3629 18149 3641
rect 18071 3573 18083 3629
rect 18139 3573 18149 3629
rect 18071 3561 18149 3573
rect 19178 3511 19378 4311
rect 19578 3511 19778 4311
rect 19178 2891 19778 3511
rect 20109 4171 20155 4182
rect 20324 4180 20420 4211
rect 20324 4134 20335 4180
rect 20409 4134 20420 4180
rect 20589 4171 21043 4311
rect 20247 4088 20293 4099
rect 20230 3804 20247 3814
rect 20451 4088 20589 4099
rect 20293 3804 20310 3814
rect 20230 3564 20242 3804
rect 20298 3564 20310 3804
rect 20230 3554 20247 3564
rect 20293 3554 20310 3564
rect 20247 3503 20293 3514
rect 20497 3514 20589 4088
rect 20451 3503 20589 3514
rect 20109 3420 20155 3431
rect 20324 3422 20335 3468
rect 20409 3422 20420 3468
rect 20324 3347 20420 3422
rect 20635 3503 20997 4171
rect 20589 3420 20635 3431
rect 21212 4180 21308 4211
rect 21212 4134 21223 4180
rect 21297 4134 21308 4180
rect 21477 4171 21523 4311
rect 21043 4088 21181 4099
rect 21043 3514 21135 4088
rect 21339 4088 21385 4099
rect 21322 3804 21339 3814
rect 21385 3804 21402 3814
rect 21322 3564 21334 3804
rect 21390 3564 21402 3804
rect 21322 3554 21339 3564
rect 21043 3503 21181 3514
rect 21385 3554 21402 3564
rect 21339 3503 21385 3514
rect 20997 3420 21043 3431
rect 21212 3422 21223 3468
rect 21297 3422 21308 3468
rect 20324 3291 20344 3347
rect 20400 3291 20420 3347
rect 20324 3073 20420 3291
rect 21212 3203 21308 3422
rect 21692 4180 21788 4211
rect 21692 4134 21703 4180
rect 21777 4134 21788 4180
rect 21957 4171 22003 4311
rect 21523 4088 21661 4099
rect 21523 3514 21615 4088
rect 21819 4088 21865 4099
rect 21802 3804 21819 3814
rect 21865 3804 21882 3814
rect 21802 3564 21814 3804
rect 21870 3564 21882 3804
rect 21802 3554 21819 3564
rect 21523 3503 21661 3514
rect 21865 3554 21882 3564
rect 21819 3503 21865 3514
rect 21477 3420 21523 3431
rect 21692 3422 21703 3468
rect 21777 3422 21788 3468
rect 21692 3281 21788 3422
rect 21957 3420 22003 3431
rect 22300 3511 23768 4311
rect 24068 3511 24268 4311
rect 28650 4311 33740 4511
rect 34412 4414 34468 5661
rect 37368 5659 37448 5661
rect 43318 5717 43400 5729
rect 43884 5717 43940 6447
rect 44776 6445 44856 6447
rect 45506 6447 46274 6503
rect 46330 6447 46342 6503
rect 44408 6353 44488 6367
rect 44195 6331 44241 6342
rect 44408 6297 44420 6353
rect 44476 6297 44488 6353
rect 44592 6353 44672 6367
rect 44592 6297 44604 6353
rect 44660 6297 44672 6353
rect 44776 6353 44856 6367
rect 44776 6297 44788 6353
rect 44844 6297 44856 6353
rect 45023 6331 45069 6342
rect 44410 6294 44421 6297
rect 44475 6294 44486 6297
rect 44594 6294 44605 6297
rect 44659 6294 44670 6297
rect 44778 6294 44789 6297
rect 44843 6294 44854 6297
rect 44333 6248 44379 6259
rect 44241 6074 44333 6248
rect 44333 6063 44379 6074
rect 44517 6248 44563 6259
rect 44517 6063 44563 6074
rect 44701 6248 44747 6259
rect 44885 6248 44931 6259
rect 44868 6221 44885 6223
rect 44931 6221 44948 6223
rect 44868 6101 44880 6221
rect 44936 6101 44948 6221
rect 44868 6099 44885 6101
rect 44701 6063 44747 6074
rect 44931 6099 44948 6101
rect 44885 6063 44931 6074
rect 44195 5846 44241 5991
rect 44410 5982 44421 6028
rect 44475 5982 44486 6028
rect 44410 5949 44486 5982
rect 44594 5982 44605 6028
rect 44659 5982 44670 6028
rect 44594 5949 44670 5982
rect 44778 5982 44789 6028
rect 44843 5982 44854 6028
rect 44778 5949 44854 5982
rect 45023 5846 45069 5991
rect 44183 5834 44263 5846
rect 44183 5778 44195 5834
rect 44251 5778 44263 5834
rect 44183 5766 44263 5778
rect 45001 5834 45079 5846
rect 45001 5778 45013 5834
rect 45069 5778 45079 5834
rect 45001 5766 45079 5778
rect 43318 5661 43332 5717
rect 43388 5661 43940 5717
rect 45506 5717 45562 6447
rect 46262 6445 46342 6447
rect 53356 6447 54260 6503
rect 54316 6447 54328 6503
rect 45894 6353 45974 6367
rect 45681 6331 45727 6342
rect 45894 6297 45906 6353
rect 45962 6297 45974 6353
rect 46078 6353 46158 6367
rect 46078 6297 46090 6353
rect 46146 6297 46158 6353
rect 46262 6353 46342 6367
rect 46262 6297 46274 6353
rect 46330 6297 46342 6353
rect 46509 6331 46555 6342
rect 45896 6294 45907 6297
rect 45961 6294 45972 6297
rect 46080 6294 46091 6297
rect 46145 6294 46156 6297
rect 46264 6294 46275 6297
rect 46329 6294 46340 6297
rect 45819 6248 45865 6259
rect 45727 6074 45819 6248
rect 45819 6063 45865 6074
rect 46003 6248 46049 6259
rect 46003 6063 46049 6074
rect 46187 6248 46233 6259
rect 46371 6248 46417 6259
rect 46354 6221 46371 6223
rect 46417 6221 46434 6223
rect 46354 6101 46366 6221
rect 46422 6101 46434 6221
rect 46354 6099 46371 6101
rect 46187 6063 46233 6074
rect 46417 6099 46434 6101
rect 46371 6063 46417 6074
rect 45681 5846 45727 5991
rect 45896 5982 45907 6028
rect 45961 5982 45972 6028
rect 45896 5949 45972 5982
rect 46080 5982 46091 6028
rect 46145 5982 46156 6028
rect 46080 5949 46156 5982
rect 46264 5982 46275 6028
rect 46329 5982 46340 6028
rect 46264 5949 46340 5982
rect 46509 5846 46555 5991
rect 45669 5834 45749 5846
rect 45669 5778 45681 5834
rect 45737 5778 45749 5834
rect 45669 5766 45749 5778
rect 46487 5834 46565 5846
rect 46487 5778 46499 5834
rect 46555 5778 46565 5834
rect 46487 5766 46565 5778
rect 46840 5717 46920 5727
rect 45506 5661 46852 5717
rect 46908 5661 46920 5717
rect 43318 5649 43400 5661
rect 35892 5606 35962 5608
rect 37192 5607 37272 5609
rect 34548 5550 35894 5606
rect 35950 5550 35962 5606
rect 34548 4530 34604 5550
rect 35892 5538 35962 5550
rect 36034 5551 37204 5607
rect 37260 5551 37272 5607
rect 35212 5499 35298 5503
rect 35212 5443 35224 5499
rect 35280 5443 35298 5499
rect 35212 5431 35298 5443
rect 34723 5286 34769 5297
rect 34938 5295 35014 5328
rect 34938 5249 34949 5295
rect 35003 5249 35014 5295
rect 35122 5295 35198 5328
rect 35122 5249 35133 5295
rect 35187 5249 35198 5295
rect 35306 5295 35382 5328
rect 35306 5249 35317 5295
rect 35371 5249 35382 5295
rect 35551 5286 35597 5297
rect 34861 5203 34907 5214
rect 34844 5176 34861 5178
rect 35045 5203 35091 5214
rect 34907 5176 34924 5178
rect 34769 5056 34856 5176
rect 34912 5056 34924 5176
rect 34844 5054 34861 5056
rect 34769 4756 34861 4876
rect 34907 5054 34924 5056
rect 35028 4876 35045 4878
rect 35229 5203 35275 5214
rect 35212 5176 35229 5178
rect 35413 5203 35459 5214
rect 35275 5176 35292 5178
rect 35212 5056 35224 5176
rect 35280 5056 35292 5176
rect 35212 5054 35229 5056
rect 35091 4876 35108 4878
rect 35028 4756 35040 4876
rect 35096 4756 35108 4876
rect 35028 4754 35045 4756
rect 34861 4718 34907 4729
rect 35091 4754 35108 4756
rect 35045 4718 35091 4729
rect 35275 5054 35292 5056
rect 35396 4876 35413 4878
rect 35534 5176 35551 5178
rect 35597 5176 35614 5178
rect 35534 5055 35546 5176
rect 35602 5055 35614 5176
rect 35534 5053 35551 5055
rect 35459 4876 35476 4878
rect 35396 4756 35408 4876
rect 35464 4756 35476 4876
rect 35396 4754 35413 4756
rect 35229 4718 35275 4729
rect 35459 4754 35476 4756
rect 35413 4718 35459 4729
rect 34938 4680 34949 4683
rect 35003 4680 35014 4683
rect 35122 4680 35133 4683
rect 35187 4680 35198 4683
rect 35306 4680 35317 4683
rect 35371 4680 35382 4683
rect 34723 4635 34769 4646
rect 34936 4624 34948 4680
rect 35004 4624 35016 4680
rect 34936 4610 35016 4624
rect 35120 4624 35132 4680
rect 35188 4624 35200 4680
rect 35120 4610 35200 4624
rect 35304 4624 35316 4680
rect 35372 4624 35384 4680
rect 35597 5053 35614 5055
rect 35551 4635 35597 4646
rect 35304 4610 35384 4624
rect 34936 4530 35016 4532
rect 34548 4474 34948 4530
rect 35004 4474 35016 4530
rect 36034 4531 36090 5551
rect 37192 5539 37272 5551
rect 36698 5500 36784 5504
rect 36698 5444 36710 5500
rect 36766 5444 36784 5500
rect 36698 5432 36784 5444
rect 36209 5287 36255 5298
rect 36424 5296 36500 5329
rect 36424 5250 36435 5296
rect 36489 5250 36500 5296
rect 36608 5296 36684 5329
rect 36608 5250 36619 5296
rect 36673 5250 36684 5296
rect 36792 5296 36868 5329
rect 36792 5250 36803 5296
rect 36857 5250 36868 5296
rect 37037 5287 37083 5298
rect 36347 5204 36393 5215
rect 36330 5177 36347 5179
rect 36531 5204 36577 5215
rect 36393 5177 36410 5179
rect 36255 5057 36342 5177
rect 36398 5057 36410 5177
rect 36330 5055 36347 5057
rect 36255 4757 36347 4877
rect 36393 5055 36410 5057
rect 36514 4877 36531 4879
rect 36715 5204 36761 5215
rect 36698 5177 36715 5179
rect 36899 5204 36945 5215
rect 36761 5177 36778 5179
rect 36698 5057 36710 5177
rect 36766 5057 36778 5177
rect 36698 5055 36715 5057
rect 36577 4877 36594 4879
rect 36514 4757 36526 4877
rect 36582 4757 36594 4877
rect 36514 4755 36531 4757
rect 36347 4719 36393 4730
rect 36577 4755 36594 4757
rect 36531 4719 36577 4730
rect 36761 5055 36778 5057
rect 36882 4877 36899 4879
rect 37020 5177 37037 5179
rect 37083 5177 37100 5179
rect 37020 5056 37032 5177
rect 37088 5056 37100 5177
rect 37020 5054 37037 5056
rect 36945 4877 36962 4879
rect 36882 4757 36894 4877
rect 36950 4757 36962 4877
rect 36882 4755 36899 4757
rect 36715 4719 36761 4730
rect 36945 4755 36962 4757
rect 36899 4719 36945 4730
rect 36424 4681 36435 4684
rect 36489 4681 36500 4684
rect 36608 4681 36619 4684
rect 36673 4681 36684 4684
rect 36792 4681 36803 4684
rect 36857 4681 36868 4684
rect 36209 4636 36255 4647
rect 36422 4625 36434 4681
rect 36490 4625 36502 4681
rect 36422 4611 36502 4625
rect 36606 4625 36618 4681
rect 36674 4625 36686 4681
rect 36606 4611 36686 4625
rect 36790 4625 36802 4681
rect 36858 4625 36870 4681
rect 37083 5054 37100 5056
rect 37037 4636 37083 4647
rect 36790 4611 36870 4625
rect 36422 4531 36502 4533
rect 36034 4475 36434 4531
rect 36490 4475 36502 4531
rect 34936 4472 35016 4474
rect 36422 4473 36502 4475
rect 35120 4414 35200 4416
rect 34412 4358 35132 4414
rect 35188 4358 35200 4414
rect 35120 4356 35200 4358
rect 35449 4414 35529 4416
rect 35716 4415 35786 4426
rect 36606 4415 36686 4417
rect 35716 4414 36618 4415
rect 35449 4358 35461 4414
rect 35517 4358 35718 4414
rect 35774 4359 36618 4414
rect 36674 4359 36686 4415
rect 35774 4358 36034 4359
rect 35449 4356 35529 4358
rect 35716 4348 35786 4358
rect 36606 4357 36686 4359
rect 36935 4415 37015 4417
rect 37378 4415 37448 4425
rect 36935 4359 36947 4415
rect 37003 4359 37380 4415
rect 37436 4359 37448 4415
rect 36935 4357 37015 4359
rect 37378 4347 37448 4359
rect 24792 4298 24862 4310
rect 25832 4298 25912 4300
rect 27318 4299 27398 4301
rect 24792 4242 24804 4298
rect 24860 4242 25844 4298
rect 25900 4242 25912 4298
rect 24792 4230 24862 4242
rect 21144 3191 21308 3203
rect 21624 3269 21788 3281
rect 21624 3213 21636 3269
rect 21692 3213 21788 3269
rect 21624 3201 21788 3213
rect 21144 3135 21156 3191
rect 21212 3135 21308 3191
rect 21144 3123 21308 3135
rect 21212 3073 21308 3123
rect 20109 3051 20155 3062
rect 19215 2751 19261 2891
rect 19430 2760 19526 2791
rect 19430 2714 19441 2760
rect 19515 2714 19526 2760
rect 19695 2751 19741 2891
rect 19261 2668 19399 2679
rect 19261 2094 19353 2668
rect 19557 2668 19603 2679
rect 19540 2384 19557 2394
rect 19603 2384 19620 2394
rect 19540 2144 19552 2384
rect 19608 2144 19620 2384
rect 19540 2134 19557 2144
rect 19261 2083 19399 2094
rect 19603 2134 19620 2144
rect 19557 2083 19603 2094
rect 19215 2000 19261 2011
rect 19430 2002 19441 2048
rect 19515 2002 19526 2048
rect 19430 1861 19526 2002
rect 20324 3060 20624 3073
rect 20324 3014 20335 3060
rect 20409 3027 20539 3060
rect 20409 3014 20420 3027
rect 20528 3014 20539 3027
rect 20613 3014 20624 3060
rect 20793 3051 20839 3062
rect 20155 2968 20293 2979
rect 20155 2794 20247 2968
rect 20451 2968 20497 2979
rect 20434 2909 20451 2919
rect 20655 2968 20793 2979
rect 20497 2909 20514 2919
rect 20434 2853 20446 2909
rect 20502 2853 20514 2909
rect 20434 2843 20451 2853
rect 20155 2783 20293 2794
rect 20497 2843 20514 2853
rect 20451 2783 20497 2794
rect 20701 2794 20793 2968
rect 20655 2783 20793 2794
rect 20109 2571 20155 2711
rect 20324 2702 20335 2748
rect 20409 2702 20420 2748
rect 20324 2671 20420 2702
rect 20528 2702 20539 2748
rect 20613 2702 20624 2748
rect 20528 2671 20624 2702
rect 21008 3060 21308 3073
rect 21008 3014 21019 3060
rect 21093 3027 21223 3060
rect 21093 3014 21104 3027
rect 21212 3014 21223 3027
rect 21297 3014 21308 3060
rect 21477 3051 21523 3062
rect 20931 2968 20977 2979
rect 20914 2909 20931 2919
rect 21135 2968 21181 2979
rect 20977 2909 20994 2919
rect 20914 2853 20926 2909
rect 20982 2853 20994 2909
rect 20914 2843 20931 2853
rect 20977 2843 20994 2853
rect 21118 2909 21135 2919
rect 21339 2968 21385 2979
rect 21181 2909 21198 2919
rect 21118 2853 21130 2909
rect 21186 2853 21198 2909
rect 21118 2843 21135 2853
rect 20931 2783 20977 2794
rect 21181 2843 21198 2853
rect 21322 2909 21339 2919
rect 21385 2909 21402 2919
rect 21322 2853 21334 2909
rect 21390 2853 21402 2909
rect 21322 2843 21339 2853
rect 21135 2783 21181 2794
rect 21385 2843 21402 2853
rect 21339 2783 21385 2794
rect 20793 2571 20839 2711
rect 21008 2702 21019 2748
rect 21093 2702 21104 2748
rect 21008 2671 21104 2702
rect 21212 2702 21223 2748
rect 21297 2702 21308 2748
rect 21212 2671 21308 2702
rect 21692 3060 21788 3201
rect 22300 3315 24268 3511
rect 25076 3511 25132 4242
rect 25832 4240 25912 4242
rect 26562 4243 27330 4299
rect 27386 4243 27398 4299
rect 25464 4148 25544 4162
rect 25251 4126 25297 4137
rect 25464 4092 25476 4148
rect 25532 4092 25544 4148
rect 25648 4148 25728 4162
rect 25648 4092 25660 4148
rect 25716 4092 25728 4148
rect 25832 4148 25912 4162
rect 25832 4092 25844 4148
rect 25900 4092 25912 4148
rect 26079 4126 26125 4137
rect 25466 4089 25477 4092
rect 25531 4089 25542 4092
rect 25650 4089 25661 4092
rect 25715 4089 25726 4092
rect 25834 4089 25845 4092
rect 25899 4089 25910 4092
rect 25389 4043 25435 4054
rect 25297 3869 25389 4043
rect 25389 3858 25435 3869
rect 25573 4043 25619 4054
rect 25573 3858 25619 3869
rect 25757 4043 25803 4054
rect 25941 4043 25987 4054
rect 25924 4016 25941 4018
rect 25987 4016 26004 4018
rect 25924 3896 25936 4016
rect 25992 3896 26004 4016
rect 25924 3894 25941 3896
rect 25757 3858 25803 3869
rect 25987 3894 26004 3896
rect 25941 3858 25987 3869
rect 25251 3641 25297 3786
rect 25466 3777 25477 3823
rect 25531 3777 25542 3823
rect 25466 3744 25542 3777
rect 25650 3777 25661 3823
rect 25715 3777 25726 3823
rect 25650 3744 25726 3777
rect 25834 3777 25845 3823
rect 25899 3777 25910 3823
rect 25834 3744 25910 3777
rect 26079 3641 26125 3786
rect 25239 3629 25319 3641
rect 25239 3573 25251 3629
rect 25307 3573 25319 3629
rect 25239 3561 25319 3573
rect 26057 3629 26135 3641
rect 26057 3573 26069 3629
rect 26125 3573 26135 3629
rect 26057 3561 26135 3573
rect 26410 3511 26490 3521
rect 25076 3455 26422 3511
rect 26478 3455 26490 3511
rect 26410 3453 26490 3455
rect 26244 3402 26314 3404
rect 22300 3175 22400 3315
rect 24168 3175 24268 3315
rect 22300 3135 24268 3175
rect 25076 3401 26314 3402
rect 25076 3347 26246 3401
rect 26302 3347 26314 3401
rect 25076 3346 26314 3347
rect 21692 3014 21703 3060
rect 21777 3014 21788 3060
rect 21957 3051 22003 3062
rect 21523 2968 21661 2979
rect 21523 2794 21615 2968
rect 21819 2968 21865 2979
rect 21802 2909 21819 2919
rect 21865 2909 21882 2919
rect 21802 2853 21814 2909
rect 21870 2853 21882 2909
rect 21802 2843 21819 2853
rect 21523 2783 21661 2794
rect 21865 2843 21882 2853
rect 21819 2783 21865 2794
rect 21477 2571 21523 2711
rect 21692 2702 21703 2748
rect 21777 2702 21788 2748
rect 21692 2671 21788 2702
rect 21957 2571 22003 2711
rect 22337 2995 22383 3135
rect 20072 2541 22040 2571
rect 20072 2401 21340 2541
rect 21940 2401 22040 2541
rect 20072 2371 22040 2401
rect 22552 3004 22648 3035
rect 22552 2958 22563 3004
rect 22637 2958 22648 3004
rect 22756 3004 22852 3035
rect 22756 2958 22767 3004
rect 22841 2958 22852 3004
rect 23021 2995 23067 3135
rect 22383 2912 22521 2923
rect 22679 2912 22725 2923
rect 22883 2912 23021 2923
rect 22383 2338 22475 2912
rect 22662 2672 22674 2912
rect 22730 2672 22742 2912
rect 22383 2327 22521 2338
rect 22679 2327 22725 2338
rect 22929 2338 23021 2912
rect 22883 2327 23021 2338
rect 22337 2244 22383 2255
rect 22552 2246 22563 2292
rect 22637 2272 22648 2292
rect 22756 2272 22767 2292
rect 22637 2246 22767 2272
rect 22841 2246 22852 2292
rect 22552 2219 22852 2246
rect 23236 3004 23332 3035
rect 23236 2958 23247 3004
rect 23321 2958 23332 3004
rect 23440 3004 23536 3035
rect 23440 2958 23451 3004
rect 23525 2958 23536 3004
rect 23705 2995 23751 3135
rect 23159 2912 23205 2923
rect 23363 2912 23409 2923
rect 23567 2912 23613 2923
rect 23346 2672 23358 2912
rect 23414 2672 23426 2912
rect 23142 2338 23154 2578
rect 23210 2338 23222 2578
rect 23550 2338 23562 2578
rect 23618 2338 23630 2578
rect 23159 2327 23205 2338
rect 23363 2327 23409 2338
rect 23567 2327 23613 2338
rect 23021 2244 23067 2255
rect 23236 2246 23247 2292
rect 23321 2272 23332 2292
rect 23440 2272 23451 2292
rect 23321 2246 23451 2272
rect 23525 2246 23536 2292
rect 23236 2219 23536 2246
rect 23920 3004 24016 3035
rect 23920 2958 23931 3004
rect 24005 2958 24016 3004
rect 24185 2995 24231 3135
rect 23751 2912 23889 2923
rect 23751 2338 23843 2912
rect 24047 2912 24093 2923
rect 24030 2628 24047 2638
rect 24093 2628 24110 2638
rect 24030 2388 24042 2628
rect 24098 2388 24110 2628
rect 24030 2378 24047 2388
rect 23751 2327 23889 2338
rect 24093 2378 24110 2388
rect 24047 2327 24093 2338
rect 23705 2244 23751 2255
rect 23920 2246 23931 2292
rect 24005 2246 24016 2292
rect 22552 2171 22648 2219
rect 19695 2000 19741 2011
rect 20072 2141 22040 2171
rect 20072 2001 21340 2141
rect 21940 2001 22040 2141
rect 20072 1971 22040 2001
rect 22552 2115 22572 2171
rect 22628 2115 22648 2171
rect 19362 1849 19526 1861
rect 19362 1793 19374 1849
rect 19430 1793 19526 1849
rect 19362 1781 19526 1793
rect 15001 1249 15013 1305
rect 15069 1249 15196 1305
rect 15252 1249 17146 1305
rect 19215 1631 19261 1642
rect 19430 1640 19526 1781
rect 20109 1831 20155 1842
rect 19430 1594 19441 1640
rect 19515 1594 19526 1640
rect 19695 1631 19741 1642
rect 19261 1548 19399 1559
rect 19261 1374 19353 1548
rect 19557 1548 19603 1559
rect 19540 1489 19557 1499
rect 19603 1489 19620 1499
rect 19540 1433 19552 1489
rect 19608 1433 19620 1489
rect 19540 1423 19557 1433
rect 19261 1363 19399 1374
rect 19603 1423 19620 1433
rect 19557 1363 19603 1374
rect 15001 1237 15087 1249
rect 15194 1237 15254 1249
rect 11672 850 11836 862
rect 12152 928 12316 940
rect 12152 872 12164 928
rect 12220 872 12316 928
rect 12152 860 12316 872
rect 11672 794 11684 850
rect 11740 794 11836 850
rect 11672 782 11836 794
rect 11740 732 11836 782
rect 5124 230 10306 430
rect 10637 710 10683 721
rect 10852 719 11152 732
rect 10852 673 10863 719
rect 10937 686 11067 719
rect 10937 673 10948 686
rect 11056 673 11067 686
rect 11141 673 11152 719
rect 11321 710 11367 721
rect 10683 627 10821 638
rect 10683 453 10775 627
rect 10979 627 11025 638
rect 10962 568 10979 578
rect 11183 627 11321 638
rect 11025 568 11042 578
rect 10962 512 10974 568
rect 11030 512 11042 568
rect 10962 502 10979 512
rect 10683 442 10821 453
rect 11025 502 11042 512
rect 10979 442 11025 453
rect 11229 453 11321 627
rect 11183 442 11321 453
rect 10637 230 10683 370
rect 10852 361 10863 407
rect 10937 361 10948 407
rect 10852 330 10948 361
rect 11056 361 11067 407
rect 11141 361 11152 407
rect 11056 330 11152 361
rect 11536 719 11836 732
rect 11536 673 11547 719
rect 11621 686 11751 719
rect 11621 673 11632 686
rect 11740 673 11751 686
rect 11825 673 11836 719
rect 12005 710 12051 721
rect 11459 627 11505 638
rect 11442 568 11459 578
rect 11663 627 11709 638
rect 11505 568 11522 578
rect 11442 512 11454 568
rect 11510 512 11522 568
rect 11442 502 11459 512
rect 11505 502 11522 512
rect 11646 568 11663 578
rect 11867 627 11913 638
rect 11709 568 11726 578
rect 11646 512 11658 568
rect 11714 512 11726 568
rect 11646 502 11663 512
rect 11459 442 11505 453
rect 11709 502 11726 512
rect 11850 568 11867 578
rect 11913 568 11930 578
rect 11850 512 11862 568
rect 11918 512 11930 568
rect 11850 502 11867 512
rect 11663 442 11709 453
rect 11913 502 11930 512
rect 11867 442 11913 453
rect 11321 230 11367 370
rect 11536 361 11547 407
rect 11621 361 11632 407
rect 11536 330 11632 361
rect 11740 361 11751 407
rect 11825 361 11836 407
rect 11740 330 11836 361
rect 12220 719 12316 860
rect 12828 1030 14796 1214
rect 19215 1151 19261 1291
rect 19430 1282 19441 1328
rect 19515 1282 19526 1328
rect 19430 1251 19526 1282
rect 19695 1151 19741 1291
rect 12220 673 12231 719
rect 12305 673 12316 719
rect 12485 710 12531 721
rect 12051 627 12189 638
rect 12051 453 12143 627
rect 12347 627 12393 638
rect 12330 568 12347 578
rect 12393 568 12410 578
rect 12330 512 12342 568
rect 12398 512 12410 568
rect 12330 502 12347 512
rect 12051 442 12189 453
rect 12393 502 12410 512
rect 12347 442 12393 453
rect 12005 230 12051 370
rect 12220 361 12231 407
rect 12305 361 12316 407
rect 12220 330 12316 361
rect 12485 230 12531 370
rect 12828 230 14296 1030
rect 14596 430 14796 1030
rect 19178 430 19778 1151
rect 20324 1840 20420 1871
rect 20324 1794 20335 1840
rect 20409 1794 20420 1840
rect 20589 1831 21043 1971
rect 20247 1748 20293 1759
rect 20230 1464 20247 1474
rect 20451 1748 20589 1759
rect 20293 1464 20310 1474
rect 20230 1224 20242 1464
rect 20298 1224 20310 1464
rect 20230 1214 20247 1224
rect 20293 1214 20310 1224
rect 20247 1163 20293 1174
rect 20497 1174 20589 1748
rect 20451 1163 20589 1174
rect 20109 1080 20155 1091
rect 20324 1082 20335 1128
rect 20409 1082 20420 1128
rect 20324 1007 20420 1082
rect 20635 1163 20997 1831
rect 20589 1080 20635 1091
rect 21212 1840 21308 1871
rect 21212 1794 21223 1840
rect 21297 1794 21308 1840
rect 21477 1831 21523 1971
rect 21043 1748 21181 1759
rect 21043 1174 21135 1748
rect 21339 1748 21385 1759
rect 21322 1464 21339 1474
rect 21385 1464 21402 1474
rect 21322 1224 21334 1464
rect 21390 1224 21402 1464
rect 21322 1214 21339 1224
rect 21043 1163 21181 1174
rect 21385 1214 21402 1224
rect 21339 1163 21385 1174
rect 20997 1080 21043 1091
rect 21212 1082 21223 1128
rect 21297 1082 21308 1128
rect 20324 951 20344 1007
rect 20400 951 20420 1007
rect 20324 733 20420 951
rect 21212 863 21308 1082
rect 21692 1840 21788 1871
rect 21692 1794 21703 1840
rect 21777 1794 21788 1840
rect 21957 1831 22003 1971
rect 21523 1748 21661 1759
rect 21523 1174 21615 1748
rect 21819 1748 21865 1759
rect 21802 1464 21819 1474
rect 21865 1464 21882 1474
rect 21802 1224 21814 1464
rect 21870 1224 21882 1464
rect 21802 1214 21819 1224
rect 21523 1163 21661 1174
rect 21865 1214 21882 1224
rect 21819 1163 21865 1174
rect 21477 1080 21523 1091
rect 21692 1082 21703 1128
rect 21777 1082 21788 1128
rect 21692 941 21788 1082
rect 22337 1875 22383 1886
rect 22552 1884 22648 2115
rect 23236 2015 23332 2219
rect 23920 2105 24016 2246
rect 25076 2325 25132 3346
rect 26244 3338 26314 3346
rect 25740 3294 25826 3298
rect 25740 3238 25752 3294
rect 25808 3238 25826 3294
rect 25740 3226 25826 3238
rect 25251 3081 25297 3092
rect 25466 3090 25542 3123
rect 25466 3044 25477 3090
rect 25531 3044 25542 3090
rect 25650 3090 25726 3123
rect 25650 3044 25661 3090
rect 25715 3044 25726 3090
rect 25834 3090 25910 3123
rect 25834 3044 25845 3090
rect 25899 3044 25910 3090
rect 26079 3081 26125 3092
rect 25389 2998 25435 3009
rect 25372 2971 25389 2973
rect 25573 2998 25619 3009
rect 25435 2971 25452 2973
rect 25297 2851 25384 2971
rect 25440 2851 25452 2971
rect 25372 2849 25389 2851
rect 25297 2551 25389 2671
rect 25435 2849 25452 2851
rect 25556 2671 25573 2673
rect 25757 2998 25803 3009
rect 25740 2971 25757 2973
rect 25941 2998 25987 3009
rect 25803 2971 25820 2973
rect 25740 2851 25752 2971
rect 25808 2851 25820 2971
rect 25740 2849 25757 2851
rect 25619 2671 25636 2673
rect 25556 2551 25568 2671
rect 25624 2551 25636 2671
rect 25556 2549 25573 2551
rect 25389 2513 25435 2524
rect 25619 2549 25636 2551
rect 25573 2513 25619 2524
rect 25803 2849 25820 2851
rect 25924 2671 25941 2673
rect 26062 2971 26079 2973
rect 26125 2971 26142 2973
rect 26062 2850 26074 2971
rect 26130 2850 26142 2971
rect 26062 2848 26079 2850
rect 25987 2671 26004 2673
rect 25924 2551 25936 2671
rect 25992 2551 26004 2671
rect 25924 2549 25941 2551
rect 25757 2513 25803 2524
rect 25987 2549 26004 2551
rect 25941 2513 25987 2524
rect 25466 2475 25477 2478
rect 25531 2475 25542 2478
rect 25650 2475 25661 2478
rect 25715 2475 25726 2478
rect 25834 2475 25845 2478
rect 25899 2475 25910 2478
rect 25251 2430 25297 2441
rect 25464 2419 25476 2475
rect 25532 2419 25544 2475
rect 25464 2405 25544 2419
rect 25648 2419 25660 2475
rect 25716 2419 25728 2475
rect 25648 2405 25728 2419
rect 25832 2419 25844 2475
rect 25900 2419 25912 2475
rect 26125 2848 26142 2850
rect 26079 2430 26125 2441
rect 25832 2405 25912 2419
rect 25464 2325 25544 2327
rect 25076 2269 25476 2325
rect 25532 2269 25544 2325
rect 25464 2267 25544 2269
rect 24185 2244 24231 2255
rect 24656 2209 24726 2223
rect 25648 2209 25728 2211
rect 24656 2153 24668 2209
rect 24724 2153 25660 2209
rect 25716 2153 25728 2209
rect 24656 2141 24726 2153
rect 25648 2151 25728 2153
rect 25977 2209 26057 2211
rect 26420 2209 26480 2221
rect 25977 2153 25989 2209
rect 26045 2153 26422 2209
rect 26478 2153 26480 2209
rect 25977 2151 26057 2153
rect 26420 2141 26480 2153
rect 23852 2093 24016 2105
rect 23852 2037 23864 2093
rect 23920 2037 24016 2093
rect 23852 2025 24016 2037
rect 24422 2093 24500 2104
rect 25832 2093 25912 2095
rect 24422 2092 25844 2093
rect 24422 2038 24434 2092
rect 24488 2038 25844 2092
rect 24422 2037 25844 2038
rect 25900 2037 25912 2093
rect 24422 2026 24500 2037
rect 25832 2035 25912 2037
rect 23236 1959 23256 2015
rect 23312 1959 23332 2015
rect 22552 1838 22563 1884
rect 22637 1838 22648 1884
rect 22817 1875 23067 1886
rect 22475 1792 22521 1803
rect 22458 1733 22475 1743
rect 22679 1792 22817 1803
rect 22521 1733 22538 1743
rect 22458 1677 22470 1733
rect 22526 1677 22538 1733
rect 22458 1667 22475 1677
rect 22521 1667 22538 1677
rect 22475 1607 22521 1618
rect 22725 1618 22817 1792
rect 22679 1607 22817 1618
rect 22337 1395 22383 1535
rect 22552 1526 22563 1572
rect 22637 1526 22648 1572
rect 22552 1495 22648 1526
rect 22863 1535 23021 1875
rect 23236 1884 23332 1959
rect 23236 1838 23247 1884
rect 23321 1838 23332 1884
rect 23501 1875 23547 1886
rect 23067 1792 23205 1803
rect 23067 1618 23159 1792
rect 23363 1792 23409 1803
rect 23346 1733 23363 1743
rect 23409 1733 23426 1743
rect 23346 1677 23358 1733
rect 23414 1677 23426 1733
rect 23346 1667 23363 1677
rect 23067 1607 23205 1618
rect 23409 1667 23426 1677
rect 23363 1607 23409 1618
rect 22817 1524 23067 1535
rect 23236 1526 23247 1572
rect 23321 1526 23332 1572
rect 22863 1395 23021 1524
rect 23236 1495 23332 1526
rect 23501 1395 23547 1535
rect 23705 1875 23751 1886
rect 23920 1884 24016 2025
rect 25464 1943 25544 1957
rect 25251 1921 25297 1932
rect 23920 1838 23931 1884
rect 24005 1838 24016 1884
rect 24185 1875 24231 1886
rect 23751 1792 23889 1803
rect 23751 1618 23843 1792
rect 24047 1792 24093 1803
rect 24030 1733 24047 1743
rect 24093 1733 24110 1743
rect 24030 1677 24042 1733
rect 24098 1677 24110 1733
rect 24030 1667 24047 1677
rect 23751 1607 23889 1618
rect 24093 1667 24110 1677
rect 24047 1607 24093 1618
rect 23705 1395 23751 1535
rect 23920 1526 23931 1572
rect 24005 1526 24016 1572
rect 23920 1495 24016 1526
rect 24185 1395 24231 1535
rect 25464 1887 25476 1943
rect 25532 1887 25544 1943
rect 25648 1943 25728 1957
rect 25648 1887 25660 1943
rect 25716 1887 25728 1943
rect 25832 1943 25912 1957
rect 25832 1887 25844 1943
rect 25900 1887 25912 1943
rect 26079 1921 26125 1932
rect 25466 1884 25477 1887
rect 25531 1884 25542 1887
rect 25650 1884 25661 1887
rect 25715 1884 25726 1887
rect 25834 1884 25845 1887
rect 25899 1884 25910 1887
rect 25389 1838 25435 1849
rect 25297 1664 25389 1838
rect 25389 1653 25435 1664
rect 25573 1838 25619 1849
rect 25573 1653 25619 1664
rect 25757 1838 25803 1849
rect 25941 1838 25987 1849
rect 25924 1811 25941 1813
rect 25987 1811 26004 1813
rect 25924 1691 25936 1811
rect 25992 1691 26004 1811
rect 25924 1689 25941 1691
rect 25757 1653 25803 1664
rect 25987 1689 26004 1691
rect 25941 1653 25987 1664
rect 25251 1436 25297 1581
rect 25466 1572 25477 1618
rect 25531 1572 25542 1618
rect 25466 1539 25542 1572
rect 25650 1572 25661 1618
rect 25715 1572 25726 1618
rect 25650 1539 25726 1572
rect 25834 1572 25845 1618
rect 25899 1572 25910 1618
rect 25834 1539 25910 1572
rect 26079 1436 26125 1581
rect 25239 1424 25319 1436
rect 21957 1080 22003 1091
rect 22300 1355 24268 1395
rect 25239 1368 25251 1424
rect 25307 1368 25319 1424
rect 25239 1356 25319 1368
rect 26057 1424 26137 1436
rect 26057 1368 26069 1424
rect 26125 1368 26137 1424
rect 26057 1356 26137 1368
rect 22300 1215 22400 1355
rect 24168 1215 24268 1355
rect 24473 1306 24559 1318
rect 24666 1306 24726 1310
rect 26562 1306 26618 4243
rect 27318 4241 27398 4243
rect 26950 4149 27030 4163
rect 26737 4127 26783 4138
rect 26950 4093 26962 4149
rect 27018 4093 27030 4149
rect 27134 4149 27214 4163
rect 27134 4093 27146 4149
rect 27202 4093 27214 4149
rect 27318 4149 27398 4163
rect 27318 4093 27330 4149
rect 27386 4093 27398 4149
rect 27565 4127 27611 4138
rect 26952 4090 26963 4093
rect 27017 4090 27028 4093
rect 27136 4090 27147 4093
rect 27201 4090 27212 4093
rect 27320 4090 27331 4093
rect 27385 4090 27396 4093
rect 26875 4044 26921 4055
rect 26783 3870 26875 4044
rect 26875 3859 26921 3870
rect 27059 4044 27105 4055
rect 27059 3859 27105 3870
rect 27243 4044 27289 4055
rect 27427 4044 27473 4055
rect 27410 4017 27427 4019
rect 27473 4017 27490 4019
rect 27410 3897 27422 4017
rect 27478 3897 27490 4017
rect 27410 3895 27427 3897
rect 27243 3859 27289 3870
rect 27473 3895 27490 3897
rect 27427 3859 27473 3870
rect 26737 3642 26783 3787
rect 26952 3778 26963 3824
rect 27017 3778 27028 3824
rect 26952 3745 27028 3778
rect 27136 3778 27147 3824
rect 27201 3778 27212 3824
rect 27136 3745 27212 3778
rect 27320 3778 27331 3824
rect 27385 3778 27396 3824
rect 27320 3745 27396 3778
rect 27565 3642 27611 3787
rect 26725 3630 26805 3642
rect 26725 3574 26737 3630
rect 26793 3574 26805 3630
rect 26725 3562 26805 3574
rect 27543 3630 27621 3642
rect 27543 3574 27555 3630
rect 27611 3574 27621 3630
rect 27543 3562 27621 3574
rect 28650 3511 28850 4311
rect 29050 3511 29250 4311
rect 28650 2891 29250 3511
rect 29581 4171 29627 4182
rect 29796 4180 29892 4211
rect 29796 4134 29807 4180
rect 29881 4134 29892 4180
rect 30061 4171 30515 4311
rect 29719 4088 29765 4099
rect 29702 3804 29719 3814
rect 29923 4088 30061 4099
rect 29765 3804 29782 3814
rect 29702 3564 29714 3804
rect 29770 3564 29782 3804
rect 29702 3554 29719 3564
rect 29765 3554 29782 3564
rect 29719 3503 29765 3514
rect 29969 3514 30061 4088
rect 29923 3503 30061 3514
rect 29581 3420 29627 3431
rect 29796 3422 29807 3468
rect 29881 3422 29892 3468
rect 29796 3347 29892 3422
rect 30107 3503 30469 4171
rect 30061 3420 30107 3431
rect 30684 4180 30780 4211
rect 30684 4134 30695 4180
rect 30769 4134 30780 4180
rect 30949 4171 30995 4311
rect 30515 4088 30653 4099
rect 30515 3514 30607 4088
rect 30811 4088 30857 4099
rect 30794 3804 30811 3814
rect 30857 3804 30874 3814
rect 30794 3564 30806 3804
rect 30862 3564 30874 3804
rect 30794 3554 30811 3564
rect 30515 3503 30653 3514
rect 30857 3554 30874 3564
rect 30811 3503 30857 3514
rect 30469 3420 30515 3431
rect 30684 3422 30695 3468
rect 30769 3422 30780 3468
rect 29796 3291 29816 3347
rect 29872 3291 29892 3347
rect 29796 3073 29892 3291
rect 30684 3203 30780 3422
rect 31164 4180 31260 4211
rect 31164 4134 31175 4180
rect 31249 4134 31260 4180
rect 31429 4171 31475 4311
rect 30995 4088 31133 4099
rect 30995 3514 31087 4088
rect 31291 4088 31337 4099
rect 31274 3804 31291 3814
rect 31337 3804 31354 3814
rect 31274 3564 31286 3804
rect 31342 3564 31354 3804
rect 31274 3554 31291 3564
rect 30995 3503 31133 3514
rect 31337 3554 31354 3564
rect 31291 3503 31337 3514
rect 30949 3420 30995 3431
rect 31164 3422 31175 3468
rect 31249 3422 31260 3468
rect 31164 3281 31260 3422
rect 31429 3420 31475 3431
rect 31772 3511 33240 4311
rect 33540 3511 33740 4311
rect 38122 4311 43212 4511
rect 43884 4414 43940 5661
rect 46840 5659 46920 5661
rect 52790 5717 52872 5729
rect 53356 5717 53412 6447
rect 54248 6445 54328 6447
rect 54978 6447 55746 6503
rect 55802 6447 55814 6503
rect 53880 6353 53960 6367
rect 53667 6331 53713 6342
rect 53880 6297 53892 6353
rect 53948 6297 53960 6353
rect 54064 6353 54144 6367
rect 54064 6297 54076 6353
rect 54132 6297 54144 6353
rect 54248 6353 54328 6367
rect 54248 6297 54260 6353
rect 54316 6297 54328 6353
rect 54495 6331 54541 6342
rect 53882 6294 53893 6297
rect 53947 6294 53958 6297
rect 54066 6294 54077 6297
rect 54131 6294 54142 6297
rect 54250 6294 54261 6297
rect 54315 6294 54326 6297
rect 53805 6248 53851 6259
rect 53713 6074 53805 6248
rect 53805 6063 53851 6074
rect 53989 6248 54035 6259
rect 53989 6063 54035 6074
rect 54173 6248 54219 6259
rect 54357 6248 54403 6259
rect 54340 6221 54357 6223
rect 54403 6221 54420 6223
rect 54340 6101 54352 6221
rect 54408 6101 54420 6221
rect 54340 6099 54357 6101
rect 54173 6063 54219 6074
rect 54403 6099 54420 6101
rect 54357 6063 54403 6074
rect 53667 5846 53713 5991
rect 53882 5982 53893 6028
rect 53947 5982 53958 6028
rect 53882 5949 53958 5982
rect 54066 5982 54077 6028
rect 54131 5982 54142 6028
rect 54066 5949 54142 5982
rect 54250 5982 54261 6028
rect 54315 5982 54326 6028
rect 54250 5949 54326 5982
rect 54495 5846 54541 5991
rect 53655 5834 53735 5846
rect 53655 5778 53667 5834
rect 53723 5778 53735 5834
rect 53655 5766 53735 5778
rect 54473 5834 54551 5846
rect 54473 5778 54485 5834
rect 54541 5778 54551 5834
rect 54473 5766 54551 5778
rect 52790 5661 52804 5717
rect 52860 5661 53412 5717
rect 54978 5717 55034 6447
rect 55734 6445 55814 6447
rect 55366 6353 55446 6367
rect 55153 6331 55199 6342
rect 55366 6297 55378 6353
rect 55434 6297 55446 6353
rect 55550 6353 55630 6367
rect 55550 6297 55562 6353
rect 55618 6297 55630 6353
rect 55734 6353 55814 6367
rect 55734 6297 55746 6353
rect 55802 6297 55814 6353
rect 55981 6331 56027 6342
rect 55368 6294 55379 6297
rect 55433 6294 55444 6297
rect 55552 6294 55563 6297
rect 55617 6294 55628 6297
rect 55736 6294 55747 6297
rect 55801 6294 55812 6297
rect 55291 6248 55337 6259
rect 55199 6074 55291 6248
rect 55291 6063 55337 6074
rect 55475 6248 55521 6259
rect 55475 6063 55521 6074
rect 55659 6248 55705 6259
rect 55843 6248 55889 6259
rect 55826 6221 55843 6223
rect 55889 6221 55906 6223
rect 55826 6101 55838 6221
rect 55894 6101 55906 6221
rect 55826 6099 55843 6101
rect 55659 6063 55705 6074
rect 55889 6099 55906 6101
rect 55843 6063 55889 6074
rect 55153 5846 55199 5991
rect 55368 5982 55379 6028
rect 55433 5982 55444 6028
rect 55368 5949 55444 5982
rect 55552 5982 55563 6028
rect 55617 5982 55628 6028
rect 55552 5949 55628 5982
rect 55736 5982 55747 6028
rect 55801 5982 55812 6028
rect 55736 5949 55812 5982
rect 55981 5846 56027 5991
rect 55141 5834 55221 5846
rect 55141 5778 55153 5834
rect 55209 5778 55221 5834
rect 55141 5766 55221 5778
rect 55959 5834 56037 5846
rect 55959 5778 55971 5834
rect 56027 5778 56037 5834
rect 55959 5766 56037 5778
rect 56312 5717 56392 5727
rect 54978 5661 56324 5717
rect 56380 5661 56392 5717
rect 52790 5649 52872 5661
rect 45364 5606 45434 5608
rect 46664 5607 46744 5609
rect 44020 5550 45366 5606
rect 45422 5550 45434 5606
rect 44020 4530 44076 5550
rect 45364 5538 45434 5550
rect 45506 5551 46676 5607
rect 46732 5551 46744 5607
rect 44684 5499 44770 5503
rect 44684 5443 44696 5499
rect 44752 5443 44770 5499
rect 44684 5431 44770 5443
rect 44195 5286 44241 5297
rect 44410 5295 44486 5328
rect 44410 5249 44421 5295
rect 44475 5249 44486 5295
rect 44594 5295 44670 5328
rect 44594 5249 44605 5295
rect 44659 5249 44670 5295
rect 44778 5295 44854 5328
rect 44778 5249 44789 5295
rect 44843 5249 44854 5295
rect 45023 5286 45069 5297
rect 44333 5203 44379 5214
rect 44316 5176 44333 5178
rect 44517 5203 44563 5214
rect 44379 5176 44396 5178
rect 44241 5056 44328 5176
rect 44384 5056 44396 5176
rect 44316 5054 44333 5056
rect 44241 4756 44333 4876
rect 44379 5054 44396 5056
rect 44500 4876 44517 4878
rect 44701 5203 44747 5214
rect 44684 5176 44701 5178
rect 44885 5203 44931 5214
rect 44747 5176 44764 5178
rect 44684 5056 44696 5176
rect 44752 5056 44764 5176
rect 44684 5054 44701 5056
rect 44563 4876 44580 4878
rect 44500 4756 44512 4876
rect 44568 4756 44580 4876
rect 44500 4754 44517 4756
rect 44333 4718 44379 4729
rect 44563 4754 44580 4756
rect 44517 4718 44563 4729
rect 44747 5054 44764 5056
rect 44868 4876 44885 4878
rect 45006 5176 45023 5178
rect 45069 5176 45086 5178
rect 45006 5055 45018 5176
rect 45074 5055 45086 5176
rect 45006 5053 45023 5055
rect 44931 4876 44948 4878
rect 44868 4756 44880 4876
rect 44936 4756 44948 4876
rect 44868 4754 44885 4756
rect 44701 4718 44747 4729
rect 44931 4754 44948 4756
rect 44885 4718 44931 4729
rect 44410 4680 44421 4683
rect 44475 4680 44486 4683
rect 44594 4680 44605 4683
rect 44659 4680 44670 4683
rect 44778 4680 44789 4683
rect 44843 4680 44854 4683
rect 44195 4635 44241 4646
rect 44408 4624 44420 4680
rect 44476 4624 44488 4680
rect 44408 4610 44488 4624
rect 44592 4624 44604 4680
rect 44660 4624 44672 4680
rect 44592 4610 44672 4624
rect 44776 4624 44788 4680
rect 44844 4624 44856 4680
rect 45069 5053 45086 5055
rect 45023 4635 45069 4646
rect 44776 4610 44856 4624
rect 44408 4530 44488 4532
rect 44020 4474 44420 4530
rect 44476 4474 44488 4530
rect 45506 4531 45562 5551
rect 46664 5539 46744 5551
rect 46170 5500 46256 5504
rect 46170 5444 46182 5500
rect 46238 5444 46256 5500
rect 46170 5432 46256 5444
rect 45681 5287 45727 5298
rect 45896 5296 45972 5329
rect 45896 5250 45907 5296
rect 45961 5250 45972 5296
rect 46080 5296 46156 5329
rect 46080 5250 46091 5296
rect 46145 5250 46156 5296
rect 46264 5296 46340 5329
rect 46264 5250 46275 5296
rect 46329 5250 46340 5296
rect 46509 5287 46555 5298
rect 45819 5204 45865 5215
rect 45802 5177 45819 5179
rect 46003 5204 46049 5215
rect 45865 5177 45882 5179
rect 45727 5057 45814 5177
rect 45870 5057 45882 5177
rect 45802 5055 45819 5057
rect 45727 4757 45819 4877
rect 45865 5055 45882 5057
rect 45986 4877 46003 4879
rect 46187 5204 46233 5215
rect 46170 5177 46187 5179
rect 46371 5204 46417 5215
rect 46233 5177 46250 5179
rect 46170 5057 46182 5177
rect 46238 5057 46250 5177
rect 46170 5055 46187 5057
rect 46049 4877 46066 4879
rect 45986 4757 45998 4877
rect 46054 4757 46066 4877
rect 45986 4755 46003 4757
rect 45819 4719 45865 4730
rect 46049 4755 46066 4757
rect 46003 4719 46049 4730
rect 46233 5055 46250 5057
rect 46354 4877 46371 4879
rect 46492 5177 46509 5179
rect 46555 5177 46572 5179
rect 46492 5056 46504 5177
rect 46560 5056 46572 5177
rect 46492 5054 46509 5056
rect 46417 4877 46434 4879
rect 46354 4757 46366 4877
rect 46422 4757 46434 4877
rect 46354 4755 46371 4757
rect 46187 4719 46233 4730
rect 46417 4755 46434 4757
rect 46371 4719 46417 4730
rect 45896 4681 45907 4684
rect 45961 4681 45972 4684
rect 46080 4681 46091 4684
rect 46145 4681 46156 4684
rect 46264 4681 46275 4684
rect 46329 4681 46340 4684
rect 45681 4636 45727 4647
rect 45894 4625 45906 4681
rect 45962 4625 45974 4681
rect 45894 4611 45974 4625
rect 46078 4625 46090 4681
rect 46146 4625 46158 4681
rect 46078 4611 46158 4625
rect 46262 4625 46274 4681
rect 46330 4625 46342 4681
rect 46555 5054 46572 5056
rect 46509 4636 46555 4647
rect 46262 4611 46342 4625
rect 45894 4531 45974 4533
rect 45506 4475 45906 4531
rect 45962 4475 45974 4531
rect 44408 4472 44488 4474
rect 45894 4473 45974 4475
rect 44592 4414 44672 4416
rect 43884 4358 44604 4414
rect 44660 4358 44672 4414
rect 44592 4356 44672 4358
rect 44921 4414 45001 4416
rect 45188 4415 45258 4426
rect 46078 4415 46158 4417
rect 45188 4414 46090 4415
rect 44921 4358 44933 4414
rect 44989 4358 45190 4414
rect 45246 4359 46090 4414
rect 46146 4359 46158 4415
rect 45246 4358 45506 4359
rect 44921 4356 45001 4358
rect 45188 4348 45258 4358
rect 46078 4357 46158 4359
rect 46407 4415 46487 4417
rect 46850 4415 46920 4425
rect 46407 4359 46419 4415
rect 46475 4359 46852 4415
rect 46908 4359 46920 4415
rect 46407 4357 46487 4359
rect 46850 4347 46920 4359
rect 34264 4298 34334 4310
rect 35304 4298 35384 4300
rect 36790 4299 36870 4301
rect 34264 4242 34276 4298
rect 34332 4242 35316 4298
rect 35372 4242 35384 4298
rect 34264 4230 34334 4242
rect 30616 3191 30780 3203
rect 31096 3269 31260 3281
rect 31096 3213 31108 3269
rect 31164 3213 31260 3269
rect 31096 3201 31260 3213
rect 30616 3135 30628 3191
rect 30684 3135 30780 3191
rect 30616 3123 30780 3135
rect 30684 3073 30780 3123
rect 29581 3051 29627 3062
rect 28687 2751 28733 2891
rect 28902 2760 28998 2791
rect 28902 2714 28913 2760
rect 28987 2714 28998 2760
rect 29167 2751 29213 2891
rect 28733 2668 28871 2679
rect 28733 2094 28825 2668
rect 29029 2668 29075 2679
rect 29012 2384 29029 2394
rect 29075 2384 29092 2394
rect 29012 2144 29024 2384
rect 29080 2144 29092 2384
rect 29012 2134 29029 2144
rect 28733 2083 28871 2094
rect 29075 2134 29092 2144
rect 29029 2083 29075 2094
rect 28687 2000 28733 2011
rect 28902 2002 28913 2048
rect 28987 2002 28998 2048
rect 28902 1861 28998 2002
rect 29796 3060 30096 3073
rect 29796 3014 29807 3060
rect 29881 3027 30011 3060
rect 29881 3014 29892 3027
rect 30000 3014 30011 3027
rect 30085 3014 30096 3060
rect 30265 3051 30311 3062
rect 29627 2968 29765 2979
rect 29627 2794 29719 2968
rect 29923 2968 29969 2979
rect 29906 2909 29923 2919
rect 30127 2968 30265 2979
rect 29969 2909 29986 2919
rect 29906 2853 29918 2909
rect 29974 2853 29986 2909
rect 29906 2843 29923 2853
rect 29627 2783 29765 2794
rect 29969 2843 29986 2853
rect 29923 2783 29969 2794
rect 30173 2794 30265 2968
rect 30127 2783 30265 2794
rect 29581 2571 29627 2711
rect 29796 2702 29807 2748
rect 29881 2702 29892 2748
rect 29796 2671 29892 2702
rect 30000 2702 30011 2748
rect 30085 2702 30096 2748
rect 30000 2671 30096 2702
rect 30480 3060 30780 3073
rect 30480 3014 30491 3060
rect 30565 3027 30695 3060
rect 30565 3014 30576 3027
rect 30684 3014 30695 3027
rect 30769 3014 30780 3060
rect 30949 3051 30995 3062
rect 30403 2968 30449 2979
rect 30386 2909 30403 2919
rect 30607 2968 30653 2979
rect 30449 2909 30466 2919
rect 30386 2853 30398 2909
rect 30454 2853 30466 2909
rect 30386 2843 30403 2853
rect 30449 2843 30466 2853
rect 30590 2909 30607 2919
rect 30811 2968 30857 2979
rect 30653 2909 30670 2919
rect 30590 2853 30602 2909
rect 30658 2853 30670 2909
rect 30590 2843 30607 2853
rect 30403 2783 30449 2794
rect 30653 2843 30670 2853
rect 30794 2909 30811 2919
rect 30857 2909 30874 2919
rect 30794 2853 30806 2909
rect 30862 2853 30874 2909
rect 30794 2843 30811 2853
rect 30607 2783 30653 2794
rect 30857 2843 30874 2853
rect 30811 2783 30857 2794
rect 30265 2571 30311 2711
rect 30480 2702 30491 2748
rect 30565 2702 30576 2748
rect 30480 2671 30576 2702
rect 30684 2702 30695 2748
rect 30769 2702 30780 2748
rect 30684 2671 30780 2702
rect 31164 3060 31260 3201
rect 31772 3315 33740 3511
rect 34548 3511 34604 4242
rect 35304 4240 35384 4242
rect 36034 4243 36802 4299
rect 36858 4243 36870 4299
rect 34936 4148 35016 4162
rect 34723 4126 34769 4137
rect 34936 4092 34948 4148
rect 35004 4092 35016 4148
rect 35120 4148 35200 4162
rect 35120 4092 35132 4148
rect 35188 4092 35200 4148
rect 35304 4148 35384 4162
rect 35304 4092 35316 4148
rect 35372 4092 35384 4148
rect 35551 4126 35597 4137
rect 34938 4089 34949 4092
rect 35003 4089 35014 4092
rect 35122 4089 35133 4092
rect 35187 4089 35198 4092
rect 35306 4089 35317 4092
rect 35371 4089 35382 4092
rect 34861 4043 34907 4054
rect 34769 3869 34861 4043
rect 34861 3858 34907 3869
rect 35045 4043 35091 4054
rect 35045 3858 35091 3869
rect 35229 4043 35275 4054
rect 35413 4043 35459 4054
rect 35396 4016 35413 4018
rect 35459 4016 35476 4018
rect 35396 3896 35408 4016
rect 35464 3896 35476 4016
rect 35396 3894 35413 3896
rect 35229 3858 35275 3869
rect 35459 3894 35476 3896
rect 35413 3858 35459 3869
rect 34723 3641 34769 3786
rect 34938 3777 34949 3823
rect 35003 3777 35014 3823
rect 34938 3744 35014 3777
rect 35122 3777 35133 3823
rect 35187 3777 35198 3823
rect 35122 3744 35198 3777
rect 35306 3777 35317 3823
rect 35371 3777 35382 3823
rect 35306 3744 35382 3777
rect 35551 3641 35597 3786
rect 34711 3629 34791 3641
rect 34711 3573 34723 3629
rect 34779 3573 34791 3629
rect 34711 3561 34791 3573
rect 35529 3629 35607 3641
rect 35529 3573 35541 3629
rect 35597 3573 35607 3629
rect 35529 3561 35607 3573
rect 35882 3511 35962 3521
rect 34548 3455 35894 3511
rect 35950 3455 35962 3511
rect 35882 3453 35962 3455
rect 35716 3402 35786 3404
rect 31772 3175 31872 3315
rect 33640 3175 33740 3315
rect 31772 3135 33740 3175
rect 34548 3401 35786 3402
rect 34548 3347 35718 3401
rect 35774 3347 35786 3401
rect 34548 3346 35786 3347
rect 31164 3014 31175 3060
rect 31249 3014 31260 3060
rect 31429 3051 31475 3062
rect 30995 2968 31133 2979
rect 30995 2794 31087 2968
rect 31291 2968 31337 2979
rect 31274 2909 31291 2919
rect 31337 2909 31354 2919
rect 31274 2853 31286 2909
rect 31342 2853 31354 2909
rect 31274 2843 31291 2853
rect 30995 2783 31133 2794
rect 31337 2843 31354 2853
rect 31291 2783 31337 2794
rect 30949 2571 30995 2711
rect 31164 2702 31175 2748
rect 31249 2702 31260 2748
rect 31164 2671 31260 2702
rect 31429 2571 31475 2711
rect 31809 2995 31855 3135
rect 29544 2541 31512 2571
rect 29544 2401 30812 2541
rect 31412 2401 31512 2541
rect 29544 2371 31512 2401
rect 32024 3004 32120 3035
rect 32024 2958 32035 3004
rect 32109 2958 32120 3004
rect 32228 3004 32324 3035
rect 32228 2958 32239 3004
rect 32313 2958 32324 3004
rect 32493 2995 32539 3135
rect 31855 2912 31993 2923
rect 32151 2912 32197 2923
rect 32355 2912 32493 2923
rect 31855 2338 31947 2912
rect 32134 2672 32146 2912
rect 32202 2672 32214 2912
rect 31855 2327 31993 2338
rect 32151 2327 32197 2338
rect 32401 2338 32493 2912
rect 32355 2327 32493 2338
rect 31809 2244 31855 2255
rect 32024 2246 32035 2292
rect 32109 2272 32120 2292
rect 32228 2272 32239 2292
rect 32109 2246 32239 2272
rect 32313 2246 32324 2292
rect 32024 2219 32324 2246
rect 32708 3004 32804 3035
rect 32708 2958 32719 3004
rect 32793 2958 32804 3004
rect 32912 3004 33008 3035
rect 32912 2958 32923 3004
rect 32997 2958 33008 3004
rect 33177 2995 33223 3135
rect 32631 2912 32677 2923
rect 32835 2912 32881 2923
rect 33039 2912 33085 2923
rect 32818 2672 32830 2912
rect 32886 2672 32898 2912
rect 32614 2338 32626 2578
rect 32682 2338 32694 2578
rect 33022 2338 33034 2578
rect 33090 2338 33102 2578
rect 32631 2327 32677 2338
rect 32835 2327 32881 2338
rect 33039 2327 33085 2338
rect 32493 2244 32539 2255
rect 32708 2246 32719 2292
rect 32793 2272 32804 2292
rect 32912 2272 32923 2292
rect 32793 2246 32923 2272
rect 32997 2246 33008 2292
rect 32708 2219 33008 2246
rect 33392 3004 33488 3035
rect 33392 2958 33403 3004
rect 33477 2958 33488 3004
rect 33657 2995 33703 3135
rect 33223 2912 33361 2923
rect 33223 2338 33315 2912
rect 33519 2912 33565 2923
rect 33502 2628 33519 2638
rect 33565 2628 33582 2638
rect 33502 2388 33514 2628
rect 33570 2388 33582 2628
rect 33502 2378 33519 2388
rect 33223 2327 33361 2338
rect 33565 2378 33582 2388
rect 33519 2327 33565 2338
rect 33177 2244 33223 2255
rect 33392 2246 33403 2292
rect 33477 2246 33488 2292
rect 32024 2171 32120 2219
rect 29167 2000 29213 2011
rect 29544 2141 31512 2171
rect 29544 2001 30812 2141
rect 31412 2001 31512 2141
rect 29544 1971 31512 2001
rect 32024 2115 32044 2171
rect 32100 2115 32120 2171
rect 28834 1849 28998 1861
rect 28834 1793 28846 1849
rect 28902 1793 28998 1849
rect 28834 1781 28998 1793
rect 24473 1250 24485 1306
rect 24541 1250 24668 1306
rect 24724 1250 26618 1306
rect 28687 1631 28733 1642
rect 28902 1640 28998 1781
rect 29581 1831 29627 1842
rect 28902 1594 28913 1640
rect 28987 1594 28998 1640
rect 29167 1631 29213 1642
rect 28733 1548 28871 1559
rect 28733 1374 28825 1548
rect 29029 1548 29075 1559
rect 29012 1489 29029 1499
rect 29075 1489 29092 1499
rect 29012 1433 29024 1489
rect 29080 1433 29092 1489
rect 29012 1423 29029 1433
rect 28733 1363 28871 1374
rect 29075 1423 29092 1433
rect 29029 1363 29075 1374
rect 24473 1238 24559 1250
rect 24666 1238 24726 1250
rect 21144 851 21308 863
rect 21624 929 21788 941
rect 21624 873 21636 929
rect 21692 873 21788 929
rect 21624 861 21788 873
rect 21144 795 21156 851
rect 21212 795 21308 851
rect 21144 783 21308 795
rect 21212 733 21308 783
rect 14596 231 19778 430
rect 20109 711 20155 722
rect 20324 720 20624 733
rect 20324 674 20335 720
rect 20409 687 20539 720
rect 20409 674 20420 687
rect 20528 674 20539 687
rect 20613 674 20624 720
rect 20793 711 20839 722
rect 20155 628 20293 639
rect 20155 454 20247 628
rect 20451 628 20497 639
rect 20434 569 20451 579
rect 20655 628 20793 639
rect 20497 569 20514 579
rect 20434 513 20446 569
rect 20502 513 20514 569
rect 20434 503 20451 513
rect 20155 443 20293 454
rect 20497 503 20514 513
rect 20451 443 20497 454
rect 20701 454 20793 628
rect 20655 443 20793 454
rect 20109 231 20155 371
rect 20324 362 20335 408
rect 20409 362 20420 408
rect 20324 331 20420 362
rect 20528 362 20539 408
rect 20613 362 20624 408
rect 20528 331 20624 362
rect 21008 720 21308 733
rect 21008 674 21019 720
rect 21093 687 21223 720
rect 21093 674 21104 687
rect 21212 674 21223 687
rect 21297 674 21308 720
rect 21477 711 21523 722
rect 20931 628 20977 639
rect 20914 569 20931 579
rect 21135 628 21181 639
rect 20977 569 20994 579
rect 20914 513 20926 569
rect 20982 513 20994 569
rect 20914 503 20931 513
rect 20977 503 20994 513
rect 21118 569 21135 579
rect 21339 628 21385 639
rect 21181 569 21198 579
rect 21118 513 21130 569
rect 21186 513 21198 569
rect 21118 503 21135 513
rect 20931 443 20977 454
rect 21181 503 21198 513
rect 21322 569 21339 579
rect 21385 569 21402 579
rect 21322 513 21334 569
rect 21390 513 21402 569
rect 21322 503 21339 513
rect 21135 443 21181 454
rect 21385 503 21402 513
rect 21339 443 21385 454
rect 20793 231 20839 371
rect 21008 362 21019 408
rect 21093 362 21104 408
rect 21008 331 21104 362
rect 21212 362 21223 408
rect 21297 362 21308 408
rect 21212 331 21308 362
rect 21692 720 21788 861
rect 22300 1031 24268 1215
rect 28687 1151 28733 1291
rect 28902 1282 28913 1328
rect 28987 1282 28998 1328
rect 28902 1251 28998 1282
rect 29167 1151 29213 1291
rect 21692 674 21703 720
rect 21777 674 21788 720
rect 21957 711 22003 722
rect 21523 628 21661 639
rect 21523 454 21615 628
rect 21819 628 21865 639
rect 21802 569 21819 579
rect 21865 569 21882 579
rect 21802 513 21814 569
rect 21870 513 21882 569
rect 21802 503 21819 513
rect 21523 443 21661 454
rect 21865 503 21882 513
rect 21819 443 21865 454
rect 21477 231 21523 371
rect 21692 362 21703 408
rect 21777 362 21788 408
rect 21692 331 21788 362
rect 21957 231 22003 371
rect 22300 231 23768 1031
rect 24068 431 24268 1031
rect 28650 431 29250 1151
rect 29796 1840 29892 1871
rect 29796 1794 29807 1840
rect 29881 1794 29892 1840
rect 30061 1831 30515 1971
rect 29719 1748 29765 1759
rect 29702 1464 29719 1474
rect 29923 1748 30061 1759
rect 29765 1464 29782 1474
rect 29702 1224 29714 1464
rect 29770 1224 29782 1464
rect 29702 1214 29719 1224
rect 29765 1214 29782 1224
rect 29719 1163 29765 1174
rect 29969 1174 30061 1748
rect 29923 1163 30061 1174
rect 29581 1080 29627 1091
rect 29796 1082 29807 1128
rect 29881 1082 29892 1128
rect 29796 1007 29892 1082
rect 30107 1163 30469 1831
rect 30061 1080 30107 1091
rect 30684 1840 30780 1871
rect 30684 1794 30695 1840
rect 30769 1794 30780 1840
rect 30949 1831 30995 1971
rect 30515 1748 30653 1759
rect 30515 1174 30607 1748
rect 30811 1748 30857 1759
rect 30794 1464 30811 1474
rect 30857 1464 30874 1474
rect 30794 1224 30806 1464
rect 30862 1224 30874 1464
rect 30794 1214 30811 1224
rect 30515 1163 30653 1174
rect 30857 1214 30874 1224
rect 30811 1163 30857 1174
rect 30469 1080 30515 1091
rect 30684 1082 30695 1128
rect 30769 1082 30780 1128
rect 29796 951 29816 1007
rect 29872 951 29892 1007
rect 29796 733 29892 951
rect 30684 863 30780 1082
rect 31164 1840 31260 1871
rect 31164 1794 31175 1840
rect 31249 1794 31260 1840
rect 31429 1831 31475 1971
rect 30995 1748 31133 1759
rect 30995 1174 31087 1748
rect 31291 1748 31337 1759
rect 31274 1464 31291 1474
rect 31337 1464 31354 1474
rect 31274 1224 31286 1464
rect 31342 1224 31354 1464
rect 31274 1214 31291 1224
rect 30995 1163 31133 1174
rect 31337 1214 31354 1224
rect 31291 1163 31337 1174
rect 30949 1080 30995 1091
rect 31164 1082 31175 1128
rect 31249 1082 31260 1128
rect 31164 941 31260 1082
rect 31809 1875 31855 1886
rect 32024 1884 32120 2115
rect 32708 2015 32804 2219
rect 33392 2105 33488 2246
rect 34548 2325 34604 3346
rect 35716 3338 35786 3346
rect 35212 3294 35298 3298
rect 35212 3238 35224 3294
rect 35280 3238 35298 3294
rect 35212 3226 35298 3238
rect 34723 3081 34769 3092
rect 34938 3090 35014 3123
rect 34938 3044 34949 3090
rect 35003 3044 35014 3090
rect 35122 3090 35198 3123
rect 35122 3044 35133 3090
rect 35187 3044 35198 3090
rect 35306 3090 35382 3123
rect 35306 3044 35317 3090
rect 35371 3044 35382 3090
rect 35551 3081 35597 3092
rect 34861 2998 34907 3009
rect 34844 2971 34861 2973
rect 35045 2998 35091 3009
rect 34907 2971 34924 2973
rect 34769 2851 34856 2971
rect 34912 2851 34924 2971
rect 34844 2849 34861 2851
rect 34769 2551 34861 2671
rect 34907 2849 34924 2851
rect 35028 2671 35045 2673
rect 35229 2998 35275 3009
rect 35212 2971 35229 2973
rect 35413 2998 35459 3009
rect 35275 2971 35292 2973
rect 35212 2851 35224 2971
rect 35280 2851 35292 2971
rect 35212 2849 35229 2851
rect 35091 2671 35108 2673
rect 35028 2551 35040 2671
rect 35096 2551 35108 2671
rect 35028 2549 35045 2551
rect 34861 2513 34907 2524
rect 35091 2549 35108 2551
rect 35045 2513 35091 2524
rect 35275 2849 35292 2851
rect 35396 2671 35413 2673
rect 35534 2971 35551 2973
rect 35597 2971 35614 2973
rect 35534 2850 35546 2971
rect 35602 2850 35614 2971
rect 35534 2848 35551 2850
rect 35459 2671 35476 2673
rect 35396 2551 35408 2671
rect 35464 2551 35476 2671
rect 35396 2549 35413 2551
rect 35229 2513 35275 2524
rect 35459 2549 35476 2551
rect 35413 2513 35459 2524
rect 34938 2475 34949 2478
rect 35003 2475 35014 2478
rect 35122 2475 35133 2478
rect 35187 2475 35198 2478
rect 35306 2475 35317 2478
rect 35371 2475 35382 2478
rect 34723 2430 34769 2441
rect 34936 2419 34948 2475
rect 35004 2419 35016 2475
rect 34936 2405 35016 2419
rect 35120 2419 35132 2475
rect 35188 2419 35200 2475
rect 35120 2405 35200 2419
rect 35304 2419 35316 2475
rect 35372 2419 35384 2475
rect 35597 2848 35614 2850
rect 35551 2430 35597 2441
rect 35304 2405 35384 2419
rect 34936 2325 35016 2327
rect 34548 2269 34948 2325
rect 35004 2269 35016 2325
rect 34936 2267 35016 2269
rect 33657 2244 33703 2255
rect 34128 2209 34198 2223
rect 35120 2209 35200 2211
rect 34128 2153 34140 2209
rect 34196 2153 35132 2209
rect 35188 2153 35200 2209
rect 34128 2141 34198 2153
rect 35120 2151 35200 2153
rect 35449 2209 35529 2211
rect 35892 2209 35952 2221
rect 35449 2153 35461 2209
rect 35517 2153 35894 2209
rect 35950 2153 35952 2209
rect 35449 2151 35529 2153
rect 35892 2141 35952 2153
rect 33324 2093 33488 2105
rect 33324 2037 33336 2093
rect 33392 2037 33488 2093
rect 33324 2025 33488 2037
rect 33894 2093 33972 2104
rect 35304 2093 35384 2095
rect 33894 2092 35316 2093
rect 33894 2038 33906 2092
rect 33960 2038 35316 2092
rect 33894 2037 35316 2038
rect 35372 2037 35384 2093
rect 33894 2026 33972 2037
rect 35304 2035 35384 2037
rect 32708 1959 32728 2015
rect 32784 1959 32804 2015
rect 32024 1838 32035 1884
rect 32109 1838 32120 1884
rect 32289 1875 32539 1886
rect 31947 1792 31993 1803
rect 31930 1733 31947 1743
rect 32151 1792 32289 1803
rect 31993 1733 32010 1743
rect 31930 1677 31942 1733
rect 31998 1677 32010 1733
rect 31930 1667 31947 1677
rect 31993 1667 32010 1677
rect 31947 1607 31993 1618
rect 32197 1618 32289 1792
rect 32151 1607 32289 1618
rect 31809 1395 31855 1535
rect 32024 1526 32035 1572
rect 32109 1526 32120 1572
rect 32024 1495 32120 1526
rect 32335 1535 32493 1875
rect 32708 1884 32804 1959
rect 32708 1838 32719 1884
rect 32793 1838 32804 1884
rect 32973 1875 33019 1886
rect 32539 1792 32677 1803
rect 32539 1618 32631 1792
rect 32835 1792 32881 1803
rect 32818 1733 32835 1743
rect 32881 1733 32898 1743
rect 32818 1677 32830 1733
rect 32886 1677 32898 1733
rect 32818 1667 32835 1677
rect 32539 1607 32677 1618
rect 32881 1667 32898 1677
rect 32835 1607 32881 1618
rect 32289 1524 32539 1535
rect 32708 1526 32719 1572
rect 32793 1526 32804 1572
rect 32335 1395 32493 1524
rect 32708 1495 32804 1526
rect 32973 1395 33019 1535
rect 33177 1875 33223 1886
rect 33392 1884 33488 2025
rect 34936 1943 35016 1957
rect 34723 1921 34769 1932
rect 33392 1838 33403 1884
rect 33477 1838 33488 1884
rect 33657 1875 33703 1886
rect 33223 1792 33361 1803
rect 33223 1618 33315 1792
rect 33519 1792 33565 1803
rect 33502 1733 33519 1743
rect 33565 1733 33582 1743
rect 33502 1677 33514 1733
rect 33570 1677 33582 1733
rect 33502 1667 33519 1677
rect 33223 1607 33361 1618
rect 33565 1667 33582 1677
rect 33519 1607 33565 1618
rect 33177 1395 33223 1535
rect 33392 1526 33403 1572
rect 33477 1526 33488 1572
rect 33392 1495 33488 1526
rect 33657 1395 33703 1535
rect 34936 1887 34948 1943
rect 35004 1887 35016 1943
rect 35120 1943 35200 1957
rect 35120 1887 35132 1943
rect 35188 1887 35200 1943
rect 35304 1943 35384 1957
rect 35304 1887 35316 1943
rect 35372 1887 35384 1943
rect 35551 1921 35597 1932
rect 34938 1884 34949 1887
rect 35003 1884 35014 1887
rect 35122 1884 35133 1887
rect 35187 1884 35198 1887
rect 35306 1884 35317 1887
rect 35371 1884 35382 1887
rect 34861 1838 34907 1849
rect 34769 1664 34861 1838
rect 34861 1653 34907 1664
rect 35045 1838 35091 1849
rect 35045 1653 35091 1664
rect 35229 1838 35275 1849
rect 35413 1838 35459 1849
rect 35396 1811 35413 1813
rect 35459 1811 35476 1813
rect 35396 1691 35408 1811
rect 35464 1691 35476 1811
rect 35396 1689 35413 1691
rect 35229 1653 35275 1664
rect 35459 1689 35476 1691
rect 35413 1653 35459 1664
rect 34723 1436 34769 1581
rect 34938 1572 34949 1618
rect 35003 1572 35014 1618
rect 34938 1539 35014 1572
rect 35122 1572 35133 1618
rect 35187 1572 35198 1618
rect 35122 1539 35198 1572
rect 35306 1572 35317 1618
rect 35371 1572 35382 1618
rect 35306 1539 35382 1572
rect 35551 1436 35597 1581
rect 34711 1424 34791 1436
rect 31429 1080 31475 1091
rect 31772 1355 33740 1395
rect 34711 1368 34723 1424
rect 34779 1368 34791 1424
rect 34711 1356 34791 1368
rect 35529 1424 35609 1436
rect 35529 1368 35541 1424
rect 35597 1368 35609 1424
rect 35529 1356 35609 1368
rect 31772 1215 31872 1355
rect 33640 1215 33740 1355
rect 33945 1306 34031 1318
rect 34138 1306 34198 1310
rect 36034 1306 36090 4243
rect 36790 4241 36870 4243
rect 36422 4149 36502 4163
rect 36209 4127 36255 4138
rect 36422 4093 36434 4149
rect 36490 4093 36502 4149
rect 36606 4149 36686 4163
rect 36606 4093 36618 4149
rect 36674 4093 36686 4149
rect 36790 4149 36870 4163
rect 36790 4093 36802 4149
rect 36858 4093 36870 4149
rect 37037 4127 37083 4138
rect 36424 4090 36435 4093
rect 36489 4090 36500 4093
rect 36608 4090 36619 4093
rect 36673 4090 36684 4093
rect 36792 4090 36803 4093
rect 36857 4090 36868 4093
rect 36347 4044 36393 4055
rect 36255 3870 36347 4044
rect 36347 3859 36393 3870
rect 36531 4044 36577 4055
rect 36531 3859 36577 3870
rect 36715 4044 36761 4055
rect 36899 4044 36945 4055
rect 36882 4017 36899 4019
rect 36945 4017 36962 4019
rect 36882 3897 36894 4017
rect 36950 3897 36962 4017
rect 36882 3895 36899 3897
rect 36715 3859 36761 3870
rect 36945 3895 36962 3897
rect 36899 3859 36945 3870
rect 36209 3642 36255 3787
rect 36424 3778 36435 3824
rect 36489 3778 36500 3824
rect 36424 3745 36500 3778
rect 36608 3778 36619 3824
rect 36673 3778 36684 3824
rect 36608 3745 36684 3778
rect 36792 3778 36803 3824
rect 36857 3778 36868 3824
rect 36792 3745 36868 3778
rect 37037 3642 37083 3787
rect 36197 3630 36277 3642
rect 36197 3574 36209 3630
rect 36265 3574 36277 3630
rect 36197 3562 36277 3574
rect 37015 3630 37093 3642
rect 37015 3574 37027 3630
rect 37083 3574 37093 3630
rect 37015 3562 37093 3574
rect 38122 3511 38322 4311
rect 38522 3511 38722 4311
rect 38122 2891 38722 3511
rect 39053 4171 39099 4182
rect 39268 4180 39364 4211
rect 39268 4134 39279 4180
rect 39353 4134 39364 4180
rect 39533 4171 39987 4311
rect 39191 4088 39237 4099
rect 39174 3804 39191 3814
rect 39395 4088 39533 4099
rect 39237 3804 39254 3814
rect 39174 3564 39186 3804
rect 39242 3564 39254 3804
rect 39174 3554 39191 3564
rect 39237 3554 39254 3564
rect 39191 3503 39237 3514
rect 39441 3514 39533 4088
rect 39395 3503 39533 3514
rect 39053 3420 39099 3431
rect 39268 3422 39279 3468
rect 39353 3422 39364 3468
rect 39268 3347 39364 3422
rect 39579 3503 39941 4171
rect 39533 3420 39579 3431
rect 40156 4180 40252 4211
rect 40156 4134 40167 4180
rect 40241 4134 40252 4180
rect 40421 4171 40467 4311
rect 39987 4088 40125 4099
rect 39987 3514 40079 4088
rect 40283 4088 40329 4099
rect 40266 3804 40283 3814
rect 40329 3804 40346 3814
rect 40266 3564 40278 3804
rect 40334 3564 40346 3804
rect 40266 3554 40283 3564
rect 39987 3503 40125 3514
rect 40329 3554 40346 3564
rect 40283 3503 40329 3514
rect 39941 3420 39987 3431
rect 40156 3422 40167 3468
rect 40241 3422 40252 3468
rect 39268 3291 39288 3347
rect 39344 3291 39364 3347
rect 39268 3073 39364 3291
rect 40156 3203 40252 3422
rect 40636 4180 40732 4211
rect 40636 4134 40647 4180
rect 40721 4134 40732 4180
rect 40901 4171 40947 4311
rect 40467 4088 40605 4099
rect 40467 3514 40559 4088
rect 40763 4088 40809 4099
rect 40746 3804 40763 3814
rect 40809 3804 40826 3814
rect 40746 3564 40758 3804
rect 40814 3564 40826 3804
rect 40746 3554 40763 3564
rect 40467 3503 40605 3514
rect 40809 3554 40826 3564
rect 40763 3503 40809 3514
rect 40421 3420 40467 3431
rect 40636 3422 40647 3468
rect 40721 3422 40732 3468
rect 40636 3281 40732 3422
rect 40901 3420 40947 3431
rect 41244 3511 42712 4311
rect 43012 3511 43212 4311
rect 47594 4311 52684 4511
rect 53356 4414 53412 5661
rect 56312 5659 56392 5661
rect 54836 5606 54906 5608
rect 56136 5607 56216 5609
rect 53492 5550 54838 5606
rect 54894 5550 54906 5606
rect 53492 4530 53548 5550
rect 54836 5538 54906 5550
rect 54978 5551 56148 5607
rect 56204 5551 56216 5607
rect 54156 5499 54242 5503
rect 54156 5443 54168 5499
rect 54224 5443 54242 5499
rect 54156 5431 54242 5443
rect 53667 5286 53713 5297
rect 53882 5295 53958 5328
rect 53882 5249 53893 5295
rect 53947 5249 53958 5295
rect 54066 5295 54142 5328
rect 54066 5249 54077 5295
rect 54131 5249 54142 5295
rect 54250 5295 54326 5328
rect 54250 5249 54261 5295
rect 54315 5249 54326 5295
rect 54495 5286 54541 5297
rect 53805 5203 53851 5214
rect 53788 5176 53805 5178
rect 53989 5203 54035 5214
rect 53851 5176 53868 5178
rect 53713 5056 53800 5176
rect 53856 5056 53868 5176
rect 53788 5054 53805 5056
rect 53713 4756 53805 4876
rect 53851 5054 53868 5056
rect 53972 4876 53989 4878
rect 54173 5203 54219 5214
rect 54156 5176 54173 5178
rect 54357 5203 54403 5214
rect 54219 5176 54236 5178
rect 54156 5056 54168 5176
rect 54224 5056 54236 5176
rect 54156 5054 54173 5056
rect 54035 4876 54052 4878
rect 53972 4756 53984 4876
rect 54040 4756 54052 4876
rect 53972 4754 53989 4756
rect 53805 4718 53851 4729
rect 54035 4754 54052 4756
rect 53989 4718 54035 4729
rect 54219 5054 54236 5056
rect 54340 4876 54357 4878
rect 54478 5176 54495 5178
rect 54541 5176 54558 5178
rect 54478 5055 54490 5176
rect 54546 5055 54558 5176
rect 54478 5053 54495 5055
rect 54403 4876 54420 4878
rect 54340 4756 54352 4876
rect 54408 4756 54420 4876
rect 54340 4754 54357 4756
rect 54173 4718 54219 4729
rect 54403 4754 54420 4756
rect 54357 4718 54403 4729
rect 53882 4680 53893 4683
rect 53947 4680 53958 4683
rect 54066 4680 54077 4683
rect 54131 4680 54142 4683
rect 54250 4680 54261 4683
rect 54315 4680 54326 4683
rect 53667 4635 53713 4646
rect 53880 4624 53892 4680
rect 53948 4624 53960 4680
rect 53880 4610 53960 4624
rect 54064 4624 54076 4680
rect 54132 4624 54144 4680
rect 54064 4610 54144 4624
rect 54248 4624 54260 4680
rect 54316 4624 54328 4680
rect 54541 5053 54558 5055
rect 54495 4635 54541 4646
rect 54248 4610 54328 4624
rect 53880 4530 53960 4532
rect 53492 4474 53892 4530
rect 53948 4474 53960 4530
rect 54978 4531 55034 5551
rect 56136 5539 56216 5551
rect 55642 5500 55728 5504
rect 55642 5444 55654 5500
rect 55710 5444 55728 5500
rect 55642 5432 55728 5444
rect 55153 5287 55199 5298
rect 55368 5296 55444 5329
rect 55368 5250 55379 5296
rect 55433 5250 55444 5296
rect 55552 5296 55628 5329
rect 55552 5250 55563 5296
rect 55617 5250 55628 5296
rect 55736 5296 55812 5329
rect 55736 5250 55747 5296
rect 55801 5250 55812 5296
rect 55981 5287 56027 5298
rect 55291 5204 55337 5215
rect 55274 5177 55291 5179
rect 55475 5204 55521 5215
rect 55337 5177 55354 5179
rect 55199 5057 55286 5177
rect 55342 5057 55354 5177
rect 55274 5055 55291 5057
rect 55199 4757 55291 4877
rect 55337 5055 55354 5057
rect 55458 4877 55475 4879
rect 55659 5204 55705 5215
rect 55642 5177 55659 5179
rect 55843 5204 55889 5215
rect 55705 5177 55722 5179
rect 55642 5057 55654 5177
rect 55710 5057 55722 5177
rect 55642 5055 55659 5057
rect 55521 4877 55538 4879
rect 55458 4757 55470 4877
rect 55526 4757 55538 4877
rect 55458 4755 55475 4757
rect 55291 4719 55337 4730
rect 55521 4755 55538 4757
rect 55475 4719 55521 4730
rect 55705 5055 55722 5057
rect 55826 4877 55843 4879
rect 55964 5177 55981 5179
rect 56027 5177 56044 5179
rect 55964 5056 55976 5177
rect 56032 5056 56044 5177
rect 55964 5054 55981 5056
rect 55889 4877 55906 4879
rect 55826 4757 55838 4877
rect 55894 4757 55906 4877
rect 55826 4755 55843 4757
rect 55659 4719 55705 4730
rect 55889 4755 55906 4757
rect 55843 4719 55889 4730
rect 55368 4681 55379 4684
rect 55433 4681 55444 4684
rect 55552 4681 55563 4684
rect 55617 4681 55628 4684
rect 55736 4681 55747 4684
rect 55801 4681 55812 4684
rect 55153 4636 55199 4647
rect 55366 4625 55378 4681
rect 55434 4625 55446 4681
rect 55366 4611 55446 4625
rect 55550 4625 55562 4681
rect 55618 4625 55630 4681
rect 55550 4611 55630 4625
rect 55734 4625 55746 4681
rect 55802 4625 55814 4681
rect 56027 5054 56044 5056
rect 55981 4636 56027 4647
rect 55734 4611 55814 4625
rect 55366 4531 55446 4533
rect 54978 4475 55378 4531
rect 55434 4475 55446 4531
rect 53880 4472 53960 4474
rect 55366 4473 55446 4475
rect 54064 4414 54144 4416
rect 53356 4358 54076 4414
rect 54132 4358 54144 4414
rect 54064 4356 54144 4358
rect 54393 4414 54473 4416
rect 54660 4415 54730 4426
rect 55550 4415 55630 4417
rect 54660 4414 55562 4415
rect 54393 4358 54405 4414
rect 54461 4358 54662 4414
rect 54718 4359 55562 4414
rect 55618 4359 55630 4415
rect 54718 4358 54978 4359
rect 54393 4356 54473 4358
rect 54660 4348 54730 4358
rect 55550 4357 55630 4359
rect 55879 4415 55959 4417
rect 56322 4415 56392 4425
rect 55879 4359 55891 4415
rect 55947 4359 56324 4415
rect 56380 4359 56392 4415
rect 55879 4357 55959 4359
rect 56322 4347 56392 4359
rect 43736 4298 43806 4310
rect 44776 4298 44856 4300
rect 46262 4299 46342 4301
rect 43736 4242 43748 4298
rect 43804 4242 44788 4298
rect 44844 4242 44856 4298
rect 43736 4230 43806 4242
rect 40088 3191 40252 3203
rect 40568 3269 40732 3281
rect 40568 3213 40580 3269
rect 40636 3213 40732 3269
rect 40568 3201 40732 3213
rect 40088 3135 40100 3191
rect 40156 3135 40252 3191
rect 40088 3123 40252 3135
rect 40156 3073 40252 3123
rect 39053 3051 39099 3062
rect 38159 2751 38205 2891
rect 38374 2760 38470 2791
rect 38374 2714 38385 2760
rect 38459 2714 38470 2760
rect 38639 2751 38685 2891
rect 38205 2668 38343 2679
rect 38205 2094 38297 2668
rect 38501 2668 38547 2679
rect 38484 2384 38501 2394
rect 38547 2384 38564 2394
rect 38484 2144 38496 2384
rect 38552 2144 38564 2384
rect 38484 2134 38501 2144
rect 38205 2083 38343 2094
rect 38547 2134 38564 2144
rect 38501 2083 38547 2094
rect 38159 2000 38205 2011
rect 38374 2002 38385 2048
rect 38459 2002 38470 2048
rect 38374 1861 38470 2002
rect 39268 3060 39568 3073
rect 39268 3014 39279 3060
rect 39353 3027 39483 3060
rect 39353 3014 39364 3027
rect 39472 3014 39483 3027
rect 39557 3014 39568 3060
rect 39737 3051 39783 3062
rect 39099 2968 39237 2979
rect 39099 2794 39191 2968
rect 39395 2968 39441 2979
rect 39378 2909 39395 2919
rect 39599 2968 39737 2979
rect 39441 2909 39458 2919
rect 39378 2853 39390 2909
rect 39446 2853 39458 2909
rect 39378 2843 39395 2853
rect 39099 2783 39237 2794
rect 39441 2843 39458 2853
rect 39395 2783 39441 2794
rect 39645 2794 39737 2968
rect 39599 2783 39737 2794
rect 39053 2571 39099 2711
rect 39268 2702 39279 2748
rect 39353 2702 39364 2748
rect 39268 2671 39364 2702
rect 39472 2702 39483 2748
rect 39557 2702 39568 2748
rect 39472 2671 39568 2702
rect 39952 3060 40252 3073
rect 39952 3014 39963 3060
rect 40037 3027 40167 3060
rect 40037 3014 40048 3027
rect 40156 3014 40167 3027
rect 40241 3014 40252 3060
rect 40421 3051 40467 3062
rect 39875 2968 39921 2979
rect 39858 2909 39875 2919
rect 40079 2968 40125 2979
rect 39921 2909 39938 2919
rect 39858 2853 39870 2909
rect 39926 2853 39938 2909
rect 39858 2843 39875 2853
rect 39921 2843 39938 2853
rect 40062 2909 40079 2919
rect 40283 2968 40329 2979
rect 40125 2909 40142 2919
rect 40062 2853 40074 2909
rect 40130 2853 40142 2909
rect 40062 2843 40079 2853
rect 39875 2783 39921 2794
rect 40125 2843 40142 2853
rect 40266 2909 40283 2919
rect 40329 2909 40346 2919
rect 40266 2853 40278 2909
rect 40334 2853 40346 2909
rect 40266 2843 40283 2853
rect 40079 2783 40125 2794
rect 40329 2843 40346 2853
rect 40283 2783 40329 2794
rect 39737 2571 39783 2711
rect 39952 2702 39963 2748
rect 40037 2702 40048 2748
rect 39952 2671 40048 2702
rect 40156 2702 40167 2748
rect 40241 2702 40252 2748
rect 40156 2671 40252 2702
rect 40636 3060 40732 3201
rect 41244 3315 43212 3511
rect 44020 3511 44076 4242
rect 44776 4240 44856 4242
rect 45506 4243 46274 4299
rect 46330 4243 46342 4299
rect 44408 4148 44488 4162
rect 44195 4126 44241 4137
rect 44408 4092 44420 4148
rect 44476 4092 44488 4148
rect 44592 4148 44672 4162
rect 44592 4092 44604 4148
rect 44660 4092 44672 4148
rect 44776 4148 44856 4162
rect 44776 4092 44788 4148
rect 44844 4092 44856 4148
rect 45023 4126 45069 4137
rect 44410 4089 44421 4092
rect 44475 4089 44486 4092
rect 44594 4089 44605 4092
rect 44659 4089 44670 4092
rect 44778 4089 44789 4092
rect 44843 4089 44854 4092
rect 44333 4043 44379 4054
rect 44241 3869 44333 4043
rect 44333 3858 44379 3869
rect 44517 4043 44563 4054
rect 44517 3858 44563 3869
rect 44701 4043 44747 4054
rect 44885 4043 44931 4054
rect 44868 4016 44885 4018
rect 44931 4016 44948 4018
rect 44868 3896 44880 4016
rect 44936 3896 44948 4016
rect 44868 3894 44885 3896
rect 44701 3858 44747 3869
rect 44931 3894 44948 3896
rect 44885 3858 44931 3869
rect 44195 3641 44241 3786
rect 44410 3777 44421 3823
rect 44475 3777 44486 3823
rect 44410 3744 44486 3777
rect 44594 3777 44605 3823
rect 44659 3777 44670 3823
rect 44594 3744 44670 3777
rect 44778 3777 44789 3823
rect 44843 3777 44854 3823
rect 44778 3744 44854 3777
rect 45023 3641 45069 3786
rect 44183 3629 44263 3641
rect 44183 3573 44195 3629
rect 44251 3573 44263 3629
rect 44183 3561 44263 3573
rect 45001 3629 45079 3641
rect 45001 3573 45013 3629
rect 45069 3573 45079 3629
rect 45001 3561 45079 3573
rect 45354 3511 45434 3521
rect 44020 3455 45366 3511
rect 45422 3455 45434 3511
rect 45354 3453 45434 3455
rect 45188 3402 45258 3404
rect 41244 3175 41344 3315
rect 43112 3175 43212 3315
rect 41244 3135 43212 3175
rect 44020 3401 45258 3402
rect 44020 3347 45190 3401
rect 45246 3347 45258 3401
rect 44020 3346 45258 3347
rect 40636 3014 40647 3060
rect 40721 3014 40732 3060
rect 40901 3051 40947 3062
rect 40467 2968 40605 2979
rect 40467 2794 40559 2968
rect 40763 2968 40809 2979
rect 40746 2909 40763 2919
rect 40809 2909 40826 2919
rect 40746 2853 40758 2909
rect 40814 2853 40826 2909
rect 40746 2843 40763 2853
rect 40467 2783 40605 2794
rect 40809 2843 40826 2853
rect 40763 2783 40809 2794
rect 40421 2571 40467 2711
rect 40636 2702 40647 2748
rect 40721 2702 40732 2748
rect 40636 2671 40732 2702
rect 40901 2571 40947 2711
rect 41281 2995 41327 3135
rect 39016 2541 40984 2571
rect 39016 2401 40284 2541
rect 40884 2401 40984 2541
rect 39016 2371 40984 2401
rect 41496 3004 41592 3035
rect 41496 2958 41507 3004
rect 41581 2958 41592 3004
rect 41700 3004 41796 3035
rect 41700 2958 41711 3004
rect 41785 2958 41796 3004
rect 41965 2995 42011 3135
rect 41327 2912 41465 2923
rect 41623 2912 41669 2923
rect 41827 2912 41965 2923
rect 41327 2338 41419 2912
rect 41606 2672 41618 2912
rect 41674 2672 41686 2912
rect 41327 2327 41465 2338
rect 41623 2327 41669 2338
rect 41873 2338 41965 2912
rect 41827 2327 41965 2338
rect 41281 2244 41327 2255
rect 41496 2246 41507 2292
rect 41581 2272 41592 2292
rect 41700 2272 41711 2292
rect 41581 2246 41711 2272
rect 41785 2246 41796 2292
rect 41496 2219 41796 2246
rect 42180 3004 42276 3035
rect 42180 2958 42191 3004
rect 42265 2958 42276 3004
rect 42384 3004 42480 3035
rect 42384 2958 42395 3004
rect 42469 2958 42480 3004
rect 42649 2995 42695 3135
rect 42103 2912 42149 2923
rect 42307 2912 42353 2923
rect 42511 2912 42557 2923
rect 42290 2672 42302 2912
rect 42358 2672 42370 2912
rect 42086 2338 42098 2578
rect 42154 2338 42166 2578
rect 42494 2338 42506 2578
rect 42562 2338 42574 2578
rect 42103 2327 42149 2338
rect 42307 2327 42353 2338
rect 42511 2327 42557 2338
rect 41965 2244 42011 2255
rect 42180 2246 42191 2292
rect 42265 2272 42276 2292
rect 42384 2272 42395 2292
rect 42265 2246 42395 2272
rect 42469 2246 42480 2292
rect 42180 2219 42480 2246
rect 42864 3004 42960 3035
rect 42864 2958 42875 3004
rect 42949 2958 42960 3004
rect 43129 2995 43175 3135
rect 42695 2912 42833 2923
rect 42695 2338 42787 2912
rect 42991 2912 43037 2923
rect 42974 2628 42991 2638
rect 43037 2628 43054 2638
rect 42974 2388 42986 2628
rect 43042 2388 43054 2628
rect 42974 2378 42991 2388
rect 42695 2327 42833 2338
rect 43037 2378 43054 2388
rect 42991 2327 43037 2338
rect 42649 2244 42695 2255
rect 42864 2246 42875 2292
rect 42949 2246 42960 2292
rect 41496 2171 41592 2219
rect 38639 2000 38685 2011
rect 39016 2141 40984 2171
rect 39016 2001 40284 2141
rect 40884 2001 40984 2141
rect 39016 1971 40984 2001
rect 41496 2115 41516 2171
rect 41572 2115 41592 2171
rect 38306 1849 38470 1861
rect 38306 1793 38318 1849
rect 38374 1793 38470 1849
rect 38306 1781 38470 1793
rect 33945 1250 33957 1306
rect 34013 1250 34140 1306
rect 34196 1250 36090 1306
rect 38159 1631 38205 1642
rect 38374 1640 38470 1781
rect 39053 1831 39099 1842
rect 38374 1594 38385 1640
rect 38459 1594 38470 1640
rect 38639 1631 38685 1642
rect 38205 1548 38343 1559
rect 38205 1374 38297 1548
rect 38501 1548 38547 1559
rect 38484 1489 38501 1499
rect 38547 1489 38564 1499
rect 38484 1433 38496 1489
rect 38552 1433 38564 1489
rect 38484 1423 38501 1433
rect 38205 1363 38343 1374
rect 38547 1423 38564 1433
rect 38501 1363 38547 1374
rect 33945 1238 34031 1250
rect 34138 1238 34198 1250
rect 30616 851 30780 863
rect 31096 929 31260 941
rect 31096 873 31108 929
rect 31164 873 31260 929
rect 31096 861 31260 873
rect 30616 795 30628 851
rect 30684 795 30780 851
rect 30616 783 30780 795
rect 30684 733 30780 783
rect 24068 231 29250 431
rect 29581 711 29627 722
rect 29796 720 30096 733
rect 29796 674 29807 720
rect 29881 687 30011 720
rect 29881 674 29892 687
rect 30000 674 30011 687
rect 30085 674 30096 720
rect 30265 711 30311 722
rect 29627 628 29765 639
rect 29627 454 29719 628
rect 29923 628 29969 639
rect 29906 569 29923 579
rect 30127 628 30265 639
rect 29969 569 29986 579
rect 29906 513 29918 569
rect 29974 513 29986 569
rect 29906 503 29923 513
rect 29627 443 29765 454
rect 29969 503 29986 513
rect 29923 443 29969 454
rect 30173 454 30265 628
rect 30127 443 30265 454
rect 29581 231 29627 371
rect 29796 362 29807 408
rect 29881 362 29892 408
rect 29796 331 29892 362
rect 30000 362 30011 408
rect 30085 362 30096 408
rect 30000 331 30096 362
rect 30480 720 30780 733
rect 30480 674 30491 720
rect 30565 687 30695 720
rect 30565 674 30576 687
rect 30684 674 30695 687
rect 30769 674 30780 720
rect 30949 711 30995 722
rect 30403 628 30449 639
rect 30386 569 30403 579
rect 30607 628 30653 639
rect 30449 569 30466 579
rect 30386 513 30398 569
rect 30454 513 30466 569
rect 30386 503 30403 513
rect 30449 503 30466 513
rect 30590 569 30607 579
rect 30811 628 30857 639
rect 30653 569 30670 579
rect 30590 513 30602 569
rect 30658 513 30670 569
rect 30590 503 30607 513
rect 30403 443 30449 454
rect 30653 503 30670 513
rect 30794 569 30811 579
rect 30857 569 30874 579
rect 30794 513 30806 569
rect 30862 513 30874 569
rect 30794 503 30811 513
rect 30607 443 30653 454
rect 30857 503 30874 513
rect 30811 443 30857 454
rect 30265 231 30311 371
rect 30480 362 30491 408
rect 30565 362 30576 408
rect 30480 331 30576 362
rect 30684 362 30695 408
rect 30769 362 30780 408
rect 30684 331 30780 362
rect 31164 720 31260 861
rect 31772 1031 33740 1215
rect 38159 1151 38205 1291
rect 38374 1282 38385 1328
rect 38459 1282 38470 1328
rect 38374 1251 38470 1282
rect 38639 1151 38685 1291
rect 31164 674 31175 720
rect 31249 674 31260 720
rect 31429 711 31475 722
rect 30995 628 31133 639
rect 30995 454 31087 628
rect 31291 628 31337 639
rect 31274 569 31291 579
rect 31337 569 31354 579
rect 31274 513 31286 569
rect 31342 513 31354 569
rect 31274 503 31291 513
rect 30995 443 31133 454
rect 31337 503 31354 513
rect 31291 443 31337 454
rect 30949 231 30995 371
rect 31164 362 31175 408
rect 31249 362 31260 408
rect 31164 331 31260 362
rect 31429 231 31475 371
rect 31772 231 33240 1031
rect 33540 431 33740 1031
rect 38122 431 38722 1151
rect 39268 1840 39364 1871
rect 39268 1794 39279 1840
rect 39353 1794 39364 1840
rect 39533 1831 39987 1971
rect 39191 1748 39237 1759
rect 39174 1464 39191 1474
rect 39395 1748 39533 1759
rect 39237 1464 39254 1474
rect 39174 1224 39186 1464
rect 39242 1224 39254 1464
rect 39174 1214 39191 1224
rect 39237 1214 39254 1224
rect 39191 1163 39237 1174
rect 39441 1174 39533 1748
rect 39395 1163 39533 1174
rect 39053 1080 39099 1091
rect 39268 1082 39279 1128
rect 39353 1082 39364 1128
rect 39268 1007 39364 1082
rect 39579 1163 39941 1831
rect 39533 1080 39579 1091
rect 40156 1840 40252 1871
rect 40156 1794 40167 1840
rect 40241 1794 40252 1840
rect 40421 1831 40467 1971
rect 39987 1748 40125 1759
rect 39987 1174 40079 1748
rect 40283 1748 40329 1759
rect 40266 1464 40283 1474
rect 40329 1464 40346 1474
rect 40266 1224 40278 1464
rect 40334 1224 40346 1464
rect 40266 1214 40283 1224
rect 39987 1163 40125 1174
rect 40329 1214 40346 1224
rect 40283 1163 40329 1174
rect 39941 1080 39987 1091
rect 40156 1082 40167 1128
rect 40241 1082 40252 1128
rect 39268 951 39288 1007
rect 39344 951 39364 1007
rect 39268 733 39364 951
rect 40156 863 40252 1082
rect 40636 1840 40732 1871
rect 40636 1794 40647 1840
rect 40721 1794 40732 1840
rect 40901 1831 40947 1971
rect 40467 1748 40605 1759
rect 40467 1174 40559 1748
rect 40763 1748 40809 1759
rect 40746 1464 40763 1474
rect 40809 1464 40826 1474
rect 40746 1224 40758 1464
rect 40814 1224 40826 1464
rect 40746 1214 40763 1224
rect 40467 1163 40605 1174
rect 40809 1214 40826 1224
rect 40763 1163 40809 1174
rect 40421 1080 40467 1091
rect 40636 1082 40647 1128
rect 40721 1082 40732 1128
rect 40636 941 40732 1082
rect 41281 1875 41327 1886
rect 41496 1884 41592 2115
rect 42180 2015 42276 2219
rect 42864 2105 42960 2246
rect 44020 2325 44076 3346
rect 45188 3338 45258 3346
rect 44684 3294 44770 3298
rect 44684 3238 44696 3294
rect 44752 3238 44770 3294
rect 44684 3226 44770 3238
rect 44195 3081 44241 3092
rect 44410 3090 44486 3123
rect 44410 3044 44421 3090
rect 44475 3044 44486 3090
rect 44594 3090 44670 3123
rect 44594 3044 44605 3090
rect 44659 3044 44670 3090
rect 44778 3090 44854 3123
rect 44778 3044 44789 3090
rect 44843 3044 44854 3090
rect 45023 3081 45069 3092
rect 44333 2998 44379 3009
rect 44316 2971 44333 2973
rect 44517 2998 44563 3009
rect 44379 2971 44396 2973
rect 44241 2851 44328 2971
rect 44384 2851 44396 2971
rect 44316 2849 44333 2851
rect 44241 2551 44333 2671
rect 44379 2849 44396 2851
rect 44500 2671 44517 2673
rect 44701 2998 44747 3009
rect 44684 2971 44701 2973
rect 44885 2998 44931 3009
rect 44747 2971 44764 2973
rect 44684 2851 44696 2971
rect 44752 2851 44764 2971
rect 44684 2849 44701 2851
rect 44563 2671 44580 2673
rect 44500 2551 44512 2671
rect 44568 2551 44580 2671
rect 44500 2549 44517 2551
rect 44333 2513 44379 2524
rect 44563 2549 44580 2551
rect 44517 2513 44563 2524
rect 44747 2849 44764 2851
rect 44868 2671 44885 2673
rect 45006 2971 45023 2973
rect 45069 2971 45086 2973
rect 45006 2850 45018 2971
rect 45074 2850 45086 2971
rect 45006 2848 45023 2850
rect 44931 2671 44948 2673
rect 44868 2551 44880 2671
rect 44936 2551 44948 2671
rect 44868 2549 44885 2551
rect 44701 2513 44747 2524
rect 44931 2549 44948 2551
rect 44885 2513 44931 2524
rect 44410 2475 44421 2478
rect 44475 2475 44486 2478
rect 44594 2475 44605 2478
rect 44659 2475 44670 2478
rect 44778 2475 44789 2478
rect 44843 2475 44854 2478
rect 44195 2430 44241 2441
rect 44408 2419 44420 2475
rect 44476 2419 44488 2475
rect 44408 2405 44488 2419
rect 44592 2419 44604 2475
rect 44660 2419 44672 2475
rect 44592 2405 44672 2419
rect 44776 2419 44788 2475
rect 44844 2419 44856 2475
rect 45069 2848 45086 2850
rect 45023 2430 45069 2441
rect 44776 2405 44856 2419
rect 44408 2325 44488 2327
rect 44020 2269 44420 2325
rect 44476 2269 44488 2325
rect 44408 2267 44488 2269
rect 43129 2244 43175 2255
rect 43600 2209 43670 2223
rect 44592 2209 44672 2211
rect 43600 2153 43612 2209
rect 43668 2153 44604 2209
rect 44660 2153 44672 2209
rect 43600 2141 43670 2153
rect 44592 2151 44672 2153
rect 44921 2209 45001 2211
rect 45364 2209 45424 2221
rect 44921 2153 44933 2209
rect 44989 2153 45366 2209
rect 45422 2153 45424 2209
rect 44921 2151 45001 2153
rect 45364 2141 45424 2153
rect 42796 2093 42960 2105
rect 42796 2037 42808 2093
rect 42864 2037 42960 2093
rect 42796 2025 42960 2037
rect 43366 2093 43444 2104
rect 44776 2093 44856 2095
rect 43366 2092 44788 2093
rect 43366 2038 43378 2092
rect 43432 2038 44788 2092
rect 43366 2037 44788 2038
rect 44844 2037 44856 2093
rect 43366 2026 43444 2037
rect 44776 2035 44856 2037
rect 42180 1959 42200 2015
rect 42256 1959 42276 2015
rect 41496 1838 41507 1884
rect 41581 1838 41592 1884
rect 41761 1875 42011 1886
rect 41419 1792 41465 1803
rect 41402 1733 41419 1743
rect 41623 1792 41761 1803
rect 41465 1733 41482 1743
rect 41402 1677 41414 1733
rect 41470 1677 41482 1733
rect 41402 1667 41419 1677
rect 41465 1667 41482 1677
rect 41419 1607 41465 1618
rect 41669 1618 41761 1792
rect 41623 1607 41761 1618
rect 41281 1395 41327 1535
rect 41496 1526 41507 1572
rect 41581 1526 41592 1572
rect 41496 1495 41592 1526
rect 41807 1535 41965 1875
rect 42180 1884 42276 1959
rect 42180 1838 42191 1884
rect 42265 1838 42276 1884
rect 42445 1875 42491 1886
rect 42011 1792 42149 1803
rect 42011 1618 42103 1792
rect 42307 1792 42353 1803
rect 42290 1733 42307 1743
rect 42353 1733 42370 1743
rect 42290 1677 42302 1733
rect 42358 1677 42370 1733
rect 42290 1667 42307 1677
rect 42011 1607 42149 1618
rect 42353 1667 42370 1677
rect 42307 1607 42353 1618
rect 41761 1524 42011 1535
rect 42180 1526 42191 1572
rect 42265 1526 42276 1572
rect 41807 1395 41965 1524
rect 42180 1495 42276 1526
rect 42445 1395 42491 1535
rect 42649 1875 42695 1886
rect 42864 1884 42960 2025
rect 44408 1943 44488 1957
rect 44195 1921 44241 1932
rect 42864 1838 42875 1884
rect 42949 1838 42960 1884
rect 43129 1875 43175 1886
rect 42695 1792 42833 1803
rect 42695 1618 42787 1792
rect 42991 1792 43037 1803
rect 42974 1733 42991 1743
rect 43037 1733 43054 1743
rect 42974 1677 42986 1733
rect 43042 1677 43054 1733
rect 42974 1667 42991 1677
rect 42695 1607 42833 1618
rect 43037 1667 43054 1677
rect 42991 1607 43037 1618
rect 42649 1395 42695 1535
rect 42864 1526 42875 1572
rect 42949 1526 42960 1572
rect 42864 1495 42960 1526
rect 43129 1395 43175 1535
rect 44408 1887 44420 1943
rect 44476 1887 44488 1943
rect 44592 1943 44672 1957
rect 44592 1887 44604 1943
rect 44660 1887 44672 1943
rect 44776 1943 44856 1957
rect 44776 1887 44788 1943
rect 44844 1887 44856 1943
rect 45023 1921 45069 1932
rect 44410 1884 44421 1887
rect 44475 1884 44486 1887
rect 44594 1884 44605 1887
rect 44659 1884 44670 1887
rect 44778 1884 44789 1887
rect 44843 1884 44854 1887
rect 44333 1838 44379 1849
rect 44241 1664 44333 1838
rect 44333 1653 44379 1664
rect 44517 1838 44563 1849
rect 44517 1653 44563 1664
rect 44701 1838 44747 1849
rect 44885 1838 44931 1849
rect 44868 1811 44885 1813
rect 44931 1811 44948 1813
rect 44868 1691 44880 1811
rect 44936 1691 44948 1811
rect 44868 1689 44885 1691
rect 44701 1653 44747 1664
rect 44931 1689 44948 1691
rect 44885 1653 44931 1664
rect 44195 1436 44241 1581
rect 44410 1572 44421 1618
rect 44475 1572 44486 1618
rect 44410 1539 44486 1572
rect 44594 1572 44605 1618
rect 44659 1572 44670 1618
rect 44594 1539 44670 1572
rect 44778 1572 44789 1618
rect 44843 1572 44854 1618
rect 44778 1539 44854 1572
rect 45023 1436 45069 1581
rect 44183 1424 44263 1436
rect 40901 1080 40947 1091
rect 41244 1355 43212 1395
rect 44183 1368 44195 1424
rect 44251 1368 44263 1424
rect 44183 1356 44263 1368
rect 45001 1424 45081 1436
rect 45001 1368 45013 1424
rect 45069 1368 45081 1424
rect 45001 1356 45081 1368
rect 41244 1215 41344 1355
rect 43112 1215 43212 1355
rect 43417 1306 43503 1318
rect 43610 1306 43670 1310
rect 45506 1306 45562 4243
rect 46262 4241 46342 4243
rect 45894 4149 45974 4163
rect 45681 4127 45727 4138
rect 45894 4093 45906 4149
rect 45962 4093 45974 4149
rect 46078 4149 46158 4163
rect 46078 4093 46090 4149
rect 46146 4093 46158 4149
rect 46262 4149 46342 4163
rect 46262 4093 46274 4149
rect 46330 4093 46342 4149
rect 46509 4127 46555 4138
rect 45896 4090 45907 4093
rect 45961 4090 45972 4093
rect 46080 4090 46091 4093
rect 46145 4090 46156 4093
rect 46264 4090 46275 4093
rect 46329 4090 46340 4093
rect 45819 4044 45865 4055
rect 45727 3870 45819 4044
rect 45819 3859 45865 3870
rect 46003 4044 46049 4055
rect 46003 3859 46049 3870
rect 46187 4044 46233 4055
rect 46371 4044 46417 4055
rect 46354 4017 46371 4019
rect 46417 4017 46434 4019
rect 46354 3897 46366 4017
rect 46422 3897 46434 4017
rect 46354 3895 46371 3897
rect 46187 3859 46233 3870
rect 46417 3895 46434 3897
rect 46371 3859 46417 3870
rect 45681 3642 45727 3787
rect 45896 3778 45907 3824
rect 45961 3778 45972 3824
rect 45896 3745 45972 3778
rect 46080 3778 46091 3824
rect 46145 3778 46156 3824
rect 46080 3745 46156 3778
rect 46264 3778 46275 3824
rect 46329 3778 46340 3824
rect 46264 3745 46340 3778
rect 46509 3642 46555 3787
rect 45669 3630 45749 3642
rect 45669 3574 45681 3630
rect 45737 3574 45749 3630
rect 45669 3562 45749 3574
rect 46487 3630 46565 3642
rect 46487 3574 46499 3630
rect 46555 3574 46565 3630
rect 46487 3562 46565 3574
rect 47594 3511 47794 4311
rect 47994 3511 48194 4311
rect 47594 2891 48194 3511
rect 48525 4171 48571 4182
rect 48740 4180 48836 4211
rect 48740 4134 48751 4180
rect 48825 4134 48836 4180
rect 49005 4171 49459 4311
rect 48663 4088 48709 4099
rect 48646 3804 48663 3814
rect 48867 4088 49005 4099
rect 48709 3804 48726 3814
rect 48646 3564 48658 3804
rect 48714 3564 48726 3804
rect 48646 3554 48663 3564
rect 48709 3554 48726 3564
rect 48663 3503 48709 3514
rect 48913 3514 49005 4088
rect 48867 3503 49005 3514
rect 48525 3420 48571 3431
rect 48740 3422 48751 3468
rect 48825 3422 48836 3468
rect 48740 3347 48836 3422
rect 49051 3503 49413 4171
rect 49005 3420 49051 3431
rect 49628 4180 49724 4211
rect 49628 4134 49639 4180
rect 49713 4134 49724 4180
rect 49893 4171 49939 4311
rect 49459 4088 49597 4099
rect 49459 3514 49551 4088
rect 49755 4088 49801 4099
rect 49738 3804 49755 3814
rect 49801 3804 49818 3814
rect 49738 3564 49750 3804
rect 49806 3564 49818 3804
rect 49738 3554 49755 3564
rect 49459 3503 49597 3514
rect 49801 3554 49818 3564
rect 49755 3503 49801 3514
rect 49413 3420 49459 3431
rect 49628 3422 49639 3468
rect 49713 3422 49724 3468
rect 48740 3291 48760 3347
rect 48816 3291 48836 3347
rect 48740 3073 48836 3291
rect 49628 3203 49724 3422
rect 50108 4180 50204 4211
rect 50108 4134 50119 4180
rect 50193 4134 50204 4180
rect 50373 4171 50419 4311
rect 49939 4088 50077 4099
rect 49939 3514 50031 4088
rect 50235 4088 50281 4099
rect 50218 3804 50235 3814
rect 50281 3804 50298 3814
rect 50218 3564 50230 3804
rect 50286 3564 50298 3804
rect 50218 3554 50235 3564
rect 49939 3503 50077 3514
rect 50281 3554 50298 3564
rect 50235 3503 50281 3514
rect 49893 3420 49939 3431
rect 50108 3422 50119 3468
rect 50193 3422 50204 3468
rect 50108 3281 50204 3422
rect 50373 3420 50419 3431
rect 50716 3511 52184 4311
rect 52484 3511 52684 4311
rect 53208 4298 53278 4310
rect 54248 4298 54328 4300
rect 55734 4299 55814 4301
rect 53208 4242 53220 4298
rect 53276 4242 54260 4298
rect 54316 4242 54328 4298
rect 53208 4230 53278 4242
rect 49560 3191 49724 3203
rect 50040 3269 50204 3281
rect 50040 3213 50052 3269
rect 50108 3213 50204 3269
rect 50040 3201 50204 3213
rect 49560 3135 49572 3191
rect 49628 3135 49724 3191
rect 49560 3123 49724 3135
rect 49628 3073 49724 3123
rect 48525 3051 48571 3062
rect 47631 2751 47677 2891
rect 47846 2760 47942 2791
rect 47846 2714 47857 2760
rect 47931 2714 47942 2760
rect 48111 2751 48157 2891
rect 47677 2668 47815 2679
rect 47677 2094 47769 2668
rect 47973 2668 48019 2679
rect 47956 2384 47973 2394
rect 48019 2384 48036 2394
rect 47956 2144 47968 2384
rect 48024 2144 48036 2384
rect 47956 2134 47973 2144
rect 47677 2083 47815 2094
rect 48019 2134 48036 2144
rect 47973 2083 48019 2094
rect 47631 2000 47677 2011
rect 47846 2002 47857 2048
rect 47931 2002 47942 2048
rect 47846 1861 47942 2002
rect 48740 3060 49040 3073
rect 48740 3014 48751 3060
rect 48825 3027 48955 3060
rect 48825 3014 48836 3027
rect 48944 3014 48955 3027
rect 49029 3014 49040 3060
rect 49209 3051 49255 3062
rect 48571 2968 48709 2979
rect 48571 2794 48663 2968
rect 48867 2968 48913 2979
rect 48850 2909 48867 2919
rect 49071 2968 49209 2979
rect 48913 2909 48930 2919
rect 48850 2853 48862 2909
rect 48918 2853 48930 2909
rect 48850 2843 48867 2853
rect 48571 2783 48709 2794
rect 48913 2843 48930 2853
rect 48867 2783 48913 2794
rect 49117 2794 49209 2968
rect 49071 2783 49209 2794
rect 48525 2571 48571 2711
rect 48740 2702 48751 2748
rect 48825 2702 48836 2748
rect 48740 2671 48836 2702
rect 48944 2702 48955 2748
rect 49029 2702 49040 2748
rect 48944 2671 49040 2702
rect 49424 3060 49724 3073
rect 49424 3014 49435 3060
rect 49509 3027 49639 3060
rect 49509 3014 49520 3027
rect 49628 3014 49639 3027
rect 49713 3014 49724 3060
rect 49893 3051 49939 3062
rect 49347 2968 49393 2979
rect 49330 2909 49347 2919
rect 49551 2968 49597 2979
rect 49393 2909 49410 2919
rect 49330 2853 49342 2909
rect 49398 2853 49410 2909
rect 49330 2843 49347 2853
rect 49393 2843 49410 2853
rect 49534 2909 49551 2919
rect 49755 2968 49801 2979
rect 49597 2909 49614 2919
rect 49534 2853 49546 2909
rect 49602 2853 49614 2909
rect 49534 2843 49551 2853
rect 49347 2783 49393 2794
rect 49597 2843 49614 2853
rect 49738 2909 49755 2919
rect 49801 2909 49818 2919
rect 49738 2853 49750 2909
rect 49806 2853 49818 2909
rect 49738 2843 49755 2853
rect 49551 2783 49597 2794
rect 49801 2843 49818 2853
rect 49755 2783 49801 2794
rect 49209 2571 49255 2711
rect 49424 2702 49435 2748
rect 49509 2702 49520 2748
rect 49424 2671 49520 2702
rect 49628 2702 49639 2748
rect 49713 2702 49724 2748
rect 49628 2671 49724 2702
rect 50108 3060 50204 3201
rect 50716 3315 52684 3511
rect 53492 3511 53548 4242
rect 54248 4240 54328 4242
rect 54978 4243 55746 4299
rect 55802 4243 55814 4299
rect 53880 4148 53960 4162
rect 53667 4126 53713 4137
rect 53880 4092 53892 4148
rect 53948 4092 53960 4148
rect 54064 4148 54144 4162
rect 54064 4092 54076 4148
rect 54132 4092 54144 4148
rect 54248 4148 54328 4162
rect 54248 4092 54260 4148
rect 54316 4092 54328 4148
rect 54495 4126 54541 4137
rect 53882 4089 53893 4092
rect 53947 4089 53958 4092
rect 54066 4089 54077 4092
rect 54131 4089 54142 4092
rect 54250 4089 54261 4092
rect 54315 4089 54326 4092
rect 53805 4043 53851 4054
rect 53713 3869 53805 4043
rect 53805 3858 53851 3869
rect 53989 4043 54035 4054
rect 53989 3858 54035 3869
rect 54173 4043 54219 4054
rect 54357 4043 54403 4054
rect 54340 4016 54357 4018
rect 54403 4016 54420 4018
rect 54340 3896 54352 4016
rect 54408 3896 54420 4016
rect 54340 3894 54357 3896
rect 54173 3858 54219 3869
rect 54403 3894 54420 3896
rect 54357 3858 54403 3869
rect 53667 3641 53713 3786
rect 53882 3777 53893 3823
rect 53947 3777 53958 3823
rect 53882 3744 53958 3777
rect 54066 3777 54077 3823
rect 54131 3777 54142 3823
rect 54066 3744 54142 3777
rect 54250 3777 54261 3823
rect 54315 3777 54326 3823
rect 54250 3744 54326 3777
rect 54495 3641 54541 3786
rect 53655 3629 53735 3641
rect 53655 3573 53667 3629
rect 53723 3573 53735 3629
rect 53655 3561 53735 3573
rect 54473 3629 54551 3641
rect 54473 3573 54485 3629
rect 54541 3573 54551 3629
rect 54473 3561 54551 3573
rect 54826 3511 54906 3521
rect 53492 3455 54838 3511
rect 54894 3455 54906 3511
rect 54826 3453 54906 3455
rect 54660 3402 54730 3404
rect 50716 3175 50816 3315
rect 52584 3175 52684 3315
rect 50716 3135 52684 3175
rect 53492 3401 54730 3402
rect 53492 3347 54662 3401
rect 54718 3347 54730 3401
rect 53492 3346 54730 3347
rect 50108 3014 50119 3060
rect 50193 3014 50204 3060
rect 50373 3051 50419 3062
rect 49939 2968 50077 2979
rect 49939 2794 50031 2968
rect 50235 2968 50281 2979
rect 50218 2909 50235 2919
rect 50281 2909 50298 2919
rect 50218 2853 50230 2909
rect 50286 2853 50298 2909
rect 50218 2843 50235 2853
rect 49939 2783 50077 2794
rect 50281 2843 50298 2853
rect 50235 2783 50281 2794
rect 49893 2571 49939 2711
rect 50108 2702 50119 2748
rect 50193 2702 50204 2748
rect 50108 2671 50204 2702
rect 50373 2571 50419 2711
rect 50753 2995 50799 3135
rect 48488 2541 50456 2571
rect 48488 2401 49756 2541
rect 50356 2401 50456 2541
rect 48488 2371 50456 2401
rect 50968 3004 51064 3035
rect 50968 2958 50979 3004
rect 51053 2958 51064 3004
rect 51172 3004 51268 3035
rect 51172 2958 51183 3004
rect 51257 2958 51268 3004
rect 51437 2995 51483 3135
rect 50799 2912 50937 2923
rect 51095 2912 51141 2923
rect 51299 2912 51437 2923
rect 50799 2338 50891 2912
rect 51078 2672 51090 2912
rect 51146 2672 51158 2912
rect 50799 2327 50937 2338
rect 51095 2327 51141 2338
rect 51345 2338 51437 2912
rect 51299 2327 51437 2338
rect 50753 2244 50799 2255
rect 50968 2246 50979 2292
rect 51053 2272 51064 2292
rect 51172 2272 51183 2292
rect 51053 2246 51183 2272
rect 51257 2246 51268 2292
rect 50968 2219 51268 2246
rect 51652 3004 51748 3035
rect 51652 2958 51663 3004
rect 51737 2958 51748 3004
rect 51856 3004 51952 3035
rect 51856 2958 51867 3004
rect 51941 2958 51952 3004
rect 52121 2995 52167 3135
rect 51575 2912 51621 2923
rect 51779 2912 51825 2923
rect 51983 2912 52029 2923
rect 51762 2672 51774 2912
rect 51830 2672 51842 2912
rect 51558 2338 51570 2578
rect 51626 2338 51638 2578
rect 51966 2338 51978 2578
rect 52034 2338 52046 2578
rect 51575 2327 51621 2338
rect 51779 2327 51825 2338
rect 51983 2327 52029 2338
rect 51437 2244 51483 2255
rect 51652 2246 51663 2292
rect 51737 2272 51748 2292
rect 51856 2272 51867 2292
rect 51737 2246 51867 2272
rect 51941 2246 51952 2292
rect 51652 2219 51952 2246
rect 52336 3004 52432 3035
rect 52336 2958 52347 3004
rect 52421 2958 52432 3004
rect 52601 2995 52647 3135
rect 52167 2912 52305 2923
rect 52167 2338 52259 2912
rect 52463 2912 52509 2923
rect 52446 2628 52463 2638
rect 52509 2628 52526 2638
rect 52446 2388 52458 2628
rect 52514 2388 52526 2628
rect 52446 2378 52463 2388
rect 52167 2327 52305 2338
rect 52509 2378 52526 2388
rect 52463 2327 52509 2338
rect 52121 2244 52167 2255
rect 52336 2246 52347 2292
rect 52421 2246 52432 2292
rect 50968 2171 51064 2219
rect 48111 2000 48157 2011
rect 48488 2141 50456 2171
rect 48488 2001 49756 2141
rect 50356 2001 50456 2141
rect 48488 1971 50456 2001
rect 50968 2115 50988 2171
rect 51044 2115 51064 2171
rect 47778 1849 47942 1861
rect 47778 1793 47790 1849
rect 47846 1793 47942 1849
rect 47778 1781 47942 1793
rect 43417 1250 43429 1306
rect 43485 1250 43612 1306
rect 43668 1250 45562 1306
rect 47631 1631 47677 1642
rect 47846 1640 47942 1781
rect 48525 1831 48571 1842
rect 47846 1594 47857 1640
rect 47931 1594 47942 1640
rect 48111 1631 48157 1642
rect 47677 1548 47815 1559
rect 47677 1374 47769 1548
rect 47973 1548 48019 1559
rect 47956 1489 47973 1499
rect 48019 1489 48036 1499
rect 47956 1433 47968 1489
rect 48024 1433 48036 1489
rect 47956 1423 47973 1433
rect 47677 1363 47815 1374
rect 48019 1423 48036 1433
rect 47973 1363 48019 1374
rect 43417 1238 43503 1250
rect 43610 1238 43670 1250
rect 40088 851 40252 863
rect 40568 929 40732 941
rect 40568 873 40580 929
rect 40636 873 40732 929
rect 40568 861 40732 873
rect 40088 795 40100 851
rect 40156 795 40252 851
rect 40088 783 40252 795
rect 40156 733 40252 783
rect 33540 231 38722 431
rect 39053 711 39099 722
rect 39268 720 39568 733
rect 39268 674 39279 720
rect 39353 687 39483 720
rect 39353 674 39364 687
rect 39472 674 39483 687
rect 39557 674 39568 720
rect 39737 711 39783 722
rect 39099 628 39237 639
rect 39099 454 39191 628
rect 39395 628 39441 639
rect 39378 569 39395 579
rect 39599 628 39737 639
rect 39441 569 39458 579
rect 39378 513 39390 569
rect 39446 513 39458 569
rect 39378 503 39395 513
rect 39099 443 39237 454
rect 39441 503 39458 513
rect 39395 443 39441 454
rect 39645 454 39737 628
rect 39599 443 39737 454
rect 39053 231 39099 371
rect 39268 362 39279 408
rect 39353 362 39364 408
rect 39268 331 39364 362
rect 39472 362 39483 408
rect 39557 362 39568 408
rect 39472 331 39568 362
rect 39952 720 40252 733
rect 39952 674 39963 720
rect 40037 687 40167 720
rect 40037 674 40048 687
rect 40156 674 40167 687
rect 40241 674 40252 720
rect 40421 711 40467 722
rect 39875 628 39921 639
rect 39858 569 39875 579
rect 40079 628 40125 639
rect 39921 569 39938 579
rect 39858 513 39870 569
rect 39926 513 39938 569
rect 39858 503 39875 513
rect 39921 503 39938 513
rect 40062 569 40079 579
rect 40283 628 40329 639
rect 40125 569 40142 579
rect 40062 513 40074 569
rect 40130 513 40142 569
rect 40062 503 40079 513
rect 39875 443 39921 454
rect 40125 503 40142 513
rect 40266 569 40283 579
rect 40329 569 40346 579
rect 40266 513 40278 569
rect 40334 513 40346 569
rect 40266 503 40283 513
rect 40079 443 40125 454
rect 40329 503 40346 513
rect 40283 443 40329 454
rect 39737 231 39783 371
rect 39952 362 39963 408
rect 40037 362 40048 408
rect 39952 331 40048 362
rect 40156 362 40167 408
rect 40241 362 40252 408
rect 40156 331 40252 362
rect 40636 720 40732 861
rect 41244 1031 43212 1215
rect 47631 1151 47677 1291
rect 47846 1282 47857 1328
rect 47931 1282 47942 1328
rect 47846 1251 47942 1282
rect 48111 1151 48157 1291
rect 40636 674 40647 720
rect 40721 674 40732 720
rect 40901 711 40947 722
rect 40467 628 40605 639
rect 40467 454 40559 628
rect 40763 628 40809 639
rect 40746 569 40763 579
rect 40809 569 40826 579
rect 40746 513 40758 569
rect 40814 513 40826 569
rect 40746 503 40763 513
rect 40467 443 40605 454
rect 40809 503 40826 513
rect 40763 443 40809 454
rect 40421 231 40467 371
rect 40636 362 40647 408
rect 40721 362 40732 408
rect 40636 331 40732 362
rect 40901 231 40947 371
rect 41244 231 42712 1031
rect 43012 431 43212 1031
rect 47594 431 48194 1151
rect 48740 1840 48836 1871
rect 48740 1794 48751 1840
rect 48825 1794 48836 1840
rect 49005 1831 49459 1971
rect 48663 1748 48709 1759
rect 48646 1464 48663 1474
rect 48867 1748 49005 1759
rect 48709 1464 48726 1474
rect 48646 1224 48658 1464
rect 48714 1224 48726 1464
rect 48646 1214 48663 1224
rect 48709 1214 48726 1224
rect 48663 1163 48709 1174
rect 48913 1174 49005 1748
rect 48867 1163 49005 1174
rect 48525 1080 48571 1091
rect 48740 1082 48751 1128
rect 48825 1082 48836 1128
rect 48740 1007 48836 1082
rect 49051 1163 49413 1831
rect 49005 1080 49051 1091
rect 49628 1840 49724 1871
rect 49628 1794 49639 1840
rect 49713 1794 49724 1840
rect 49893 1831 49939 1971
rect 49459 1748 49597 1759
rect 49459 1174 49551 1748
rect 49755 1748 49801 1759
rect 49738 1464 49755 1474
rect 49801 1464 49818 1474
rect 49738 1224 49750 1464
rect 49806 1224 49818 1464
rect 49738 1214 49755 1224
rect 49459 1163 49597 1174
rect 49801 1214 49818 1224
rect 49755 1163 49801 1174
rect 49413 1080 49459 1091
rect 49628 1082 49639 1128
rect 49713 1082 49724 1128
rect 48740 951 48760 1007
rect 48816 951 48836 1007
rect 48740 733 48836 951
rect 49628 863 49724 1082
rect 50108 1840 50204 1871
rect 50108 1794 50119 1840
rect 50193 1794 50204 1840
rect 50373 1831 50419 1971
rect 49939 1748 50077 1759
rect 49939 1174 50031 1748
rect 50235 1748 50281 1759
rect 50218 1464 50235 1474
rect 50281 1464 50298 1474
rect 50218 1224 50230 1464
rect 50286 1224 50298 1464
rect 50218 1214 50235 1224
rect 49939 1163 50077 1174
rect 50281 1214 50298 1224
rect 50235 1163 50281 1174
rect 49893 1080 49939 1091
rect 50108 1082 50119 1128
rect 50193 1082 50204 1128
rect 50108 941 50204 1082
rect 50753 1875 50799 1886
rect 50968 1884 51064 2115
rect 51652 2015 51748 2219
rect 52336 2105 52432 2246
rect 53492 2325 53548 3346
rect 54660 3338 54730 3346
rect 54156 3294 54242 3298
rect 54156 3238 54168 3294
rect 54224 3238 54242 3294
rect 54156 3226 54242 3238
rect 53667 3081 53713 3092
rect 53882 3090 53958 3123
rect 53882 3044 53893 3090
rect 53947 3044 53958 3090
rect 54066 3090 54142 3123
rect 54066 3044 54077 3090
rect 54131 3044 54142 3090
rect 54250 3090 54326 3123
rect 54250 3044 54261 3090
rect 54315 3044 54326 3090
rect 54495 3081 54541 3092
rect 53805 2998 53851 3009
rect 53788 2971 53805 2973
rect 53989 2998 54035 3009
rect 53851 2971 53868 2973
rect 53713 2851 53800 2971
rect 53856 2851 53868 2971
rect 53788 2849 53805 2851
rect 53713 2551 53805 2671
rect 53851 2849 53868 2851
rect 53972 2671 53989 2673
rect 54173 2998 54219 3009
rect 54156 2971 54173 2973
rect 54357 2998 54403 3009
rect 54219 2971 54236 2973
rect 54156 2851 54168 2971
rect 54224 2851 54236 2971
rect 54156 2849 54173 2851
rect 54035 2671 54052 2673
rect 53972 2551 53984 2671
rect 54040 2551 54052 2671
rect 53972 2549 53989 2551
rect 53805 2513 53851 2524
rect 54035 2549 54052 2551
rect 53989 2513 54035 2524
rect 54219 2849 54236 2851
rect 54340 2671 54357 2673
rect 54478 2971 54495 2973
rect 54541 2971 54558 2973
rect 54478 2850 54490 2971
rect 54546 2850 54558 2971
rect 54478 2848 54495 2850
rect 54403 2671 54420 2673
rect 54340 2551 54352 2671
rect 54408 2551 54420 2671
rect 54340 2549 54357 2551
rect 54173 2513 54219 2524
rect 54403 2549 54420 2551
rect 54357 2513 54403 2524
rect 53882 2475 53893 2478
rect 53947 2475 53958 2478
rect 54066 2475 54077 2478
rect 54131 2475 54142 2478
rect 54250 2475 54261 2478
rect 54315 2475 54326 2478
rect 53667 2430 53713 2441
rect 53880 2419 53892 2475
rect 53948 2419 53960 2475
rect 53880 2405 53960 2419
rect 54064 2419 54076 2475
rect 54132 2419 54144 2475
rect 54064 2405 54144 2419
rect 54248 2419 54260 2475
rect 54316 2419 54328 2475
rect 54541 2848 54558 2850
rect 54495 2430 54541 2441
rect 54248 2405 54328 2419
rect 53880 2325 53960 2327
rect 53492 2269 53892 2325
rect 53948 2269 53960 2325
rect 53880 2267 53960 2269
rect 52601 2244 52647 2255
rect 53072 2209 53142 2223
rect 54064 2209 54144 2211
rect 53072 2153 53084 2209
rect 53140 2153 54076 2209
rect 54132 2153 54144 2209
rect 53072 2141 53142 2153
rect 54064 2151 54144 2153
rect 54393 2209 54473 2211
rect 54836 2209 54896 2221
rect 54393 2153 54405 2209
rect 54461 2153 54838 2209
rect 54894 2153 54896 2209
rect 54393 2151 54473 2153
rect 54836 2141 54896 2153
rect 52268 2093 52432 2105
rect 52268 2037 52280 2093
rect 52336 2037 52432 2093
rect 52268 2025 52432 2037
rect 52838 2093 52916 2104
rect 54248 2093 54328 2095
rect 52838 2092 54260 2093
rect 52838 2038 52850 2092
rect 52904 2038 54260 2092
rect 52838 2037 54260 2038
rect 54316 2037 54328 2093
rect 52838 2026 52916 2037
rect 54248 2035 54328 2037
rect 51652 1959 51672 2015
rect 51728 1959 51748 2015
rect 50968 1838 50979 1884
rect 51053 1838 51064 1884
rect 51233 1875 51483 1886
rect 50891 1792 50937 1803
rect 50874 1733 50891 1743
rect 51095 1792 51233 1803
rect 50937 1733 50954 1743
rect 50874 1677 50886 1733
rect 50942 1677 50954 1733
rect 50874 1667 50891 1677
rect 50937 1667 50954 1677
rect 50891 1607 50937 1618
rect 51141 1618 51233 1792
rect 51095 1607 51233 1618
rect 50753 1395 50799 1535
rect 50968 1526 50979 1572
rect 51053 1526 51064 1572
rect 50968 1495 51064 1526
rect 51279 1535 51437 1875
rect 51652 1884 51748 1959
rect 51652 1838 51663 1884
rect 51737 1838 51748 1884
rect 51917 1875 51963 1886
rect 51483 1792 51621 1803
rect 51483 1618 51575 1792
rect 51779 1792 51825 1803
rect 51762 1733 51779 1743
rect 51825 1733 51842 1743
rect 51762 1677 51774 1733
rect 51830 1677 51842 1733
rect 51762 1667 51779 1677
rect 51483 1607 51621 1618
rect 51825 1667 51842 1677
rect 51779 1607 51825 1618
rect 51233 1524 51483 1535
rect 51652 1526 51663 1572
rect 51737 1526 51748 1572
rect 51279 1395 51437 1524
rect 51652 1495 51748 1526
rect 51917 1395 51963 1535
rect 52121 1875 52167 1886
rect 52336 1884 52432 2025
rect 53880 1943 53960 1957
rect 53667 1921 53713 1932
rect 52336 1838 52347 1884
rect 52421 1838 52432 1884
rect 52601 1875 52647 1886
rect 52167 1792 52305 1803
rect 52167 1618 52259 1792
rect 52463 1792 52509 1803
rect 52446 1733 52463 1743
rect 52509 1733 52526 1743
rect 52446 1677 52458 1733
rect 52514 1677 52526 1733
rect 52446 1667 52463 1677
rect 52167 1607 52305 1618
rect 52509 1667 52526 1677
rect 52463 1607 52509 1618
rect 52121 1395 52167 1535
rect 52336 1526 52347 1572
rect 52421 1526 52432 1572
rect 52336 1495 52432 1526
rect 52601 1395 52647 1535
rect 53880 1887 53892 1943
rect 53948 1887 53960 1943
rect 54064 1943 54144 1957
rect 54064 1887 54076 1943
rect 54132 1887 54144 1943
rect 54248 1943 54328 1957
rect 54248 1887 54260 1943
rect 54316 1887 54328 1943
rect 54495 1921 54541 1932
rect 53882 1884 53893 1887
rect 53947 1884 53958 1887
rect 54066 1884 54077 1887
rect 54131 1884 54142 1887
rect 54250 1884 54261 1887
rect 54315 1884 54326 1887
rect 53805 1838 53851 1849
rect 53713 1664 53805 1838
rect 53805 1653 53851 1664
rect 53989 1838 54035 1849
rect 53989 1653 54035 1664
rect 54173 1838 54219 1849
rect 54357 1838 54403 1849
rect 54340 1811 54357 1813
rect 54403 1811 54420 1813
rect 54340 1691 54352 1811
rect 54408 1691 54420 1811
rect 54340 1689 54357 1691
rect 54173 1653 54219 1664
rect 54403 1689 54420 1691
rect 54357 1653 54403 1664
rect 53667 1436 53713 1581
rect 53882 1572 53893 1618
rect 53947 1572 53958 1618
rect 53882 1539 53958 1572
rect 54066 1572 54077 1618
rect 54131 1572 54142 1618
rect 54066 1539 54142 1572
rect 54250 1572 54261 1618
rect 54315 1572 54326 1618
rect 54250 1539 54326 1572
rect 54495 1436 54541 1581
rect 53655 1424 53735 1436
rect 50373 1080 50419 1091
rect 50716 1355 52684 1395
rect 53655 1368 53667 1424
rect 53723 1368 53735 1424
rect 53655 1356 53735 1368
rect 54473 1424 54553 1436
rect 54473 1368 54485 1424
rect 54541 1368 54553 1424
rect 54473 1356 54553 1368
rect 50716 1215 50816 1355
rect 52584 1215 52684 1355
rect 52889 1306 52975 1318
rect 53082 1306 53142 1310
rect 54978 1306 55034 4243
rect 55734 4241 55814 4243
rect 55366 4149 55446 4163
rect 55153 4127 55199 4138
rect 55366 4093 55378 4149
rect 55434 4093 55446 4149
rect 55550 4149 55630 4163
rect 55550 4093 55562 4149
rect 55618 4093 55630 4149
rect 55734 4149 55814 4163
rect 55734 4093 55746 4149
rect 55802 4093 55814 4149
rect 55981 4127 56027 4138
rect 55368 4090 55379 4093
rect 55433 4090 55444 4093
rect 55552 4090 55563 4093
rect 55617 4090 55628 4093
rect 55736 4090 55747 4093
rect 55801 4090 55812 4093
rect 55291 4044 55337 4055
rect 55199 3870 55291 4044
rect 55291 3859 55337 3870
rect 55475 4044 55521 4055
rect 55475 3859 55521 3870
rect 55659 4044 55705 4055
rect 55843 4044 55889 4055
rect 55826 4017 55843 4019
rect 55889 4017 55906 4019
rect 55826 3897 55838 4017
rect 55894 3897 55906 4017
rect 55826 3895 55843 3897
rect 55659 3859 55705 3870
rect 55889 3895 55906 3897
rect 55843 3859 55889 3870
rect 55153 3642 55199 3787
rect 55368 3778 55379 3824
rect 55433 3778 55444 3824
rect 55368 3745 55444 3778
rect 55552 3778 55563 3824
rect 55617 3778 55628 3824
rect 55552 3745 55628 3778
rect 55736 3778 55747 3824
rect 55801 3778 55812 3824
rect 55736 3745 55812 3778
rect 55981 3642 56027 3787
rect 55141 3630 55221 3642
rect 55141 3574 55153 3630
rect 55209 3574 55221 3630
rect 55141 3562 55221 3574
rect 55959 3630 56037 3642
rect 55959 3574 55971 3630
rect 56027 3574 56037 3630
rect 55959 3562 56037 3574
rect 52889 1250 52901 1306
rect 52957 1250 53084 1306
rect 53140 1250 55034 1306
rect 52889 1238 52975 1250
rect 53082 1238 53142 1250
rect 49560 851 49724 863
rect 50040 929 50204 941
rect 50040 873 50052 929
rect 50108 873 50204 929
rect 50040 861 50204 873
rect 49560 795 49572 851
rect 49628 795 49724 851
rect 49560 783 49724 795
rect 49628 733 49724 783
rect 43012 231 48194 431
rect 48525 711 48571 722
rect 48740 720 49040 733
rect 48740 674 48751 720
rect 48825 687 48955 720
rect 48825 674 48836 687
rect 48944 674 48955 687
rect 49029 674 49040 720
rect 49209 711 49255 722
rect 48571 628 48709 639
rect 48571 454 48663 628
rect 48867 628 48913 639
rect 48850 569 48867 579
rect 49071 628 49209 639
rect 48913 569 48930 579
rect 48850 513 48862 569
rect 48918 513 48930 569
rect 48850 503 48867 513
rect 48571 443 48709 454
rect 48913 503 48930 513
rect 48867 443 48913 454
rect 49117 454 49209 628
rect 49071 443 49209 454
rect 48525 231 48571 371
rect 48740 362 48751 408
rect 48825 362 48836 408
rect 48740 331 48836 362
rect 48944 362 48955 408
rect 49029 362 49040 408
rect 48944 331 49040 362
rect 49424 720 49724 733
rect 49424 674 49435 720
rect 49509 687 49639 720
rect 49509 674 49520 687
rect 49628 674 49639 687
rect 49713 674 49724 720
rect 49893 711 49939 722
rect 49347 628 49393 639
rect 49330 569 49347 579
rect 49551 628 49597 639
rect 49393 569 49410 579
rect 49330 513 49342 569
rect 49398 513 49410 569
rect 49330 503 49347 513
rect 49393 503 49410 513
rect 49534 569 49551 579
rect 49755 628 49801 639
rect 49597 569 49614 579
rect 49534 513 49546 569
rect 49602 513 49614 569
rect 49534 503 49551 513
rect 49347 443 49393 454
rect 49597 503 49614 513
rect 49738 569 49755 579
rect 49801 569 49818 579
rect 49738 513 49750 569
rect 49806 513 49818 569
rect 49738 503 49755 513
rect 49551 443 49597 454
rect 49801 503 49818 513
rect 49755 443 49801 454
rect 49209 231 49255 371
rect 49424 362 49435 408
rect 49509 362 49520 408
rect 49424 331 49520 362
rect 49628 362 49639 408
rect 49713 362 49724 408
rect 49628 331 49724 362
rect 50108 720 50204 861
rect 50716 1031 52684 1215
rect 50108 674 50119 720
rect 50193 674 50204 720
rect 50373 711 50419 722
rect 49939 628 50077 639
rect 49939 454 50031 628
rect 50235 628 50281 639
rect 50218 569 50235 579
rect 50281 569 50298 579
rect 50218 513 50230 569
rect 50286 513 50298 569
rect 50218 503 50235 513
rect 49939 443 50077 454
rect 50281 503 50298 513
rect 50235 443 50281 454
rect 49893 231 49939 371
rect 50108 362 50119 408
rect 50193 362 50204 408
rect 50108 331 50204 362
rect 50373 231 50419 371
rect 50716 231 52184 1031
rect 52484 231 52684 1031
rect 14596 230 52684 231
rect 230 31 52684 230
rect 230 30 19178 31
<< via1 >>
rect 6808 9852 6864 9908
rect 6440 9465 6445 9585
rect 6445 9465 6491 9585
rect 6491 9465 6496 9585
rect 6808 9465 6813 9585
rect 6813 9465 6859 9585
rect 6859 9465 6864 9585
rect 6624 9165 6629 9285
rect 6629 9165 6675 9285
rect 6675 9165 6680 9285
rect 7130 9464 7135 9585
rect 7135 9464 7181 9585
rect 7181 9464 7186 9585
rect 6992 9165 6997 9285
rect 6997 9165 7043 9285
rect 7043 9165 7048 9285
rect 6532 9046 6533 9089
rect 6533 9046 6587 9089
rect 6587 9046 6588 9089
rect 6532 9033 6588 9046
rect 6716 9046 6717 9089
rect 6717 9046 6771 9089
rect 6771 9046 6772 9089
rect 6716 9033 6772 9046
rect 6900 9046 6901 9089
rect 6901 9046 6955 9089
rect 6955 9046 6956 9089
rect 6900 9033 6956 9046
rect 5644 8883 5700 8939
rect 6532 8883 6588 8939
rect 5860 8767 5916 8823
rect 6716 8767 6772 8823
rect 7045 8767 7101 8823
rect 7302 8767 7358 8823
rect 6900 8651 6956 8707
rect 6532 8544 6588 8557
rect 6532 8501 6533 8544
rect 6533 8501 6587 8544
rect 6587 8501 6588 8544
rect 6716 8544 6772 8557
rect 6716 8501 6717 8544
rect 6717 8501 6771 8544
rect 6771 8501 6772 8544
rect 6900 8544 6956 8557
rect 6900 8501 6901 8544
rect 6901 8501 6955 8544
rect 6955 8501 6956 8544
rect 6992 8305 6997 8425
rect 6997 8305 7043 8425
rect 7043 8305 7048 8425
rect 6307 7982 6363 8038
rect 7125 7982 7181 8038
rect 7478 7864 7534 7920
rect 7302 7756 7358 7810
rect 6808 7647 6864 7703
rect 6440 7260 6445 7380
rect 6445 7260 6491 7380
rect 6491 7260 6496 7380
rect 6808 7260 6813 7380
rect 6813 7260 6859 7380
rect 6859 7260 6864 7380
rect 6624 6960 6629 7080
rect 6629 6960 6675 7080
rect 6675 6960 6680 7080
rect 7130 7259 7135 7380
rect 7135 7259 7181 7380
rect 7181 7259 7186 7380
rect 6992 6960 6997 7080
rect 6997 6960 7043 7080
rect 7043 6960 7048 7080
rect 6532 6841 6533 6884
rect 6533 6841 6587 6884
rect 6587 6841 6588 6884
rect 6532 6828 6588 6841
rect 6716 6841 6717 6884
rect 6717 6841 6771 6884
rect 6771 6841 6772 6884
rect 6716 6828 6772 6841
rect 6900 6841 6901 6884
rect 6901 6841 6955 6884
rect 6955 6841 6956 6884
rect 6900 6828 6956 6841
rect 6532 6678 6588 6734
rect 16280 9852 16336 9908
rect 15912 9465 15917 9585
rect 15917 9465 15963 9585
rect 15963 9465 15968 9585
rect 16280 9465 16285 9585
rect 16285 9465 16331 9585
rect 16331 9465 16336 9585
rect 16096 9165 16101 9285
rect 16101 9165 16147 9285
rect 16147 9165 16152 9285
rect 16602 9464 16607 9585
rect 16607 9464 16653 9585
rect 16653 9464 16658 9585
rect 16464 9165 16469 9285
rect 16469 9165 16515 9285
rect 16515 9165 16520 9285
rect 16004 9046 16005 9089
rect 16005 9046 16059 9089
rect 16059 9046 16060 9089
rect 16004 9033 16060 9046
rect 16188 9046 16189 9089
rect 16189 9046 16243 9089
rect 16243 9046 16244 9089
rect 16188 9033 16244 9046
rect 16372 9046 16373 9089
rect 16373 9046 16427 9089
rect 16427 9046 16428 9089
rect 16372 9033 16428 9046
rect 15116 8883 15172 8939
rect 16004 8883 16060 8939
rect 15332 8767 15388 8823
rect 16188 8767 16244 8823
rect 16517 8767 16573 8823
rect 16774 8767 16830 8823
rect 16372 8651 16428 8707
rect 16004 8544 16060 8557
rect 16004 8501 16005 8544
rect 16005 8501 16059 8544
rect 16059 8501 16060 8544
rect 16188 8544 16244 8557
rect 16188 8501 16189 8544
rect 16189 8501 16243 8544
rect 16243 8501 16244 8544
rect 16372 8544 16428 8557
rect 16372 8501 16373 8544
rect 16373 8501 16427 8544
rect 16427 8501 16428 8544
rect 16464 8305 16469 8425
rect 16469 8305 16515 8425
rect 16515 8305 16520 8425
rect 15779 7982 15835 8038
rect 16597 7982 16653 8038
rect 16950 7864 17006 7920
rect 16774 7756 16830 7810
rect 8294 7647 8350 7703
rect 7926 7260 7931 7380
rect 7931 7260 7977 7380
rect 7977 7260 7982 7380
rect 8294 7260 8299 7380
rect 8299 7260 8345 7380
rect 8345 7260 8350 7380
rect 8110 6960 8115 7080
rect 8115 6960 8161 7080
rect 8161 6960 8166 7080
rect 8616 7259 8621 7380
rect 8621 7259 8667 7380
rect 8667 7259 8672 7380
rect 8478 6960 8483 7080
rect 8483 6960 8529 7080
rect 8529 6960 8534 7080
rect 8018 6841 8019 6884
rect 8019 6841 8073 6884
rect 8073 6841 8074 6884
rect 8018 6828 8074 6841
rect 8202 6841 8203 6884
rect 8203 6841 8257 6884
rect 8257 6841 8258 6884
rect 8202 6828 8258 6841
rect 8386 6841 8387 6884
rect 8387 6841 8441 6884
rect 8441 6841 8442 6884
rect 8386 6828 8442 6841
rect 8018 6678 8074 6734
rect 16280 7647 16336 7703
rect 15912 7260 15917 7380
rect 15917 7260 15963 7380
rect 15963 7260 15968 7380
rect 16280 7260 16285 7380
rect 16285 7260 16331 7380
rect 16331 7260 16336 7380
rect 16096 6960 16101 7080
rect 16101 6960 16147 7080
rect 16147 6960 16152 7080
rect 16602 7259 16607 7380
rect 16607 7259 16653 7380
rect 16653 7259 16658 7380
rect 16464 6960 16469 7080
rect 16469 6960 16515 7080
rect 16515 6960 16520 7080
rect 16004 6841 16005 6884
rect 16005 6841 16059 6884
rect 16059 6841 16060 6884
rect 16004 6828 16060 6841
rect 16188 6841 16189 6884
rect 16189 6841 16243 6884
rect 16243 6841 16244 6884
rect 16188 6828 16244 6841
rect 16372 6841 16373 6884
rect 16373 6841 16427 6884
rect 16427 6841 16428 6884
rect 16372 6828 16428 6841
rect 16004 6678 16060 6734
rect 25752 9853 25808 9909
rect 25384 9466 25389 9586
rect 25389 9466 25435 9586
rect 25435 9466 25440 9586
rect 25752 9466 25757 9586
rect 25757 9466 25803 9586
rect 25803 9466 25808 9586
rect 25568 9166 25573 9286
rect 25573 9166 25619 9286
rect 25619 9166 25624 9286
rect 26074 9465 26079 9586
rect 26079 9465 26125 9586
rect 26125 9465 26130 9586
rect 25936 9166 25941 9286
rect 25941 9166 25987 9286
rect 25987 9166 25992 9286
rect 25476 9047 25477 9090
rect 25477 9047 25531 9090
rect 25531 9047 25532 9090
rect 25476 9034 25532 9047
rect 25660 9047 25661 9090
rect 25661 9047 25715 9090
rect 25715 9047 25716 9090
rect 25660 9034 25716 9047
rect 25844 9047 25845 9090
rect 25845 9047 25899 9090
rect 25899 9047 25900 9090
rect 25844 9034 25900 9047
rect 24588 8884 24644 8940
rect 25476 8884 25532 8940
rect 24804 8768 24860 8824
rect 25660 8768 25716 8824
rect 25989 8768 26045 8824
rect 26246 8768 26302 8824
rect 25844 8652 25900 8708
rect 25476 8545 25532 8558
rect 25476 8502 25477 8545
rect 25477 8502 25531 8545
rect 25531 8502 25532 8545
rect 25660 8545 25716 8558
rect 25660 8502 25661 8545
rect 25661 8502 25715 8545
rect 25715 8502 25716 8545
rect 25844 8545 25900 8558
rect 25844 8502 25845 8545
rect 25845 8502 25899 8545
rect 25899 8502 25900 8545
rect 25936 8306 25941 8426
rect 25941 8306 25987 8426
rect 25987 8306 25992 8426
rect 25251 7983 25307 8039
rect 26069 7983 26125 8039
rect 26422 7865 26478 7921
rect 26246 7757 26302 7811
rect 17766 7647 17822 7703
rect 17398 7260 17403 7380
rect 17403 7260 17449 7380
rect 17449 7260 17454 7380
rect 17766 7260 17771 7380
rect 17771 7260 17817 7380
rect 17817 7260 17822 7380
rect 17582 6960 17587 7080
rect 17587 6960 17633 7080
rect 17633 6960 17638 7080
rect 18088 7259 18093 7380
rect 18093 7259 18139 7380
rect 18139 7259 18144 7380
rect 17950 6960 17955 7080
rect 17955 6960 18001 7080
rect 18001 6960 18006 7080
rect 17490 6841 17491 6884
rect 17491 6841 17545 6884
rect 17545 6841 17546 6884
rect 17490 6828 17546 6841
rect 17674 6841 17675 6884
rect 17675 6841 17729 6884
rect 17729 6841 17730 6884
rect 17674 6828 17730 6841
rect 17858 6841 17859 6884
rect 17859 6841 17913 6884
rect 17913 6841 17914 6884
rect 17858 6828 17914 6841
rect 17490 6678 17546 6734
rect 25752 7648 25808 7704
rect 25384 7261 25389 7381
rect 25389 7261 25435 7381
rect 25435 7261 25440 7381
rect 25752 7261 25757 7381
rect 25757 7261 25803 7381
rect 25803 7261 25808 7381
rect 25568 6961 25573 7081
rect 25573 6961 25619 7081
rect 25619 6961 25624 7081
rect 26074 7260 26079 7381
rect 26079 7260 26125 7381
rect 26125 7260 26130 7381
rect 25936 6961 25941 7081
rect 25941 6961 25987 7081
rect 25987 6961 25992 7081
rect 25476 6842 25477 6885
rect 25477 6842 25531 6885
rect 25531 6842 25532 6885
rect 25476 6829 25532 6842
rect 25660 6842 25661 6885
rect 25661 6842 25715 6885
rect 25715 6842 25716 6885
rect 25660 6829 25716 6842
rect 25844 6842 25845 6885
rect 25845 6842 25899 6885
rect 25899 6842 25900 6885
rect 25844 6829 25900 6842
rect 25476 6679 25532 6735
rect 35224 9853 35280 9909
rect 34856 9466 34861 9586
rect 34861 9466 34907 9586
rect 34907 9466 34912 9586
rect 35224 9466 35229 9586
rect 35229 9466 35275 9586
rect 35275 9466 35280 9586
rect 35040 9166 35045 9286
rect 35045 9166 35091 9286
rect 35091 9166 35096 9286
rect 35546 9465 35551 9586
rect 35551 9465 35597 9586
rect 35597 9465 35602 9586
rect 35408 9166 35413 9286
rect 35413 9166 35459 9286
rect 35459 9166 35464 9286
rect 34948 9047 34949 9090
rect 34949 9047 35003 9090
rect 35003 9047 35004 9090
rect 34948 9034 35004 9047
rect 35132 9047 35133 9090
rect 35133 9047 35187 9090
rect 35187 9047 35188 9090
rect 35132 9034 35188 9047
rect 35316 9047 35317 9090
rect 35317 9047 35371 9090
rect 35371 9047 35372 9090
rect 35316 9034 35372 9047
rect 34060 8884 34116 8940
rect 34948 8884 35004 8940
rect 34276 8768 34332 8824
rect 35132 8768 35188 8824
rect 35461 8768 35517 8824
rect 35718 8768 35774 8824
rect 35316 8652 35372 8708
rect 34948 8545 35004 8558
rect 34948 8502 34949 8545
rect 34949 8502 35003 8545
rect 35003 8502 35004 8545
rect 35132 8545 35188 8558
rect 35132 8502 35133 8545
rect 35133 8502 35187 8545
rect 35187 8502 35188 8545
rect 35316 8545 35372 8558
rect 35316 8502 35317 8545
rect 35317 8502 35371 8545
rect 35371 8502 35372 8545
rect 35408 8306 35413 8426
rect 35413 8306 35459 8426
rect 35459 8306 35464 8426
rect 34723 7983 34779 8039
rect 35541 7983 35597 8039
rect 35894 7865 35950 7921
rect 35718 7757 35774 7811
rect 27238 7648 27294 7704
rect 26870 7261 26875 7381
rect 26875 7261 26921 7381
rect 26921 7261 26926 7381
rect 27238 7261 27243 7381
rect 27243 7261 27289 7381
rect 27289 7261 27294 7381
rect 27054 6961 27059 7081
rect 27059 6961 27105 7081
rect 27105 6961 27110 7081
rect 27560 7260 27565 7381
rect 27565 7260 27611 7381
rect 27611 7260 27616 7381
rect 27422 6961 27427 7081
rect 27427 6961 27473 7081
rect 27473 6961 27478 7081
rect 26962 6842 26963 6885
rect 26963 6842 27017 6885
rect 27017 6842 27018 6885
rect 26962 6829 27018 6842
rect 27146 6842 27147 6885
rect 27147 6842 27201 6885
rect 27201 6842 27202 6885
rect 27146 6829 27202 6842
rect 27330 6842 27331 6885
rect 27331 6842 27385 6885
rect 27385 6842 27386 6885
rect 27330 6829 27386 6842
rect 26962 6679 27018 6735
rect 35224 7648 35280 7704
rect 34856 7261 34861 7381
rect 34861 7261 34907 7381
rect 34907 7261 34912 7381
rect 35224 7261 35229 7381
rect 35229 7261 35275 7381
rect 35275 7261 35280 7381
rect 35040 6961 35045 7081
rect 35045 6961 35091 7081
rect 35091 6961 35096 7081
rect 35546 7260 35551 7381
rect 35551 7260 35597 7381
rect 35597 7260 35602 7381
rect 35408 6961 35413 7081
rect 35413 6961 35459 7081
rect 35459 6961 35464 7081
rect 34948 6842 34949 6885
rect 34949 6842 35003 6885
rect 35003 6842 35004 6885
rect 34948 6829 35004 6842
rect 35132 6842 35133 6885
rect 35133 6842 35187 6885
rect 35187 6842 35188 6885
rect 35132 6829 35188 6842
rect 35316 6842 35317 6885
rect 35317 6842 35371 6885
rect 35371 6842 35372 6885
rect 35316 6829 35372 6842
rect 34948 6679 35004 6735
rect 44696 9853 44752 9909
rect 44328 9466 44333 9586
rect 44333 9466 44379 9586
rect 44379 9466 44384 9586
rect 44696 9466 44701 9586
rect 44701 9466 44747 9586
rect 44747 9466 44752 9586
rect 44512 9166 44517 9286
rect 44517 9166 44563 9286
rect 44563 9166 44568 9286
rect 45018 9465 45023 9586
rect 45023 9465 45069 9586
rect 45069 9465 45074 9586
rect 44880 9166 44885 9286
rect 44885 9166 44931 9286
rect 44931 9166 44936 9286
rect 44420 9047 44421 9090
rect 44421 9047 44475 9090
rect 44475 9047 44476 9090
rect 44420 9034 44476 9047
rect 44604 9047 44605 9090
rect 44605 9047 44659 9090
rect 44659 9047 44660 9090
rect 44604 9034 44660 9047
rect 44788 9047 44789 9090
rect 44789 9047 44843 9090
rect 44843 9047 44844 9090
rect 44788 9034 44844 9047
rect 43532 8884 43588 8940
rect 44420 8884 44476 8940
rect 43748 8768 43804 8824
rect 44604 8768 44660 8824
rect 44933 8768 44989 8824
rect 45190 8768 45246 8824
rect 44788 8652 44844 8708
rect 44420 8545 44476 8558
rect 44420 8502 44421 8545
rect 44421 8502 44475 8545
rect 44475 8502 44476 8545
rect 44604 8545 44660 8558
rect 44604 8502 44605 8545
rect 44605 8502 44659 8545
rect 44659 8502 44660 8545
rect 44788 8545 44844 8558
rect 44788 8502 44789 8545
rect 44789 8502 44843 8545
rect 44843 8502 44844 8545
rect 44880 8306 44885 8426
rect 44885 8306 44931 8426
rect 44931 8306 44936 8426
rect 44195 7983 44251 8039
rect 45013 7983 45069 8039
rect 45366 7865 45422 7921
rect 45190 7757 45246 7811
rect 36710 7648 36766 7704
rect 36342 7261 36347 7381
rect 36347 7261 36393 7381
rect 36393 7261 36398 7381
rect 36710 7261 36715 7381
rect 36715 7261 36761 7381
rect 36761 7261 36766 7381
rect 36526 6961 36531 7081
rect 36531 6961 36577 7081
rect 36577 6961 36582 7081
rect 37032 7260 37037 7381
rect 37037 7260 37083 7381
rect 37083 7260 37088 7381
rect 36894 6961 36899 7081
rect 36899 6961 36945 7081
rect 36945 6961 36950 7081
rect 36434 6842 36435 6885
rect 36435 6842 36489 6885
rect 36489 6842 36490 6885
rect 36434 6829 36490 6842
rect 36618 6842 36619 6885
rect 36619 6842 36673 6885
rect 36673 6842 36674 6885
rect 36618 6829 36674 6842
rect 36802 6842 36803 6885
rect 36803 6842 36857 6885
rect 36857 6842 36858 6885
rect 36802 6829 36858 6842
rect 36434 6679 36490 6735
rect 44696 7648 44752 7704
rect 44328 7261 44333 7381
rect 44333 7261 44379 7381
rect 44379 7261 44384 7381
rect 44696 7261 44701 7381
rect 44701 7261 44747 7381
rect 44747 7261 44752 7381
rect 44512 6961 44517 7081
rect 44517 6961 44563 7081
rect 44563 6961 44568 7081
rect 45018 7260 45023 7381
rect 45023 7260 45069 7381
rect 45069 7260 45074 7381
rect 44880 6961 44885 7081
rect 44885 6961 44931 7081
rect 44931 6961 44936 7081
rect 44420 6842 44421 6885
rect 44421 6842 44475 6885
rect 44475 6842 44476 6885
rect 44420 6829 44476 6842
rect 44604 6842 44605 6885
rect 44605 6842 44659 6885
rect 44659 6842 44660 6885
rect 44604 6829 44660 6842
rect 44788 6842 44789 6885
rect 44789 6842 44843 6885
rect 44843 6842 44844 6885
rect 44788 6829 44844 6842
rect 44420 6679 44476 6735
rect 54168 9853 54224 9909
rect 53800 9466 53805 9586
rect 53805 9466 53851 9586
rect 53851 9466 53856 9586
rect 54168 9466 54173 9586
rect 54173 9466 54219 9586
rect 54219 9466 54224 9586
rect 53984 9166 53989 9286
rect 53989 9166 54035 9286
rect 54035 9166 54040 9286
rect 54490 9465 54495 9586
rect 54495 9465 54541 9586
rect 54541 9465 54546 9586
rect 54352 9166 54357 9286
rect 54357 9166 54403 9286
rect 54403 9166 54408 9286
rect 53892 9047 53893 9090
rect 53893 9047 53947 9090
rect 53947 9047 53948 9090
rect 53892 9034 53948 9047
rect 54076 9047 54077 9090
rect 54077 9047 54131 9090
rect 54131 9047 54132 9090
rect 54076 9034 54132 9047
rect 54260 9047 54261 9090
rect 54261 9047 54315 9090
rect 54315 9047 54316 9090
rect 54260 9034 54316 9047
rect 53004 8884 53060 8940
rect 53892 8884 53948 8940
rect 53220 8768 53276 8824
rect 54076 8768 54132 8824
rect 54405 8768 54461 8824
rect 54662 8768 54718 8824
rect 54260 8652 54316 8708
rect 53892 8545 53948 8558
rect 53892 8502 53893 8545
rect 53893 8502 53947 8545
rect 53947 8502 53948 8545
rect 54076 8545 54132 8558
rect 54076 8502 54077 8545
rect 54077 8502 54131 8545
rect 54131 8502 54132 8545
rect 54260 8545 54316 8558
rect 54260 8502 54261 8545
rect 54261 8502 54315 8545
rect 54315 8502 54316 8545
rect 54352 8306 54357 8426
rect 54357 8306 54403 8426
rect 54403 8306 54408 8426
rect 53667 7983 53723 8039
rect 54485 7983 54541 8039
rect 54838 7865 54894 7921
rect 54662 7757 54718 7811
rect 46182 7648 46238 7704
rect 45814 7261 45819 7381
rect 45819 7261 45865 7381
rect 45865 7261 45870 7381
rect 46182 7261 46187 7381
rect 46187 7261 46233 7381
rect 46233 7261 46238 7381
rect 45998 6961 46003 7081
rect 46003 6961 46049 7081
rect 46049 6961 46054 7081
rect 46504 7260 46509 7381
rect 46509 7260 46555 7381
rect 46555 7260 46560 7381
rect 46366 6961 46371 7081
rect 46371 6961 46417 7081
rect 46417 6961 46422 7081
rect 45906 6842 45907 6885
rect 45907 6842 45961 6885
rect 45961 6842 45962 6885
rect 45906 6829 45962 6842
rect 46090 6842 46091 6885
rect 46091 6842 46145 6885
rect 46145 6842 46146 6885
rect 46090 6829 46146 6842
rect 46274 6842 46275 6885
rect 46275 6842 46329 6885
rect 46329 6842 46330 6885
rect 46274 6829 46330 6842
rect 45906 6679 45962 6735
rect 54168 7648 54224 7704
rect 53800 7261 53805 7381
rect 53805 7261 53851 7381
rect 53851 7261 53856 7381
rect 54168 7261 54173 7381
rect 54173 7261 54219 7381
rect 54219 7261 54224 7381
rect 53984 6961 53989 7081
rect 53989 6961 54035 7081
rect 54035 6961 54040 7081
rect 54490 7260 54495 7381
rect 54495 7260 54541 7381
rect 54541 7260 54546 7381
rect 54352 6961 54357 7081
rect 54357 6961 54403 7081
rect 54403 6961 54408 7081
rect 53892 6842 53893 6885
rect 53893 6842 53947 6885
rect 53947 6842 53948 6885
rect 53892 6829 53948 6842
rect 54076 6842 54077 6885
rect 54077 6842 54131 6885
rect 54131 6842 54132 6885
rect 54076 6829 54132 6842
rect 54260 6842 54261 6885
rect 54261 6842 54315 6885
rect 54315 6842 54316 6885
rect 54260 6829 54316 6842
rect 53892 6679 53948 6735
rect 55654 7648 55710 7704
rect 55286 7261 55291 7381
rect 55291 7261 55337 7381
rect 55337 7261 55342 7381
rect 55654 7261 55659 7381
rect 55659 7261 55705 7381
rect 55705 7261 55710 7381
rect 55470 6961 55475 7081
rect 55475 6961 55521 7081
rect 55521 6961 55526 7081
rect 55976 7260 55981 7381
rect 55981 7260 56027 7381
rect 56027 7260 56032 7381
rect 55838 6961 55843 7081
rect 55843 6961 55889 7081
rect 55889 6961 55894 7081
rect 55378 6842 55379 6885
rect 55379 6842 55433 6885
rect 55433 6842 55434 6885
rect 55378 6829 55434 6842
rect 55562 6842 55563 6885
rect 55563 6842 55617 6885
rect 55617 6842 55618 6885
rect 55562 6829 55618 6842
rect 55746 6842 55747 6885
rect 55747 6842 55801 6885
rect 55801 6842 55802 6885
rect 55746 6829 55802 6842
rect 55378 6679 55434 6735
rect 5724 6562 5780 6618
rect 6716 6562 6772 6618
rect 7045 6562 7101 6618
rect 7478 6562 7534 6618
rect 8202 6562 8258 6618
rect 8531 6562 8587 6618
rect 8788 6562 8844 6618
rect 15196 6562 15252 6618
rect 16188 6562 16244 6618
rect 16517 6562 16573 6618
rect 16950 6562 17006 6618
rect 17674 6562 17730 6618
rect 18003 6562 18059 6618
rect 18260 6562 18316 6618
rect 24668 6563 24724 6619
rect 25660 6563 25716 6619
rect 25989 6563 26045 6619
rect 26422 6563 26478 6619
rect 27146 6563 27202 6619
rect 27475 6563 27531 6619
rect 27732 6563 27788 6619
rect 34140 6563 34196 6619
rect 35132 6563 35188 6619
rect 35461 6563 35517 6619
rect 35894 6563 35950 6619
rect 36618 6563 36674 6619
rect 36947 6563 37003 6619
rect 37204 6563 37260 6619
rect 43612 6563 43668 6619
rect 44604 6563 44660 6619
rect 44933 6563 44989 6619
rect 45366 6563 45422 6619
rect 46090 6563 46146 6619
rect 46419 6563 46475 6619
rect 46676 6563 46732 6619
rect 53084 6563 53140 6619
rect 54076 6563 54132 6619
rect 54405 6563 54461 6619
rect 54838 6563 54894 6619
rect 55562 6563 55618 6619
rect 55891 6563 55947 6619
rect 56148 6563 56204 6619
rect 6900 6446 6956 6502
rect 8386 6446 8442 6502
rect 6532 6339 6588 6352
rect 6532 6296 6533 6339
rect 6533 6296 6587 6339
rect 6587 6296 6588 6339
rect 6716 6339 6772 6352
rect 6716 6296 6717 6339
rect 6717 6296 6771 6339
rect 6771 6296 6772 6339
rect 6900 6339 6956 6352
rect 6900 6296 6901 6339
rect 6901 6296 6955 6339
rect 6955 6296 6956 6339
rect 6992 6100 6997 6220
rect 6997 6100 7043 6220
rect 7043 6100 7048 6220
rect 6307 5777 6363 5833
rect 7125 5777 7181 5833
rect 5444 5660 5500 5716
rect 16372 6446 16428 6502
rect 8018 6339 8074 6352
rect 8018 6296 8019 6339
rect 8019 6296 8073 6339
rect 8073 6296 8074 6339
rect 8202 6339 8258 6352
rect 8202 6296 8203 6339
rect 8203 6296 8257 6339
rect 8257 6296 8258 6339
rect 8386 6339 8442 6352
rect 8386 6296 8387 6339
rect 8387 6296 8441 6339
rect 8441 6296 8442 6339
rect 8478 6100 8483 6220
rect 8483 6100 8529 6220
rect 8529 6100 8534 6220
rect 7793 5777 7849 5833
rect 8611 5777 8667 5833
rect 8964 5660 9020 5716
rect 17858 6446 17914 6502
rect 16004 6339 16060 6352
rect 16004 6296 16005 6339
rect 16005 6296 16059 6339
rect 16059 6296 16060 6339
rect 16188 6339 16244 6352
rect 16188 6296 16189 6339
rect 16189 6296 16243 6339
rect 16243 6296 16244 6339
rect 16372 6339 16428 6352
rect 16372 6296 16373 6339
rect 16373 6296 16427 6339
rect 16427 6296 16428 6339
rect 16464 6100 16469 6220
rect 16469 6100 16515 6220
rect 16515 6100 16520 6220
rect 15779 5777 15835 5833
rect 16597 5777 16653 5833
rect 14916 5660 14972 5716
rect 25844 6447 25900 6503
rect 17490 6339 17546 6352
rect 17490 6296 17491 6339
rect 17491 6296 17545 6339
rect 17545 6296 17546 6339
rect 17674 6339 17730 6352
rect 17674 6296 17675 6339
rect 17675 6296 17729 6339
rect 17729 6296 17730 6339
rect 17858 6339 17914 6352
rect 17858 6296 17859 6339
rect 17859 6296 17913 6339
rect 17913 6296 17914 6339
rect 17950 6100 17955 6220
rect 17955 6100 18001 6220
rect 18001 6100 18006 6220
rect 17265 5777 17321 5833
rect 18083 5777 18139 5833
rect 18436 5660 18492 5716
rect 7478 5549 7534 5605
rect 8788 5550 8844 5606
rect 6808 5442 6864 5498
rect 6440 5055 6445 5175
rect 6445 5055 6491 5175
rect 6491 5055 6496 5175
rect 6808 5055 6813 5175
rect 6813 5055 6859 5175
rect 6859 5055 6864 5175
rect 6624 4755 6629 4875
rect 6629 4755 6675 4875
rect 6675 4755 6680 4875
rect 7130 5054 7135 5175
rect 7135 5054 7181 5175
rect 7181 5054 7186 5175
rect 6992 4755 6997 4875
rect 6997 4755 7043 4875
rect 7043 4755 7048 4875
rect 6532 4636 6533 4679
rect 6533 4636 6587 4679
rect 6587 4636 6588 4679
rect 6532 4623 6588 4636
rect 6716 4636 6717 4679
rect 6717 4636 6771 4679
rect 6771 4636 6772 4679
rect 6716 4623 6772 4636
rect 6900 4636 6901 4679
rect 6901 4636 6955 4679
rect 6955 4636 6956 4679
rect 6900 4623 6956 4636
rect 6532 4473 6588 4529
rect 8294 5443 8350 5499
rect 7926 5056 7931 5176
rect 7931 5056 7977 5176
rect 7977 5056 7982 5176
rect 8294 5056 8299 5176
rect 8299 5056 8345 5176
rect 8345 5056 8350 5176
rect 8110 4756 8115 4876
rect 8115 4756 8161 4876
rect 8161 4756 8166 4876
rect 8616 5055 8621 5176
rect 8621 5055 8667 5176
rect 8667 5055 8672 5176
rect 8478 4756 8483 4876
rect 8483 4756 8529 4876
rect 8529 4756 8534 4876
rect 8018 4637 8019 4680
rect 8019 4637 8073 4680
rect 8073 4637 8074 4680
rect 8018 4624 8074 4637
rect 8202 4637 8203 4680
rect 8203 4637 8257 4680
rect 8257 4637 8258 4680
rect 8202 4624 8258 4637
rect 8386 4637 8387 4680
rect 8387 4637 8441 4680
rect 8441 4637 8442 4680
rect 8386 4624 8442 4637
rect 8018 4474 8074 4530
rect 6716 4357 6772 4413
rect 7045 4357 7101 4413
rect 7302 4357 7358 4413
rect 8202 4358 8258 4414
rect 8531 4358 8587 4414
rect 8964 4358 9020 4414
rect 1298 3563 1303 3803
rect 1303 3563 1349 3803
rect 1349 3563 1354 3803
rect 952 3290 1008 3346
rect 2390 3563 2395 3803
rect 2395 3563 2441 3803
rect 2441 3563 2446 3803
rect 1400 3290 1456 3346
rect 2870 3563 2875 3803
rect 2875 3563 2921 3803
rect 2921 3563 2926 3803
rect 4824 3510 5124 4310
rect 27330 6447 27386 6503
rect 25476 6340 25532 6353
rect 25476 6297 25477 6340
rect 25477 6297 25531 6340
rect 25531 6297 25532 6340
rect 25660 6340 25716 6353
rect 25660 6297 25661 6340
rect 25661 6297 25715 6340
rect 25715 6297 25716 6340
rect 25844 6340 25900 6353
rect 25844 6297 25845 6340
rect 25845 6297 25899 6340
rect 25899 6297 25900 6340
rect 25936 6101 25941 6221
rect 25941 6101 25987 6221
rect 25987 6101 25992 6221
rect 25251 5778 25307 5834
rect 26069 5778 26125 5834
rect 24388 5661 24444 5717
rect 35316 6447 35372 6503
rect 26962 6340 27018 6353
rect 26962 6297 26963 6340
rect 26963 6297 27017 6340
rect 27017 6297 27018 6340
rect 27146 6340 27202 6353
rect 27146 6297 27147 6340
rect 27147 6297 27201 6340
rect 27201 6297 27202 6340
rect 27330 6340 27386 6353
rect 27330 6297 27331 6340
rect 27331 6297 27385 6340
rect 27385 6297 27386 6340
rect 27422 6101 27427 6221
rect 27427 6101 27473 6221
rect 27473 6101 27478 6221
rect 26737 5778 26793 5834
rect 27555 5778 27611 5834
rect 27908 5661 27964 5717
rect 16950 5549 17006 5605
rect 18260 5550 18316 5606
rect 16280 5442 16336 5498
rect 15912 5055 15917 5175
rect 15917 5055 15963 5175
rect 15963 5055 15968 5175
rect 16280 5055 16285 5175
rect 16285 5055 16331 5175
rect 16331 5055 16336 5175
rect 16096 4755 16101 4875
rect 16101 4755 16147 4875
rect 16147 4755 16152 4875
rect 16602 5054 16607 5175
rect 16607 5054 16653 5175
rect 16653 5054 16658 5175
rect 16464 4755 16469 4875
rect 16469 4755 16515 4875
rect 16515 4755 16520 4875
rect 16004 4636 16005 4679
rect 16005 4636 16059 4679
rect 16059 4636 16060 4679
rect 16004 4623 16060 4636
rect 16188 4636 16189 4679
rect 16189 4636 16243 4679
rect 16243 4636 16244 4679
rect 16188 4623 16244 4636
rect 16372 4636 16373 4679
rect 16373 4636 16427 4679
rect 16427 4636 16428 4679
rect 16372 4623 16428 4636
rect 16004 4473 16060 4529
rect 17766 5443 17822 5499
rect 17398 5056 17403 5176
rect 17403 5056 17449 5176
rect 17449 5056 17454 5176
rect 17766 5056 17771 5176
rect 17771 5056 17817 5176
rect 17817 5056 17822 5176
rect 17582 4756 17587 4876
rect 17587 4756 17633 4876
rect 17633 4756 17638 4876
rect 18088 5055 18093 5176
rect 18093 5055 18139 5176
rect 18139 5055 18144 5176
rect 17950 4756 17955 4876
rect 17955 4756 18001 4876
rect 18001 4756 18006 4876
rect 17490 4637 17491 4680
rect 17491 4637 17545 4680
rect 17545 4637 17546 4680
rect 17490 4624 17546 4637
rect 17674 4637 17675 4680
rect 17675 4637 17729 4680
rect 17729 4637 17730 4680
rect 17674 4624 17730 4637
rect 17858 4637 17859 4680
rect 17859 4637 17913 4680
rect 17913 4637 17914 4680
rect 17858 4624 17914 4637
rect 17490 4474 17546 4530
rect 16188 4357 16244 4413
rect 16517 4357 16573 4413
rect 16774 4357 16830 4413
rect 17674 4358 17730 4414
rect 18003 4358 18059 4414
rect 18436 4358 18492 4414
rect 5860 4241 5916 4297
rect 6900 4241 6956 4297
rect 2692 3212 2748 3268
rect 2212 3134 2268 3190
rect 608 2143 613 2383
rect 613 2143 659 2383
rect 659 2143 664 2383
rect 1502 2852 1507 2908
rect 1507 2852 1553 2908
rect 1553 2852 1558 2908
rect 1982 2852 1987 2908
rect 1987 2852 2033 2908
rect 2033 2852 2038 2908
rect 2186 2852 2191 2908
rect 2191 2852 2237 2908
rect 2237 2852 2242 2908
rect 2390 2852 2395 2908
rect 2395 2852 2441 2908
rect 2441 2852 2446 2908
rect 8386 4242 8442 4298
rect 6532 4134 6588 4147
rect 6532 4091 6533 4134
rect 6533 4091 6587 4134
rect 6587 4091 6588 4134
rect 6716 4134 6772 4147
rect 6716 4091 6717 4134
rect 6717 4091 6771 4134
rect 6771 4091 6772 4134
rect 6900 4134 6956 4147
rect 6900 4091 6901 4134
rect 6901 4091 6955 4134
rect 6955 4091 6956 4134
rect 6992 3895 6997 4015
rect 6997 3895 7043 4015
rect 7043 3895 7048 4015
rect 6307 3572 6363 3628
rect 7125 3572 7181 3628
rect 7478 3454 7534 3510
rect 3456 3174 5224 3314
rect 7302 3346 7358 3400
rect 2870 2852 2875 2908
rect 2875 2852 2921 2908
rect 2921 2852 2926 2908
rect 1166 2431 1246 2507
rect 2396 2400 2996 2540
rect 3730 2671 3735 2911
rect 3735 2671 3781 2911
rect 3781 2671 3786 2911
rect 4414 2671 4419 2911
rect 4419 2671 4465 2911
rect 4465 2671 4470 2911
rect 4210 2337 4215 2577
rect 4215 2337 4261 2577
rect 4261 2337 4266 2577
rect 4618 2337 4623 2577
rect 4623 2337 4669 2577
rect 4669 2337 4674 2577
rect 5098 2387 5103 2627
rect 5103 2387 5149 2627
rect 5149 2387 5154 2627
rect 2396 2000 2996 2140
rect 3628 2114 3684 2170
rect 430 1792 486 1848
rect 608 1432 613 1488
rect 613 1432 659 1488
rect 659 1432 664 1488
rect 1298 1223 1303 1463
rect 1303 1223 1349 1463
rect 1349 1223 1354 1463
rect 2390 1223 2395 1463
rect 2395 1223 2441 1463
rect 2441 1223 2446 1463
rect 1400 950 1456 1006
rect 2870 1223 2875 1463
rect 2875 1223 2921 1463
rect 2921 1223 2926 1463
rect 6808 3237 6864 3293
rect 6440 2850 6445 2970
rect 6445 2850 6491 2970
rect 6491 2850 6496 2970
rect 6808 2850 6813 2970
rect 6813 2850 6859 2970
rect 6859 2850 6864 2970
rect 6624 2550 6629 2670
rect 6629 2550 6675 2670
rect 6675 2550 6680 2670
rect 7130 2849 7135 2970
rect 7135 2849 7181 2970
rect 7181 2849 7186 2970
rect 6992 2550 6997 2670
rect 6997 2550 7043 2670
rect 7043 2550 7048 2670
rect 6532 2431 6533 2474
rect 6533 2431 6587 2474
rect 6587 2431 6588 2474
rect 6532 2418 6588 2431
rect 6716 2431 6717 2474
rect 6717 2431 6771 2474
rect 6771 2431 6772 2474
rect 6716 2418 6772 2431
rect 6900 2431 6901 2474
rect 6901 2431 6955 2474
rect 6955 2431 6956 2474
rect 6900 2418 6956 2431
rect 6532 2268 6588 2324
rect 5724 2152 5780 2208
rect 6716 2152 6772 2208
rect 7045 2152 7101 2208
rect 7478 2152 7534 2208
rect 4920 2036 4976 2092
rect 5490 2037 5544 2091
rect 6900 2036 6956 2092
rect 4312 1958 4368 2014
rect 3526 1676 3531 1732
rect 3531 1676 3577 1732
rect 3577 1676 3582 1732
rect 4414 1676 4419 1732
rect 4419 1676 4465 1732
rect 4465 1676 4470 1732
rect 5098 1676 5103 1732
rect 5103 1676 5149 1732
rect 5149 1676 5154 1732
rect 6532 1929 6588 1942
rect 6532 1886 6533 1929
rect 6533 1886 6587 1929
rect 6587 1886 6588 1929
rect 6716 1929 6772 1942
rect 6716 1886 6717 1929
rect 6717 1886 6771 1929
rect 6771 1886 6772 1929
rect 6900 1929 6956 1942
rect 6900 1886 6901 1929
rect 6901 1886 6955 1929
rect 6955 1886 6956 1929
rect 6992 1690 6997 1810
rect 6997 1690 7043 1810
rect 7043 1690 7048 1810
rect 6307 1367 6363 1423
rect 7125 1367 7181 1423
rect 3456 1214 5224 1354
rect 8018 4135 8074 4148
rect 8018 4092 8019 4135
rect 8019 4092 8073 4135
rect 8073 4092 8074 4135
rect 8202 4135 8258 4148
rect 8202 4092 8203 4135
rect 8203 4092 8257 4135
rect 8257 4092 8258 4135
rect 8386 4135 8442 4148
rect 8386 4092 8387 4135
rect 8387 4092 8441 4135
rect 8441 4092 8442 4135
rect 8478 3896 8483 4016
rect 8483 3896 8529 4016
rect 8529 3896 8534 4016
rect 7793 3573 7849 3629
rect 8611 3573 8667 3629
rect 9906 3510 10106 4310
rect 10770 3563 10775 3803
rect 10775 3563 10821 3803
rect 10821 3563 10826 3803
rect 11862 3563 11867 3803
rect 11867 3563 11913 3803
rect 11913 3563 11918 3803
rect 10872 3290 10928 3346
rect 12342 3563 12347 3803
rect 12347 3563 12393 3803
rect 12393 3563 12398 3803
rect 14296 3510 14596 4310
rect 36802 6447 36858 6503
rect 34948 6340 35004 6353
rect 34948 6297 34949 6340
rect 34949 6297 35003 6340
rect 35003 6297 35004 6340
rect 35132 6340 35188 6353
rect 35132 6297 35133 6340
rect 35133 6297 35187 6340
rect 35187 6297 35188 6340
rect 35316 6340 35372 6353
rect 35316 6297 35317 6340
rect 35317 6297 35371 6340
rect 35371 6297 35372 6340
rect 35408 6101 35413 6221
rect 35413 6101 35459 6221
rect 35459 6101 35464 6221
rect 34723 5778 34779 5834
rect 35541 5778 35597 5834
rect 33860 5661 33916 5717
rect 44788 6447 44844 6503
rect 36434 6340 36490 6353
rect 36434 6297 36435 6340
rect 36435 6297 36489 6340
rect 36489 6297 36490 6340
rect 36618 6340 36674 6353
rect 36618 6297 36619 6340
rect 36619 6297 36673 6340
rect 36673 6297 36674 6340
rect 36802 6340 36858 6353
rect 36802 6297 36803 6340
rect 36803 6297 36857 6340
rect 36857 6297 36858 6340
rect 36894 6101 36899 6221
rect 36899 6101 36945 6221
rect 36945 6101 36950 6221
rect 36209 5778 36265 5834
rect 37027 5778 37083 5834
rect 37380 5661 37436 5717
rect 26422 5550 26478 5606
rect 27732 5551 27788 5607
rect 25752 5443 25808 5499
rect 25384 5056 25389 5176
rect 25389 5056 25435 5176
rect 25435 5056 25440 5176
rect 25752 5056 25757 5176
rect 25757 5056 25803 5176
rect 25803 5056 25808 5176
rect 25568 4756 25573 4876
rect 25573 4756 25619 4876
rect 25619 4756 25624 4876
rect 26074 5055 26079 5176
rect 26079 5055 26125 5176
rect 26125 5055 26130 5176
rect 25936 4756 25941 4876
rect 25941 4756 25987 4876
rect 25987 4756 25992 4876
rect 25476 4637 25477 4680
rect 25477 4637 25531 4680
rect 25531 4637 25532 4680
rect 25476 4624 25532 4637
rect 25660 4637 25661 4680
rect 25661 4637 25715 4680
rect 25715 4637 25716 4680
rect 25660 4624 25716 4637
rect 25844 4637 25845 4680
rect 25845 4637 25899 4680
rect 25899 4637 25900 4680
rect 25844 4624 25900 4637
rect 25476 4474 25532 4530
rect 27238 5444 27294 5500
rect 26870 5057 26875 5177
rect 26875 5057 26921 5177
rect 26921 5057 26926 5177
rect 27238 5057 27243 5177
rect 27243 5057 27289 5177
rect 27289 5057 27294 5177
rect 27054 4757 27059 4877
rect 27059 4757 27105 4877
rect 27105 4757 27110 4877
rect 27560 5056 27565 5177
rect 27565 5056 27611 5177
rect 27611 5056 27616 5177
rect 27422 4757 27427 4877
rect 27427 4757 27473 4877
rect 27473 4757 27478 4877
rect 26962 4638 26963 4681
rect 26963 4638 27017 4681
rect 27017 4638 27018 4681
rect 26962 4625 27018 4638
rect 27146 4638 27147 4681
rect 27147 4638 27201 4681
rect 27201 4638 27202 4681
rect 27146 4625 27202 4638
rect 27330 4638 27331 4681
rect 27331 4638 27385 4681
rect 27385 4638 27386 4681
rect 27330 4625 27386 4638
rect 26962 4475 27018 4531
rect 25660 4358 25716 4414
rect 25989 4358 26045 4414
rect 26246 4358 26302 4414
rect 27146 4359 27202 4415
rect 27475 4359 27531 4415
rect 27908 4359 27964 4415
rect 15332 4241 15388 4297
rect 16372 4241 16428 4297
rect 12164 3212 12220 3268
rect 11684 3134 11740 3190
rect 10080 2143 10085 2383
rect 10085 2143 10131 2383
rect 10131 2143 10136 2383
rect 10974 2852 10979 2908
rect 10979 2852 11025 2908
rect 11025 2852 11030 2908
rect 11454 2852 11459 2908
rect 11459 2852 11505 2908
rect 11505 2852 11510 2908
rect 11658 2852 11663 2908
rect 11663 2852 11709 2908
rect 11709 2852 11714 2908
rect 11862 2852 11867 2908
rect 11867 2852 11913 2908
rect 11913 2852 11918 2908
rect 17858 4242 17914 4298
rect 16004 4134 16060 4147
rect 16004 4091 16005 4134
rect 16005 4091 16059 4134
rect 16059 4091 16060 4134
rect 16188 4134 16244 4147
rect 16188 4091 16189 4134
rect 16189 4091 16243 4134
rect 16243 4091 16244 4134
rect 16372 4134 16428 4147
rect 16372 4091 16373 4134
rect 16373 4091 16427 4134
rect 16427 4091 16428 4134
rect 16464 3895 16469 4015
rect 16469 3895 16515 4015
rect 16515 3895 16520 4015
rect 15779 3572 15835 3628
rect 16597 3572 16653 3628
rect 16950 3454 17006 3510
rect 12928 3174 14696 3314
rect 16774 3346 16830 3400
rect 12342 2852 12347 2908
rect 12347 2852 12393 2908
rect 12393 2852 12398 2908
rect 11868 2400 12468 2540
rect 13202 2671 13207 2911
rect 13207 2671 13253 2911
rect 13253 2671 13258 2911
rect 13886 2671 13891 2911
rect 13891 2671 13937 2911
rect 13937 2671 13942 2911
rect 13682 2337 13687 2577
rect 13687 2337 13733 2577
rect 13733 2337 13738 2577
rect 14090 2337 14095 2577
rect 14095 2337 14141 2577
rect 14141 2337 14146 2577
rect 14570 2387 14575 2627
rect 14575 2387 14621 2627
rect 14621 2387 14626 2627
rect 11868 2000 12468 2140
rect 13100 2114 13156 2170
rect 9902 1792 9958 1848
rect 5541 1249 5597 1305
rect 5724 1249 5780 1305
rect 10080 1432 10085 1488
rect 10085 1432 10131 1488
rect 10131 1432 10136 1488
rect 2692 872 2748 928
rect 2212 794 2268 850
rect 1502 512 1507 568
rect 1507 512 1553 568
rect 1553 512 1558 568
rect 1982 512 1987 568
rect 1987 512 2033 568
rect 2033 512 2038 568
rect 2186 512 2191 568
rect 2191 512 2237 568
rect 2237 512 2242 568
rect 2390 512 2395 568
rect 2395 512 2441 568
rect 2441 512 2446 568
rect 2870 512 2875 568
rect 2875 512 2921 568
rect 2921 512 2926 568
rect 4824 230 5124 1030
rect 10770 1223 10775 1463
rect 10775 1223 10821 1463
rect 10821 1223 10826 1463
rect 11862 1223 11867 1463
rect 11867 1223 11913 1463
rect 11913 1223 11918 1463
rect 10872 950 10928 1006
rect 12342 1223 12347 1463
rect 12347 1223 12393 1463
rect 12393 1223 12398 1463
rect 16280 3237 16336 3293
rect 15912 2850 15917 2970
rect 15917 2850 15963 2970
rect 15963 2850 15968 2970
rect 16280 2850 16285 2970
rect 16285 2850 16331 2970
rect 16331 2850 16336 2970
rect 16096 2550 16101 2670
rect 16101 2550 16147 2670
rect 16147 2550 16152 2670
rect 16602 2849 16607 2970
rect 16607 2849 16653 2970
rect 16653 2849 16658 2970
rect 16464 2550 16469 2670
rect 16469 2550 16515 2670
rect 16515 2550 16520 2670
rect 16004 2431 16005 2474
rect 16005 2431 16059 2474
rect 16059 2431 16060 2474
rect 16004 2418 16060 2431
rect 16188 2431 16189 2474
rect 16189 2431 16243 2474
rect 16243 2431 16244 2474
rect 16188 2418 16244 2431
rect 16372 2431 16373 2474
rect 16373 2431 16427 2474
rect 16427 2431 16428 2474
rect 16372 2418 16428 2431
rect 16004 2268 16060 2324
rect 15196 2152 15252 2208
rect 16188 2152 16244 2208
rect 16517 2152 16573 2208
rect 16950 2152 17006 2208
rect 14392 2036 14448 2092
rect 14962 2037 15016 2091
rect 16372 2036 16428 2092
rect 13784 1958 13840 2014
rect 12998 1676 13003 1732
rect 13003 1676 13049 1732
rect 13049 1676 13054 1732
rect 13886 1676 13891 1732
rect 13891 1676 13937 1732
rect 13937 1676 13942 1732
rect 14570 1676 14575 1732
rect 14575 1676 14621 1732
rect 14621 1676 14626 1732
rect 16004 1929 16060 1942
rect 16004 1886 16005 1929
rect 16005 1886 16059 1929
rect 16059 1886 16060 1929
rect 16188 1929 16244 1942
rect 16188 1886 16189 1929
rect 16189 1886 16243 1929
rect 16243 1886 16244 1929
rect 16372 1929 16428 1942
rect 16372 1886 16373 1929
rect 16373 1886 16427 1929
rect 16427 1886 16428 1929
rect 16464 1690 16469 1810
rect 16469 1690 16515 1810
rect 16515 1690 16520 1810
rect 15779 1367 15835 1423
rect 16597 1367 16653 1423
rect 12928 1214 14696 1354
rect 17490 4135 17546 4148
rect 17490 4092 17491 4135
rect 17491 4092 17545 4135
rect 17545 4092 17546 4135
rect 17674 4135 17730 4148
rect 17674 4092 17675 4135
rect 17675 4092 17729 4135
rect 17729 4092 17730 4135
rect 17858 4135 17914 4148
rect 17858 4092 17859 4135
rect 17859 4092 17913 4135
rect 17913 4092 17914 4135
rect 17950 3896 17955 4016
rect 17955 3896 18001 4016
rect 18001 3896 18006 4016
rect 17265 3573 17321 3629
rect 18083 3573 18139 3629
rect 19378 3511 19578 4311
rect 20242 3564 20247 3804
rect 20247 3564 20293 3804
rect 20293 3564 20298 3804
rect 21334 3564 21339 3804
rect 21339 3564 21385 3804
rect 21385 3564 21390 3804
rect 20344 3291 20400 3347
rect 21814 3564 21819 3804
rect 21819 3564 21865 3804
rect 21865 3564 21870 3804
rect 23768 3511 24068 4311
rect 46274 6447 46330 6503
rect 44420 6340 44476 6353
rect 44420 6297 44421 6340
rect 44421 6297 44475 6340
rect 44475 6297 44476 6340
rect 44604 6340 44660 6353
rect 44604 6297 44605 6340
rect 44605 6297 44659 6340
rect 44659 6297 44660 6340
rect 44788 6340 44844 6353
rect 44788 6297 44789 6340
rect 44789 6297 44843 6340
rect 44843 6297 44844 6340
rect 44880 6101 44885 6221
rect 44885 6101 44931 6221
rect 44931 6101 44936 6221
rect 44195 5778 44251 5834
rect 45013 5778 45069 5834
rect 43332 5661 43388 5717
rect 54260 6447 54316 6503
rect 45906 6340 45962 6353
rect 45906 6297 45907 6340
rect 45907 6297 45961 6340
rect 45961 6297 45962 6340
rect 46090 6340 46146 6353
rect 46090 6297 46091 6340
rect 46091 6297 46145 6340
rect 46145 6297 46146 6340
rect 46274 6340 46330 6353
rect 46274 6297 46275 6340
rect 46275 6297 46329 6340
rect 46329 6297 46330 6340
rect 46366 6101 46371 6221
rect 46371 6101 46417 6221
rect 46417 6101 46422 6221
rect 45681 5778 45737 5834
rect 46499 5778 46555 5834
rect 46852 5661 46908 5717
rect 35894 5550 35950 5606
rect 37204 5551 37260 5607
rect 35224 5443 35280 5499
rect 34856 5056 34861 5176
rect 34861 5056 34907 5176
rect 34907 5056 34912 5176
rect 35224 5056 35229 5176
rect 35229 5056 35275 5176
rect 35275 5056 35280 5176
rect 35040 4756 35045 4876
rect 35045 4756 35091 4876
rect 35091 4756 35096 4876
rect 35546 5055 35551 5176
rect 35551 5055 35597 5176
rect 35597 5055 35602 5176
rect 35408 4756 35413 4876
rect 35413 4756 35459 4876
rect 35459 4756 35464 4876
rect 34948 4637 34949 4680
rect 34949 4637 35003 4680
rect 35003 4637 35004 4680
rect 34948 4624 35004 4637
rect 35132 4637 35133 4680
rect 35133 4637 35187 4680
rect 35187 4637 35188 4680
rect 35132 4624 35188 4637
rect 35316 4637 35317 4680
rect 35317 4637 35371 4680
rect 35371 4637 35372 4680
rect 35316 4624 35372 4637
rect 34948 4474 35004 4530
rect 36710 5444 36766 5500
rect 36342 5057 36347 5177
rect 36347 5057 36393 5177
rect 36393 5057 36398 5177
rect 36710 5057 36715 5177
rect 36715 5057 36761 5177
rect 36761 5057 36766 5177
rect 36526 4757 36531 4877
rect 36531 4757 36577 4877
rect 36577 4757 36582 4877
rect 37032 5056 37037 5177
rect 37037 5056 37083 5177
rect 37083 5056 37088 5177
rect 36894 4757 36899 4877
rect 36899 4757 36945 4877
rect 36945 4757 36950 4877
rect 36434 4638 36435 4681
rect 36435 4638 36489 4681
rect 36489 4638 36490 4681
rect 36434 4625 36490 4638
rect 36618 4638 36619 4681
rect 36619 4638 36673 4681
rect 36673 4638 36674 4681
rect 36618 4625 36674 4638
rect 36802 4638 36803 4681
rect 36803 4638 36857 4681
rect 36857 4638 36858 4681
rect 36802 4625 36858 4638
rect 36434 4475 36490 4531
rect 35132 4358 35188 4414
rect 35461 4358 35517 4414
rect 35718 4358 35774 4414
rect 36618 4359 36674 4415
rect 36947 4359 37003 4415
rect 37380 4359 37436 4415
rect 24804 4242 24860 4298
rect 25844 4242 25900 4298
rect 21636 3213 21692 3269
rect 21156 3135 21212 3191
rect 19552 2144 19557 2384
rect 19557 2144 19603 2384
rect 19603 2144 19608 2384
rect 20446 2853 20451 2909
rect 20451 2853 20497 2909
rect 20497 2853 20502 2909
rect 20926 2853 20931 2909
rect 20931 2853 20977 2909
rect 20977 2853 20982 2909
rect 21130 2853 21135 2909
rect 21135 2853 21181 2909
rect 21181 2853 21186 2909
rect 21334 2853 21339 2909
rect 21339 2853 21385 2909
rect 21385 2853 21390 2909
rect 27330 4243 27386 4299
rect 25476 4135 25532 4148
rect 25476 4092 25477 4135
rect 25477 4092 25531 4135
rect 25531 4092 25532 4135
rect 25660 4135 25716 4148
rect 25660 4092 25661 4135
rect 25661 4092 25715 4135
rect 25715 4092 25716 4135
rect 25844 4135 25900 4148
rect 25844 4092 25845 4135
rect 25845 4092 25899 4135
rect 25899 4092 25900 4135
rect 25936 3896 25941 4016
rect 25941 3896 25987 4016
rect 25987 3896 25992 4016
rect 25251 3573 25307 3629
rect 26069 3573 26125 3629
rect 26422 3455 26478 3511
rect 22400 3175 24168 3315
rect 26246 3347 26302 3401
rect 21814 2853 21819 2909
rect 21819 2853 21865 2909
rect 21865 2853 21870 2909
rect 21340 2401 21940 2541
rect 22674 2672 22679 2912
rect 22679 2672 22725 2912
rect 22725 2672 22730 2912
rect 23358 2672 23363 2912
rect 23363 2672 23409 2912
rect 23409 2672 23414 2912
rect 23154 2338 23159 2578
rect 23159 2338 23205 2578
rect 23205 2338 23210 2578
rect 23562 2338 23567 2578
rect 23567 2338 23613 2578
rect 23613 2338 23618 2578
rect 24042 2388 24047 2628
rect 24047 2388 24093 2628
rect 24093 2388 24098 2628
rect 21340 2001 21940 2141
rect 22572 2115 22628 2171
rect 19374 1793 19430 1849
rect 15013 1249 15069 1305
rect 15196 1249 15252 1305
rect 19552 1433 19557 1489
rect 19557 1433 19603 1489
rect 19603 1433 19608 1489
rect 12164 872 12220 928
rect 11684 794 11740 850
rect 10974 512 10979 568
rect 10979 512 11025 568
rect 11025 512 11030 568
rect 11454 512 11459 568
rect 11459 512 11505 568
rect 11505 512 11510 568
rect 11658 512 11663 568
rect 11663 512 11709 568
rect 11709 512 11714 568
rect 11862 512 11867 568
rect 11867 512 11913 568
rect 11913 512 11918 568
rect 12342 512 12347 568
rect 12347 512 12393 568
rect 12393 512 12398 568
rect 14296 230 14596 1030
rect 20242 1224 20247 1464
rect 20247 1224 20293 1464
rect 20293 1224 20298 1464
rect 21334 1224 21339 1464
rect 21339 1224 21385 1464
rect 21385 1224 21390 1464
rect 20344 951 20400 1007
rect 21814 1224 21819 1464
rect 21819 1224 21865 1464
rect 21865 1224 21870 1464
rect 25752 3238 25808 3294
rect 25384 2851 25389 2971
rect 25389 2851 25435 2971
rect 25435 2851 25440 2971
rect 25752 2851 25757 2971
rect 25757 2851 25803 2971
rect 25803 2851 25808 2971
rect 25568 2551 25573 2671
rect 25573 2551 25619 2671
rect 25619 2551 25624 2671
rect 26074 2850 26079 2971
rect 26079 2850 26125 2971
rect 26125 2850 26130 2971
rect 25936 2551 25941 2671
rect 25941 2551 25987 2671
rect 25987 2551 25992 2671
rect 25476 2432 25477 2475
rect 25477 2432 25531 2475
rect 25531 2432 25532 2475
rect 25476 2419 25532 2432
rect 25660 2432 25661 2475
rect 25661 2432 25715 2475
rect 25715 2432 25716 2475
rect 25660 2419 25716 2432
rect 25844 2432 25845 2475
rect 25845 2432 25899 2475
rect 25899 2432 25900 2475
rect 25844 2419 25900 2432
rect 25476 2269 25532 2325
rect 24668 2153 24724 2209
rect 25660 2153 25716 2209
rect 25989 2153 26045 2209
rect 26422 2153 26478 2209
rect 23864 2037 23920 2093
rect 24434 2038 24488 2092
rect 25844 2037 25900 2093
rect 23256 1959 23312 2015
rect 22470 1677 22475 1733
rect 22475 1677 22521 1733
rect 22521 1677 22526 1733
rect 23358 1677 23363 1733
rect 23363 1677 23409 1733
rect 23409 1677 23414 1733
rect 24042 1677 24047 1733
rect 24047 1677 24093 1733
rect 24093 1677 24098 1733
rect 25476 1930 25532 1943
rect 25476 1887 25477 1930
rect 25477 1887 25531 1930
rect 25531 1887 25532 1930
rect 25660 1930 25716 1943
rect 25660 1887 25661 1930
rect 25661 1887 25715 1930
rect 25715 1887 25716 1930
rect 25844 1930 25900 1943
rect 25844 1887 25845 1930
rect 25845 1887 25899 1930
rect 25899 1887 25900 1930
rect 25936 1691 25941 1811
rect 25941 1691 25987 1811
rect 25987 1691 25992 1811
rect 25251 1368 25307 1424
rect 26069 1368 26125 1424
rect 22400 1215 24168 1355
rect 26962 4136 27018 4149
rect 26962 4093 26963 4136
rect 26963 4093 27017 4136
rect 27017 4093 27018 4136
rect 27146 4136 27202 4149
rect 27146 4093 27147 4136
rect 27147 4093 27201 4136
rect 27201 4093 27202 4136
rect 27330 4136 27386 4149
rect 27330 4093 27331 4136
rect 27331 4093 27385 4136
rect 27385 4093 27386 4136
rect 27422 3897 27427 4017
rect 27427 3897 27473 4017
rect 27473 3897 27478 4017
rect 26737 3574 26793 3630
rect 27555 3574 27611 3630
rect 28850 3511 29050 4311
rect 29714 3564 29719 3804
rect 29719 3564 29765 3804
rect 29765 3564 29770 3804
rect 30806 3564 30811 3804
rect 30811 3564 30857 3804
rect 30857 3564 30862 3804
rect 29816 3291 29872 3347
rect 31286 3564 31291 3804
rect 31291 3564 31337 3804
rect 31337 3564 31342 3804
rect 33240 3511 33540 4311
rect 55746 6447 55802 6503
rect 53892 6340 53948 6353
rect 53892 6297 53893 6340
rect 53893 6297 53947 6340
rect 53947 6297 53948 6340
rect 54076 6340 54132 6353
rect 54076 6297 54077 6340
rect 54077 6297 54131 6340
rect 54131 6297 54132 6340
rect 54260 6340 54316 6353
rect 54260 6297 54261 6340
rect 54261 6297 54315 6340
rect 54315 6297 54316 6340
rect 54352 6101 54357 6221
rect 54357 6101 54403 6221
rect 54403 6101 54408 6221
rect 53667 5778 53723 5834
rect 54485 5778 54541 5834
rect 52804 5661 52860 5717
rect 55378 6340 55434 6353
rect 55378 6297 55379 6340
rect 55379 6297 55433 6340
rect 55433 6297 55434 6340
rect 55562 6340 55618 6353
rect 55562 6297 55563 6340
rect 55563 6297 55617 6340
rect 55617 6297 55618 6340
rect 55746 6340 55802 6353
rect 55746 6297 55747 6340
rect 55747 6297 55801 6340
rect 55801 6297 55802 6340
rect 55838 6101 55843 6221
rect 55843 6101 55889 6221
rect 55889 6101 55894 6221
rect 55153 5778 55209 5834
rect 55971 5778 56027 5834
rect 56324 5661 56380 5717
rect 45366 5550 45422 5606
rect 46676 5551 46732 5607
rect 44696 5443 44752 5499
rect 44328 5056 44333 5176
rect 44333 5056 44379 5176
rect 44379 5056 44384 5176
rect 44696 5056 44701 5176
rect 44701 5056 44747 5176
rect 44747 5056 44752 5176
rect 44512 4756 44517 4876
rect 44517 4756 44563 4876
rect 44563 4756 44568 4876
rect 45018 5055 45023 5176
rect 45023 5055 45069 5176
rect 45069 5055 45074 5176
rect 44880 4756 44885 4876
rect 44885 4756 44931 4876
rect 44931 4756 44936 4876
rect 44420 4637 44421 4680
rect 44421 4637 44475 4680
rect 44475 4637 44476 4680
rect 44420 4624 44476 4637
rect 44604 4637 44605 4680
rect 44605 4637 44659 4680
rect 44659 4637 44660 4680
rect 44604 4624 44660 4637
rect 44788 4637 44789 4680
rect 44789 4637 44843 4680
rect 44843 4637 44844 4680
rect 44788 4624 44844 4637
rect 44420 4474 44476 4530
rect 46182 5444 46238 5500
rect 45814 5057 45819 5177
rect 45819 5057 45865 5177
rect 45865 5057 45870 5177
rect 46182 5057 46187 5177
rect 46187 5057 46233 5177
rect 46233 5057 46238 5177
rect 45998 4757 46003 4877
rect 46003 4757 46049 4877
rect 46049 4757 46054 4877
rect 46504 5056 46509 5177
rect 46509 5056 46555 5177
rect 46555 5056 46560 5177
rect 46366 4757 46371 4877
rect 46371 4757 46417 4877
rect 46417 4757 46422 4877
rect 45906 4638 45907 4681
rect 45907 4638 45961 4681
rect 45961 4638 45962 4681
rect 45906 4625 45962 4638
rect 46090 4638 46091 4681
rect 46091 4638 46145 4681
rect 46145 4638 46146 4681
rect 46090 4625 46146 4638
rect 46274 4638 46275 4681
rect 46275 4638 46329 4681
rect 46329 4638 46330 4681
rect 46274 4625 46330 4638
rect 45906 4475 45962 4531
rect 44604 4358 44660 4414
rect 44933 4358 44989 4414
rect 45190 4358 45246 4414
rect 46090 4359 46146 4415
rect 46419 4359 46475 4415
rect 46852 4359 46908 4415
rect 34276 4242 34332 4298
rect 35316 4242 35372 4298
rect 31108 3213 31164 3269
rect 30628 3135 30684 3191
rect 29024 2144 29029 2384
rect 29029 2144 29075 2384
rect 29075 2144 29080 2384
rect 29918 2853 29923 2909
rect 29923 2853 29969 2909
rect 29969 2853 29974 2909
rect 30398 2853 30403 2909
rect 30403 2853 30449 2909
rect 30449 2853 30454 2909
rect 30602 2853 30607 2909
rect 30607 2853 30653 2909
rect 30653 2853 30658 2909
rect 30806 2853 30811 2909
rect 30811 2853 30857 2909
rect 30857 2853 30862 2909
rect 36802 4243 36858 4299
rect 34948 4135 35004 4148
rect 34948 4092 34949 4135
rect 34949 4092 35003 4135
rect 35003 4092 35004 4135
rect 35132 4135 35188 4148
rect 35132 4092 35133 4135
rect 35133 4092 35187 4135
rect 35187 4092 35188 4135
rect 35316 4135 35372 4148
rect 35316 4092 35317 4135
rect 35317 4092 35371 4135
rect 35371 4092 35372 4135
rect 35408 3896 35413 4016
rect 35413 3896 35459 4016
rect 35459 3896 35464 4016
rect 34723 3573 34779 3629
rect 35541 3573 35597 3629
rect 35894 3455 35950 3511
rect 31872 3175 33640 3315
rect 35718 3347 35774 3401
rect 31286 2853 31291 2909
rect 31291 2853 31337 2909
rect 31337 2853 31342 2909
rect 30812 2401 31412 2541
rect 32146 2672 32151 2912
rect 32151 2672 32197 2912
rect 32197 2672 32202 2912
rect 32830 2672 32835 2912
rect 32835 2672 32881 2912
rect 32881 2672 32886 2912
rect 32626 2338 32631 2578
rect 32631 2338 32677 2578
rect 32677 2338 32682 2578
rect 33034 2338 33039 2578
rect 33039 2338 33085 2578
rect 33085 2338 33090 2578
rect 33514 2388 33519 2628
rect 33519 2388 33565 2628
rect 33565 2388 33570 2628
rect 30812 2001 31412 2141
rect 32044 2115 32100 2171
rect 28846 1793 28902 1849
rect 24485 1250 24541 1306
rect 24668 1250 24724 1306
rect 29024 1433 29029 1489
rect 29029 1433 29075 1489
rect 29075 1433 29080 1489
rect 21636 873 21692 929
rect 21156 795 21212 851
rect 20446 513 20451 569
rect 20451 513 20497 569
rect 20497 513 20502 569
rect 20926 513 20931 569
rect 20931 513 20977 569
rect 20977 513 20982 569
rect 21130 513 21135 569
rect 21135 513 21181 569
rect 21181 513 21186 569
rect 21334 513 21339 569
rect 21339 513 21385 569
rect 21385 513 21390 569
rect 21814 513 21819 569
rect 21819 513 21865 569
rect 21865 513 21870 569
rect 23768 231 24068 1031
rect 29714 1224 29719 1464
rect 29719 1224 29765 1464
rect 29765 1224 29770 1464
rect 30806 1224 30811 1464
rect 30811 1224 30857 1464
rect 30857 1224 30862 1464
rect 29816 951 29872 1007
rect 31286 1224 31291 1464
rect 31291 1224 31337 1464
rect 31337 1224 31342 1464
rect 35224 3238 35280 3294
rect 34856 2851 34861 2971
rect 34861 2851 34907 2971
rect 34907 2851 34912 2971
rect 35224 2851 35229 2971
rect 35229 2851 35275 2971
rect 35275 2851 35280 2971
rect 35040 2551 35045 2671
rect 35045 2551 35091 2671
rect 35091 2551 35096 2671
rect 35546 2850 35551 2971
rect 35551 2850 35597 2971
rect 35597 2850 35602 2971
rect 35408 2551 35413 2671
rect 35413 2551 35459 2671
rect 35459 2551 35464 2671
rect 34948 2432 34949 2475
rect 34949 2432 35003 2475
rect 35003 2432 35004 2475
rect 34948 2419 35004 2432
rect 35132 2432 35133 2475
rect 35133 2432 35187 2475
rect 35187 2432 35188 2475
rect 35132 2419 35188 2432
rect 35316 2432 35317 2475
rect 35317 2432 35371 2475
rect 35371 2432 35372 2475
rect 35316 2419 35372 2432
rect 34948 2269 35004 2325
rect 34140 2153 34196 2209
rect 35132 2153 35188 2209
rect 35461 2153 35517 2209
rect 35894 2153 35950 2209
rect 33336 2037 33392 2093
rect 33906 2038 33960 2092
rect 35316 2037 35372 2093
rect 32728 1959 32784 2015
rect 31942 1677 31947 1733
rect 31947 1677 31993 1733
rect 31993 1677 31998 1733
rect 32830 1677 32835 1733
rect 32835 1677 32881 1733
rect 32881 1677 32886 1733
rect 33514 1677 33519 1733
rect 33519 1677 33565 1733
rect 33565 1677 33570 1733
rect 34948 1930 35004 1943
rect 34948 1887 34949 1930
rect 34949 1887 35003 1930
rect 35003 1887 35004 1930
rect 35132 1930 35188 1943
rect 35132 1887 35133 1930
rect 35133 1887 35187 1930
rect 35187 1887 35188 1930
rect 35316 1930 35372 1943
rect 35316 1887 35317 1930
rect 35317 1887 35371 1930
rect 35371 1887 35372 1930
rect 35408 1691 35413 1811
rect 35413 1691 35459 1811
rect 35459 1691 35464 1811
rect 34723 1368 34779 1424
rect 35541 1368 35597 1424
rect 31872 1215 33640 1355
rect 36434 4136 36490 4149
rect 36434 4093 36435 4136
rect 36435 4093 36489 4136
rect 36489 4093 36490 4136
rect 36618 4136 36674 4149
rect 36618 4093 36619 4136
rect 36619 4093 36673 4136
rect 36673 4093 36674 4136
rect 36802 4136 36858 4149
rect 36802 4093 36803 4136
rect 36803 4093 36857 4136
rect 36857 4093 36858 4136
rect 36894 3897 36899 4017
rect 36899 3897 36945 4017
rect 36945 3897 36950 4017
rect 36209 3574 36265 3630
rect 37027 3574 37083 3630
rect 38322 3511 38522 4311
rect 39186 3564 39191 3804
rect 39191 3564 39237 3804
rect 39237 3564 39242 3804
rect 40278 3564 40283 3804
rect 40283 3564 40329 3804
rect 40329 3564 40334 3804
rect 39288 3291 39344 3347
rect 40758 3564 40763 3804
rect 40763 3564 40809 3804
rect 40809 3564 40814 3804
rect 42712 3511 43012 4311
rect 54838 5550 54894 5606
rect 56148 5551 56204 5607
rect 54168 5443 54224 5499
rect 53800 5056 53805 5176
rect 53805 5056 53851 5176
rect 53851 5056 53856 5176
rect 54168 5056 54173 5176
rect 54173 5056 54219 5176
rect 54219 5056 54224 5176
rect 53984 4756 53989 4876
rect 53989 4756 54035 4876
rect 54035 4756 54040 4876
rect 54490 5055 54495 5176
rect 54495 5055 54541 5176
rect 54541 5055 54546 5176
rect 54352 4756 54357 4876
rect 54357 4756 54403 4876
rect 54403 4756 54408 4876
rect 53892 4637 53893 4680
rect 53893 4637 53947 4680
rect 53947 4637 53948 4680
rect 53892 4624 53948 4637
rect 54076 4637 54077 4680
rect 54077 4637 54131 4680
rect 54131 4637 54132 4680
rect 54076 4624 54132 4637
rect 54260 4637 54261 4680
rect 54261 4637 54315 4680
rect 54315 4637 54316 4680
rect 54260 4624 54316 4637
rect 53892 4474 53948 4530
rect 55654 5444 55710 5500
rect 55286 5057 55291 5177
rect 55291 5057 55337 5177
rect 55337 5057 55342 5177
rect 55654 5057 55659 5177
rect 55659 5057 55705 5177
rect 55705 5057 55710 5177
rect 55470 4757 55475 4877
rect 55475 4757 55521 4877
rect 55521 4757 55526 4877
rect 55976 5056 55981 5177
rect 55981 5056 56027 5177
rect 56027 5056 56032 5177
rect 55838 4757 55843 4877
rect 55843 4757 55889 4877
rect 55889 4757 55894 4877
rect 55378 4638 55379 4681
rect 55379 4638 55433 4681
rect 55433 4638 55434 4681
rect 55378 4625 55434 4638
rect 55562 4638 55563 4681
rect 55563 4638 55617 4681
rect 55617 4638 55618 4681
rect 55562 4625 55618 4638
rect 55746 4638 55747 4681
rect 55747 4638 55801 4681
rect 55801 4638 55802 4681
rect 55746 4625 55802 4638
rect 55378 4475 55434 4531
rect 54076 4358 54132 4414
rect 54405 4358 54461 4414
rect 54662 4358 54718 4414
rect 55562 4359 55618 4415
rect 55891 4359 55947 4415
rect 56324 4359 56380 4415
rect 43748 4242 43804 4298
rect 44788 4242 44844 4298
rect 40580 3213 40636 3269
rect 40100 3135 40156 3191
rect 38496 2144 38501 2384
rect 38501 2144 38547 2384
rect 38547 2144 38552 2384
rect 39390 2853 39395 2909
rect 39395 2853 39441 2909
rect 39441 2853 39446 2909
rect 39870 2853 39875 2909
rect 39875 2853 39921 2909
rect 39921 2853 39926 2909
rect 40074 2853 40079 2909
rect 40079 2853 40125 2909
rect 40125 2853 40130 2909
rect 40278 2853 40283 2909
rect 40283 2853 40329 2909
rect 40329 2853 40334 2909
rect 46274 4243 46330 4299
rect 44420 4135 44476 4148
rect 44420 4092 44421 4135
rect 44421 4092 44475 4135
rect 44475 4092 44476 4135
rect 44604 4135 44660 4148
rect 44604 4092 44605 4135
rect 44605 4092 44659 4135
rect 44659 4092 44660 4135
rect 44788 4135 44844 4148
rect 44788 4092 44789 4135
rect 44789 4092 44843 4135
rect 44843 4092 44844 4135
rect 44880 3896 44885 4016
rect 44885 3896 44931 4016
rect 44931 3896 44936 4016
rect 44195 3573 44251 3629
rect 45013 3573 45069 3629
rect 45366 3455 45422 3511
rect 41344 3175 43112 3315
rect 45190 3347 45246 3401
rect 40758 2853 40763 2909
rect 40763 2853 40809 2909
rect 40809 2853 40814 2909
rect 40284 2401 40884 2541
rect 41618 2672 41623 2912
rect 41623 2672 41669 2912
rect 41669 2672 41674 2912
rect 42302 2672 42307 2912
rect 42307 2672 42353 2912
rect 42353 2672 42358 2912
rect 42098 2338 42103 2578
rect 42103 2338 42149 2578
rect 42149 2338 42154 2578
rect 42506 2338 42511 2578
rect 42511 2338 42557 2578
rect 42557 2338 42562 2578
rect 42986 2388 42991 2628
rect 42991 2388 43037 2628
rect 43037 2388 43042 2628
rect 40284 2001 40884 2141
rect 41516 2115 41572 2171
rect 38318 1793 38374 1849
rect 33957 1250 34013 1306
rect 34140 1250 34196 1306
rect 38496 1433 38501 1489
rect 38501 1433 38547 1489
rect 38547 1433 38552 1489
rect 31108 873 31164 929
rect 30628 795 30684 851
rect 29918 513 29923 569
rect 29923 513 29969 569
rect 29969 513 29974 569
rect 30398 513 30403 569
rect 30403 513 30449 569
rect 30449 513 30454 569
rect 30602 513 30607 569
rect 30607 513 30653 569
rect 30653 513 30658 569
rect 30806 513 30811 569
rect 30811 513 30857 569
rect 30857 513 30862 569
rect 31286 513 31291 569
rect 31291 513 31337 569
rect 31337 513 31342 569
rect 33240 231 33540 1031
rect 39186 1224 39191 1464
rect 39191 1224 39237 1464
rect 39237 1224 39242 1464
rect 40278 1224 40283 1464
rect 40283 1224 40329 1464
rect 40329 1224 40334 1464
rect 39288 951 39344 1007
rect 40758 1224 40763 1464
rect 40763 1224 40809 1464
rect 40809 1224 40814 1464
rect 44696 3238 44752 3294
rect 44328 2851 44333 2971
rect 44333 2851 44379 2971
rect 44379 2851 44384 2971
rect 44696 2851 44701 2971
rect 44701 2851 44747 2971
rect 44747 2851 44752 2971
rect 44512 2551 44517 2671
rect 44517 2551 44563 2671
rect 44563 2551 44568 2671
rect 45018 2850 45023 2971
rect 45023 2850 45069 2971
rect 45069 2850 45074 2971
rect 44880 2551 44885 2671
rect 44885 2551 44931 2671
rect 44931 2551 44936 2671
rect 44420 2432 44421 2475
rect 44421 2432 44475 2475
rect 44475 2432 44476 2475
rect 44420 2419 44476 2432
rect 44604 2432 44605 2475
rect 44605 2432 44659 2475
rect 44659 2432 44660 2475
rect 44604 2419 44660 2432
rect 44788 2432 44789 2475
rect 44789 2432 44843 2475
rect 44843 2432 44844 2475
rect 44788 2419 44844 2432
rect 44420 2269 44476 2325
rect 43612 2153 43668 2209
rect 44604 2153 44660 2209
rect 44933 2153 44989 2209
rect 45366 2153 45422 2209
rect 42808 2037 42864 2093
rect 43378 2038 43432 2092
rect 44788 2037 44844 2093
rect 42200 1959 42256 2015
rect 41414 1677 41419 1733
rect 41419 1677 41465 1733
rect 41465 1677 41470 1733
rect 42302 1677 42307 1733
rect 42307 1677 42353 1733
rect 42353 1677 42358 1733
rect 42986 1677 42991 1733
rect 42991 1677 43037 1733
rect 43037 1677 43042 1733
rect 44420 1930 44476 1943
rect 44420 1887 44421 1930
rect 44421 1887 44475 1930
rect 44475 1887 44476 1930
rect 44604 1930 44660 1943
rect 44604 1887 44605 1930
rect 44605 1887 44659 1930
rect 44659 1887 44660 1930
rect 44788 1930 44844 1943
rect 44788 1887 44789 1930
rect 44789 1887 44843 1930
rect 44843 1887 44844 1930
rect 44880 1691 44885 1811
rect 44885 1691 44931 1811
rect 44931 1691 44936 1811
rect 44195 1368 44251 1424
rect 45013 1368 45069 1424
rect 41344 1215 43112 1355
rect 45906 4136 45962 4149
rect 45906 4093 45907 4136
rect 45907 4093 45961 4136
rect 45961 4093 45962 4136
rect 46090 4136 46146 4149
rect 46090 4093 46091 4136
rect 46091 4093 46145 4136
rect 46145 4093 46146 4136
rect 46274 4136 46330 4149
rect 46274 4093 46275 4136
rect 46275 4093 46329 4136
rect 46329 4093 46330 4136
rect 46366 3897 46371 4017
rect 46371 3897 46417 4017
rect 46417 3897 46422 4017
rect 45681 3574 45737 3630
rect 46499 3574 46555 3630
rect 47794 3511 47994 4311
rect 48658 3564 48663 3804
rect 48663 3564 48709 3804
rect 48709 3564 48714 3804
rect 49750 3564 49755 3804
rect 49755 3564 49801 3804
rect 49801 3564 49806 3804
rect 48760 3291 48816 3347
rect 50230 3564 50235 3804
rect 50235 3564 50281 3804
rect 50281 3564 50286 3804
rect 52184 3511 52484 4311
rect 53220 4242 53276 4298
rect 54260 4242 54316 4298
rect 50052 3213 50108 3269
rect 49572 3135 49628 3191
rect 47968 2144 47973 2384
rect 47973 2144 48019 2384
rect 48019 2144 48024 2384
rect 48862 2853 48867 2909
rect 48867 2853 48913 2909
rect 48913 2853 48918 2909
rect 49342 2853 49347 2909
rect 49347 2853 49393 2909
rect 49393 2853 49398 2909
rect 49546 2853 49551 2909
rect 49551 2853 49597 2909
rect 49597 2853 49602 2909
rect 49750 2853 49755 2909
rect 49755 2853 49801 2909
rect 49801 2853 49806 2909
rect 55746 4243 55802 4299
rect 53892 4135 53948 4148
rect 53892 4092 53893 4135
rect 53893 4092 53947 4135
rect 53947 4092 53948 4135
rect 54076 4135 54132 4148
rect 54076 4092 54077 4135
rect 54077 4092 54131 4135
rect 54131 4092 54132 4135
rect 54260 4135 54316 4148
rect 54260 4092 54261 4135
rect 54261 4092 54315 4135
rect 54315 4092 54316 4135
rect 54352 3896 54357 4016
rect 54357 3896 54403 4016
rect 54403 3896 54408 4016
rect 53667 3573 53723 3629
rect 54485 3573 54541 3629
rect 54838 3455 54894 3511
rect 50816 3175 52584 3315
rect 54662 3347 54718 3401
rect 50230 2853 50235 2909
rect 50235 2853 50281 2909
rect 50281 2853 50286 2909
rect 49756 2401 50356 2541
rect 51090 2672 51095 2912
rect 51095 2672 51141 2912
rect 51141 2672 51146 2912
rect 51774 2672 51779 2912
rect 51779 2672 51825 2912
rect 51825 2672 51830 2912
rect 51570 2338 51575 2578
rect 51575 2338 51621 2578
rect 51621 2338 51626 2578
rect 51978 2338 51983 2578
rect 51983 2338 52029 2578
rect 52029 2338 52034 2578
rect 52458 2388 52463 2628
rect 52463 2388 52509 2628
rect 52509 2388 52514 2628
rect 49756 2001 50356 2141
rect 50988 2115 51044 2171
rect 47790 1793 47846 1849
rect 43429 1250 43485 1306
rect 43612 1250 43668 1306
rect 47968 1433 47973 1489
rect 47973 1433 48019 1489
rect 48019 1433 48024 1489
rect 40580 873 40636 929
rect 40100 795 40156 851
rect 39390 513 39395 569
rect 39395 513 39441 569
rect 39441 513 39446 569
rect 39870 513 39875 569
rect 39875 513 39921 569
rect 39921 513 39926 569
rect 40074 513 40079 569
rect 40079 513 40125 569
rect 40125 513 40130 569
rect 40278 513 40283 569
rect 40283 513 40329 569
rect 40329 513 40334 569
rect 40758 513 40763 569
rect 40763 513 40809 569
rect 40809 513 40814 569
rect 42712 231 43012 1031
rect 48658 1224 48663 1464
rect 48663 1224 48709 1464
rect 48709 1224 48714 1464
rect 49750 1224 49755 1464
rect 49755 1224 49801 1464
rect 49801 1224 49806 1464
rect 48760 951 48816 1007
rect 50230 1224 50235 1464
rect 50235 1224 50281 1464
rect 50281 1224 50286 1464
rect 54168 3238 54224 3294
rect 53800 2851 53805 2971
rect 53805 2851 53851 2971
rect 53851 2851 53856 2971
rect 54168 2851 54173 2971
rect 54173 2851 54219 2971
rect 54219 2851 54224 2971
rect 53984 2551 53989 2671
rect 53989 2551 54035 2671
rect 54035 2551 54040 2671
rect 54490 2850 54495 2971
rect 54495 2850 54541 2971
rect 54541 2850 54546 2971
rect 54352 2551 54357 2671
rect 54357 2551 54403 2671
rect 54403 2551 54408 2671
rect 53892 2432 53893 2475
rect 53893 2432 53947 2475
rect 53947 2432 53948 2475
rect 53892 2419 53948 2432
rect 54076 2432 54077 2475
rect 54077 2432 54131 2475
rect 54131 2432 54132 2475
rect 54076 2419 54132 2432
rect 54260 2432 54261 2475
rect 54261 2432 54315 2475
rect 54315 2432 54316 2475
rect 54260 2419 54316 2432
rect 53892 2269 53948 2325
rect 53084 2153 53140 2209
rect 54076 2153 54132 2209
rect 54405 2153 54461 2209
rect 54838 2153 54894 2209
rect 52280 2037 52336 2093
rect 52850 2038 52904 2092
rect 54260 2037 54316 2093
rect 51672 1959 51728 2015
rect 50886 1677 50891 1733
rect 50891 1677 50937 1733
rect 50937 1677 50942 1733
rect 51774 1677 51779 1733
rect 51779 1677 51825 1733
rect 51825 1677 51830 1733
rect 52458 1677 52463 1733
rect 52463 1677 52509 1733
rect 52509 1677 52514 1733
rect 53892 1930 53948 1943
rect 53892 1887 53893 1930
rect 53893 1887 53947 1930
rect 53947 1887 53948 1930
rect 54076 1930 54132 1943
rect 54076 1887 54077 1930
rect 54077 1887 54131 1930
rect 54131 1887 54132 1930
rect 54260 1930 54316 1943
rect 54260 1887 54261 1930
rect 54261 1887 54315 1930
rect 54315 1887 54316 1930
rect 54352 1691 54357 1811
rect 54357 1691 54403 1811
rect 54403 1691 54408 1811
rect 53667 1368 53723 1424
rect 54485 1368 54541 1424
rect 50816 1215 52584 1355
rect 55378 4136 55434 4149
rect 55378 4093 55379 4136
rect 55379 4093 55433 4136
rect 55433 4093 55434 4136
rect 55562 4136 55618 4149
rect 55562 4093 55563 4136
rect 55563 4093 55617 4136
rect 55617 4093 55618 4136
rect 55746 4136 55802 4149
rect 55746 4093 55747 4136
rect 55747 4093 55801 4136
rect 55801 4093 55802 4136
rect 55838 3897 55843 4017
rect 55843 3897 55889 4017
rect 55889 3897 55894 4017
rect 55153 3574 55209 3630
rect 55971 3574 56027 3630
rect 52901 1250 52957 1306
rect 53084 1250 53140 1306
rect 50052 873 50108 929
rect 49572 795 49628 851
rect 48862 513 48867 569
rect 48867 513 48913 569
rect 48913 513 48918 569
rect 49342 513 49347 569
rect 49347 513 49393 569
rect 49393 513 49398 569
rect 49546 513 49551 569
rect 49551 513 49597 569
rect 49597 513 49602 569
rect 49750 513 49755 569
rect 49755 513 49801 569
rect 49801 513 49806 569
rect 50230 513 50235 569
rect 50235 513 50281 569
rect 50281 513 50286 569
rect 52184 231 52484 1031
<< metal2 >>
rect 6440 9908 7186 9920
rect 6440 9852 6808 9908
rect 6864 9852 7186 9908
rect 6440 9840 7186 9852
rect 6440 9587 6496 9840
rect 6808 9587 6864 9840
rect 7130 9587 7186 9840
rect 15912 9908 16658 9920
rect 15912 9852 16280 9908
rect 16336 9852 16658 9908
rect 15912 9840 16658 9852
rect 15912 9587 15968 9840
rect 16280 9587 16336 9840
rect 16602 9587 16658 9840
rect 25384 9909 26130 9921
rect 25384 9853 25752 9909
rect 25808 9853 26130 9909
rect 25384 9841 26130 9853
rect 25384 9588 25440 9841
rect 25752 9588 25808 9841
rect 26074 9588 26130 9841
rect 34856 9909 35602 9921
rect 34856 9853 35224 9909
rect 35280 9853 35602 9909
rect 34856 9841 35602 9853
rect 34856 9588 34912 9841
rect 35224 9588 35280 9841
rect 35546 9588 35602 9841
rect 44328 9909 45074 9921
rect 44328 9853 44696 9909
rect 44752 9853 45074 9909
rect 44328 9841 45074 9853
rect 44328 9588 44384 9841
rect 44696 9588 44752 9841
rect 45018 9588 45074 9841
rect 53800 9909 54546 9921
rect 53800 9853 54168 9909
rect 54224 9853 54546 9909
rect 53800 9841 54546 9853
rect 53800 9588 53856 9841
rect 54168 9588 54224 9841
rect 54490 9588 54546 9841
rect 6428 9585 6508 9587
rect 6428 9465 6440 9585
rect 6496 9465 6508 9585
rect 6428 9463 6508 9465
rect 6796 9585 6876 9587
rect 6796 9465 6808 9585
rect 6864 9465 6876 9585
rect 6796 9463 6876 9465
rect 7118 9585 7198 9587
rect 7118 9464 7130 9585
rect 7186 9464 7198 9585
rect 6440 9455 6496 9463
rect 6808 9455 6864 9463
rect 7118 9462 7198 9464
rect 15900 9585 15980 9587
rect 15900 9465 15912 9585
rect 15968 9465 15980 9585
rect 15900 9463 15980 9465
rect 16268 9585 16348 9587
rect 16268 9465 16280 9585
rect 16336 9465 16348 9585
rect 16268 9463 16348 9465
rect 16590 9585 16670 9587
rect 16590 9464 16602 9585
rect 16658 9464 16670 9585
rect 25372 9586 25452 9588
rect 25372 9466 25384 9586
rect 25440 9466 25452 9586
rect 25372 9464 25452 9466
rect 25740 9586 25820 9588
rect 25740 9466 25752 9586
rect 25808 9466 25820 9586
rect 25740 9464 25820 9466
rect 26062 9586 26142 9588
rect 26062 9465 26074 9586
rect 26130 9465 26142 9586
rect 7130 9454 7186 9462
rect 15912 9455 15968 9463
rect 16280 9455 16336 9463
rect 16590 9462 16670 9464
rect 16602 9454 16658 9462
rect 25384 9456 25440 9464
rect 25752 9456 25808 9464
rect 26062 9463 26142 9465
rect 34844 9586 34924 9588
rect 34844 9466 34856 9586
rect 34912 9466 34924 9586
rect 34844 9464 34924 9466
rect 35212 9586 35292 9588
rect 35212 9466 35224 9586
rect 35280 9466 35292 9586
rect 35212 9464 35292 9466
rect 35534 9586 35614 9588
rect 35534 9465 35546 9586
rect 35602 9465 35614 9586
rect 26074 9455 26130 9463
rect 34856 9456 34912 9464
rect 35224 9456 35280 9464
rect 35534 9463 35614 9465
rect 44316 9586 44396 9588
rect 44316 9466 44328 9586
rect 44384 9466 44396 9586
rect 44316 9464 44396 9466
rect 44684 9586 44764 9588
rect 44684 9466 44696 9586
rect 44752 9466 44764 9586
rect 44684 9464 44764 9466
rect 45006 9586 45086 9588
rect 45006 9465 45018 9586
rect 45074 9465 45086 9586
rect 35546 9455 35602 9463
rect 44328 9456 44384 9464
rect 44696 9456 44752 9464
rect 45006 9463 45086 9465
rect 53788 9586 53868 9588
rect 53788 9466 53800 9586
rect 53856 9466 53868 9586
rect 53788 9464 53868 9466
rect 54156 9586 54236 9588
rect 54156 9466 54168 9586
rect 54224 9466 54236 9586
rect 54156 9464 54236 9466
rect 54478 9586 54558 9588
rect 54478 9465 54490 9586
rect 54546 9465 54558 9586
rect 45018 9455 45074 9463
rect 53800 9456 53856 9464
rect 54168 9456 54224 9464
rect 54478 9463 54558 9465
rect 54490 9455 54546 9463
rect 6624 9287 6680 9295
rect 6992 9287 7048 9295
rect 16096 9287 16152 9295
rect 16464 9287 16520 9295
rect 25568 9288 25624 9296
rect 25936 9288 25992 9296
rect 35040 9288 35096 9296
rect 35408 9288 35464 9296
rect 44512 9288 44568 9296
rect 44880 9288 44936 9296
rect 53984 9288 54040 9296
rect 54352 9288 54408 9296
rect 6612 9285 7101 9287
rect 6612 9165 6624 9285
rect 6680 9165 6992 9285
rect 7048 9165 7101 9285
rect 6612 9163 7101 9165
rect 16084 9285 16573 9287
rect 16084 9165 16096 9285
rect 16152 9165 16464 9285
rect 16520 9165 16573 9285
rect 16084 9163 16573 9165
rect 25556 9286 26045 9288
rect 25556 9166 25568 9286
rect 25624 9166 25936 9286
rect 25992 9166 26045 9286
rect 25556 9164 26045 9166
rect 35028 9286 35517 9288
rect 35028 9166 35040 9286
rect 35096 9166 35408 9286
rect 35464 9166 35517 9286
rect 35028 9164 35517 9166
rect 44500 9286 44989 9288
rect 44500 9166 44512 9286
rect 44568 9166 44880 9286
rect 44936 9166 44989 9286
rect 44500 9164 44989 9166
rect 53972 9286 54461 9288
rect 53972 9166 53984 9286
rect 54040 9166 54352 9286
rect 54408 9166 54461 9286
rect 53972 9164 54461 9166
rect 6624 9155 6680 9163
rect 6992 9155 7101 9163
rect 16096 9155 16152 9163
rect 16464 9155 16573 9163
rect 25568 9156 25624 9164
rect 25936 9156 26045 9164
rect 35040 9156 35096 9164
rect 35408 9156 35517 9164
rect 44512 9156 44568 9164
rect 44880 9156 44989 9164
rect 53984 9156 54040 9164
rect 54352 9156 54461 9164
rect 6520 9089 6600 9099
rect 6520 9033 6532 9089
rect 6588 9033 6600 9089
rect 6520 9023 6600 9033
rect 6704 9089 6784 9099
rect 6704 9033 6716 9089
rect 6772 9033 6784 9089
rect 6704 9023 6784 9033
rect 6888 9089 6968 9099
rect 6888 9033 6900 9089
rect 6956 9033 6968 9089
rect 6888 9023 6968 9033
rect 5630 8939 5718 8951
rect 6532 8941 6588 9023
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 6520 8939 6600 8941
rect 6520 8883 6532 8939
rect 6588 8883 6600 8939
rect 6520 8881 6600 8883
rect 5848 8823 5918 8835
rect 5848 8767 5860 8823
rect 5916 8767 5918 8823
rect 5848 8755 5918 8767
rect 5712 6618 5782 6632
rect 5712 6562 5724 6618
rect 5780 6562 5782 6618
rect 5712 6550 5782 6562
rect 5430 5716 5512 5728
rect 5430 5660 5444 5716
rect 5500 5660 5512 5716
rect 5430 5648 5512 5660
rect 4814 4310 5134 4320
rect 1286 3803 2458 3813
rect 1286 3563 1298 3803
rect 1354 3563 2390 3803
rect 2446 3563 2458 3803
rect 1286 3553 2458 3563
rect 940 3346 1020 3356
rect 1380 3346 1458 3358
rect 10 3290 952 3346
rect 1008 3290 1400 3346
rect 1456 3290 1458 3346
rect 940 3280 1020 3290
rect 1380 3278 1458 3290
rect 2378 3268 2458 3553
rect 2858 3803 2938 3813
rect 2858 3563 2870 3803
rect 2926 3563 2938 3803
rect 2680 3268 2750 3280
rect 2378 3212 2692 3268
rect 2748 3212 2750 3268
rect 2200 3190 2270 3202
rect 10 3134 2212 3190
rect 2268 3134 2270 3190
rect 122 1848 178 3134
rect 2200 3122 2270 3134
rect 1490 2908 1570 2918
rect 1490 2852 1502 2908
rect 1558 2852 1570 2908
rect 1490 2666 1570 2852
rect 1970 2908 2050 2918
rect 1970 2852 1982 2908
rect 2038 2852 2050 2908
rect 1970 2842 2050 2852
rect 2174 2908 2254 2918
rect 2174 2852 2186 2908
rect 2242 2852 2254 2908
rect 2174 2666 2254 2852
rect 2378 2908 2458 3212
rect 2680 3200 2750 3212
rect 2858 3268 2938 3563
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 4814 3500 5134 3510
rect 3444 3314 5236 3326
rect 2858 3212 3215 3268
rect 2378 2852 2390 2908
rect 2446 2852 2458 2908
rect 2378 2842 2458 2852
rect 2858 2908 2938 3212
rect 2858 2852 2870 2908
rect 2926 2852 2938 2908
rect 2858 2842 2938 2852
rect 1490 2594 2254 2666
rect 2384 2540 3008 2552
rect 1156 2507 1256 2517
rect 1156 2431 1166 2507
rect 1246 2431 1256 2507
rect 1156 2421 1256 2431
rect 2384 2400 2396 2540
rect 2996 2400 3008 2540
rect 596 2383 676 2393
rect 2384 2388 3008 2400
rect 596 2143 608 2383
rect 664 2143 676 2383
rect 3159 2170 3215 3212
rect 3444 3174 3456 3314
rect 5224 3174 5236 3314
rect 3444 3162 5236 3174
rect 3718 2911 4482 2921
rect 3718 2671 3730 2911
rect 3786 2671 4414 2911
rect 4470 2671 4482 2911
rect 3718 2661 4482 2671
rect 5086 2627 5166 2637
rect 4198 2577 4686 2587
rect 4198 2337 4210 2577
rect 4266 2337 4618 2577
rect 4674 2337 4686 2577
rect 4198 2327 4686 2337
rect 3608 2170 3704 2182
rect 418 1848 488 1860
rect -446 1792 430 1848
rect 486 1792 488 1848
rect -441 -51 -385 1792
rect 418 1780 488 1792
rect 596 1848 676 2143
rect 2384 2140 3008 2152
rect 2384 2000 2396 2140
rect 2996 2000 3008 2140
rect 3159 2114 3628 2170
rect 3684 2114 3704 2170
rect 3608 2102 3704 2114
rect 4606 2092 4686 2327
rect 5086 2387 5098 2627
rect 5154 2387 5166 2627
rect 4908 2092 4978 2104
rect 4606 2036 4920 2092
rect 4976 2036 4978 2092
rect 4292 2014 4388 2024
rect 2384 1988 3008 2000
rect 3159 1958 4312 2014
rect 4368 1958 4388 2014
rect 596 1792 1034 1848
rect 596 1488 676 1792
rect 596 1432 608 1488
rect 664 1432 676 1488
rect 596 1422 676 1432
rect 978 1006 1034 1792
rect 1286 1463 2458 1473
rect 1286 1223 1298 1463
rect 1354 1223 2390 1463
rect 2446 1223 2458 1463
rect 1286 1213 2458 1223
rect 1380 1006 1458 1018
rect 978 950 1400 1006
rect 1456 950 1458 1006
rect 1380 938 1458 950
rect 2378 928 2458 1213
rect 2858 1463 2938 1473
rect 2858 1223 2870 1463
rect 2926 1223 2938 1463
rect 2680 928 2750 940
rect 2378 872 2692 928
rect 2748 872 2750 928
rect 2200 850 2270 862
rect -441 -181 -385 -171
rect 10 794 2212 850
rect 2268 794 2270 850
rect 10 -370 66 794
rect 2200 782 2270 794
rect 1490 568 1570 578
rect 1490 512 1502 568
rect 1558 512 1570 568
rect 1490 326 1570 512
rect 1970 568 2050 578
rect 1970 512 1982 568
rect 2038 512 2050 568
rect 1970 502 2050 512
rect 2174 568 2254 578
rect 2174 512 2186 568
rect 2242 512 2254 568
rect 2174 326 2254 512
rect 2378 568 2458 872
rect 2680 860 2750 872
rect 2858 928 2938 1223
rect 3159 928 3215 1958
rect 4292 1948 4388 1958
rect 4606 1742 4686 2036
rect 4908 2024 4978 2036
rect 5086 2092 5166 2387
rect 5724 2222 5780 6550
rect 5860 4309 5916 8755
rect 6532 8567 6588 8881
rect 6716 8825 6772 9023
rect 6704 8823 6784 8825
rect 6704 8767 6716 8823
rect 6772 8767 6784 8823
rect 6704 8765 6784 8767
rect 6716 8567 6772 8765
rect 6900 8709 6956 9023
rect 7033 8825 7101 9155
rect 15992 9089 16072 9099
rect 15992 9033 16004 9089
rect 16060 9033 16072 9089
rect 15992 9023 16072 9033
rect 16176 9089 16256 9099
rect 16176 9033 16188 9089
rect 16244 9033 16256 9089
rect 16176 9023 16256 9033
rect 16360 9089 16440 9099
rect 16360 9033 16372 9089
rect 16428 9033 16440 9089
rect 16360 9023 16440 9033
rect 15102 8939 15190 8951
rect 16004 8941 16060 9023
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 15992 8939 16072 8941
rect 15992 8883 16004 8939
rect 16060 8883 16072 8939
rect 15992 8881 16072 8883
rect 7033 8823 7113 8825
rect 7033 8767 7045 8823
rect 7101 8767 7113 8823
rect 7033 8765 7113 8767
rect 7300 8823 7370 8835
rect 7300 8767 7302 8823
rect 7358 8767 7370 8823
rect 6888 8707 6968 8709
rect 6888 8651 6900 8707
rect 6956 8651 6968 8707
rect 6888 8649 6968 8651
rect 6900 8567 6956 8649
rect 6520 8557 6600 8567
rect 6520 8501 6532 8557
rect 6588 8501 6600 8557
rect 6520 8491 6600 8501
rect 6704 8557 6784 8567
rect 6704 8501 6716 8557
rect 6772 8501 6784 8557
rect 6704 8491 6784 8501
rect 6888 8557 6968 8567
rect 6888 8501 6900 8557
rect 6956 8501 6968 8557
rect 6888 8491 6968 8501
rect 7033 8435 7101 8765
rect 7300 8757 7370 8767
rect 15320 8823 15390 8835
rect 15320 8767 15332 8823
rect 15388 8767 15390 8823
rect 6992 8427 7101 8435
rect 6980 8425 7101 8427
rect 6980 8305 6992 8425
rect 7048 8305 7101 8425
rect 6980 8303 7101 8305
rect 6992 8295 7048 8303
rect 6295 8038 7193 8050
rect 6295 7982 6307 8038
rect 6363 7982 7125 8038
rect 7181 7982 7193 8038
rect 6295 7970 7193 7982
rect 7302 7813 7358 8757
rect 15320 8755 15390 8767
rect 7466 7920 7546 7930
rect 7466 7864 7478 7920
rect 7534 7864 7546 7920
rect 7466 7862 7546 7864
rect 7300 7810 7370 7813
rect 7300 7756 7302 7810
rect 7358 7756 7370 7810
rect 7300 7744 7370 7756
rect 6440 7703 7186 7715
rect 6440 7647 6808 7703
rect 6864 7647 7186 7703
rect 6440 7635 7186 7647
rect 6440 7382 6496 7635
rect 6808 7382 6864 7635
rect 7130 7382 7186 7635
rect 6428 7380 6508 7382
rect 6428 7260 6440 7380
rect 6496 7260 6508 7380
rect 6428 7258 6508 7260
rect 6796 7380 6876 7382
rect 6796 7260 6808 7380
rect 6864 7260 6876 7380
rect 6796 7258 6876 7260
rect 7118 7380 7198 7382
rect 7118 7259 7130 7380
rect 7186 7259 7198 7380
rect 6440 7250 6496 7258
rect 6808 7250 6864 7258
rect 7118 7257 7198 7259
rect 7130 7249 7186 7257
rect 6624 7082 6680 7090
rect 6992 7082 7048 7090
rect 6612 7080 7101 7082
rect 6612 6960 6624 7080
rect 6680 6960 6992 7080
rect 7048 6960 7101 7080
rect 6612 6958 7101 6960
rect 6624 6950 6680 6958
rect 6992 6950 7101 6958
rect 6520 6884 6600 6894
rect 6520 6828 6532 6884
rect 6588 6828 6600 6884
rect 6520 6818 6600 6828
rect 6704 6884 6784 6894
rect 6704 6828 6716 6884
rect 6772 6828 6784 6884
rect 6704 6818 6784 6828
rect 6888 6884 6968 6894
rect 6888 6828 6900 6884
rect 6956 6828 6968 6884
rect 6888 6818 6968 6828
rect 6532 6736 6588 6818
rect 6520 6734 6600 6736
rect 6520 6678 6532 6734
rect 6588 6678 6600 6734
rect 6520 6676 6600 6678
rect 6532 6362 6588 6676
rect 6716 6620 6772 6818
rect 6704 6618 6784 6620
rect 6704 6562 6716 6618
rect 6772 6562 6784 6618
rect 6704 6560 6784 6562
rect 6716 6362 6772 6560
rect 6900 6504 6956 6818
rect 7033 6620 7101 6950
rect 7478 6628 7534 7862
rect 7926 7703 8672 7715
rect 7926 7647 8294 7703
rect 8350 7647 8672 7703
rect 7926 7635 8672 7647
rect 7926 7382 7982 7635
rect 8294 7382 8350 7635
rect 8616 7382 8672 7635
rect 7914 7380 7994 7382
rect 7914 7260 7926 7380
rect 7982 7260 7994 7380
rect 7914 7258 7994 7260
rect 8282 7380 8362 7382
rect 8282 7260 8294 7380
rect 8350 7260 8362 7380
rect 8282 7258 8362 7260
rect 8604 7380 8684 7382
rect 8604 7259 8616 7380
rect 8672 7259 8684 7380
rect 7926 7250 7982 7258
rect 8294 7250 8350 7258
rect 8604 7257 8684 7259
rect 8616 7249 8672 7257
rect 8110 7082 8166 7090
rect 8478 7082 8534 7090
rect 8098 7080 8587 7082
rect 8098 6960 8110 7080
rect 8166 6960 8478 7080
rect 8534 6960 8587 7080
rect 8098 6958 8587 6960
rect 8110 6950 8166 6958
rect 8478 6950 8587 6958
rect 8006 6884 8086 6894
rect 8006 6828 8018 6884
rect 8074 6828 8086 6884
rect 8006 6818 8086 6828
rect 8190 6884 8270 6894
rect 8190 6828 8202 6884
rect 8258 6828 8270 6884
rect 8190 6818 8270 6828
rect 8374 6884 8454 6894
rect 8374 6828 8386 6884
rect 8442 6828 8454 6884
rect 8374 6818 8454 6828
rect 8018 6736 8074 6818
rect 8006 6734 8086 6736
rect 8006 6678 8018 6734
rect 8074 6678 8086 6734
rect 8006 6676 8086 6678
rect 7033 6618 7113 6620
rect 7033 6562 7045 6618
rect 7101 6562 7113 6618
rect 7033 6560 7113 6562
rect 7476 6618 7536 6628
rect 7476 6562 7478 6618
rect 7534 6562 7536 6618
rect 6888 6502 6968 6504
rect 6888 6446 6900 6502
rect 6956 6446 6968 6502
rect 6888 6444 6968 6446
rect 6900 6362 6956 6444
rect 6520 6352 6600 6362
rect 6520 6296 6532 6352
rect 6588 6296 6600 6352
rect 6520 6286 6600 6296
rect 6704 6352 6784 6362
rect 6704 6296 6716 6352
rect 6772 6296 6784 6352
rect 6704 6286 6784 6296
rect 6888 6352 6968 6362
rect 6888 6296 6900 6352
rect 6956 6296 6968 6352
rect 6888 6286 6968 6296
rect 7033 6230 7101 6560
rect 7476 6550 7536 6562
rect 6992 6222 7101 6230
rect 6980 6220 7101 6222
rect 6980 6100 6992 6220
rect 7048 6100 7101 6220
rect 6980 6098 7101 6100
rect 6992 6090 7048 6098
rect 6295 5833 7191 5845
rect 6295 5777 6307 5833
rect 6363 5777 7125 5833
rect 7181 5777 7191 5833
rect 6295 5765 7191 5777
rect 7478 5607 7534 6550
rect 8018 6362 8074 6676
rect 8202 6620 8258 6818
rect 8190 6618 8270 6620
rect 8190 6562 8202 6618
rect 8258 6562 8270 6618
rect 8190 6560 8270 6562
rect 8202 6362 8258 6560
rect 8386 6504 8442 6818
rect 8519 6620 8587 6950
rect 8519 6618 8599 6620
rect 8519 6562 8531 6618
rect 8587 6562 8599 6618
rect 8519 6560 8599 6562
rect 8786 6618 8856 6630
rect 15184 6618 15254 6632
rect 8786 6562 8788 6618
rect 8844 6562 9542 6618
rect 8374 6502 8454 6504
rect 8374 6446 8386 6502
rect 8442 6446 8454 6502
rect 8374 6444 8454 6446
rect 8386 6362 8442 6444
rect 8006 6352 8086 6362
rect 8006 6296 8018 6352
rect 8074 6296 8086 6352
rect 8006 6286 8086 6296
rect 8190 6352 8270 6362
rect 8190 6296 8202 6352
rect 8258 6296 8270 6352
rect 8190 6286 8270 6296
rect 8374 6352 8454 6362
rect 8374 6296 8386 6352
rect 8442 6296 8454 6352
rect 8374 6286 8454 6296
rect 8519 6230 8587 6560
rect 8786 6552 8856 6562
rect 8478 6222 8587 6230
rect 8466 6220 8587 6222
rect 8466 6100 8478 6220
rect 8534 6100 8587 6220
rect 8466 6098 8587 6100
rect 8478 6090 8534 6098
rect 7781 5833 8677 5845
rect 7781 5777 7793 5833
rect 7849 5777 8611 5833
rect 8667 5777 8677 5833
rect 7781 5765 8677 5777
rect 8788 5608 8844 6552
rect 8952 5716 9032 5726
rect 8952 5660 8964 5716
rect 9020 5660 9032 5716
rect 8952 5658 9032 5660
rect 7476 5605 7546 5607
rect 7476 5549 7478 5605
rect 7534 5549 7546 5605
rect 7476 5537 7546 5549
rect 8776 5606 8856 5608
rect 8776 5550 8788 5606
rect 8844 5550 8856 5606
rect 8776 5538 8856 5550
rect 6440 5498 7186 5510
rect 6440 5442 6808 5498
rect 6864 5442 7186 5498
rect 6440 5430 7186 5442
rect 6440 5177 6496 5430
rect 6808 5177 6864 5430
rect 7130 5177 7186 5430
rect 7926 5499 8672 5511
rect 7926 5443 8294 5499
rect 8350 5443 8672 5499
rect 7926 5431 8672 5443
rect 7926 5178 7982 5431
rect 8294 5178 8350 5431
rect 8616 5178 8672 5431
rect 6428 5175 6508 5177
rect 6428 5055 6440 5175
rect 6496 5055 6508 5175
rect 6428 5053 6508 5055
rect 6796 5175 6876 5177
rect 6796 5055 6808 5175
rect 6864 5055 6876 5175
rect 6796 5053 6876 5055
rect 7118 5175 7198 5177
rect 7118 5054 7130 5175
rect 7186 5054 7198 5175
rect 7914 5176 7994 5178
rect 7914 5056 7926 5176
rect 7982 5056 7994 5176
rect 7914 5054 7994 5056
rect 8282 5176 8362 5178
rect 8282 5056 8294 5176
rect 8350 5056 8362 5176
rect 8282 5054 8362 5056
rect 8604 5176 8684 5178
rect 8604 5055 8616 5176
rect 8672 5055 8684 5176
rect 6440 5045 6496 5053
rect 6808 5045 6864 5053
rect 7118 5052 7198 5054
rect 7130 5044 7186 5052
rect 7926 5046 7982 5054
rect 8294 5046 8350 5054
rect 8604 5053 8684 5055
rect 8616 5045 8672 5053
rect 6624 4877 6680 4885
rect 6992 4877 7048 4885
rect 8110 4878 8166 4886
rect 8478 4878 8534 4886
rect 6612 4875 7101 4877
rect 6612 4755 6624 4875
rect 6680 4755 6992 4875
rect 7048 4755 7101 4875
rect 6612 4753 7101 4755
rect 8098 4876 8587 4878
rect 8098 4756 8110 4876
rect 8166 4756 8478 4876
rect 8534 4756 8587 4876
rect 8098 4754 8587 4756
rect 6624 4745 6680 4753
rect 6992 4745 7101 4753
rect 8110 4746 8166 4754
rect 8478 4746 8587 4754
rect 6520 4679 6600 4689
rect 6520 4623 6532 4679
rect 6588 4623 6600 4679
rect 6520 4613 6600 4623
rect 6704 4679 6784 4689
rect 6704 4623 6716 4679
rect 6772 4623 6784 4679
rect 6704 4613 6784 4623
rect 6888 4679 6968 4689
rect 6888 4623 6900 4679
rect 6956 4623 6968 4679
rect 6888 4613 6968 4623
rect 6532 4531 6588 4613
rect 6520 4529 6600 4531
rect 6520 4473 6532 4529
rect 6588 4473 6600 4529
rect 6520 4471 6600 4473
rect 5848 4297 5918 4309
rect 5848 4241 5860 4297
rect 5916 4241 5918 4297
rect 5848 4229 5918 4241
rect 6532 4157 6588 4471
rect 6716 4415 6772 4613
rect 6704 4413 6784 4415
rect 6704 4357 6716 4413
rect 6772 4357 6784 4413
rect 6704 4355 6784 4357
rect 6716 4157 6772 4355
rect 6900 4299 6956 4613
rect 7033 4415 7101 4745
rect 8006 4680 8086 4690
rect 8006 4624 8018 4680
rect 8074 4624 8086 4680
rect 8006 4614 8086 4624
rect 8190 4680 8270 4690
rect 8190 4624 8202 4680
rect 8258 4624 8270 4680
rect 8190 4614 8270 4624
rect 8374 4680 8454 4690
rect 8374 4624 8386 4680
rect 8442 4624 8454 4680
rect 8374 4614 8454 4624
rect 8018 4532 8074 4614
rect 8006 4530 8086 4532
rect 8006 4474 8018 4530
rect 8074 4474 8086 4530
rect 8006 4472 8086 4474
rect 7033 4413 7113 4415
rect 7033 4357 7045 4413
rect 7101 4357 7113 4413
rect 7033 4355 7113 4357
rect 7300 4413 7370 4425
rect 7300 4357 7302 4413
rect 7358 4357 7370 4413
rect 6888 4297 6968 4299
rect 6888 4241 6900 4297
rect 6956 4241 6968 4297
rect 6888 4239 6968 4241
rect 6900 4157 6956 4239
rect 6520 4147 6600 4157
rect 6520 4091 6532 4147
rect 6588 4091 6600 4147
rect 6520 4081 6600 4091
rect 6704 4147 6784 4157
rect 6704 4091 6716 4147
rect 6772 4091 6784 4147
rect 6704 4081 6784 4091
rect 6888 4147 6968 4157
rect 6888 4091 6900 4147
rect 6956 4091 6968 4147
rect 6888 4081 6968 4091
rect 7033 4025 7101 4355
rect 7300 4347 7370 4357
rect 6992 4017 7101 4025
rect 6980 4015 7101 4017
rect 6980 3895 6992 4015
rect 7048 3895 7101 4015
rect 6980 3893 7101 3895
rect 6992 3885 7048 3893
rect 6295 3628 7191 3640
rect 6295 3572 6307 3628
rect 6363 3572 7125 3628
rect 7181 3572 7191 3628
rect 6295 3560 7191 3572
rect 7302 3403 7358 4347
rect 8018 4158 8074 4472
rect 8202 4416 8258 4614
rect 8190 4414 8270 4416
rect 8190 4358 8202 4414
rect 8258 4358 8270 4414
rect 8190 4356 8270 4358
rect 8202 4158 8258 4356
rect 8386 4300 8442 4614
rect 8519 4416 8587 4746
rect 8964 4424 9020 5658
rect 8519 4414 8599 4416
rect 8519 4358 8531 4414
rect 8587 4358 8599 4414
rect 8519 4356 8599 4358
rect 8962 4414 9032 4424
rect 8962 4358 8964 4414
rect 9020 4358 9112 4414
rect 8374 4298 8454 4300
rect 8374 4242 8386 4298
rect 8442 4242 8454 4298
rect 8374 4240 8454 4242
rect 8386 4158 8442 4240
rect 8006 4148 8086 4158
rect 8006 4092 8018 4148
rect 8074 4092 8086 4148
rect 8006 4082 8086 4092
rect 8190 4148 8270 4158
rect 8190 4092 8202 4148
rect 8258 4092 8270 4148
rect 8190 4082 8270 4092
rect 8374 4148 8454 4158
rect 8374 4092 8386 4148
rect 8442 4092 8454 4148
rect 8374 4082 8454 4092
rect 8519 4026 8587 4356
rect 8962 4346 9032 4358
rect 8478 4018 8587 4026
rect 8466 4016 8587 4018
rect 8466 3896 8478 4016
rect 8534 3896 8587 4016
rect 8466 3894 8587 3896
rect 8478 3886 8534 3894
rect 7781 3629 8677 3641
rect 7781 3573 7793 3629
rect 7849 3573 8611 3629
rect 8667 3573 8677 3629
rect 7781 3561 8677 3573
rect 7466 3510 7546 3520
rect 7466 3454 7478 3510
rect 7534 3454 7546 3510
rect 7466 3452 7546 3454
rect 7300 3400 7370 3403
rect 7300 3346 7302 3400
rect 7358 3346 7370 3400
rect 7300 3334 7370 3346
rect 6440 3293 7186 3305
rect 6440 3237 6808 3293
rect 6864 3237 7186 3293
rect 6440 3225 7186 3237
rect 6440 2972 6496 3225
rect 6808 2972 6864 3225
rect 7130 2972 7186 3225
rect 6428 2970 6508 2972
rect 6428 2850 6440 2970
rect 6496 2850 6508 2970
rect 6428 2848 6508 2850
rect 6796 2970 6876 2972
rect 6796 2850 6808 2970
rect 6864 2850 6876 2970
rect 6796 2848 6876 2850
rect 7118 2970 7198 2972
rect 7118 2849 7130 2970
rect 7186 2849 7198 2970
rect 6440 2840 6496 2848
rect 6808 2840 6864 2848
rect 7118 2847 7198 2849
rect 7130 2839 7186 2847
rect 6624 2672 6680 2680
rect 6992 2672 7048 2680
rect 6612 2670 7101 2672
rect 6612 2550 6624 2670
rect 6680 2550 6992 2670
rect 7048 2550 7101 2670
rect 6612 2548 7101 2550
rect 6624 2540 6680 2548
rect 6992 2540 7101 2548
rect 6520 2474 6600 2484
rect 6520 2418 6532 2474
rect 6588 2418 6600 2474
rect 6520 2408 6600 2418
rect 6704 2474 6784 2484
rect 6704 2418 6716 2474
rect 6772 2418 6784 2474
rect 6704 2408 6784 2418
rect 6888 2474 6968 2484
rect 6888 2418 6900 2474
rect 6956 2418 6968 2474
rect 6888 2408 6968 2418
rect 6532 2326 6588 2408
rect 6520 2324 6600 2326
rect 6520 2268 6532 2324
rect 6588 2268 6600 2324
rect 6520 2266 6600 2268
rect 5712 2208 5782 2222
rect 5712 2152 5724 2208
rect 5780 2152 5782 2208
rect 5712 2140 5782 2152
rect 5478 2092 5556 2103
rect 5086 2091 5556 2092
rect 5086 2037 5490 2091
rect 5544 2037 5556 2091
rect 5086 2036 5556 2037
rect 3514 1732 4686 1742
rect 3514 1676 3526 1732
rect 3582 1676 4414 1732
rect 4470 1676 4686 1732
rect 3514 1666 4686 1676
rect 5086 1732 5166 2036
rect 5478 2025 5556 2036
rect 5086 1676 5098 1732
rect 5154 1676 5166 1732
rect 5086 1666 5166 1676
rect 3444 1354 5236 1366
rect 3444 1214 3456 1354
rect 5224 1214 5236 1354
rect 5529 1305 5615 1317
rect 5724 1309 5780 2140
rect 6532 1952 6588 2266
rect 6716 2210 6772 2408
rect 6704 2208 6784 2210
rect 6704 2152 6716 2208
rect 6772 2152 6784 2208
rect 6704 2150 6784 2152
rect 6716 1952 6772 2150
rect 6900 2094 6956 2408
rect 7033 2210 7101 2540
rect 7478 2220 7534 3452
rect 9486 3346 9542 6562
rect 15184 6562 15196 6618
rect 15252 6562 15254 6618
rect 15184 6550 15254 6562
rect 14902 5716 14984 5728
rect 14902 5660 14916 5716
rect 14972 5660 14984 5716
rect 14902 5648 14984 5660
rect 9896 4310 10116 4320
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 14286 4310 14606 4320
rect 10758 3803 11930 3813
rect 10758 3563 10770 3803
rect 10826 3563 11862 3803
rect 11918 3563 11930 3803
rect 10758 3553 11930 3563
rect 9896 3500 10116 3510
rect 10852 3346 10930 3358
rect 9482 3290 10872 3346
rect 10928 3290 10930 3346
rect 10852 3278 10930 3290
rect 11850 3268 11930 3553
rect 12330 3803 12410 3813
rect 12330 3563 12342 3803
rect 12398 3563 12410 3803
rect 12152 3268 12222 3280
rect 11850 3212 12164 3268
rect 12220 3212 12222 3268
rect 11672 3190 11742 3202
rect 9482 3134 11684 3190
rect 11740 3134 11742 3190
rect 7033 2208 7113 2210
rect 7033 2152 7045 2208
rect 7101 2152 7113 2208
rect 7033 2150 7113 2152
rect 7476 2208 7536 2220
rect 7476 2152 7478 2208
rect 7534 2152 7536 2208
rect 6888 2092 6968 2094
rect 6888 2036 6900 2092
rect 6956 2036 6968 2092
rect 6888 2034 6968 2036
rect 6900 1952 6956 2034
rect 6520 1942 6600 1952
rect 6520 1886 6532 1942
rect 6588 1886 6600 1942
rect 6520 1876 6600 1886
rect 6704 1942 6784 1952
rect 6704 1886 6716 1942
rect 6772 1886 6784 1942
rect 6704 1876 6784 1886
rect 6888 1942 6968 1952
rect 6888 1886 6900 1942
rect 6956 1886 6968 1942
rect 6888 1876 6968 1886
rect 7033 1820 7101 2150
rect 7476 2140 7536 2152
rect 9594 1849 9650 3134
rect 11672 3122 11742 3134
rect 10962 2908 11042 2918
rect 10962 2852 10974 2908
rect 11030 2852 11042 2908
rect 10962 2666 11042 2852
rect 11442 2908 11522 2918
rect 11442 2852 11454 2908
rect 11510 2852 11522 2908
rect 11442 2842 11522 2852
rect 11646 2908 11726 2918
rect 11646 2852 11658 2908
rect 11714 2852 11726 2908
rect 11646 2666 11726 2852
rect 11850 2908 11930 3212
rect 12152 3200 12222 3212
rect 12330 3268 12410 3563
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 14286 3500 14606 3510
rect 12916 3314 14708 3326
rect 12330 3212 12687 3268
rect 11850 2852 11862 2908
rect 11918 2852 11930 2908
rect 11850 2842 11930 2852
rect 12330 2908 12410 3212
rect 12330 2852 12342 2908
rect 12398 2852 12410 2908
rect 12330 2842 12410 2852
rect 10962 2594 11726 2666
rect 11856 2540 12480 2552
rect 11856 2400 11868 2540
rect 12468 2400 12480 2540
rect 10068 2383 10148 2393
rect 11856 2388 12480 2400
rect 10068 2143 10080 2383
rect 10136 2143 10148 2383
rect 12631 2170 12687 3212
rect 12916 3174 12928 3314
rect 14696 3174 14708 3314
rect 12916 3162 14708 3174
rect 13190 2911 13954 2921
rect 13190 2671 13202 2911
rect 13258 2671 13886 2911
rect 13942 2671 13954 2911
rect 13190 2661 13954 2671
rect 14558 2627 14638 2637
rect 13670 2577 14158 2587
rect 13670 2337 13682 2577
rect 13738 2337 14090 2577
rect 14146 2337 14158 2577
rect 13670 2327 14158 2337
rect 13080 2170 13176 2182
rect 6992 1812 7101 1820
rect 6980 1810 7101 1812
rect 6980 1690 6992 1810
rect 7048 1690 7101 1810
rect 9082 1848 9650 1849
rect 9890 1848 9960 1860
rect 9082 1793 9902 1848
rect 6980 1688 7101 1690
rect 6992 1680 7048 1688
rect 6295 1423 7193 1435
rect 6295 1367 6307 1423
rect 6363 1367 7125 1423
rect 7181 1367 7193 1423
rect 6295 1355 7193 1367
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 5722 1305 5782 1309
rect 5722 1249 5724 1305
rect 5780 1249 5782 1305
rect 5722 1237 5782 1249
rect 3444 1202 5236 1214
rect 2858 872 3215 928
rect 4814 1030 5134 1040
rect 2378 512 2390 568
rect 2446 512 2458 568
rect 2378 502 2458 512
rect 2858 568 2938 872
rect 2858 512 2870 568
rect 2926 512 2938 568
rect 2858 502 2938 512
rect 1490 254 2254 326
rect 4814 230 4824 1030
rect 5124 230 5134 1030
rect 4814 220 5134 230
rect 9087 -50 9143 1793
rect 9594 1792 9902 1793
rect 9958 1792 9960 1848
rect 9890 1780 9960 1792
rect 10068 1848 10148 2143
rect 11856 2140 12480 2152
rect 11856 2000 11868 2140
rect 12468 2000 12480 2140
rect 12631 2114 13100 2170
rect 13156 2114 13176 2170
rect 13080 2102 13176 2114
rect 14078 2092 14158 2327
rect 14558 2387 14570 2627
rect 14626 2387 14638 2627
rect 14380 2092 14450 2104
rect 14078 2036 14392 2092
rect 14448 2036 14450 2092
rect 13764 2014 13860 2024
rect 11856 1988 12480 2000
rect 12631 1958 13784 2014
rect 13840 1958 13860 2014
rect 10068 1792 10506 1848
rect 10068 1488 10148 1792
rect 10068 1432 10080 1488
rect 10136 1432 10148 1488
rect 10068 1422 10148 1432
rect 10450 1006 10506 1792
rect 10758 1463 11930 1473
rect 10758 1223 10770 1463
rect 10826 1223 11862 1463
rect 11918 1223 11930 1463
rect 10758 1213 11930 1223
rect 10852 1006 10930 1018
rect 10450 950 10872 1006
rect 10928 950 10930 1006
rect 10852 938 10930 950
rect 11850 928 11930 1213
rect 12330 1463 12410 1473
rect 12330 1223 12342 1463
rect 12398 1223 12410 1463
rect 12152 928 12222 940
rect 11850 872 12164 928
rect 12220 872 12222 928
rect 11672 850 11742 862
rect 9087 -180 9143 -170
rect 9482 794 11684 850
rect 11740 794 11742 850
rect 9482 -370 9538 794
rect 11672 782 11742 794
rect 10962 568 11042 578
rect 10962 512 10974 568
rect 11030 512 11042 568
rect 10962 326 11042 512
rect 11442 568 11522 578
rect 11442 512 11454 568
rect 11510 512 11522 568
rect 11442 502 11522 512
rect 11646 568 11726 578
rect 11646 512 11658 568
rect 11714 512 11726 568
rect 11646 326 11726 512
rect 11850 568 11930 872
rect 12152 860 12222 872
rect 12330 928 12410 1223
rect 12631 928 12687 1958
rect 13764 1948 13860 1958
rect 14078 1742 14158 2036
rect 14380 2024 14450 2036
rect 14558 2092 14638 2387
rect 15196 2222 15252 6550
rect 15332 4309 15388 8755
rect 16004 8567 16060 8881
rect 16188 8825 16244 9023
rect 16176 8823 16256 8825
rect 16176 8767 16188 8823
rect 16244 8767 16256 8823
rect 16176 8765 16256 8767
rect 16188 8567 16244 8765
rect 16372 8709 16428 9023
rect 16505 8825 16573 9155
rect 25464 9090 25544 9100
rect 25464 9034 25476 9090
rect 25532 9034 25544 9090
rect 25464 9024 25544 9034
rect 25648 9090 25728 9100
rect 25648 9034 25660 9090
rect 25716 9034 25728 9090
rect 25648 9024 25728 9034
rect 25832 9090 25912 9100
rect 25832 9034 25844 9090
rect 25900 9034 25912 9090
rect 25832 9024 25912 9034
rect 24574 8940 24662 8952
rect 25476 8942 25532 9024
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 25464 8940 25544 8942
rect 25464 8884 25476 8940
rect 25532 8884 25544 8940
rect 25464 8882 25544 8884
rect 16505 8823 16585 8825
rect 16505 8767 16517 8823
rect 16573 8767 16585 8823
rect 16505 8765 16585 8767
rect 16772 8823 16842 8835
rect 16772 8767 16774 8823
rect 16830 8767 16842 8823
rect 16360 8707 16440 8709
rect 16360 8651 16372 8707
rect 16428 8651 16440 8707
rect 16360 8649 16440 8651
rect 16372 8567 16428 8649
rect 15992 8557 16072 8567
rect 15992 8501 16004 8557
rect 16060 8501 16072 8557
rect 15992 8491 16072 8501
rect 16176 8557 16256 8567
rect 16176 8501 16188 8557
rect 16244 8501 16256 8557
rect 16176 8491 16256 8501
rect 16360 8557 16440 8567
rect 16360 8501 16372 8557
rect 16428 8501 16440 8557
rect 16360 8491 16440 8501
rect 16505 8435 16573 8765
rect 16772 8757 16842 8767
rect 24792 8824 24862 8836
rect 24792 8768 24804 8824
rect 24860 8768 24862 8824
rect 16464 8427 16573 8435
rect 16452 8425 16573 8427
rect 16452 8305 16464 8425
rect 16520 8305 16573 8425
rect 16452 8303 16573 8305
rect 16464 8295 16520 8303
rect 15767 8038 16665 8050
rect 15767 7982 15779 8038
rect 15835 7982 16597 8038
rect 16653 7982 16665 8038
rect 15767 7970 16665 7982
rect 16774 7813 16830 8757
rect 24792 8756 24862 8768
rect 16938 7920 17018 7930
rect 16938 7864 16950 7920
rect 17006 7864 17018 7920
rect 16938 7862 17018 7864
rect 16772 7810 16842 7813
rect 16772 7756 16774 7810
rect 16830 7756 16842 7810
rect 16772 7744 16842 7756
rect 15912 7703 16658 7715
rect 15912 7647 16280 7703
rect 16336 7647 16658 7703
rect 15912 7635 16658 7647
rect 15912 7382 15968 7635
rect 16280 7382 16336 7635
rect 16602 7382 16658 7635
rect 15900 7380 15980 7382
rect 15900 7260 15912 7380
rect 15968 7260 15980 7380
rect 15900 7258 15980 7260
rect 16268 7380 16348 7382
rect 16268 7260 16280 7380
rect 16336 7260 16348 7380
rect 16268 7258 16348 7260
rect 16590 7380 16670 7382
rect 16590 7259 16602 7380
rect 16658 7259 16670 7380
rect 15912 7250 15968 7258
rect 16280 7250 16336 7258
rect 16590 7257 16670 7259
rect 16602 7249 16658 7257
rect 16096 7082 16152 7090
rect 16464 7082 16520 7090
rect 16084 7080 16573 7082
rect 16084 6960 16096 7080
rect 16152 6960 16464 7080
rect 16520 6960 16573 7080
rect 16084 6958 16573 6960
rect 16096 6950 16152 6958
rect 16464 6950 16573 6958
rect 15992 6884 16072 6894
rect 15992 6828 16004 6884
rect 16060 6828 16072 6884
rect 15992 6818 16072 6828
rect 16176 6884 16256 6894
rect 16176 6828 16188 6884
rect 16244 6828 16256 6884
rect 16176 6818 16256 6828
rect 16360 6884 16440 6894
rect 16360 6828 16372 6884
rect 16428 6828 16440 6884
rect 16360 6818 16440 6828
rect 16004 6736 16060 6818
rect 15992 6734 16072 6736
rect 15992 6678 16004 6734
rect 16060 6678 16072 6734
rect 15992 6676 16072 6678
rect 16004 6362 16060 6676
rect 16188 6620 16244 6818
rect 16176 6618 16256 6620
rect 16176 6562 16188 6618
rect 16244 6562 16256 6618
rect 16176 6560 16256 6562
rect 16188 6362 16244 6560
rect 16372 6504 16428 6818
rect 16505 6620 16573 6950
rect 16950 6628 17006 7862
rect 17398 7703 18144 7715
rect 17398 7647 17766 7703
rect 17822 7647 18144 7703
rect 17398 7635 18144 7647
rect 17398 7382 17454 7635
rect 17766 7382 17822 7635
rect 18088 7382 18144 7635
rect 17386 7380 17466 7382
rect 17386 7260 17398 7380
rect 17454 7260 17466 7380
rect 17386 7258 17466 7260
rect 17754 7380 17834 7382
rect 17754 7260 17766 7380
rect 17822 7260 17834 7380
rect 17754 7258 17834 7260
rect 18076 7380 18156 7382
rect 18076 7259 18088 7380
rect 18144 7259 18156 7380
rect 17398 7250 17454 7258
rect 17766 7250 17822 7258
rect 18076 7257 18156 7259
rect 18088 7249 18144 7257
rect 17582 7082 17638 7090
rect 17950 7082 18006 7090
rect 17570 7080 18059 7082
rect 17570 6960 17582 7080
rect 17638 6960 17950 7080
rect 18006 6960 18059 7080
rect 17570 6958 18059 6960
rect 17582 6950 17638 6958
rect 17950 6950 18059 6958
rect 17478 6884 17558 6894
rect 17478 6828 17490 6884
rect 17546 6828 17558 6884
rect 17478 6818 17558 6828
rect 17662 6884 17742 6894
rect 17662 6828 17674 6884
rect 17730 6828 17742 6884
rect 17662 6818 17742 6828
rect 17846 6884 17926 6894
rect 17846 6828 17858 6884
rect 17914 6828 17926 6884
rect 17846 6818 17926 6828
rect 17490 6736 17546 6818
rect 17478 6734 17558 6736
rect 17478 6678 17490 6734
rect 17546 6678 17558 6734
rect 17478 6676 17558 6678
rect 16505 6618 16585 6620
rect 16505 6562 16517 6618
rect 16573 6562 16585 6618
rect 16505 6560 16585 6562
rect 16948 6618 17008 6628
rect 16948 6562 16950 6618
rect 17006 6562 17008 6618
rect 16360 6502 16440 6504
rect 16360 6446 16372 6502
rect 16428 6446 16440 6502
rect 16360 6444 16440 6446
rect 16372 6362 16428 6444
rect 15992 6352 16072 6362
rect 15992 6296 16004 6352
rect 16060 6296 16072 6352
rect 15992 6286 16072 6296
rect 16176 6352 16256 6362
rect 16176 6296 16188 6352
rect 16244 6296 16256 6352
rect 16176 6286 16256 6296
rect 16360 6352 16440 6362
rect 16360 6296 16372 6352
rect 16428 6296 16440 6352
rect 16360 6286 16440 6296
rect 16505 6230 16573 6560
rect 16948 6550 17008 6562
rect 16464 6222 16573 6230
rect 16452 6220 16573 6222
rect 16452 6100 16464 6220
rect 16520 6100 16573 6220
rect 16452 6098 16573 6100
rect 16464 6090 16520 6098
rect 15767 5833 16663 5845
rect 15767 5777 15779 5833
rect 15835 5777 16597 5833
rect 16653 5777 16663 5833
rect 15767 5765 16663 5777
rect 16950 5607 17006 6550
rect 17490 6362 17546 6676
rect 17674 6620 17730 6818
rect 17662 6618 17742 6620
rect 17662 6562 17674 6618
rect 17730 6562 17742 6618
rect 17662 6560 17742 6562
rect 17674 6362 17730 6560
rect 17858 6504 17914 6818
rect 17991 6620 18059 6950
rect 17991 6618 18071 6620
rect 17991 6562 18003 6618
rect 18059 6562 18071 6618
rect 17991 6560 18071 6562
rect 18258 6618 18328 6630
rect 24656 6619 24726 6633
rect 18258 6562 18260 6618
rect 18316 6562 19014 6618
rect 17846 6502 17926 6504
rect 17846 6446 17858 6502
rect 17914 6446 17926 6502
rect 17846 6444 17926 6446
rect 17858 6362 17914 6444
rect 17478 6352 17558 6362
rect 17478 6296 17490 6352
rect 17546 6296 17558 6352
rect 17478 6286 17558 6296
rect 17662 6352 17742 6362
rect 17662 6296 17674 6352
rect 17730 6296 17742 6352
rect 17662 6286 17742 6296
rect 17846 6352 17926 6362
rect 17846 6296 17858 6352
rect 17914 6296 17926 6352
rect 17846 6286 17926 6296
rect 17991 6230 18059 6560
rect 18258 6552 18328 6562
rect 17950 6222 18059 6230
rect 17938 6220 18059 6222
rect 17938 6100 17950 6220
rect 18006 6100 18059 6220
rect 17938 6098 18059 6100
rect 17950 6090 18006 6098
rect 17253 5833 18149 5845
rect 17253 5777 17265 5833
rect 17321 5777 18083 5833
rect 18139 5777 18149 5833
rect 17253 5765 18149 5777
rect 18260 5608 18316 6552
rect 18424 5716 18504 5726
rect 18424 5660 18436 5716
rect 18492 5660 18504 5716
rect 18424 5658 18504 5660
rect 16948 5605 17018 5607
rect 16948 5549 16950 5605
rect 17006 5549 17018 5605
rect 16948 5537 17018 5549
rect 18248 5606 18328 5608
rect 18248 5550 18260 5606
rect 18316 5550 18328 5606
rect 18248 5538 18328 5550
rect 15912 5498 16658 5510
rect 15912 5442 16280 5498
rect 16336 5442 16658 5498
rect 15912 5430 16658 5442
rect 15912 5177 15968 5430
rect 16280 5177 16336 5430
rect 16602 5177 16658 5430
rect 17398 5499 18144 5511
rect 17398 5443 17766 5499
rect 17822 5443 18144 5499
rect 17398 5431 18144 5443
rect 17398 5178 17454 5431
rect 17766 5178 17822 5431
rect 18088 5178 18144 5431
rect 15900 5175 15980 5177
rect 15900 5055 15912 5175
rect 15968 5055 15980 5175
rect 15900 5053 15980 5055
rect 16268 5175 16348 5177
rect 16268 5055 16280 5175
rect 16336 5055 16348 5175
rect 16268 5053 16348 5055
rect 16590 5175 16670 5177
rect 16590 5054 16602 5175
rect 16658 5054 16670 5175
rect 17386 5176 17466 5178
rect 17386 5056 17398 5176
rect 17454 5056 17466 5176
rect 17386 5054 17466 5056
rect 17754 5176 17834 5178
rect 17754 5056 17766 5176
rect 17822 5056 17834 5176
rect 17754 5054 17834 5056
rect 18076 5176 18156 5178
rect 18076 5055 18088 5176
rect 18144 5055 18156 5176
rect 15912 5045 15968 5053
rect 16280 5045 16336 5053
rect 16590 5052 16670 5054
rect 16602 5044 16658 5052
rect 17398 5046 17454 5054
rect 17766 5046 17822 5054
rect 18076 5053 18156 5055
rect 18088 5045 18144 5053
rect 16096 4877 16152 4885
rect 16464 4877 16520 4885
rect 17582 4878 17638 4886
rect 17950 4878 18006 4886
rect 16084 4875 16573 4877
rect 16084 4755 16096 4875
rect 16152 4755 16464 4875
rect 16520 4755 16573 4875
rect 16084 4753 16573 4755
rect 17570 4876 18059 4878
rect 17570 4756 17582 4876
rect 17638 4756 17950 4876
rect 18006 4756 18059 4876
rect 17570 4754 18059 4756
rect 16096 4745 16152 4753
rect 16464 4745 16573 4753
rect 17582 4746 17638 4754
rect 17950 4746 18059 4754
rect 15992 4679 16072 4689
rect 15992 4623 16004 4679
rect 16060 4623 16072 4679
rect 15992 4613 16072 4623
rect 16176 4679 16256 4689
rect 16176 4623 16188 4679
rect 16244 4623 16256 4679
rect 16176 4613 16256 4623
rect 16360 4679 16440 4689
rect 16360 4623 16372 4679
rect 16428 4623 16440 4679
rect 16360 4613 16440 4623
rect 16004 4531 16060 4613
rect 15992 4529 16072 4531
rect 15992 4473 16004 4529
rect 16060 4473 16072 4529
rect 15992 4471 16072 4473
rect 15320 4297 15390 4309
rect 15320 4241 15332 4297
rect 15388 4241 15390 4297
rect 15320 4229 15390 4241
rect 16004 4157 16060 4471
rect 16188 4415 16244 4613
rect 16176 4413 16256 4415
rect 16176 4357 16188 4413
rect 16244 4357 16256 4413
rect 16176 4355 16256 4357
rect 16188 4157 16244 4355
rect 16372 4299 16428 4613
rect 16505 4415 16573 4745
rect 17478 4680 17558 4690
rect 17478 4624 17490 4680
rect 17546 4624 17558 4680
rect 17478 4614 17558 4624
rect 17662 4680 17742 4690
rect 17662 4624 17674 4680
rect 17730 4624 17742 4680
rect 17662 4614 17742 4624
rect 17846 4680 17926 4690
rect 17846 4624 17858 4680
rect 17914 4624 17926 4680
rect 17846 4614 17926 4624
rect 17490 4532 17546 4614
rect 17478 4530 17558 4532
rect 17478 4474 17490 4530
rect 17546 4474 17558 4530
rect 17478 4472 17558 4474
rect 16505 4413 16585 4415
rect 16505 4357 16517 4413
rect 16573 4357 16585 4413
rect 16505 4355 16585 4357
rect 16772 4413 16842 4425
rect 16772 4357 16774 4413
rect 16830 4357 16842 4413
rect 16360 4297 16440 4299
rect 16360 4241 16372 4297
rect 16428 4241 16440 4297
rect 16360 4239 16440 4241
rect 16372 4157 16428 4239
rect 15992 4147 16072 4157
rect 15992 4091 16004 4147
rect 16060 4091 16072 4147
rect 15992 4081 16072 4091
rect 16176 4147 16256 4157
rect 16176 4091 16188 4147
rect 16244 4091 16256 4147
rect 16176 4081 16256 4091
rect 16360 4147 16440 4157
rect 16360 4091 16372 4147
rect 16428 4091 16440 4147
rect 16360 4081 16440 4091
rect 16505 4025 16573 4355
rect 16772 4347 16842 4357
rect 16464 4017 16573 4025
rect 16452 4015 16573 4017
rect 16452 3895 16464 4015
rect 16520 3895 16573 4015
rect 16452 3893 16573 3895
rect 16464 3885 16520 3893
rect 15767 3628 16663 3640
rect 15767 3572 15779 3628
rect 15835 3572 16597 3628
rect 16653 3572 16663 3628
rect 15767 3560 16663 3572
rect 16774 3403 16830 4347
rect 17490 4158 17546 4472
rect 17674 4416 17730 4614
rect 17662 4414 17742 4416
rect 17662 4358 17674 4414
rect 17730 4358 17742 4414
rect 17662 4356 17742 4358
rect 17674 4158 17730 4356
rect 17858 4300 17914 4614
rect 17991 4416 18059 4746
rect 18436 4424 18492 5658
rect 17991 4414 18071 4416
rect 17991 4358 18003 4414
rect 18059 4358 18071 4414
rect 17991 4356 18071 4358
rect 18434 4414 18504 4424
rect 18434 4358 18436 4414
rect 18492 4358 18584 4414
rect 17846 4298 17926 4300
rect 17846 4242 17858 4298
rect 17914 4242 17926 4298
rect 17846 4240 17926 4242
rect 17858 4158 17914 4240
rect 17478 4148 17558 4158
rect 17478 4092 17490 4148
rect 17546 4092 17558 4148
rect 17478 4082 17558 4092
rect 17662 4148 17742 4158
rect 17662 4092 17674 4148
rect 17730 4092 17742 4148
rect 17662 4082 17742 4092
rect 17846 4148 17926 4158
rect 17846 4092 17858 4148
rect 17914 4092 17926 4148
rect 17846 4082 17926 4092
rect 17991 4026 18059 4356
rect 18434 4346 18504 4358
rect 17950 4018 18059 4026
rect 17938 4016 18059 4018
rect 17938 3896 17950 4016
rect 18006 3896 18059 4016
rect 17938 3894 18059 3896
rect 17950 3886 18006 3894
rect 17253 3629 18149 3641
rect 17253 3573 17265 3629
rect 17321 3573 18083 3629
rect 18139 3573 18149 3629
rect 17253 3561 18149 3573
rect 16938 3510 17018 3520
rect 16938 3454 16950 3510
rect 17006 3454 17018 3510
rect 16938 3452 17018 3454
rect 16772 3400 16842 3403
rect 16772 3346 16774 3400
rect 16830 3346 16842 3400
rect 16772 3334 16842 3346
rect 15912 3293 16658 3305
rect 15912 3237 16280 3293
rect 16336 3237 16658 3293
rect 15912 3225 16658 3237
rect 15912 2972 15968 3225
rect 16280 2972 16336 3225
rect 16602 2972 16658 3225
rect 15900 2970 15980 2972
rect 15900 2850 15912 2970
rect 15968 2850 15980 2970
rect 15900 2848 15980 2850
rect 16268 2970 16348 2972
rect 16268 2850 16280 2970
rect 16336 2850 16348 2970
rect 16268 2848 16348 2850
rect 16590 2970 16670 2972
rect 16590 2849 16602 2970
rect 16658 2849 16670 2970
rect 15912 2840 15968 2848
rect 16280 2840 16336 2848
rect 16590 2847 16670 2849
rect 16602 2839 16658 2847
rect 16096 2672 16152 2680
rect 16464 2672 16520 2680
rect 16084 2670 16573 2672
rect 16084 2550 16096 2670
rect 16152 2550 16464 2670
rect 16520 2550 16573 2670
rect 16084 2548 16573 2550
rect 16096 2540 16152 2548
rect 16464 2540 16573 2548
rect 15992 2474 16072 2484
rect 15992 2418 16004 2474
rect 16060 2418 16072 2474
rect 15992 2408 16072 2418
rect 16176 2474 16256 2484
rect 16176 2418 16188 2474
rect 16244 2418 16256 2474
rect 16176 2408 16256 2418
rect 16360 2474 16440 2484
rect 16360 2418 16372 2474
rect 16428 2418 16440 2474
rect 16360 2408 16440 2418
rect 16004 2326 16060 2408
rect 15992 2324 16072 2326
rect 15992 2268 16004 2324
rect 16060 2268 16072 2324
rect 15992 2266 16072 2268
rect 15184 2208 15254 2222
rect 15184 2152 15196 2208
rect 15252 2152 15254 2208
rect 15184 2140 15254 2152
rect 14950 2092 15028 2103
rect 14558 2091 15028 2092
rect 14558 2037 14962 2091
rect 15016 2037 15028 2091
rect 14558 2036 15028 2037
rect 12986 1732 14158 1742
rect 12986 1676 12998 1732
rect 13054 1676 13886 1732
rect 13942 1676 14158 1732
rect 12986 1666 14158 1676
rect 14558 1732 14638 2036
rect 14950 2025 15028 2036
rect 14558 1676 14570 1732
rect 14626 1676 14638 1732
rect 14558 1666 14638 1676
rect 12916 1354 14708 1366
rect 12916 1214 12928 1354
rect 14696 1214 14708 1354
rect 15001 1305 15087 1317
rect 15196 1309 15252 2140
rect 16004 1952 16060 2266
rect 16188 2210 16244 2408
rect 16176 2208 16256 2210
rect 16176 2152 16188 2208
rect 16244 2152 16256 2208
rect 16176 2150 16256 2152
rect 16188 1952 16244 2150
rect 16372 2094 16428 2408
rect 16505 2210 16573 2540
rect 16950 2220 17006 3452
rect 18958 3347 19014 6562
rect 24656 6563 24668 6619
rect 24724 6563 24726 6619
rect 24656 6551 24726 6563
rect 24374 5717 24456 5729
rect 24374 5661 24388 5717
rect 24444 5661 24456 5717
rect 24374 5649 24456 5661
rect 19368 4311 19588 4321
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 23758 4311 24078 4321
rect 20230 3804 21402 3814
rect 20230 3564 20242 3804
rect 20298 3564 21334 3804
rect 21390 3564 21402 3804
rect 20230 3554 21402 3564
rect 19368 3501 19588 3511
rect 20324 3347 20402 3359
rect 18954 3291 20344 3347
rect 20400 3291 20402 3347
rect 18958 3290 19014 3291
rect 20324 3279 20402 3291
rect 21322 3269 21402 3554
rect 21802 3804 21882 3814
rect 21802 3564 21814 3804
rect 21870 3564 21882 3804
rect 21624 3269 21694 3281
rect 21322 3213 21636 3269
rect 21692 3213 21694 3269
rect 21144 3191 21214 3203
rect 18954 3135 21156 3191
rect 21212 3135 21214 3191
rect 16505 2208 16585 2210
rect 16505 2152 16517 2208
rect 16573 2152 16585 2208
rect 16505 2150 16585 2152
rect 16948 2208 17008 2220
rect 16948 2152 16950 2208
rect 17006 2152 17008 2208
rect 16360 2092 16440 2094
rect 16360 2036 16372 2092
rect 16428 2036 16440 2092
rect 16360 2034 16440 2036
rect 16372 1952 16428 2034
rect 15992 1942 16072 1952
rect 15992 1886 16004 1942
rect 16060 1886 16072 1942
rect 15992 1876 16072 1886
rect 16176 1942 16256 1952
rect 16176 1886 16188 1942
rect 16244 1886 16256 1942
rect 16176 1876 16256 1886
rect 16360 1942 16440 1952
rect 16360 1886 16372 1942
rect 16428 1886 16440 1942
rect 16360 1876 16440 1886
rect 16505 1820 16573 2150
rect 16948 2140 17008 2152
rect 19066 1849 19122 3135
rect 21144 3123 21214 3135
rect 20434 2909 20514 2919
rect 20434 2853 20446 2909
rect 20502 2853 20514 2909
rect 20434 2667 20514 2853
rect 20914 2909 20994 2919
rect 20914 2853 20926 2909
rect 20982 2853 20994 2909
rect 20914 2843 20994 2853
rect 21118 2909 21198 2919
rect 21118 2853 21130 2909
rect 21186 2853 21198 2909
rect 21118 2667 21198 2853
rect 21322 2909 21402 3213
rect 21624 3201 21694 3213
rect 21802 3269 21882 3564
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 23758 3501 24078 3511
rect 22388 3315 24180 3327
rect 21802 3213 22159 3269
rect 21322 2853 21334 2909
rect 21390 2853 21402 2909
rect 21322 2843 21402 2853
rect 21802 2909 21882 3213
rect 21802 2853 21814 2909
rect 21870 2853 21882 2909
rect 21802 2843 21882 2853
rect 20434 2595 21198 2667
rect 21328 2541 21952 2553
rect 21328 2401 21340 2541
rect 21940 2401 21952 2541
rect 19540 2384 19620 2394
rect 21328 2389 21952 2401
rect 19540 2144 19552 2384
rect 19608 2144 19620 2384
rect 22103 2171 22159 3213
rect 22388 3175 22400 3315
rect 24168 3175 24180 3315
rect 22388 3163 24180 3175
rect 22662 2912 23426 2922
rect 22662 2672 22674 2912
rect 22730 2672 23358 2912
rect 23414 2672 23426 2912
rect 22662 2662 23426 2672
rect 24030 2628 24110 2638
rect 23142 2578 23630 2588
rect 23142 2338 23154 2578
rect 23210 2338 23562 2578
rect 23618 2338 23630 2578
rect 23142 2328 23630 2338
rect 22552 2171 22648 2183
rect 19362 1849 19432 1861
rect 16464 1812 16573 1820
rect 16452 1810 16573 1812
rect 16452 1690 16464 1810
rect 16520 1690 16573 1810
rect 18554 1793 19374 1849
rect 19430 1793 19432 1849
rect 16452 1688 16573 1690
rect 16464 1680 16520 1688
rect 15767 1423 16665 1435
rect 15767 1367 15779 1423
rect 15835 1367 16597 1423
rect 16653 1367 16665 1423
rect 15767 1355 16665 1367
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 15194 1305 15254 1309
rect 15194 1249 15196 1305
rect 15252 1249 15254 1305
rect 15194 1237 15254 1249
rect 12916 1202 14708 1214
rect 12330 872 12687 928
rect 14286 1030 14606 1040
rect 11850 512 11862 568
rect 11918 512 11930 568
rect 11850 502 11930 512
rect 12330 568 12410 872
rect 12330 512 12342 568
rect 12398 512 12410 568
rect 12330 502 12410 512
rect 10962 254 11726 326
rect 14286 230 14296 1030
rect 14596 230 14606 1030
rect 14286 220 14606 230
rect 18559 -50 18615 1793
rect 19362 1781 19432 1793
rect 19540 1849 19620 2144
rect 21328 2141 21952 2153
rect 21328 2001 21340 2141
rect 21940 2001 21952 2141
rect 22103 2115 22572 2171
rect 22628 2115 22648 2171
rect 22552 2103 22648 2115
rect 23550 2093 23630 2328
rect 24030 2388 24042 2628
rect 24098 2388 24110 2628
rect 23852 2093 23922 2105
rect 23550 2037 23864 2093
rect 23920 2037 23922 2093
rect 23236 2015 23332 2025
rect 21328 1989 21952 2001
rect 22103 1959 23256 2015
rect 23312 1959 23332 2015
rect 19540 1793 19978 1849
rect 19540 1489 19620 1793
rect 19540 1433 19552 1489
rect 19608 1433 19620 1489
rect 19540 1423 19620 1433
rect 19922 1007 19978 1793
rect 20230 1464 21402 1474
rect 20230 1224 20242 1464
rect 20298 1224 21334 1464
rect 21390 1224 21402 1464
rect 20230 1214 21402 1224
rect 20324 1007 20402 1019
rect 19922 951 20344 1007
rect 20400 951 20402 1007
rect 20324 939 20402 951
rect 21322 929 21402 1214
rect 21802 1464 21882 1474
rect 21802 1224 21814 1464
rect 21870 1224 21882 1464
rect 21624 929 21694 941
rect 21322 873 21636 929
rect 21692 873 21694 929
rect 21144 851 21214 863
rect 18559 -180 18615 -170
rect 18954 795 21156 851
rect 21212 795 21214 851
rect 18954 -370 19010 795
rect 21144 783 21214 795
rect 20434 569 20514 579
rect 20434 513 20446 569
rect 20502 513 20514 569
rect 20434 327 20514 513
rect 20914 569 20994 579
rect 20914 513 20926 569
rect 20982 513 20994 569
rect 20914 503 20994 513
rect 21118 569 21198 579
rect 21118 513 21130 569
rect 21186 513 21198 569
rect 21118 327 21198 513
rect 21322 569 21402 873
rect 21624 861 21694 873
rect 21802 929 21882 1224
rect 22103 929 22159 1959
rect 23236 1949 23332 1959
rect 23550 1743 23630 2037
rect 23852 2025 23922 2037
rect 24030 2093 24110 2388
rect 24668 2223 24724 6551
rect 24804 4310 24860 8756
rect 25476 8568 25532 8882
rect 25660 8826 25716 9024
rect 25648 8824 25728 8826
rect 25648 8768 25660 8824
rect 25716 8768 25728 8824
rect 25648 8766 25728 8768
rect 25660 8568 25716 8766
rect 25844 8710 25900 9024
rect 25977 8826 26045 9156
rect 34936 9090 35016 9100
rect 34936 9034 34948 9090
rect 35004 9034 35016 9090
rect 34936 9024 35016 9034
rect 35120 9090 35200 9100
rect 35120 9034 35132 9090
rect 35188 9034 35200 9090
rect 35120 9024 35200 9034
rect 35304 9090 35384 9100
rect 35304 9034 35316 9090
rect 35372 9034 35384 9090
rect 35304 9024 35384 9034
rect 34046 8940 34134 8952
rect 34948 8942 35004 9024
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 34936 8940 35016 8942
rect 34936 8884 34948 8940
rect 35004 8884 35016 8940
rect 34936 8882 35016 8884
rect 25977 8824 26057 8826
rect 25977 8768 25989 8824
rect 26045 8768 26057 8824
rect 25977 8766 26057 8768
rect 26244 8824 26314 8836
rect 26244 8768 26246 8824
rect 26302 8768 26314 8824
rect 25832 8708 25912 8710
rect 25832 8652 25844 8708
rect 25900 8652 25912 8708
rect 25832 8650 25912 8652
rect 25844 8568 25900 8650
rect 25464 8558 25544 8568
rect 25464 8502 25476 8558
rect 25532 8502 25544 8558
rect 25464 8492 25544 8502
rect 25648 8558 25728 8568
rect 25648 8502 25660 8558
rect 25716 8502 25728 8558
rect 25648 8492 25728 8502
rect 25832 8558 25912 8568
rect 25832 8502 25844 8558
rect 25900 8502 25912 8558
rect 25832 8492 25912 8502
rect 25977 8436 26045 8766
rect 26244 8758 26314 8768
rect 34264 8824 34334 8836
rect 34264 8768 34276 8824
rect 34332 8768 34334 8824
rect 25936 8428 26045 8436
rect 25924 8426 26045 8428
rect 25924 8306 25936 8426
rect 25992 8306 26045 8426
rect 25924 8304 26045 8306
rect 25936 8296 25992 8304
rect 25239 8039 26137 8051
rect 25239 7983 25251 8039
rect 25307 7983 26069 8039
rect 26125 7983 26137 8039
rect 25239 7971 26137 7983
rect 26246 7814 26302 8758
rect 34264 8756 34334 8768
rect 26410 7921 26490 7931
rect 26410 7865 26422 7921
rect 26478 7865 26490 7921
rect 26410 7863 26490 7865
rect 26244 7811 26314 7814
rect 26244 7757 26246 7811
rect 26302 7757 26314 7811
rect 26244 7745 26314 7757
rect 25384 7704 26130 7716
rect 25384 7648 25752 7704
rect 25808 7648 26130 7704
rect 25384 7636 26130 7648
rect 25384 7383 25440 7636
rect 25752 7383 25808 7636
rect 26074 7383 26130 7636
rect 25372 7381 25452 7383
rect 25372 7261 25384 7381
rect 25440 7261 25452 7381
rect 25372 7259 25452 7261
rect 25740 7381 25820 7383
rect 25740 7261 25752 7381
rect 25808 7261 25820 7381
rect 25740 7259 25820 7261
rect 26062 7381 26142 7383
rect 26062 7260 26074 7381
rect 26130 7260 26142 7381
rect 25384 7251 25440 7259
rect 25752 7251 25808 7259
rect 26062 7258 26142 7260
rect 26074 7250 26130 7258
rect 25568 7083 25624 7091
rect 25936 7083 25992 7091
rect 25556 7081 26045 7083
rect 25556 6961 25568 7081
rect 25624 6961 25936 7081
rect 25992 6961 26045 7081
rect 25556 6959 26045 6961
rect 25568 6951 25624 6959
rect 25936 6951 26045 6959
rect 25464 6885 25544 6895
rect 25464 6829 25476 6885
rect 25532 6829 25544 6885
rect 25464 6819 25544 6829
rect 25648 6885 25728 6895
rect 25648 6829 25660 6885
rect 25716 6829 25728 6885
rect 25648 6819 25728 6829
rect 25832 6885 25912 6895
rect 25832 6829 25844 6885
rect 25900 6829 25912 6885
rect 25832 6819 25912 6829
rect 25476 6737 25532 6819
rect 25464 6735 25544 6737
rect 25464 6679 25476 6735
rect 25532 6679 25544 6735
rect 25464 6677 25544 6679
rect 25476 6363 25532 6677
rect 25660 6621 25716 6819
rect 25648 6619 25728 6621
rect 25648 6563 25660 6619
rect 25716 6563 25728 6619
rect 25648 6561 25728 6563
rect 25660 6363 25716 6561
rect 25844 6505 25900 6819
rect 25977 6621 26045 6951
rect 26422 6629 26478 7863
rect 26870 7704 27616 7716
rect 26870 7648 27238 7704
rect 27294 7648 27616 7704
rect 26870 7636 27616 7648
rect 26870 7383 26926 7636
rect 27238 7383 27294 7636
rect 27560 7383 27616 7636
rect 26858 7381 26938 7383
rect 26858 7261 26870 7381
rect 26926 7261 26938 7381
rect 26858 7259 26938 7261
rect 27226 7381 27306 7383
rect 27226 7261 27238 7381
rect 27294 7261 27306 7381
rect 27226 7259 27306 7261
rect 27548 7381 27628 7383
rect 27548 7260 27560 7381
rect 27616 7260 27628 7381
rect 26870 7251 26926 7259
rect 27238 7251 27294 7259
rect 27548 7258 27628 7260
rect 27560 7250 27616 7258
rect 27054 7083 27110 7091
rect 27422 7083 27478 7091
rect 27042 7081 27531 7083
rect 27042 6961 27054 7081
rect 27110 6961 27422 7081
rect 27478 6961 27531 7081
rect 27042 6959 27531 6961
rect 27054 6951 27110 6959
rect 27422 6951 27531 6959
rect 26950 6885 27030 6895
rect 26950 6829 26962 6885
rect 27018 6829 27030 6885
rect 26950 6819 27030 6829
rect 27134 6885 27214 6895
rect 27134 6829 27146 6885
rect 27202 6829 27214 6885
rect 27134 6819 27214 6829
rect 27318 6885 27398 6895
rect 27318 6829 27330 6885
rect 27386 6829 27398 6885
rect 27318 6819 27398 6829
rect 26962 6737 27018 6819
rect 26950 6735 27030 6737
rect 26950 6679 26962 6735
rect 27018 6679 27030 6735
rect 26950 6677 27030 6679
rect 25977 6619 26057 6621
rect 25977 6563 25989 6619
rect 26045 6563 26057 6619
rect 25977 6561 26057 6563
rect 26420 6619 26480 6629
rect 26420 6563 26422 6619
rect 26478 6563 26480 6619
rect 25832 6503 25912 6505
rect 25832 6447 25844 6503
rect 25900 6447 25912 6503
rect 25832 6445 25912 6447
rect 25844 6363 25900 6445
rect 25464 6353 25544 6363
rect 25464 6297 25476 6353
rect 25532 6297 25544 6353
rect 25464 6287 25544 6297
rect 25648 6353 25728 6363
rect 25648 6297 25660 6353
rect 25716 6297 25728 6353
rect 25648 6287 25728 6297
rect 25832 6353 25912 6363
rect 25832 6297 25844 6353
rect 25900 6297 25912 6353
rect 25832 6287 25912 6297
rect 25977 6231 26045 6561
rect 26420 6551 26480 6563
rect 25936 6223 26045 6231
rect 25924 6221 26045 6223
rect 25924 6101 25936 6221
rect 25992 6101 26045 6221
rect 25924 6099 26045 6101
rect 25936 6091 25992 6099
rect 25239 5834 26135 5846
rect 25239 5778 25251 5834
rect 25307 5778 26069 5834
rect 26125 5778 26135 5834
rect 25239 5766 26135 5778
rect 26422 5608 26478 6551
rect 26962 6363 27018 6677
rect 27146 6621 27202 6819
rect 27134 6619 27214 6621
rect 27134 6563 27146 6619
rect 27202 6563 27214 6619
rect 27134 6561 27214 6563
rect 27146 6363 27202 6561
rect 27330 6505 27386 6819
rect 27463 6621 27531 6951
rect 27463 6619 27543 6621
rect 27463 6563 27475 6619
rect 27531 6563 27543 6619
rect 27463 6561 27543 6563
rect 27730 6619 27800 6631
rect 34128 6619 34198 6633
rect 27730 6563 27732 6619
rect 27788 6563 28486 6619
rect 27318 6503 27398 6505
rect 27318 6447 27330 6503
rect 27386 6447 27398 6503
rect 27318 6445 27398 6447
rect 27330 6363 27386 6445
rect 26950 6353 27030 6363
rect 26950 6297 26962 6353
rect 27018 6297 27030 6353
rect 26950 6287 27030 6297
rect 27134 6353 27214 6363
rect 27134 6297 27146 6353
rect 27202 6297 27214 6353
rect 27134 6287 27214 6297
rect 27318 6353 27398 6363
rect 27318 6297 27330 6353
rect 27386 6297 27398 6353
rect 27318 6287 27398 6297
rect 27463 6231 27531 6561
rect 27730 6553 27800 6563
rect 27422 6223 27531 6231
rect 27410 6221 27531 6223
rect 27410 6101 27422 6221
rect 27478 6101 27531 6221
rect 27410 6099 27531 6101
rect 27422 6091 27478 6099
rect 26725 5834 27621 5846
rect 26725 5778 26737 5834
rect 26793 5778 27555 5834
rect 27611 5778 27621 5834
rect 26725 5766 27621 5778
rect 27732 5609 27788 6553
rect 27896 5717 27976 5727
rect 27896 5661 27908 5717
rect 27964 5661 27976 5717
rect 27896 5659 27976 5661
rect 26420 5606 26490 5608
rect 26420 5550 26422 5606
rect 26478 5550 26490 5606
rect 26420 5538 26490 5550
rect 27720 5607 27800 5609
rect 27720 5551 27732 5607
rect 27788 5551 27800 5607
rect 27720 5539 27800 5551
rect 25384 5499 26130 5511
rect 25384 5443 25752 5499
rect 25808 5443 26130 5499
rect 25384 5431 26130 5443
rect 25384 5178 25440 5431
rect 25752 5178 25808 5431
rect 26074 5178 26130 5431
rect 26870 5500 27616 5512
rect 26870 5444 27238 5500
rect 27294 5444 27616 5500
rect 26870 5432 27616 5444
rect 26870 5179 26926 5432
rect 27238 5179 27294 5432
rect 27560 5179 27616 5432
rect 25372 5176 25452 5178
rect 25372 5056 25384 5176
rect 25440 5056 25452 5176
rect 25372 5054 25452 5056
rect 25740 5176 25820 5178
rect 25740 5056 25752 5176
rect 25808 5056 25820 5176
rect 25740 5054 25820 5056
rect 26062 5176 26142 5178
rect 26062 5055 26074 5176
rect 26130 5055 26142 5176
rect 26858 5177 26938 5179
rect 26858 5057 26870 5177
rect 26926 5057 26938 5177
rect 26858 5055 26938 5057
rect 27226 5177 27306 5179
rect 27226 5057 27238 5177
rect 27294 5057 27306 5177
rect 27226 5055 27306 5057
rect 27548 5177 27628 5179
rect 27548 5056 27560 5177
rect 27616 5056 27628 5177
rect 25384 5046 25440 5054
rect 25752 5046 25808 5054
rect 26062 5053 26142 5055
rect 26074 5045 26130 5053
rect 26870 5047 26926 5055
rect 27238 5047 27294 5055
rect 27548 5054 27628 5056
rect 27560 5046 27616 5054
rect 25568 4878 25624 4886
rect 25936 4878 25992 4886
rect 27054 4879 27110 4887
rect 27422 4879 27478 4887
rect 25556 4876 26045 4878
rect 25556 4756 25568 4876
rect 25624 4756 25936 4876
rect 25992 4756 26045 4876
rect 25556 4754 26045 4756
rect 27042 4877 27531 4879
rect 27042 4757 27054 4877
rect 27110 4757 27422 4877
rect 27478 4757 27531 4877
rect 27042 4755 27531 4757
rect 25568 4746 25624 4754
rect 25936 4746 26045 4754
rect 27054 4747 27110 4755
rect 27422 4747 27531 4755
rect 25464 4680 25544 4690
rect 25464 4624 25476 4680
rect 25532 4624 25544 4680
rect 25464 4614 25544 4624
rect 25648 4680 25728 4690
rect 25648 4624 25660 4680
rect 25716 4624 25728 4680
rect 25648 4614 25728 4624
rect 25832 4680 25912 4690
rect 25832 4624 25844 4680
rect 25900 4624 25912 4680
rect 25832 4614 25912 4624
rect 25476 4532 25532 4614
rect 25464 4530 25544 4532
rect 25464 4474 25476 4530
rect 25532 4474 25544 4530
rect 25464 4472 25544 4474
rect 24792 4298 24862 4310
rect 24792 4242 24804 4298
rect 24860 4242 24862 4298
rect 24792 4230 24862 4242
rect 25476 4158 25532 4472
rect 25660 4416 25716 4614
rect 25648 4414 25728 4416
rect 25648 4358 25660 4414
rect 25716 4358 25728 4414
rect 25648 4356 25728 4358
rect 25660 4158 25716 4356
rect 25844 4300 25900 4614
rect 25977 4416 26045 4746
rect 26950 4681 27030 4691
rect 26950 4625 26962 4681
rect 27018 4625 27030 4681
rect 26950 4615 27030 4625
rect 27134 4681 27214 4691
rect 27134 4625 27146 4681
rect 27202 4625 27214 4681
rect 27134 4615 27214 4625
rect 27318 4681 27398 4691
rect 27318 4625 27330 4681
rect 27386 4625 27398 4681
rect 27318 4615 27398 4625
rect 26962 4533 27018 4615
rect 26950 4531 27030 4533
rect 26950 4475 26962 4531
rect 27018 4475 27030 4531
rect 26950 4473 27030 4475
rect 25977 4414 26057 4416
rect 25977 4358 25989 4414
rect 26045 4358 26057 4414
rect 25977 4356 26057 4358
rect 26244 4414 26314 4426
rect 26244 4358 26246 4414
rect 26302 4358 26314 4414
rect 25832 4298 25912 4300
rect 25832 4242 25844 4298
rect 25900 4242 25912 4298
rect 25832 4240 25912 4242
rect 25844 4158 25900 4240
rect 25464 4148 25544 4158
rect 25464 4092 25476 4148
rect 25532 4092 25544 4148
rect 25464 4082 25544 4092
rect 25648 4148 25728 4158
rect 25648 4092 25660 4148
rect 25716 4092 25728 4148
rect 25648 4082 25728 4092
rect 25832 4148 25912 4158
rect 25832 4092 25844 4148
rect 25900 4092 25912 4148
rect 25832 4082 25912 4092
rect 25977 4026 26045 4356
rect 26244 4348 26314 4358
rect 25936 4018 26045 4026
rect 25924 4016 26045 4018
rect 25924 3896 25936 4016
rect 25992 3896 26045 4016
rect 25924 3894 26045 3896
rect 25936 3886 25992 3894
rect 25239 3629 26135 3641
rect 25239 3573 25251 3629
rect 25307 3573 26069 3629
rect 26125 3573 26135 3629
rect 25239 3561 26135 3573
rect 26246 3404 26302 4348
rect 26962 4159 27018 4473
rect 27146 4417 27202 4615
rect 27134 4415 27214 4417
rect 27134 4359 27146 4415
rect 27202 4359 27214 4415
rect 27134 4357 27214 4359
rect 27146 4159 27202 4357
rect 27330 4301 27386 4615
rect 27463 4417 27531 4747
rect 27908 4425 27964 5659
rect 27463 4415 27543 4417
rect 27463 4359 27475 4415
rect 27531 4359 27543 4415
rect 27463 4357 27543 4359
rect 27906 4415 27976 4425
rect 27906 4359 27908 4415
rect 27964 4359 28056 4415
rect 27318 4299 27398 4301
rect 27318 4243 27330 4299
rect 27386 4243 27398 4299
rect 27318 4241 27398 4243
rect 27330 4159 27386 4241
rect 26950 4149 27030 4159
rect 26950 4093 26962 4149
rect 27018 4093 27030 4149
rect 26950 4083 27030 4093
rect 27134 4149 27214 4159
rect 27134 4093 27146 4149
rect 27202 4093 27214 4149
rect 27134 4083 27214 4093
rect 27318 4149 27398 4159
rect 27318 4093 27330 4149
rect 27386 4093 27398 4149
rect 27318 4083 27398 4093
rect 27463 4027 27531 4357
rect 27906 4347 27976 4359
rect 27422 4019 27531 4027
rect 27410 4017 27531 4019
rect 27410 3897 27422 4017
rect 27478 3897 27531 4017
rect 27410 3895 27531 3897
rect 27422 3887 27478 3895
rect 26725 3630 27621 3642
rect 26725 3574 26737 3630
rect 26793 3574 27555 3630
rect 27611 3574 27621 3630
rect 26725 3562 27621 3574
rect 26410 3511 26490 3521
rect 26410 3455 26422 3511
rect 26478 3455 26490 3511
rect 26410 3453 26490 3455
rect 26244 3401 26314 3404
rect 26244 3347 26246 3401
rect 26302 3347 26314 3401
rect 26244 3335 26314 3347
rect 25384 3294 26130 3306
rect 25384 3238 25752 3294
rect 25808 3238 26130 3294
rect 25384 3226 26130 3238
rect 25384 2973 25440 3226
rect 25752 2973 25808 3226
rect 26074 2973 26130 3226
rect 25372 2971 25452 2973
rect 25372 2851 25384 2971
rect 25440 2851 25452 2971
rect 25372 2849 25452 2851
rect 25740 2971 25820 2973
rect 25740 2851 25752 2971
rect 25808 2851 25820 2971
rect 25740 2849 25820 2851
rect 26062 2971 26142 2973
rect 26062 2850 26074 2971
rect 26130 2850 26142 2971
rect 25384 2841 25440 2849
rect 25752 2841 25808 2849
rect 26062 2848 26142 2850
rect 26074 2840 26130 2848
rect 25568 2673 25624 2681
rect 25936 2673 25992 2681
rect 25556 2671 26045 2673
rect 25556 2551 25568 2671
rect 25624 2551 25936 2671
rect 25992 2551 26045 2671
rect 25556 2549 26045 2551
rect 25568 2541 25624 2549
rect 25936 2541 26045 2549
rect 25464 2475 25544 2485
rect 25464 2419 25476 2475
rect 25532 2419 25544 2475
rect 25464 2409 25544 2419
rect 25648 2475 25728 2485
rect 25648 2419 25660 2475
rect 25716 2419 25728 2475
rect 25648 2409 25728 2419
rect 25832 2475 25912 2485
rect 25832 2419 25844 2475
rect 25900 2419 25912 2475
rect 25832 2409 25912 2419
rect 25476 2327 25532 2409
rect 25464 2325 25544 2327
rect 25464 2269 25476 2325
rect 25532 2269 25544 2325
rect 25464 2267 25544 2269
rect 24656 2209 24726 2223
rect 24656 2153 24668 2209
rect 24724 2153 24726 2209
rect 24656 2141 24726 2153
rect 24422 2093 24500 2104
rect 24030 2092 24500 2093
rect 24030 2038 24434 2092
rect 24488 2038 24500 2092
rect 24030 2037 24500 2038
rect 22458 1733 23630 1743
rect 22458 1677 22470 1733
rect 22526 1677 23358 1733
rect 23414 1677 23630 1733
rect 22458 1667 23630 1677
rect 24030 1733 24110 2037
rect 24422 2026 24500 2037
rect 24030 1677 24042 1733
rect 24098 1677 24110 1733
rect 24030 1667 24110 1677
rect 22388 1355 24180 1367
rect 22388 1215 22400 1355
rect 24168 1215 24180 1355
rect 24473 1306 24559 1318
rect 24668 1310 24724 2141
rect 25476 1953 25532 2267
rect 25660 2211 25716 2409
rect 25648 2209 25728 2211
rect 25648 2153 25660 2209
rect 25716 2153 25728 2209
rect 25648 2151 25728 2153
rect 25660 1953 25716 2151
rect 25844 2095 25900 2409
rect 25977 2211 26045 2541
rect 26422 2221 26478 3453
rect 28430 3347 28486 6563
rect 34128 6563 34140 6619
rect 34196 6563 34198 6619
rect 34128 6551 34198 6563
rect 33846 5717 33928 5729
rect 33846 5661 33860 5717
rect 33916 5661 33928 5717
rect 33846 5649 33928 5661
rect 28840 4311 29060 4321
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 33230 4311 33550 4321
rect 29702 3804 30874 3814
rect 29702 3564 29714 3804
rect 29770 3564 30806 3804
rect 30862 3564 30874 3804
rect 29702 3554 30874 3564
rect 28840 3501 29060 3511
rect 29796 3347 29874 3359
rect 28426 3291 29816 3347
rect 29872 3291 29874 3347
rect 29796 3279 29874 3291
rect 30794 3269 30874 3554
rect 31274 3804 31354 3814
rect 31274 3564 31286 3804
rect 31342 3564 31354 3804
rect 31096 3269 31166 3281
rect 30794 3213 31108 3269
rect 31164 3213 31166 3269
rect 30616 3191 30686 3203
rect 28426 3135 30628 3191
rect 30684 3135 30686 3191
rect 25977 2209 26057 2211
rect 25977 2153 25989 2209
rect 26045 2153 26057 2209
rect 25977 2151 26057 2153
rect 26420 2209 26480 2221
rect 26420 2153 26422 2209
rect 26478 2153 26480 2209
rect 25832 2093 25912 2095
rect 25832 2037 25844 2093
rect 25900 2037 25912 2093
rect 25832 2035 25912 2037
rect 25844 1953 25900 2035
rect 25464 1943 25544 1953
rect 25464 1887 25476 1943
rect 25532 1887 25544 1943
rect 25464 1877 25544 1887
rect 25648 1943 25728 1953
rect 25648 1887 25660 1943
rect 25716 1887 25728 1943
rect 25648 1877 25728 1887
rect 25832 1943 25912 1953
rect 25832 1887 25844 1943
rect 25900 1887 25912 1943
rect 25832 1877 25912 1887
rect 25977 1821 26045 2151
rect 26420 2141 26480 2153
rect 28538 1850 28594 3135
rect 30616 3123 30686 3135
rect 29906 2909 29986 2919
rect 29906 2853 29918 2909
rect 29974 2853 29986 2909
rect 29906 2667 29986 2853
rect 30386 2909 30466 2919
rect 30386 2853 30398 2909
rect 30454 2853 30466 2909
rect 30386 2843 30466 2853
rect 30590 2909 30670 2919
rect 30590 2853 30602 2909
rect 30658 2853 30670 2909
rect 30590 2667 30670 2853
rect 30794 2909 30874 3213
rect 31096 3201 31166 3213
rect 31274 3269 31354 3564
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 33230 3501 33550 3511
rect 31860 3315 33652 3327
rect 31274 3213 31631 3269
rect 30794 2853 30806 2909
rect 30862 2853 30874 2909
rect 30794 2843 30874 2853
rect 31274 2909 31354 3213
rect 31274 2853 31286 2909
rect 31342 2853 31354 2909
rect 31274 2843 31354 2853
rect 29906 2595 30670 2667
rect 30800 2541 31424 2553
rect 30800 2401 30812 2541
rect 31412 2401 31424 2541
rect 29012 2384 29092 2394
rect 30800 2389 31424 2401
rect 29012 2144 29024 2384
rect 29080 2144 29092 2384
rect 31575 2171 31631 3213
rect 31860 3175 31872 3315
rect 33640 3175 33652 3315
rect 31860 3163 33652 3175
rect 32134 2912 32898 2922
rect 32134 2672 32146 2912
rect 32202 2672 32830 2912
rect 32886 2672 32898 2912
rect 32134 2662 32898 2672
rect 33502 2628 33582 2638
rect 32614 2578 33102 2588
rect 32614 2338 32626 2578
rect 32682 2338 33034 2578
rect 33090 2338 33102 2578
rect 32614 2328 33102 2338
rect 32024 2171 32120 2183
rect 25936 1813 26045 1821
rect 25924 1811 26045 1813
rect 25924 1691 25936 1811
rect 25992 1691 26045 1811
rect 28026 1849 28594 1850
rect 28834 1849 28904 1861
rect 28026 1794 28846 1849
rect 25924 1689 26045 1691
rect 25936 1681 25992 1689
rect 25239 1424 26137 1436
rect 25239 1368 25251 1424
rect 25307 1368 26069 1424
rect 26125 1368 26137 1424
rect 25239 1356 26137 1368
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 24666 1306 24726 1310
rect 24666 1250 24668 1306
rect 24724 1250 24726 1306
rect 24666 1238 24726 1250
rect 22388 1203 24180 1215
rect 21802 873 22159 929
rect 23758 1031 24078 1041
rect 21322 513 21334 569
rect 21390 513 21402 569
rect 21322 503 21402 513
rect 21802 569 21882 873
rect 21802 513 21814 569
rect 21870 513 21882 569
rect 21802 503 21882 513
rect 20434 255 21198 327
rect 23758 231 23768 1031
rect 24068 231 24078 1031
rect 23758 221 24078 231
rect 28031 -49 28087 1794
rect 28538 1793 28846 1794
rect 28902 1793 28904 1849
rect 28834 1781 28904 1793
rect 29012 1849 29092 2144
rect 30800 2141 31424 2153
rect 30800 2001 30812 2141
rect 31412 2001 31424 2141
rect 31575 2115 32044 2171
rect 32100 2115 32120 2171
rect 32024 2103 32120 2115
rect 33022 2093 33102 2328
rect 33502 2388 33514 2628
rect 33570 2388 33582 2628
rect 33324 2093 33394 2105
rect 33022 2037 33336 2093
rect 33392 2037 33394 2093
rect 32708 2015 32804 2025
rect 30800 1989 31424 2001
rect 31575 1959 32728 2015
rect 32784 1959 32804 2015
rect 29012 1793 29450 1849
rect 29012 1489 29092 1793
rect 29012 1433 29024 1489
rect 29080 1433 29092 1489
rect 29012 1423 29092 1433
rect 29394 1007 29450 1793
rect 29702 1464 30874 1474
rect 29702 1224 29714 1464
rect 29770 1224 30806 1464
rect 30862 1224 30874 1464
rect 29702 1214 30874 1224
rect 29796 1007 29874 1019
rect 29394 951 29816 1007
rect 29872 951 29874 1007
rect 29796 939 29874 951
rect 30794 929 30874 1214
rect 31274 1464 31354 1474
rect 31274 1224 31286 1464
rect 31342 1224 31354 1464
rect 31096 929 31166 941
rect 30794 873 31108 929
rect 31164 873 31166 929
rect 30616 851 30686 863
rect 28031 -179 28087 -169
rect 28426 795 30628 851
rect 30684 795 30686 851
rect 28426 -369 28482 795
rect 30616 783 30686 795
rect 29906 569 29986 579
rect 29906 513 29918 569
rect 29974 513 29986 569
rect 29906 327 29986 513
rect 30386 569 30466 579
rect 30386 513 30398 569
rect 30454 513 30466 569
rect 30386 503 30466 513
rect 30590 569 30670 579
rect 30590 513 30602 569
rect 30658 513 30670 569
rect 30590 327 30670 513
rect 30794 569 30874 873
rect 31096 861 31166 873
rect 31274 929 31354 1224
rect 31575 929 31631 1959
rect 32708 1949 32804 1959
rect 33022 1743 33102 2037
rect 33324 2025 33394 2037
rect 33502 2093 33582 2388
rect 34140 2223 34196 6551
rect 34276 4310 34332 8756
rect 34948 8568 35004 8882
rect 35132 8826 35188 9024
rect 35120 8824 35200 8826
rect 35120 8768 35132 8824
rect 35188 8768 35200 8824
rect 35120 8766 35200 8768
rect 35132 8568 35188 8766
rect 35316 8710 35372 9024
rect 35449 8826 35517 9156
rect 44408 9090 44488 9100
rect 44408 9034 44420 9090
rect 44476 9034 44488 9090
rect 44408 9024 44488 9034
rect 44592 9090 44672 9100
rect 44592 9034 44604 9090
rect 44660 9034 44672 9090
rect 44592 9024 44672 9034
rect 44776 9090 44856 9100
rect 44776 9034 44788 9090
rect 44844 9034 44856 9090
rect 44776 9024 44856 9034
rect 43518 8940 43606 8952
rect 44420 8942 44476 9024
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 44408 8940 44488 8942
rect 44408 8884 44420 8940
rect 44476 8884 44488 8940
rect 44408 8882 44488 8884
rect 35449 8824 35529 8826
rect 35449 8768 35461 8824
rect 35517 8768 35529 8824
rect 35449 8766 35529 8768
rect 35716 8824 35786 8836
rect 35716 8768 35718 8824
rect 35774 8768 35786 8824
rect 35304 8708 35384 8710
rect 35304 8652 35316 8708
rect 35372 8652 35384 8708
rect 35304 8650 35384 8652
rect 35316 8568 35372 8650
rect 34936 8558 35016 8568
rect 34936 8502 34948 8558
rect 35004 8502 35016 8558
rect 34936 8492 35016 8502
rect 35120 8558 35200 8568
rect 35120 8502 35132 8558
rect 35188 8502 35200 8558
rect 35120 8492 35200 8502
rect 35304 8558 35384 8568
rect 35304 8502 35316 8558
rect 35372 8502 35384 8558
rect 35304 8492 35384 8502
rect 35449 8436 35517 8766
rect 35716 8758 35786 8768
rect 43736 8824 43806 8836
rect 43736 8768 43748 8824
rect 43804 8768 43806 8824
rect 35408 8428 35517 8436
rect 35396 8426 35517 8428
rect 35396 8306 35408 8426
rect 35464 8306 35517 8426
rect 35396 8304 35517 8306
rect 35408 8296 35464 8304
rect 34711 8039 35609 8051
rect 34711 7983 34723 8039
rect 34779 7983 35541 8039
rect 35597 7983 35609 8039
rect 34711 7971 35609 7983
rect 35718 7814 35774 8758
rect 43736 8756 43806 8768
rect 35882 7921 35962 7931
rect 35882 7865 35894 7921
rect 35950 7865 35962 7921
rect 35882 7863 35962 7865
rect 35716 7811 35786 7814
rect 35716 7757 35718 7811
rect 35774 7757 35786 7811
rect 35716 7745 35786 7757
rect 34856 7704 35602 7716
rect 34856 7648 35224 7704
rect 35280 7648 35602 7704
rect 34856 7636 35602 7648
rect 34856 7383 34912 7636
rect 35224 7383 35280 7636
rect 35546 7383 35602 7636
rect 34844 7381 34924 7383
rect 34844 7261 34856 7381
rect 34912 7261 34924 7381
rect 34844 7259 34924 7261
rect 35212 7381 35292 7383
rect 35212 7261 35224 7381
rect 35280 7261 35292 7381
rect 35212 7259 35292 7261
rect 35534 7381 35614 7383
rect 35534 7260 35546 7381
rect 35602 7260 35614 7381
rect 34856 7251 34912 7259
rect 35224 7251 35280 7259
rect 35534 7258 35614 7260
rect 35546 7250 35602 7258
rect 35040 7083 35096 7091
rect 35408 7083 35464 7091
rect 35028 7081 35517 7083
rect 35028 6961 35040 7081
rect 35096 6961 35408 7081
rect 35464 6961 35517 7081
rect 35028 6959 35517 6961
rect 35040 6951 35096 6959
rect 35408 6951 35517 6959
rect 34936 6885 35016 6895
rect 34936 6829 34948 6885
rect 35004 6829 35016 6885
rect 34936 6819 35016 6829
rect 35120 6885 35200 6895
rect 35120 6829 35132 6885
rect 35188 6829 35200 6885
rect 35120 6819 35200 6829
rect 35304 6885 35384 6895
rect 35304 6829 35316 6885
rect 35372 6829 35384 6885
rect 35304 6819 35384 6829
rect 34948 6737 35004 6819
rect 34936 6735 35016 6737
rect 34936 6679 34948 6735
rect 35004 6679 35016 6735
rect 34936 6677 35016 6679
rect 34948 6363 35004 6677
rect 35132 6621 35188 6819
rect 35120 6619 35200 6621
rect 35120 6563 35132 6619
rect 35188 6563 35200 6619
rect 35120 6561 35200 6563
rect 35132 6363 35188 6561
rect 35316 6505 35372 6819
rect 35449 6621 35517 6951
rect 35894 6629 35950 7863
rect 36342 7704 37088 7716
rect 36342 7648 36710 7704
rect 36766 7648 37088 7704
rect 36342 7636 37088 7648
rect 36342 7383 36398 7636
rect 36710 7383 36766 7636
rect 37032 7383 37088 7636
rect 36330 7381 36410 7383
rect 36330 7261 36342 7381
rect 36398 7261 36410 7381
rect 36330 7259 36410 7261
rect 36698 7381 36778 7383
rect 36698 7261 36710 7381
rect 36766 7261 36778 7381
rect 36698 7259 36778 7261
rect 37020 7381 37100 7383
rect 37020 7260 37032 7381
rect 37088 7260 37100 7381
rect 36342 7251 36398 7259
rect 36710 7251 36766 7259
rect 37020 7258 37100 7260
rect 37032 7250 37088 7258
rect 36526 7083 36582 7091
rect 36894 7083 36950 7091
rect 36514 7081 37003 7083
rect 36514 6961 36526 7081
rect 36582 6961 36894 7081
rect 36950 6961 37003 7081
rect 36514 6959 37003 6961
rect 36526 6951 36582 6959
rect 36894 6951 37003 6959
rect 36422 6885 36502 6895
rect 36422 6829 36434 6885
rect 36490 6829 36502 6885
rect 36422 6819 36502 6829
rect 36606 6885 36686 6895
rect 36606 6829 36618 6885
rect 36674 6829 36686 6885
rect 36606 6819 36686 6829
rect 36790 6885 36870 6895
rect 36790 6829 36802 6885
rect 36858 6829 36870 6885
rect 36790 6819 36870 6829
rect 36434 6737 36490 6819
rect 36422 6735 36502 6737
rect 36422 6679 36434 6735
rect 36490 6679 36502 6735
rect 36422 6677 36502 6679
rect 35449 6619 35529 6621
rect 35449 6563 35461 6619
rect 35517 6563 35529 6619
rect 35449 6561 35529 6563
rect 35892 6619 35952 6629
rect 35892 6563 35894 6619
rect 35950 6563 35952 6619
rect 35304 6503 35384 6505
rect 35304 6447 35316 6503
rect 35372 6447 35384 6503
rect 35304 6445 35384 6447
rect 35316 6363 35372 6445
rect 34936 6353 35016 6363
rect 34936 6297 34948 6353
rect 35004 6297 35016 6353
rect 34936 6287 35016 6297
rect 35120 6353 35200 6363
rect 35120 6297 35132 6353
rect 35188 6297 35200 6353
rect 35120 6287 35200 6297
rect 35304 6353 35384 6363
rect 35304 6297 35316 6353
rect 35372 6297 35384 6353
rect 35304 6287 35384 6297
rect 35449 6231 35517 6561
rect 35892 6551 35952 6563
rect 35408 6223 35517 6231
rect 35396 6221 35517 6223
rect 35396 6101 35408 6221
rect 35464 6101 35517 6221
rect 35396 6099 35517 6101
rect 35408 6091 35464 6099
rect 34711 5834 35607 5846
rect 34711 5778 34723 5834
rect 34779 5778 35541 5834
rect 35597 5778 35607 5834
rect 34711 5766 35607 5778
rect 35894 5608 35950 6551
rect 36434 6363 36490 6677
rect 36618 6621 36674 6819
rect 36606 6619 36686 6621
rect 36606 6563 36618 6619
rect 36674 6563 36686 6619
rect 36606 6561 36686 6563
rect 36618 6363 36674 6561
rect 36802 6505 36858 6819
rect 36935 6621 37003 6951
rect 36935 6619 37015 6621
rect 36935 6563 36947 6619
rect 37003 6563 37015 6619
rect 36935 6561 37015 6563
rect 37202 6619 37272 6631
rect 43600 6619 43670 6633
rect 37202 6563 37204 6619
rect 37260 6563 37958 6619
rect 36790 6503 36870 6505
rect 36790 6447 36802 6503
rect 36858 6447 36870 6503
rect 36790 6445 36870 6447
rect 36802 6363 36858 6445
rect 36422 6353 36502 6363
rect 36422 6297 36434 6353
rect 36490 6297 36502 6353
rect 36422 6287 36502 6297
rect 36606 6353 36686 6363
rect 36606 6297 36618 6353
rect 36674 6297 36686 6353
rect 36606 6287 36686 6297
rect 36790 6353 36870 6363
rect 36790 6297 36802 6353
rect 36858 6297 36870 6353
rect 36790 6287 36870 6297
rect 36935 6231 37003 6561
rect 37202 6553 37272 6563
rect 36894 6223 37003 6231
rect 36882 6221 37003 6223
rect 36882 6101 36894 6221
rect 36950 6101 37003 6221
rect 36882 6099 37003 6101
rect 36894 6091 36950 6099
rect 36197 5834 37093 5846
rect 36197 5778 36209 5834
rect 36265 5778 37027 5834
rect 37083 5778 37093 5834
rect 36197 5766 37093 5778
rect 37204 5609 37260 6553
rect 37368 5717 37448 5727
rect 37368 5661 37380 5717
rect 37436 5661 37448 5717
rect 37368 5659 37448 5661
rect 35892 5606 35962 5608
rect 35892 5550 35894 5606
rect 35950 5550 35962 5606
rect 35892 5538 35962 5550
rect 37192 5607 37272 5609
rect 37192 5551 37204 5607
rect 37260 5551 37272 5607
rect 37192 5539 37272 5551
rect 34856 5499 35602 5511
rect 34856 5443 35224 5499
rect 35280 5443 35602 5499
rect 34856 5431 35602 5443
rect 34856 5178 34912 5431
rect 35224 5178 35280 5431
rect 35546 5178 35602 5431
rect 36342 5500 37088 5512
rect 36342 5444 36710 5500
rect 36766 5444 37088 5500
rect 36342 5432 37088 5444
rect 36342 5179 36398 5432
rect 36710 5179 36766 5432
rect 37032 5179 37088 5432
rect 34844 5176 34924 5178
rect 34844 5056 34856 5176
rect 34912 5056 34924 5176
rect 34844 5054 34924 5056
rect 35212 5176 35292 5178
rect 35212 5056 35224 5176
rect 35280 5056 35292 5176
rect 35212 5054 35292 5056
rect 35534 5176 35614 5178
rect 35534 5055 35546 5176
rect 35602 5055 35614 5176
rect 36330 5177 36410 5179
rect 36330 5057 36342 5177
rect 36398 5057 36410 5177
rect 36330 5055 36410 5057
rect 36698 5177 36778 5179
rect 36698 5057 36710 5177
rect 36766 5057 36778 5177
rect 36698 5055 36778 5057
rect 37020 5177 37100 5179
rect 37020 5056 37032 5177
rect 37088 5056 37100 5177
rect 34856 5046 34912 5054
rect 35224 5046 35280 5054
rect 35534 5053 35614 5055
rect 35546 5045 35602 5053
rect 36342 5047 36398 5055
rect 36710 5047 36766 5055
rect 37020 5054 37100 5056
rect 37032 5046 37088 5054
rect 35040 4878 35096 4886
rect 35408 4878 35464 4886
rect 36526 4879 36582 4887
rect 36894 4879 36950 4887
rect 35028 4876 35517 4878
rect 35028 4756 35040 4876
rect 35096 4756 35408 4876
rect 35464 4756 35517 4876
rect 35028 4754 35517 4756
rect 36514 4877 37003 4879
rect 36514 4757 36526 4877
rect 36582 4757 36894 4877
rect 36950 4757 37003 4877
rect 36514 4755 37003 4757
rect 35040 4746 35096 4754
rect 35408 4746 35517 4754
rect 36526 4747 36582 4755
rect 36894 4747 37003 4755
rect 34936 4680 35016 4690
rect 34936 4624 34948 4680
rect 35004 4624 35016 4680
rect 34936 4614 35016 4624
rect 35120 4680 35200 4690
rect 35120 4624 35132 4680
rect 35188 4624 35200 4680
rect 35120 4614 35200 4624
rect 35304 4680 35384 4690
rect 35304 4624 35316 4680
rect 35372 4624 35384 4680
rect 35304 4614 35384 4624
rect 34948 4532 35004 4614
rect 34936 4530 35016 4532
rect 34936 4474 34948 4530
rect 35004 4474 35016 4530
rect 34936 4472 35016 4474
rect 34264 4298 34334 4310
rect 34264 4242 34276 4298
rect 34332 4242 34334 4298
rect 34264 4230 34334 4242
rect 34948 4158 35004 4472
rect 35132 4416 35188 4614
rect 35120 4414 35200 4416
rect 35120 4358 35132 4414
rect 35188 4358 35200 4414
rect 35120 4356 35200 4358
rect 35132 4158 35188 4356
rect 35316 4300 35372 4614
rect 35449 4416 35517 4746
rect 36422 4681 36502 4691
rect 36422 4625 36434 4681
rect 36490 4625 36502 4681
rect 36422 4615 36502 4625
rect 36606 4681 36686 4691
rect 36606 4625 36618 4681
rect 36674 4625 36686 4681
rect 36606 4615 36686 4625
rect 36790 4681 36870 4691
rect 36790 4625 36802 4681
rect 36858 4625 36870 4681
rect 36790 4615 36870 4625
rect 36434 4533 36490 4615
rect 36422 4531 36502 4533
rect 36422 4475 36434 4531
rect 36490 4475 36502 4531
rect 36422 4473 36502 4475
rect 35449 4414 35529 4416
rect 35449 4358 35461 4414
rect 35517 4358 35529 4414
rect 35449 4356 35529 4358
rect 35716 4414 35786 4426
rect 35716 4358 35718 4414
rect 35774 4358 35786 4414
rect 35304 4298 35384 4300
rect 35304 4242 35316 4298
rect 35372 4242 35384 4298
rect 35304 4240 35384 4242
rect 35316 4158 35372 4240
rect 34936 4148 35016 4158
rect 34936 4092 34948 4148
rect 35004 4092 35016 4148
rect 34936 4082 35016 4092
rect 35120 4148 35200 4158
rect 35120 4092 35132 4148
rect 35188 4092 35200 4148
rect 35120 4082 35200 4092
rect 35304 4148 35384 4158
rect 35304 4092 35316 4148
rect 35372 4092 35384 4148
rect 35304 4082 35384 4092
rect 35449 4026 35517 4356
rect 35716 4348 35786 4358
rect 35408 4018 35517 4026
rect 35396 4016 35517 4018
rect 35396 3896 35408 4016
rect 35464 3896 35517 4016
rect 35396 3894 35517 3896
rect 35408 3886 35464 3894
rect 34711 3629 35607 3641
rect 34711 3573 34723 3629
rect 34779 3573 35541 3629
rect 35597 3573 35607 3629
rect 34711 3561 35607 3573
rect 35718 3404 35774 4348
rect 36434 4159 36490 4473
rect 36618 4417 36674 4615
rect 36606 4415 36686 4417
rect 36606 4359 36618 4415
rect 36674 4359 36686 4415
rect 36606 4357 36686 4359
rect 36618 4159 36674 4357
rect 36802 4301 36858 4615
rect 36935 4417 37003 4747
rect 37380 4425 37436 5659
rect 36935 4415 37015 4417
rect 36935 4359 36947 4415
rect 37003 4359 37015 4415
rect 36935 4357 37015 4359
rect 37378 4415 37448 4425
rect 37378 4359 37380 4415
rect 37436 4359 37528 4415
rect 36790 4299 36870 4301
rect 36790 4243 36802 4299
rect 36858 4243 36870 4299
rect 36790 4241 36870 4243
rect 36802 4159 36858 4241
rect 36422 4149 36502 4159
rect 36422 4093 36434 4149
rect 36490 4093 36502 4149
rect 36422 4083 36502 4093
rect 36606 4149 36686 4159
rect 36606 4093 36618 4149
rect 36674 4093 36686 4149
rect 36606 4083 36686 4093
rect 36790 4149 36870 4159
rect 36790 4093 36802 4149
rect 36858 4093 36870 4149
rect 36790 4083 36870 4093
rect 36935 4027 37003 4357
rect 37378 4347 37448 4359
rect 36894 4019 37003 4027
rect 36882 4017 37003 4019
rect 36882 3897 36894 4017
rect 36950 3897 37003 4017
rect 36882 3895 37003 3897
rect 36894 3887 36950 3895
rect 36197 3630 37093 3642
rect 36197 3574 36209 3630
rect 36265 3574 37027 3630
rect 37083 3574 37093 3630
rect 36197 3562 37093 3574
rect 35882 3511 35962 3521
rect 35882 3455 35894 3511
rect 35950 3455 35962 3511
rect 35882 3453 35962 3455
rect 35716 3401 35786 3404
rect 35716 3347 35718 3401
rect 35774 3347 35786 3401
rect 35716 3335 35786 3347
rect 34856 3294 35602 3306
rect 34856 3238 35224 3294
rect 35280 3238 35602 3294
rect 34856 3226 35602 3238
rect 34856 2973 34912 3226
rect 35224 2973 35280 3226
rect 35546 2973 35602 3226
rect 34844 2971 34924 2973
rect 34844 2851 34856 2971
rect 34912 2851 34924 2971
rect 34844 2849 34924 2851
rect 35212 2971 35292 2973
rect 35212 2851 35224 2971
rect 35280 2851 35292 2971
rect 35212 2849 35292 2851
rect 35534 2971 35614 2973
rect 35534 2850 35546 2971
rect 35602 2850 35614 2971
rect 34856 2841 34912 2849
rect 35224 2841 35280 2849
rect 35534 2848 35614 2850
rect 35546 2840 35602 2848
rect 35040 2673 35096 2681
rect 35408 2673 35464 2681
rect 35028 2671 35517 2673
rect 35028 2551 35040 2671
rect 35096 2551 35408 2671
rect 35464 2551 35517 2671
rect 35028 2549 35517 2551
rect 35040 2541 35096 2549
rect 35408 2541 35517 2549
rect 34936 2475 35016 2485
rect 34936 2419 34948 2475
rect 35004 2419 35016 2475
rect 34936 2409 35016 2419
rect 35120 2475 35200 2485
rect 35120 2419 35132 2475
rect 35188 2419 35200 2475
rect 35120 2409 35200 2419
rect 35304 2475 35384 2485
rect 35304 2419 35316 2475
rect 35372 2419 35384 2475
rect 35304 2409 35384 2419
rect 34948 2327 35004 2409
rect 34936 2325 35016 2327
rect 34936 2269 34948 2325
rect 35004 2269 35016 2325
rect 34936 2267 35016 2269
rect 34128 2209 34198 2223
rect 34128 2153 34140 2209
rect 34196 2153 34198 2209
rect 34128 2141 34198 2153
rect 33894 2093 33972 2104
rect 33502 2092 33972 2093
rect 33502 2038 33906 2092
rect 33960 2038 33972 2092
rect 33502 2037 33972 2038
rect 31930 1733 33102 1743
rect 31930 1677 31942 1733
rect 31998 1677 32830 1733
rect 32886 1677 33102 1733
rect 31930 1667 33102 1677
rect 33502 1733 33582 2037
rect 33894 2026 33972 2037
rect 33502 1677 33514 1733
rect 33570 1677 33582 1733
rect 33502 1667 33582 1677
rect 31860 1355 33652 1367
rect 31860 1215 31872 1355
rect 33640 1215 33652 1355
rect 33945 1306 34031 1318
rect 34140 1310 34196 2141
rect 34948 1953 35004 2267
rect 35132 2211 35188 2409
rect 35120 2209 35200 2211
rect 35120 2153 35132 2209
rect 35188 2153 35200 2209
rect 35120 2151 35200 2153
rect 35132 1953 35188 2151
rect 35316 2095 35372 2409
rect 35449 2211 35517 2541
rect 35894 2221 35950 3453
rect 37902 3347 37958 6563
rect 43600 6563 43612 6619
rect 43668 6563 43670 6619
rect 43600 6551 43670 6563
rect 43318 5717 43400 5729
rect 43318 5661 43332 5717
rect 43388 5661 43400 5717
rect 43318 5649 43400 5661
rect 38312 4311 38532 4321
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 42702 4311 43022 4321
rect 39174 3804 40346 3814
rect 39174 3564 39186 3804
rect 39242 3564 40278 3804
rect 40334 3564 40346 3804
rect 39174 3554 40346 3564
rect 38312 3501 38532 3511
rect 39268 3347 39346 3359
rect 37898 3291 39288 3347
rect 39344 3291 39346 3347
rect 39268 3279 39346 3291
rect 40266 3269 40346 3554
rect 40746 3804 40826 3814
rect 40746 3564 40758 3804
rect 40814 3564 40826 3804
rect 40568 3269 40638 3281
rect 40266 3213 40580 3269
rect 40636 3213 40638 3269
rect 40088 3191 40158 3203
rect 37898 3135 40100 3191
rect 40156 3135 40158 3191
rect 35449 2209 35529 2211
rect 35449 2153 35461 2209
rect 35517 2153 35529 2209
rect 35449 2151 35529 2153
rect 35892 2209 35952 2221
rect 35892 2153 35894 2209
rect 35950 2153 35952 2209
rect 35304 2093 35384 2095
rect 35304 2037 35316 2093
rect 35372 2037 35384 2093
rect 35304 2035 35384 2037
rect 35316 1953 35372 2035
rect 34936 1943 35016 1953
rect 34936 1887 34948 1943
rect 35004 1887 35016 1943
rect 34936 1877 35016 1887
rect 35120 1943 35200 1953
rect 35120 1887 35132 1943
rect 35188 1887 35200 1943
rect 35120 1877 35200 1887
rect 35304 1943 35384 1953
rect 35304 1887 35316 1943
rect 35372 1887 35384 1943
rect 35304 1877 35384 1887
rect 35449 1821 35517 2151
rect 35892 2141 35952 2153
rect 38010 1850 38066 3135
rect 40088 3123 40158 3135
rect 39378 2909 39458 2919
rect 39378 2853 39390 2909
rect 39446 2853 39458 2909
rect 39378 2667 39458 2853
rect 39858 2909 39938 2919
rect 39858 2853 39870 2909
rect 39926 2853 39938 2909
rect 39858 2843 39938 2853
rect 40062 2909 40142 2919
rect 40062 2853 40074 2909
rect 40130 2853 40142 2909
rect 40062 2667 40142 2853
rect 40266 2909 40346 3213
rect 40568 3201 40638 3213
rect 40746 3269 40826 3564
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 42702 3501 43022 3511
rect 41332 3315 43124 3327
rect 40746 3213 41103 3269
rect 40266 2853 40278 2909
rect 40334 2853 40346 2909
rect 40266 2843 40346 2853
rect 40746 2909 40826 3213
rect 40746 2853 40758 2909
rect 40814 2853 40826 2909
rect 40746 2843 40826 2853
rect 39378 2595 40142 2667
rect 40272 2541 40896 2553
rect 40272 2401 40284 2541
rect 40884 2401 40896 2541
rect 38484 2384 38564 2394
rect 40272 2389 40896 2401
rect 38484 2144 38496 2384
rect 38552 2144 38564 2384
rect 41047 2171 41103 3213
rect 41332 3175 41344 3315
rect 43112 3175 43124 3315
rect 41332 3163 43124 3175
rect 41606 2912 42370 2922
rect 41606 2672 41618 2912
rect 41674 2672 42302 2912
rect 42358 2672 42370 2912
rect 41606 2662 42370 2672
rect 42974 2628 43054 2638
rect 42086 2578 42574 2588
rect 42086 2338 42098 2578
rect 42154 2338 42506 2578
rect 42562 2338 42574 2578
rect 42086 2328 42574 2338
rect 41496 2171 41592 2183
rect 35408 1813 35517 1821
rect 35396 1811 35517 1813
rect 35396 1691 35408 1811
rect 35464 1691 35517 1811
rect 37498 1849 38066 1850
rect 38306 1849 38376 1861
rect 37498 1794 38318 1849
rect 35396 1689 35517 1691
rect 35408 1681 35464 1689
rect 34711 1424 35609 1436
rect 34711 1368 34723 1424
rect 34779 1368 35541 1424
rect 35597 1368 35609 1424
rect 34711 1356 35609 1368
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 34138 1306 34198 1310
rect 34138 1250 34140 1306
rect 34196 1250 34198 1306
rect 34138 1238 34198 1250
rect 31860 1203 33652 1215
rect 31274 873 31631 929
rect 33230 1031 33550 1041
rect 30794 513 30806 569
rect 30862 513 30874 569
rect 30794 503 30874 513
rect 31274 569 31354 873
rect 31274 513 31286 569
rect 31342 513 31354 569
rect 31274 503 31354 513
rect 29906 255 30670 327
rect 33230 231 33240 1031
rect 33540 231 33550 1031
rect 33230 221 33550 231
rect 37503 -49 37559 1794
rect 38010 1793 38318 1794
rect 38374 1793 38376 1849
rect 38306 1781 38376 1793
rect 38484 1849 38564 2144
rect 40272 2141 40896 2153
rect 40272 2001 40284 2141
rect 40884 2001 40896 2141
rect 41047 2115 41516 2171
rect 41572 2115 41592 2171
rect 41496 2103 41592 2115
rect 42494 2093 42574 2328
rect 42974 2388 42986 2628
rect 43042 2388 43054 2628
rect 42796 2093 42866 2105
rect 42494 2037 42808 2093
rect 42864 2037 42866 2093
rect 42180 2015 42276 2025
rect 40272 1989 40896 2001
rect 41047 1959 42200 2015
rect 42256 1959 42276 2015
rect 38484 1793 38922 1849
rect 38484 1489 38564 1793
rect 38484 1433 38496 1489
rect 38552 1433 38564 1489
rect 38484 1423 38564 1433
rect 38866 1007 38922 1793
rect 39174 1464 40346 1474
rect 39174 1224 39186 1464
rect 39242 1224 40278 1464
rect 40334 1224 40346 1464
rect 39174 1214 40346 1224
rect 39268 1007 39346 1019
rect 38866 951 39288 1007
rect 39344 951 39346 1007
rect 39268 939 39346 951
rect 40266 929 40346 1214
rect 40746 1464 40826 1474
rect 40746 1224 40758 1464
rect 40814 1224 40826 1464
rect 40568 929 40638 941
rect 40266 873 40580 929
rect 40636 873 40638 929
rect 40088 851 40158 863
rect 37503 -179 37559 -169
rect 37898 795 40100 851
rect 40156 795 40158 851
rect 37898 -369 37954 795
rect 40088 783 40158 795
rect 39378 569 39458 579
rect 39378 513 39390 569
rect 39446 513 39458 569
rect 39378 327 39458 513
rect 39858 569 39938 579
rect 39858 513 39870 569
rect 39926 513 39938 569
rect 39858 503 39938 513
rect 40062 569 40142 579
rect 40062 513 40074 569
rect 40130 513 40142 569
rect 40062 327 40142 513
rect 40266 569 40346 873
rect 40568 861 40638 873
rect 40746 929 40826 1224
rect 41047 929 41103 1959
rect 42180 1949 42276 1959
rect 42494 1743 42574 2037
rect 42796 2025 42866 2037
rect 42974 2093 43054 2388
rect 43612 2223 43668 6551
rect 43748 4310 43804 8756
rect 44420 8568 44476 8882
rect 44604 8826 44660 9024
rect 44592 8824 44672 8826
rect 44592 8768 44604 8824
rect 44660 8768 44672 8824
rect 44592 8766 44672 8768
rect 44604 8568 44660 8766
rect 44788 8710 44844 9024
rect 44921 8826 44989 9156
rect 53880 9090 53960 9100
rect 53880 9034 53892 9090
rect 53948 9034 53960 9090
rect 53880 9024 53960 9034
rect 54064 9090 54144 9100
rect 54064 9034 54076 9090
rect 54132 9034 54144 9090
rect 54064 9024 54144 9034
rect 54248 9090 54328 9100
rect 54248 9034 54260 9090
rect 54316 9034 54328 9090
rect 54248 9024 54328 9034
rect 52990 8940 53078 8952
rect 53892 8942 53948 9024
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 53880 8940 53960 8942
rect 53880 8884 53892 8940
rect 53948 8884 53960 8940
rect 53880 8882 53960 8884
rect 44921 8824 45001 8826
rect 44921 8768 44933 8824
rect 44989 8768 45001 8824
rect 44921 8766 45001 8768
rect 45188 8824 45258 8836
rect 45188 8768 45190 8824
rect 45246 8768 45258 8824
rect 44776 8708 44856 8710
rect 44776 8652 44788 8708
rect 44844 8652 44856 8708
rect 44776 8650 44856 8652
rect 44788 8568 44844 8650
rect 44408 8558 44488 8568
rect 44408 8502 44420 8558
rect 44476 8502 44488 8558
rect 44408 8492 44488 8502
rect 44592 8558 44672 8568
rect 44592 8502 44604 8558
rect 44660 8502 44672 8558
rect 44592 8492 44672 8502
rect 44776 8558 44856 8568
rect 44776 8502 44788 8558
rect 44844 8502 44856 8558
rect 44776 8492 44856 8502
rect 44921 8436 44989 8766
rect 45188 8758 45258 8768
rect 53208 8824 53278 8836
rect 53208 8768 53220 8824
rect 53276 8768 53278 8824
rect 44880 8428 44989 8436
rect 44868 8426 44989 8428
rect 44868 8306 44880 8426
rect 44936 8306 44989 8426
rect 44868 8304 44989 8306
rect 44880 8296 44936 8304
rect 44183 8039 45081 8051
rect 44183 7983 44195 8039
rect 44251 7983 45013 8039
rect 45069 7983 45081 8039
rect 44183 7971 45081 7983
rect 45190 7814 45246 8758
rect 53208 8756 53278 8768
rect 45354 7921 45434 7931
rect 45354 7865 45366 7921
rect 45422 7865 45434 7921
rect 45354 7863 45434 7865
rect 45188 7811 45258 7814
rect 45188 7757 45190 7811
rect 45246 7757 45258 7811
rect 45188 7745 45258 7757
rect 44328 7704 45074 7716
rect 44328 7648 44696 7704
rect 44752 7648 45074 7704
rect 44328 7636 45074 7648
rect 44328 7383 44384 7636
rect 44696 7383 44752 7636
rect 45018 7383 45074 7636
rect 44316 7381 44396 7383
rect 44316 7261 44328 7381
rect 44384 7261 44396 7381
rect 44316 7259 44396 7261
rect 44684 7381 44764 7383
rect 44684 7261 44696 7381
rect 44752 7261 44764 7381
rect 44684 7259 44764 7261
rect 45006 7381 45086 7383
rect 45006 7260 45018 7381
rect 45074 7260 45086 7381
rect 44328 7251 44384 7259
rect 44696 7251 44752 7259
rect 45006 7258 45086 7260
rect 45018 7250 45074 7258
rect 44512 7083 44568 7091
rect 44880 7083 44936 7091
rect 44500 7081 44989 7083
rect 44500 6961 44512 7081
rect 44568 6961 44880 7081
rect 44936 6961 44989 7081
rect 44500 6959 44989 6961
rect 44512 6951 44568 6959
rect 44880 6951 44989 6959
rect 44408 6885 44488 6895
rect 44408 6829 44420 6885
rect 44476 6829 44488 6885
rect 44408 6819 44488 6829
rect 44592 6885 44672 6895
rect 44592 6829 44604 6885
rect 44660 6829 44672 6885
rect 44592 6819 44672 6829
rect 44776 6885 44856 6895
rect 44776 6829 44788 6885
rect 44844 6829 44856 6885
rect 44776 6819 44856 6829
rect 44420 6737 44476 6819
rect 44408 6735 44488 6737
rect 44408 6679 44420 6735
rect 44476 6679 44488 6735
rect 44408 6677 44488 6679
rect 44420 6363 44476 6677
rect 44604 6621 44660 6819
rect 44592 6619 44672 6621
rect 44592 6563 44604 6619
rect 44660 6563 44672 6619
rect 44592 6561 44672 6563
rect 44604 6363 44660 6561
rect 44788 6505 44844 6819
rect 44921 6621 44989 6951
rect 45366 6629 45422 7863
rect 45814 7704 46560 7716
rect 45814 7648 46182 7704
rect 46238 7648 46560 7704
rect 45814 7636 46560 7648
rect 45814 7383 45870 7636
rect 46182 7383 46238 7636
rect 46504 7383 46560 7636
rect 45802 7381 45882 7383
rect 45802 7261 45814 7381
rect 45870 7261 45882 7381
rect 45802 7259 45882 7261
rect 46170 7381 46250 7383
rect 46170 7261 46182 7381
rect 46238 7261 46250 7381
rect 46170 7259 46250 7261
rect 46492 7381 46572 7383
rect 46492 7260 46504 7381
rect 46560 7260 46572 7381
rect 45814 7251 45870 7259
rect 46182 7251 46238 7259
rect 46492 7258 46572 7260
rect 46504 7250 46560 7258
rect 45998 7083 46054 7091
rect 46366 7083 46422 7091
rect 45986 7081 46475 7083
rect 45986 6961 45998 7081
rect 46054 6961 46366 7081
rect 46422 6961 46475 7081
rect 45986 6959 46475 6961
rect 45998 6951 46054 6959
rect 46366 6951 46475 6959
rect 45894 6885 45974 6895
rect 45894 6829 45906 6885
rect 45962 6829 45974 6885
rect 45894 6819 45974 6829
rect 46078 6885 46158 6895
rect 46078 6829 46090 6885
rect 46146 6829 46158 6885
rect 46078 6819 46158 6829
rect 46262 6885 46342 6895
rect 46262 6829 46274 6885
rect 46330 6829 46342 6885
rect 46262 6819 46342 6829
rect 45906 6737 45962 6819
rect 45894 6735 45974 6737
rect 45894 6679 45906 6735
rect 45962 6679 45974 6735
rect 45894 6677 45974 6679
rect 44921 6619 45001 6621
rect 44921 6563 44933 6619
rect 44989 6563 45001 6619
rect 44921 6561 45001 6563
rect 45364 6619 45424 6629
rect 45364 6563 45366 6619
rect 45422 6563 45424 6619
rect 44776 6503 44856 6505
rect 44776 6447 44788 6503
rect 44844 6447 44856 6503
rect 44776 6445 44856 6447
rect 44788 6363 44844 6445
rect 44408 6353 44488 6363
rect 44408 6297 44420 6353
rect 44476 6297 44488 6353
rect 44408 6287 44488 6297
rect 44592 6353 44672 6363
rect 44592 6297 44604 6353
rect 44660 6297 44672 6353
rect 44592 6287 44672 6297
rect 44776 6353 44856 6363
rect 44776 6297 44788 6353
rect 44844 6297 44856 6353
rect 44776 6287 44856 6297
rect 44921 6231 44989 6561
rect 45364 6551 45424 6563
rect 44880 6223 44989 6231
rect 44868 6221 44989 6223
rect 44868 6101 44880 6221
rect 44936 6101 44989 6221
rect 44868 6099 44989 6101
rect 44880 6091 44936 6099
rect 44183 5834 45079 5846
rect 44183 5778 44195 5834
rect 44251 5778 45013 5834
rect 45069 5778 45079 5834
rect 44183 5766 45079 5778
rect 45366 5608 45422 6551
rect 45906 6363 45962 6677
rect 46090 6621 46146 6819
rect 46078 6619 46158 6621
rect 46078 6563 46090 6619
rect 46146 6563 46158 6619
rect 46078 6561 46158 6563
rect 46090 6363 46146 6561
rect 46274 6505 46330 6819
rect 46407 6621 46475 6951
rect 46407 6619 46487 6621
rect 46407 6563 46419 6619
rect 46475 6563 46487 6619
rect 46407 6561 46487 6563
rect 46674 6619 46744 6631
rect 53072 6619 53142 6633
rect 46674 6563 46676 6619
rect 46732 6563 47430 6619
rect 46262 6503 46342 6505
rect 46262 6447 46274 6503
rect 46330 6447 46342 6503
rect 46262 6445 46342 6447
rect 46274 6363 46330 6445
rect 45894 6353 45974 6363
rect 45894 6297 45906 6353
rect 45962 6297 45974 6353
rect 45894 6287 45974 6297
rect 46078 6353 46158 6363
rect 46078 6297 46090 6353
rect 46146 6297 46158 6353
rect 46078 6287 46158 6297
rect 46262 6353 46342 6363
rect 46262 6297 46274 6353
rect 46330 6297 46342 6353
rect 46262 6287 46342 6297
rect 46407 6231 46475 6561
rect 46674 6553 46744 6563
rect 46366 6223 46475 6231
rect 46354 6221 46475 6223
rect 46354 6101 46366 6221
rect 46422 6101 46475 6221
rect 46354 6099 46475 6101
rect 46366 6091 46422 6099
rect 45669 5834 46565 5846
rect 45669 5778 45681 5834
rect 45737 5778 46499 5834
rect 46555 5778 46565 5834
rect 45669 5766 46565 5778
rect 46676 5609 46732 6553
rect 46840 5717 46920 5727
rect 46840 5661 46852 5717
rect 46908 5661 46920 5717
rect 46840 5659 46920 5661
rect 45364 5606 45434 5608
rect 45364 5550 45366 5606
rect 45422 5550 45434 5606
rect 45364 5538 45434 5550
rect 46664 5607 46744 5609
rect 46664 5551 46676 5607
rect 46732 5551 46744 5607
rect 46664 5539 46744 5551
rect 44328 5499 45074 5511
rect 44328 5443 44696 5499
rect 44752 5443 45074 5499
rect 44328 5431 45074 5443
rect 44328 5178 44384 5431
rect 44696 5178 44752 5431
rect 45018 5178 45074 5431
rect 45814 5500 46560 5512
rect 45814 5444 46182 5500
rect 46238 5444 46560 5500
rect 45814 5432 46560 5444
rect 45814 5179 45870 5432
rect 46182 5179 46238 5432
rect 46504 5179 46560 5432
rect 44316 5176 44396 5178
rect 44316 5056 44328 5176
rect 44384 5056 44396 5176
rect 44316 5054 44396 5056
rect 44684 5176 44764 5178
rect 44684 5056 44696 5176
rect 44752 5056 44764 5176
rect 44684 5054 44764 5056
rect 45006 5176 45086 5178
rect 45006 5055 45018 5176
rect 45074 5055 45086 5176
rect 45802 5177 45882 5179
rect 45802 5057 45814 5177
rect 45870 5057 45882 5177
rect 45802 5055 45882 5057
rect 46170 5177 46250 5179
rect 46170 5057 46182 5177
rect 46238 5057 46250 5177
rect 46170 5055 46250 5057
rect 46492 5177 46572 5179
rect 46492 5056 46504 5177
rect 46560 5056 46572 5177
rect 44328 5046 44384 5054
rect 44696 5046 44752 5054
rect 45006 5053 45086 5055
rect 45018 5045 45074 5053
rect 45814 5047 45870 5055
rect 46182 5047 46238 5055
rect 46492 5054 46572 5056
rect 46504 5046 46560 5054
rect 44512 4878 44568 4886
rect 44880 4878 44936 4886
rect 45998 4879 46054 4887
rect 46366 4879 46422 4887
rect 44500 4876 44989 4878
rect 44500 4756 44512 4876
rect 44568 4756 44880 4876
rect 44936 4756 44989 4876
rect 44500 4754 44989 4756
rect 45986 4877 46475 4879
rect 45986 4757 45998 4877
rect 46054 4757 46366 4877
rect 46422 4757 46475 4877
rect 45986 4755 46475 4757
rect 44512 4746 44568 4754
rect 44880 4746 44989 4754
rect 45998 4747 46054 4755
rect 46366 4747 46475 4755
rect 44408 4680 44488 4690
rect 44408 4624 44420 4680
rect 44476 4624 44488 4680
rect 44408 4614 44488 4624
rect 44592 4680 44672 4690
rect 44592 4624 44604 4680
rect 44660 4624 44672 4680
rect 44592 4614 44672 4624
rect 44776 4680 44856 4690
rect 44776 4624 44788 4680
rect 44844 4624 44856 4680
rect 44776 4614 44856 4624
rect 44420 4532 44476 4614
rect 44408 4530 44488 4532
rect 44408 4474 44420 4530
rect 44476 4474 44488 4530
rect 44408 4472 44488 4474
rect 43736 4298 43806 4310
rect 43736 4242 43748 4298
rect 43804 4242 43806 4298
rect 43736 4230 43806 4242
rect 44420 4158 44476 4472
rect 44604 4416 44660 4614
rect 44592 4414 44672 4416
rect 44592 4358 44604 4414
rect 44660 4358 44672 4414
rect 44592 4356 44672 4358
rect 44604 4158 44660 4356
rect 44788 4300 44844 4614
rect 44921 4416 44989 4746
rect 45894 4681 45974 4691
rect 45894 4625 45906 4681
rect 45962 4625 45974 4681
rect 45894 4615 45974 4625
rect 46078 4681 46158 4691
rect 46078 4625 46090 4681
rect 46146 4625 46158 4681
rect 46078 4615 46158 4625
rect 46262 4681 46342 4691
rect 46262 4625 46274 4681
rect 46330 4625 46342 4681
rect 46262 4615 46342 4625
rect 45906 4533 45962 4615
rect 45894 4531 45974 4533
rect 45894 4475 45906 4531
rect 45962 4475 45974 4531
rect 45894 4473 45974 4475
rect 44921 4414 45001 4416
rect 44921 4358 44933 4414
rect 44989 4358 45001 4414
rect 44921 4356 45001 4358
rect 45188 4414 45258 4426
rect 45188 4358 45190 4414
rect 45246 4358 45258 4414
rect 44776 4298 44856 4300
rect 44776 4242 44788 4298
rect 44844 4242 44856 4298
rect 44776 4240 44856 4242
rect 44788 4158 44844 4240
rect 44408 4148 44488 4158
rect 44408 4092 44420 4148
rect 44476 4092 44488 4148
rect 44408 4082 44488 4092
rect 44592 4148 44672 4158
rect 44592 4092 44604 4148
rect 44660 4092 44672 4148
rect 44592 4082 44672 4092
rect 44776 4148 44856 4158
rect 44776 4092 44788 4148
rect 44844 4092 44856 4148
rect 44776 4082 44856 4092
rect 44921 4026 44989 4356
rect 45188 4348 45258 4358
rect 44880 4018 44989 4026
rect 44868 4016 44989 4018
rect 44868 3896 44880 4016
rect 44936 3896 44989 4016
rect 44868 3894 44989 3896
rect 44880 3886 44936 3894
rect 44183 3629 45079 3641
rect 44183 3573 44195 3629
rect 44251 3573 45013 3629
rect 45069 3573 45079 3629
rect 44183 3561 45079 3573
rect 45190 3404 45246 4348
rect 45906 4159 45962 4473
rect 46090 4417 46146 4615
rect 46078 4415 46158 4417
rect 46078 4359 46090 4415
rect 46146 4359 46158 4415
rect 46078 4357 46158 4359
rect 46090 4159 46146 4357
rect 46274 4301 46330 4615
rect 46407 4417 46475 4747
rect 46852 4425 46908 5659
rect 46407 4415 46487 4417
rect 46407 4359 46419 4415
rect 46475 4359 46487 4415
rect 46407 4357 46487 4359
rect 46850 4415 46920 4425
rect 46850 4359 46852 4415
rect 46908 4359 47000 4415
rect 46262 4299 46342 4301
rect 46262 4243 46274 4299
rect 46330 4243 46342 4299
rect 46262 4241 46342 4243
rect 46274 4159 46330 4241
rect 45894 4149 45974 4159
rect 45894 4093 45906 4149
rect 45962 4093 45974 4149
rect 45894 4083 45974 4093
rect 46078 4149 46158 4159
rect 46078 4093 46090 4149
rect 46146 4093 46158 4149
rect 46078 4083 46158 4093
rect 46262 4149 46342 4159
rect 46262 4093 46274 4149
rect 46330 4093 46342 4149
rect 46262 4083 46342 4093
rect 46407 4027 46475 4357
rect 46850 4347 46920 4359
rect 46366 4019 46475 4027
rect 46354 4017 46475 4019
rect 46354 3897 46366 4017
rect 46422 3897 46475 4017
rect 46354 3895 46475 3897
rect 46366 3887 46422 3895
rect 45669 3630 46565 3642
rect 45669 3574 45681 3630
rect 45737 3574 46499 3630
rect 46555 3574 46565 3630
rect 45669 3562 46565 3574
rect 45354 3511 45434 3521
rect 45354 3455 45366 3511
rect 45422 3455 45434 3511
rect 45354 3453 45434 3455
rect 45188 3401 45258 3404
rect 45188 3347 45190 3401
rect 45246 3347 45258 3401
rect 45188 3335 45258 3347
rect 44328 3294 45074 3306
rect 44328 3238 44696 3294
rect 44752 3238 45074 3294
rect 44328 3226 45074 3238
rect 44328 2973 44384 3226
rect 44696 2973 44752 3226
rect 45018 2973 45074 3226
rect 44316 2971 44396 2973
rect 44316 2851 44328 2971
rect 44384 2851 44396 2971
rect 44316 2849 44396 2851
rect 44684 2971 44764 2973
rect 44684 2851 44696 2971
rect 44752 2851 44764 2971
rect 44684 2849 44764 2851
rect 45006 2971 45086 2973
rect 45006 2850 45018 2971
rect 45074 2850 45086 2971
rect 44328 2841 44384 2849
rect 44696 2841 44752 2849
rect 45006 2848 45086 2850
rect 45018 2840 45074 2848
rect 44512 2673 44568 2681
rect 44880 2673 44936 2681
rect 44500 2671 44989 2673
rect 44500 2551 44512 2671
rect 44568 2551 44880 2671
rect 44936 2551 44989 2671
rect 44500 2549 44989 2551
rect 44512 2541 44568 2549
rect 44880 2541 44989 2549
rect 44408 2475 44488 2485
rect 44408 2419 44420 2475
rect 44476 2419 44488 2475
rect 44408 2409 44488 2419
rect 44592 2475 44672 2485
rect 44592 2419 44604 2475
rect 44660 2419 44672 2475
rect 44592 2409 44672 2419
rect 44776 2475 44856 2485
rect 44776 2419 44788 2475
rect 44844 2419 44856 2475
rect 44776 2409 44856 2419
rect 44420 2327 44476 2409
rect 44408 2325 44488 2327
rect 44408 2269 44420 2325
rect 44476 2269 44488 2325
rect 44408 2267 44488 2269
rect 43600 2209 43670 2223
rect 43600 2153 43612 2209
rect 43668 2153 43670 2209
rect 43600 2141 43670 2153
rect 43366 2093 43444 2104
rect 42974 2092 43444 2093
rect 42974 2038 43378 2092
rect 43432 2038 43444 2092
rect 42974 2037 43444 2038
rect 41402 1733 42574 1743
rect 41402 1677 41414 1733
rect 41470 1677 42302 1733
rect 42358 1677 42574 1733
rect 41402 1667 42574 1677
rect 42974 1733 43054 2037
rect 43366 2026 43444 2037
rect 42974 1677 42986 1733
rect 43042 1677 43054 1733
rect 42974 1667 43054 1677
rect 41332 1355 43124 1367
rect 41332 1215 41344 1355
rect 43112 1215 43124 1355
rect 43417 1306 43503 1318
rect 43612 1310 43668 2141
rect 44420 1953 44476 2267
rect 44604 2211 44660 2409
rect 44592 2209 44672 2211
rect 44592 2153 44604 2209
rect 44660 2153 44672 2209
rect 44592 2151 44672 2153
rect 44604 1953 44660 2151
rect 44788 2095 44844 2409
rect 44921 2211 44989 2541
rect 45366 2221 45422 3453
rect 47374 3347 47430 6563
rect 53072 6563 53084 6619
rect 53140 6563 53142 6619
rect 53072 6551 53142 6563
rect 52790 5717 52872 5729
rect 52790 5661 52804 5717
rect 52860 5661 52872 5717
rect 52790 5649 52872 5661
rect 47784 4311 48004 4321
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 52174 4311 52494 4321
rect 48646 3804 49818 3814
rect 48646 3564 48658 3804
rect 48714 3564 49750 3804
rect 49806 3564 49818 3804
rect 48646 3554 49818 3564
rect 47784 3501 48004 3511
rect 48740 3347 48818 3359
rect 47370 3291 48760 3347
rect 48816 3291 48818 3347
rect 48740 3279 48818 3291
rect 49738 3269 49818 3554
rect 50218 3804 50298 3814
rect 50218 3564 50230 3804
rect 50286 3564 50298 3804
rect 50040 3269 50110 3281
rect 49738 3213 50052 3269
rect 50108 3213 50110 3269
rect 49560 3191 49630 3203
rect 47370 3135 49572 3191
rect 49628 3135 49630 3191
rect 44921 2209 45001 2211
rect 44921 2153 44933 2209
rect 44989 2153 45001 2209
rect 44921 2151 45001 2153
rect 45364 2209 45424 2221
rect 45364 2153 45366 2209
rect 45422 2153 45424 2209
rect 44776 2093 44856 2095
rect 44776 2037 44788 2093
rect 44844 2037 44856 2093
rect 44776 2035 44856 2037
rect 44788 1953 44844 2035
rect 44408 1943 44488 1953
rect 44408 1887 44420 1943
rect 44476 1887 44488 1943
rect 44408 1877 44488 1887
rect 44592 1943 44672 1953
rect 44592 1887 44604 1943
rect 44660 1887 44672 1943
rect 44592 1877 44672 1887
rect 44776 1943 44856 1953
rect 44776 1887 44788 1943
rect 44844 1887 44856 1943
rect 44776 1877 44856 1887
rect 44921 1821 44989 2151
rect 45364 2141 45424 2153
rect 47482 1850 47538 3135
rect 49560 3123 49630 3135
rect 48850 2909 48930 2919
rect 48850 2853 48862 2909
rect 48918 2853 48930 2909
rect 48850 2667 48930 2853
rect 49330 2909 49410 2919
rect 49330 2853 49342 2909
rect 49398 2853 49410 2909
rect 49330 2843 49410 2853
rect 49534 2909 49614 2919
rect 49534 2853 49546 2909
rect 49602 2853 49614 2909
rect 49534 2667 49614 2853
rect 49738 2909 49818 3213
rect 50040 3201 50110 3213
rect 50218 3269 50298 3564
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 52174 3501 52494 3511
rect 50804 3315 52596 3327
rect 50218 3213 50575 3269
rect 49738 2853 49750 2909
rect 49806 2853 49818 2909
rect 49738 2843 49818 2853
rect 50218 2909 50298 3213
rect 50218 2853 50230 2909
rect 50286 2853 50298 2909
rect 50218 2843 50298 2853
rect 48850 2595 49614 2667
rect 49744 2541 50368 2553
rect 49744 2401 49756 2541
rect 50356 2401 50368 2541
rect 47956 2384 48036 2394
rect 49744 2389 50368 2401
rect 47956 2144 47968 2384
rect 48024 2144 48036 2384
rect 50519 2171 50575 3213
rect 50804 3175 50816 3315
rect 52584 3175 52596 3315
rect 50804 3163 52596 3175
rect 51078 2912 51842 2922
rect 51078 2672 51090 2912
rect 51146 2672 51774 2912
rect 51830 2672 51842 2912
rect 51078 2662 51842 2672
rect 52446 2628 52526 2638
rect 51558 2578 52046 2588
rect 51558 2338 51570 2578
rect 51626 2338 51978 2578
rect 52034 2338 52046 2578
rect 51558 2328 52046 2338
rect 50968 2171 51064 2183
rect 44880 1813 44989 1821
rect 44868 1811 44989 1813
rect 44868 1691 44880 1811
rect 44936 1691 44989 1811
rect 46970 1849 47538 1850
rect 47778 1849 47848 1861
rect 46970 1794 47790 1849
rect 44868 1689 44989 1691
rect 44880 1681 44936 1689
rect 44183 1424 45081 1436
rect 44183 1368 44195 1424
rect 44251 1368 45013 1424
rect 45069 1368 45081 1424
rect 44183 1356 45081 1368
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 43610 1306 43670 1310
rect 43610 1250 43612 1306
rect 43668 1250 43670 1306
rect 43610 1238 43670 1250
rect 41332 1203 43124 1215
rect 40746 873 41103 929
rect 42702 1031 43022 1041
rect 40266 513 40278 569
rect 40334 513 40346 569
rect 40266 503 40346 513
rect 40746 569 40826 873
rect 40746 513 40758 569
rect 40814 513 40826 569
rect 40746 503 40826 513
rect 39378 255 40142 327
rect 42702 231 42712 1031
rect 43012 231 43022 1031
rect 42702 221 43022 231
rect 46975 -49 47031 1794
rect 47482 1793 47790 1794
rect 47846 1793 47848 1849
rect 47778 1781 47848 1793
rect 47956 1849 48036 2144
rect 49744 2141 50368 2153
rect 49744 2001 49756 2141
rect 50356 2001 50368 2141
rect 50519 2115 50988 2171
rect 51044 2115 51064 2171
rect 50968 2103 51064 2115
rect 51966 2093 52046 2328
rect 52446 2388 52458 2628
rect 52514 2388 52526 2628
rect 52268 2093 52338 2105
rect 51966 2037 52280 2093
rect 52336 2037 52338 2093
rect 51652 2015 51748 2025
rect 49744 1989 50368 2001
rect 50519 1959 51672 2015
rect 51728 1959 51748 2015
rect 47956 1793 48394 1849
rect 47956 1489 48036 1793
rect 47956 1433 47968 1489
rect 48024 1433 48036 1489
rect 47956 1423 48036 1433
rect 48338 1007 48394 1793
rect 48646 1464 49818 1474
rect 48646 1224 48658 1464
rect 48714 1224 49750 1464
rect 49806 1224 49818 1464
rect 48646 1214 49818 1224
rect 48740 1007 48818 1019
rect 48338 951 48760 1007
rect 48816 951 48818 1007
rect 48740 939 48818 951
rect 49738 929 49818 1214
rect 50218 1464 50298 1474
rect 50218 1224 50230 1464
rect 50286 1224 50298 1464
rect 50040 929 50110 941
rect 49738 873 50052 929
rect 50108 873 50110 929
rect 49560 851 49630 863
rect 46975 -179 47031 -169
rect 47370 795 49572 851
rect 49628 795 49630 851
rect 47370 -369 47426 795
rect 49560 783 49630 795
rect 48850 569 48930 579
rect 48850 513 48862 569
rect 48918 513 48930 569
rect 48850 327 48930 513
rect 49330 569 49410 579
rect 49330 513 49342 569
rect 49398 513 49410 569
rect 49330 503 49410 513
rect 49534 569 49614 579
rect 49534 513 49546 569
rect 49602 513 49614 569
rect 49534 327 49614 513
rect 49738 569 49818 873
rect 50040 861 50110 873
rect 50218 929 50298 1224
rect 50519 929 50575 1959
rect 51652 1949 51748 1959
rect 51966 1743 52046 2037
rect 52268 2025 52338 2037
rect 52446 2093 52526 2388
rect 53084 2223 53140 6551
rect 53220 4310 53276 8756
rect 53892 8568 53948 8882
rect 54076 8826 54132 9024
rect 54064 8824 54144 8826
rect 54064 8768 54076 8824
rect 54132 8768 54144 8824
rect 54064 8766 54144 8768
rect 54076 8568 54132 8766
rect 54260 8710 54316 9024
rect 54393 8826 54461 9156
rect 54393 8824 54473 8826
rect 54393 8768 54405 8824
rect 54461 8768 54473 8824
rect 54393 8766 54473 8768
rect 54660 8824 54730 8836
rect 54660 8768 54662 8824
rect 54718 8768 54730 8824
rect 54248 8708 54328 8710
rect 54248 8652 54260 8708
rect 54316 8652 54328 8708
rect 54248 8650 54328 8652
rect 54260 8568 54316 8650
rect 53880 8558 53960 8568
rect 53880 8502 53892 8558
rect 53948 8502 53960 8558
rect 53880 8492 53960 8502
rect 54064 8558 54144 8568
rect 54064 8502 54076 8558
rect 54132 8502 54144 8558
rect 54064 8492 54144 8502
rect 54248 8558 54328 8568
rect 54248 8502 54260 8558
rect 54316 8502 54328 8558
rect 54248 8492 54328 8502
rect 54393 8436 54461 8766
rect 54660 8758 54730 8768
rect 54352 8428 54461 8436
rect 54340 8426 54461 8428
rect 54340 8306 54352 8426
rect 54408 8306 54461 8426
rect 54340 8304 54461 8306
rect 54352 8296 54408 8304
rect 53655 8039 54553 8051
rect 53655 7983 53667 8039
rect 53723 7983 54485 8039
rect 54541 7983 54553 8039
rect 53655 7971 54553 7983
rect 54662 7814 54718 8758
rect 54826 7921 54906 7931
rect 54826 7865 54838 7921
rect 54894 7865 54906 7921
rect 54826 7863 54906 7865
rect 54660 7811 54730 7814
rect 54660 7757 54662 7811
rect 54718 7757 54730 7811
rect 54660 7745 54730 7757
rect 53800 7704 54546 7716
rect 53800 7648 54168 7704
rect 54224 7648 54546 7704
rect 53800 7636 54546 7648
rect 53800 7383 53856 7636
rect 54168 7383 54224 7636
rect 54490 7383 54546 7636
rect 53788 7381 53868 7383
rect 53788 7261 53800 7381
rect 53856 7261 53868 7381
rect 53788 7259 53868 7261
rect 54156 7381 54236 7383
rect 54156 7261 54168 7381
rect 54224 7261 54236 7381
rect 54156 7259 54236 7261
rect 54478 7381 54558 7383
rect 54478 7260 54490 7381
rect 54546 7260 54558 7381
rect 53800 7251 53856 7259
rect 54168 7251 54224 7259
rect 54478 7258 54558 7260
rect 54490 7250 54546 7258
rect 53984 7083 54040 7091
rect 54352 7083 54408 7091
rect 53972 7081 54461 7083
rect 53972 6961 53984 7081
rect 54040 6961 54352 7081
rect 54408 6961 54461 7081
rect 53972 6959 54461 6961
rect 53984 6951 54040 6959
rect 54352 6951 54461 6959
rect 53880 6885 53960 6895
rect 53880 6829 53892 6885
rect 53948 6829 53960 6885
rect 53880 6819 53960 6829
rect 54064 6885 54144 6895
rect 54064 6829 54076 6885
rect 54132 6829 54144 6885
rect 54064 6819 54144 6829
rect 54248 6885 54328 6895
rect 54248 6829 54260 6885
rect 54316 6829 54328 6885
rect 54248 6819 54328 6829
rect 53892 6737 53948 6819
rect 53880 6735 53960 6737
rect 53880 6679 53892 6735
rect 53948 6679 53960 6735
rect 53880 6677 53960 6679
rect 53892 6363 53948 6677
rect 54076 6621 54132 6819
rect 54064 6619 54144 6621
rect 54064 6563 54076 6619
rect 54132 6563 54144 6619
rect 54064 6561 54144 6563
rect 54076 6363 54132 6561
rect 54260 6505 54316 6819
rect 54393 6621 54461 6951
rect 54838 6629 54894 7863
rect 55286 7704 56032 7716
rect 55286 7648 55654 7704
rect 55710 7648 56032 7704
rect 55286 7636 56032 7648
rect 55286 7383 55342 7636
rect 55654 7383 55710 7636
rect 55976 7383 56032 7636
rect 55274 7381 55354 7383
rect 55274 7261 55286 7381
rect 55342 7261 55354 7381
rect 55274 7259 55354 7261
rect 55642 7381 55722 7383
rect 55642 7261 55654 7381
rect 55710 7261 55722 7381
rect 55642 7259 55722 7261
rect 55964 7381 56044 7383
rect 55964 7260 55976 7381
rect 56032 7260 56044 7381
rect 55286 7251 55342 7259
rect 55654 7251 55710 7259
rect 55964 7258 56044 7260
rect 55976 7250 56032 7258
rect 55470 7083 55526 7091
rect 55838 7083 55894 7091
rect 55458 7081 55947 7083
rect 55458 6961 55470 7081
rect 55526 6961 55838 7081
rect 55894 6961 55947 7081
rect 55458 6959 55947 6961
rect 55470 6951 55526 6959
rect 55838 6951 55947 6959
rect 55366 6885 55446 6895
rect 55366 6829 55378 6885
rect 55434 6829 55446 6885
rect 55366 6819 55446 6829
rect 55550 6885 55630 6895
rect 55550 6829 55562 6885
rect 55618 6829 55630 6885
rect 55550 6819 55630 6829
rect 55734 6885 55814 6895
rect 55734 6829 55746 6885
rect 55802 6829 55814 6885
rect 55734 6819 55814 6829
rect 55378 6737 55434 6819
rect 55366 6735 55446 6737
rect 55366 6679 55378 6735
rect 55434 6679 55446 6735
rect 55366 6677 55446 6679
rect 54393 6619 54473 6621
rect 54393 6563 54405 6619
rect 54461 6563 54473 6619
rect 54393 6561 54473 6563
rect 54836 6619 54896 6629
rect 54836 6563 54838 6619
rect 54894 6563 54896 6619
rect 54248 6503 54328 6505
rect 54248 6447 54260 6503
rect 54316 6447 54328 6503
rect 54248 6445 54328 6447
rect 54260 6363 54316 6445
rect 53880 6353 53960 6363
rect 53880 6297 53892 6353
rect 53948 6297 53960 6353
rect 53880 6287 53960 6297
rect 54064 6353 54144 6363
rect 54064 6297 54076 6353
rect 54132 6297 54144 6353
rect 54064 6287 54144 6297
rect 54248 6353 54328 6363
rect 54248 6297 54260 6353
rect 54316 6297 54328 6353
rect 54248 6287 54328 6297
rect 54393 6231 54461 6561
rect 54836 6551 54896 6563
rect 54352 6223 54461 6231
rect 54340 6221 54461 6223
rect 54340 6101 54352 6221
rect 54408 6101 54461 6221
rect 54340 6099 54461 6101
rect 54352 6091 54408 6099
rect 53655 5834 54551 5846
rect 53655 5778 53667 5834
rect 53723 5778 54485 5834
rect 54541 5778 54551 5834
rect 53655 5766 54551 5778
rect 54838 5608 54894 6551
rect 55378 6363 55434 6677
rect 55562 6621 55618 6819
rect 55550 6619 55630 6621
rect 55550 6563 55562 6619
rect 55618 6563 55630 6619
rect 55550 6561 55630 6563
rect 55562 6363 55618 6561
rect 55746 6505 55802 6819
rect 55879 6621 55947 6951
rect 55879 6619 55959 6621
rect 55879 6563 55891 6619
rect 55947 6563 55959 6619
rect 55879 6561 55959 6563
rect 56146 6619 56216 6631
rect 56846 6619 56902 9891
rect 56146 6563 56148 6619
rect 56204 6563 56902 6619
rect 55734 6503 55814 6505
rect 55734 6447 55746 6503
rect 55802 6447 55814 6503
rect 55734 6445 55814 6447
rect 55746 6363 55802 6445
rect 55366 6353 55446 6363
rect 55366 6297 55378 6353
rect 55434 6297 55446 6353
rect 55366 6287 55446 6297
rect 55550 6353 55630 6363
rect 55550 6297 55562 6353
rect 55618 6297 55630 6353
rect 55550 6287 55630 6297
rect 55734 6353 55814 6363
rect 55734 6297 55746 6353
rect 55802 6297 55814 6353
rect 55734 6287 55814 6297
rect 55879 6231 55947 6561
rect 56146 6553 56216 6563
rect 55838 6223 55947 6231
rect 55826 6221 55947 6223
rect 55826 6101 55838 6221
rect 55894 6101 55947 6221
rect 55826 6099 55947 6101
rect 55838 6091 55894 6099
rect 55141 5834 56037 5846
rect 55141 5778 55153 5834
rect 55209 5778 55971 5834
rect 56027 5778 56037 5834
rect 55141 5766 56037 5778
rect 56148 5609 56204 6553
rect 56312 5717 56392 5727
rect 56312 5661 56324 5717
rect 56380 5661 56392 5717
rect 56312 5659 56392 5661
rect 54836 5606 54906 5608
rect 54836 5550 54838 5606
rect 54894 5550 54906 5606
rect 54836 5538 54906 5550
rect 56136 5607 56216 5609
rect 56136 5551 56148 5607
rect 56204 5551 56216 5607
rect 56136 5539 56216 5551
rect 53800 5499 54546 5511
rect 53800 5443 54168 5499
rect 54224 5443 54546 5499
rect 53800 5431 54546 5443
rect 53800 5178 53856 5431
rect 54168 5178 54224 5431
rect 54490 5178 54546 5431
rect 55286 5500 56032 5512
rect 55286 5444 55654 5500
rect 55710 5444 56032 5500
rect 55286 5432 56032 5444
rect 55286 5179 55342 5432
rect 55654 5179 55710 5432
rect 55976 5179 56032 5432
rect 53788 5176 53868 5178
rect 53788 5056 53800 5176
rect 53856 5056 53868 5176
rect 53788 5054 53868 5056
rect 54156 5176 54236 5178
rect 54156 5056 54168 5176
rect 54224 5056 54236 5176
rect 54156 5054 54236 5056
rect 54478 5176 54558 5178
rect 54478 5055 54490 5176
rect 54546 5055 54558 5176
rect 55274 5177 55354 5179
rect 55274 5057 55286 5177
rect 55342 5057 55354 5177
rect 55274 5055 55354 5057
rect 55642 5177 55722 5179
rect 55642 5057 55654 5177
rect 55710 5057 55722 5177
rect 55642 5055 55722 5057
rect 55964 5177 56044 5179
rect 55964 5056 55976 5177
rect 56032 5056 56044 5177
rect 53800 5046 53856 5054
rect 54168 5046 54224 5054
rect 54478 5053 54558 5055
rect 54490 5045 54546 5053
rect 55286 5047 55342 5055
rect 55654 5047 55710 5055
rect 55964 5054 56044 5056
rect 55976 5046 56032 5054
rect 53984 4878 54040 4886
rect 54352 4878 54408 4886
rect 55470 4879 55526 4887
rect 55838 4879 55894 4887
rect 53972 4876 54461 4878
rect 53972 4756 53984 4876
rect 54040 4756 54352 4876
rect 54408 4756 54461 4876
rect 53972 4754 54461 4756
rect 55458 4877 55947 4879
rect 55458 4757 55470 4877
rect 55526 4757 55838 4877
rect 55894 4757 55947 4877
rect 55458 4755 55947 4757
rect 53984 4746 54040 4754
rect 54352 4746 54461 4754
rect 55470 4747 55526 4755
rect 55838 4747 55947 4755
rect 53880 4680 53960 4690
rect 53880 4624 53892 4680
rect 53948 4624 53960 4680
rect 53880 4614 53960 4624
rect 54064 4680 54144 4690
rect 54064 4624 54076 4680
rect 54132 4624 54144 4680
rect 54064 4614 54144 4624
rect 54248 4680 54328 4690
rect 54248 4624 54260 4680
rect 54316 4624 54328 4680
rect 54248 4614 54328 4624
rect 53892 4532 53948 4614
rect 53880 4530 53960 4532
rect 53880 4474 53892 4530
rect 53948 4474 53960 4530
rect 53880 4472 53960 4474
rect 53208 4298 53278 4310
rect 53208 4242 53220 4298
rect 53276 4242 53278 4298
rect 53208 4230 53278 4242
rect 53892 4158 53948 4472
rect 54076 4416 54132 4614
rect 54064 4414 54144 4416
rect 54064 4358 54076 4414
rect 54132 4358 54144 4414
rect 54064 4356 54144 4358
rect 54076 4158 54132 4356
rect 54260 4300 54316 4614
rect 54393 4416 54461 4746
rect 55366 4681 55446 4691
rect 55366 4625 55378 4681
rect 55434 4625 55446 4681
rect 55366 4615 55446 4625
rect 55550 4681 55630 4691
rect 55550 4625 55562 4681
rect 55618 4625 55630 4681
rect 55550 4615 55630 4625
rect 55734 4681 55814 4691
rect 55734 4625 55746 4681
rect 55802 4625 55814 4681
rect 55734 4615 55814 4625
rect 55378 4533 55434 4615
rect 55366 4531 55446 4533
rect 55366 4475 55378 4531
rect 55434 4475 55446 4531
rect 55366 4473 55446 4475
rect 54393 4414 54473 4416
rect 54393 4358 54405 4414
rect 54461 4358 54473 4414
rect 54393 4356 54473 4358
rect 54660 4414 54730 4426
rect 54660 4358 54662 4414
rect 54718 4358 54730 4414
rect 54248 4298 54328 4300
rect 54248 4242 54260 4298
rect 54316 4242 54328 4298
rect 54248 4240 54328 4242
rect 54260 4158 54316 4240
rect 53880 4148 53960 4158
rect 53880 4092 53892 4148
rect 53948 4092 53960 4148
rect 53880 4082 53960 4092
rect 54064 4148 54144 4158
rect 54064 4092 54076 4148
rect 54132 4092 54144 4148
rect 54064 4082 54144 4092
rect 54248 4148 54328 4158
rect 54248 4092 54260 4148
rect 54316 4092 54328 4148
rect 54248 4082 54328 4092
rect 54393 4026 54461 4356
rect 54660 4348 54730 4358
rect 54352 4018 54461 4026
rect 54340 4016 54461 4018
rect 54340 3896 54352 4016
rect 54408 3896 54461 4016
rect 54340 3894 54461 3896
rect 54352 3886 54408 3894
rect 53655 3629 54551 3641
rect 53655 3573 53667 3629
rect 53723 3573 54485 3629
rect 54541 3573 54551 3629
rect 53655 3561 54551 3573
rect 54662 3404 54718 4348
rect 55378 4159 55434 4473
rect 55562 4417 55618 4615
rect 55550 4415 55630 4417
rect 55550 4359 55562 4415
rect 55618 4359 55630 4415
rect 55550 4357 55630 4359
rect 55562 4159 55618 4357
rect 55746 4301 55802 4615
rect 55879 4417 55947 4747
rect 56324 4425 56380 5659
rect 55879 4415 55959 4417
rect 55879 4359 55891 4415
rect 55947 4359 55959 4415
rect 55879 4357 55959 4359
rect 56322 4415 56392 4425
rect 56322 4359 56324 4415
rect 56380 4359 56472 4415
rect 55734 4299 55814 4301
rect 55734 4243 55746 4299
rect 55802 4243 55814 4299
rect 55734 4241 55814 4243
rect 55746 4159 55802 4241
rect 55366 4149 55446 4159
rect 55366 4093 55378 4149
rect 55434 4093 55446 4149
rect 55366 4083 55446 4093
rect 55550 4149 55630 4159
rect 55550 4093 55562 4149
rect 55618 4093 55630 4149
rect 55550 4083 55630 4093
rect 55734 4149 55814 4159
rect 55734 4093 55746 4149
rect 55802 4093 55814 4149
rect 55734 4083 55814 4093
rect 55879 4027 55947 4357
rect 56322 4347 56392 4359
rect 55838 4019 55947 4027
rect 55826 4017 55947 4019
rect 55826 3897 55838 4017
rect 55894 3897 55947 4017
rect 55826 3895 55947 3897
rect 55838 3887 55894 3895
rect 55141 3630 56037 3642
rect 55141 3574 55153 3630
rect 55209 3574 55971 3630
rect 56027 3574 56037 3630
rect 55141 3562 56037 3574
rect 54826 3511 54906 3521
rect 54826 3455 54838 3511
rect 54894 3455 54906 3511
rect 54826 3453 54906 3455
rect 54660 3401 54730 3404
rect 54660 3347 54662 3401
rect 54718 3347 54730 3401
rect 54660 3335 54730 3347
rect 53800 3294 54546 3306
rect 53800 3238 54168 3294
rect 54224 3238 54546 3294
rect 53800 3226 54546 3238
rect 53800 2973 53856 3226
rect 54168 2973 54224 3226
rect 54490 2973 54546 3226
rect 53788 2971 53868 2973
rect 53788 2851 53800 2971
rect 53856 2851 53868 2971
rect 53788 2849 53868 2851
rect 54156 2971 54236 2973
rect 54156 2851 54168 2971
rect 54224 2851 54236 2971
rect 54156 2849 54236 2851
rect 54478 2971 54558 2973
rect 54478 2850 54490 2971
rect 54546 2850 54558 2971
rect 53800 2841 53856 2849
rect 54168 2841 54224 2849
rect 54478 2848 54558 2850
rect 54490 2840 54546 2848
rect 53984 2673 54040 2681
rect 54352 2673 54408 2681
rect 53972 2671 54461 2673
rect 53972 2551 53984 2671
rect 54040 2551 54352 2671
rect 54408 2551 54461 2671
rect 53972 2549 54461 2551
rect 53984 2541 54040 2549
rect 54352 2541 54461 2549
rect 53880 2475 53960 2485
rect 53880 2419 53892 2475
rect 53948 2419 53960 2475
rect 53880 2409 53960 2419
rect 54064 2475 54144 2485
rect 54064 2419 54076 2475
rect 54132 2419 54144 2475
rect 54064 2409 54144 2419
rect 54248 2475 54328 2485
rect 54248 2419 54260 2475
rect 54316 2419 54328 2475
rect 54248 2409 54328 2419
rect 53892 2327 53948 2409
rect 53880 2325 53960 2327
rect 53880 2269 53892 2325
rect 53948 2269 53960 2325
rect 53880 2267 53960 2269
rect 53072 2209 53142 2223
rect 53072 2153 53084 2209
rect 53140 2153 53142 2209
rect 53072 2141 53142 2153
rect 52838 2093 52916 2104
rect 52446 2092 52916 2093
rect 52446 2038 52850 2092
rect 52904 2038 52916 2092
rect 52446 2037 52916 2038
rect 50874 1733 52046 1743
rect 50874 1677 50886 1733
rect 50942 1677 51774 1733
rect 51830 1677 52046 1733
rect 50874 1667 52046 1677
rect 52446 1733 52526 2037
rect 52838 2026 52916 2037
rect 52446 1677 52458 1733
rect 52514 1677 52526 1733
rect 52446 1667 52526 1677
rect 50804 1355 52596 1367
rect 50804 1215 50816 1355
rect 52584 1215 52596 1355
rect 52889 1306 52975 1318
rect 53084 1310 53140 2141
rect 53892 1953 53948 2267
rect 54076 2211 54132 2409
rect 54064 2209 54144 2211
rect 54064 2153 54076 2209
rect 54132 2153 54144 2209
rect 54064 2151 54144 2153
rect 54076 1953 54132 2151
rect 54260 2095 54316 2409
rect 54393 2211 54461 2541
rect 54838 2221 54894 3453
rect 54393 2209 54473 2211
rect 54393 2153 54405 2209
rect 54461 2153 54473 2209
rect 54393 2151 54473 2153
rect 54836 2209 54896 2221
rect 54836 2153 54838 2209
rect 54894 2153 54896 2209
rect 54248 2093 54328 2095
rect 54248 2037 54260 2093
rect 54316 2037 54328 2093
rect 54248 2035 54328 2037
rect 54260 1953 54316 2035
rect 53880 1943 53960 1953
rect 53880 1887 53892 1943
rect 53948 1887 53960 1943
rect 53880 1877 53960 1887
rect 54064 1943 54144 1953
rect 54064 1887 54076 1943
rect 54132 1887 54144 1943
rect 54064 1877 54144 1887
rect 54248 1943 54328 1953
rect 54248 1887 54260 1943
rect 54316 1887 54328 1943
rect 54248 1877 54328 1887
rect 54393 1821 54461 2151
rect 54836 2141 54896 2153
rect 54352 1813 54461 1821
rect 54340 1811 54461 1813
rect 54340 1691 54352 1811
rect 54408 1691 54461 1811
rect 54340 1689 54461 1691
rect 54352 1681 54408 1689
rect 53655 1424 54553 1436
rect 53655 1368 53667 1424
rect 53723 1368 54485 1424
rect 54541 1368 54553 1424
rect 53655 1356 54553 1368
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 53082 1306 53142 1310
rect 53082 1250 53084 1306
rect 53140 1250 53142 1306
rect 53082 1238 53142 1250
rect 50804 1203 52596 1215
rect 50218 873 50575 929
rect 52174 1031 52494 1041
rect 49738 513 49750 569
rect 49806 513 49818 569
rect 49738 503 49818 513
rect 50218 569 50298 873
rect 50218 513 50230 569
rect 50286 513 50298 569
rect 50218 503 50298 513
rect 48850 255 49614 327
rect 52174 231 52184 1031
rect 52484 231 52494 1031
rect 52174 221 52494 231
<< via2 >>
rect 6808 9852 6864 9908
rect 16280 9852 16336 9908
rect 25752 9853 25808 9909
rect 35224 9853 35280 9909
rect 44696 9853 44752 9909
rect 54168 9853 54224 9909
rect 5644 8883 5700 8939
rect 5444 5660 5500 5716
rect 952 3290 1008 3346
rect 1982 2852 2038 2908
rect 4824 3510 5124 4310
rect 2390 2852 2446 2908
rect 1166 2431 1246 2507
rect 2396 2400 2996 2540
rect 3456 3174 5224 3314
rect 2396 2000 2996 2140
rect -441 -171 -385 -51
rect 1982 512 2038 568
rect 15116 8883 15172 8939
rect 6307 7982 6363 8038
rect 7125 7982 7181 8038
rect 6808 7647 6864 7703
rect 8294 7647 8350 7703
rect 6307 5777 6363 5833
rect 7125 5777 7181 5833
rect 7793 5777 7849 5833
rect 8611 5777 8667 5833
rect 6808 5442 6864 5498
rect 8294 5443 8350 5499
rect 6307 3572 6363 3628
rect 7125 3572 7181 3628
rect 7793 3573 7849 3629
rect 8611 3573 8667 3629
rect 6808 3237 6864 3293
rect 3456 1214 5224 1354
rect 14916 5660 14972 5716
rect 9906 3510 10106 4310
rect 11454 2852 11510 2908
rect 14296 3510 14596 4310
rect 11862 2852 11918 2908
rect 11868 2400 12468 2540
rect 12928 3174 14696 3314
rect 6307 1367 6363 1423
rect 7125 1367 7181 1423
rect 5541 1249 5597 1305
rect 2390 512 2446 568
rect 4824 230 5124 1030
rect 11868 2000 12468 2140
rect 9087 -170 9143 -50
rect 11454 512 11510 568
rect 24588 8884 24644 8940
rect 15779 7982 15835 8038
rect 16597 7982 16653 8038
rect 16280 7647 16336 7703
rect 17766 7647 17822 7703
rect 15779 5777 15835 5833
rect 16597 5777 16653 5833
rect 17265 5777 17321 5833
rect 18083 5777 18139 5833
rect 16280 5442 16336 5498
rect 17766 5443 17822 5499
rect 15779 3572 15835 3628
rect 16597 3572 16653 3628
rect 17265 3573 17321 3629
rect 18083 3573 18139 3629
rect 16280 3237 16336 3293
rect 12928 1214 14696 1354
rect 24388 5661 24444 5717
rect 19378 3511 19578 4311
rect 20926 2853 20982 2909
rect 23768 3511 24068 4311
rect 21334 2853 21390 2909
rect 21340 2401 21940 2541
rect 22400 3175 24168 3315
rect 15779 1367 15835 1423
rect 16597 1367 16653 1423
rect 15013 1249 15069 1305
rect 11862 512 11918 568
rect 14296 230 14596 1030
rect 21340 2001 21940 2141
rect 18559 -170 18615 -50
rect 20926 513 20982 569
rect 34060 8884 34116 8940
rect 25251 7983 25307 8039
rect 26069 7983 26125 8039
rect 25752 7648 25808 7704
rect 27238 7648 27294 7704
rect 25251 5778 25307 5834
rect 26069 5778 26125 5834
rect 26737 5778 26793 5834
rect 27555 5778 27611 5834
rect 25752 5443 25808 5499
rect 27238 5444 27294 5500
rect 25251 3573 25307 3629
rect 26069 3573 26125 3629
rect 26737 3574 26793 3630
rect 27555 3574 27611 3630
rect 25752 3238 25808 3294
rect 22400 1215 24168 1355
rect 33860 5661 33916 5717
rect 28850 3511 29050 4311
rect 30398 2853 30454 2909
rect 33240 3511 33540 4311
rect 30806 2853 30862 2909
rect 30812 2401 31412 2541
rect 31872 3175 33640 3315
rect 25251 1368 25307 1424
rect 26069 1368 26125 1424
rect 24485 1250 24541 1306
rect 21334 513 21390 569
rect 23768 231 24068 1031
rect 30812 2001 31412 2141
rect 28031 -169 28087 -49
rect 30398 513 30454 569
rect 43532 8884 43588 8940
rect 34723 7983 34779 8039
rect 35541 7983 35597 8039
rect 35224 7648 35280 7704
rect 36710 7648 36766 7704
rect 34723 5778 34779 5834
rect 35541 5778 35597 5834
rect 36209 5778 36265 5834
rect 37027 5778 37083 5834
rect 35224 5443 35280 5499
rect 36710 5444 36766 5500
rect 34723 3573 34779 3629
rect 35541 3573 35597 3629
rect 36209 3574 36265 3630
rect 37027 3574 37083 3630
rect 35224 3238 35280 3294
rect 31872 1215 33640 1355
rect 43332 5661 43388 5717
rect 38322 3511 38522 4311
rect 39870 2853 39926 2909
rect 42712 3511 43012 4311
rect 40278 2853 40334 2909
rect 40284 2401 40884 2541
rect 41344 3175 43112 3315
rect 34723 1368 34779 1424
rect 35541 1368 35597 1424
rect 33957 1250 34013 1306
rect 30806 513 30862 569
rect 33240 231 33540 1031
rect 40284 2001 40884 2141
rect 37503 -169 37559 -49
rect 39870 513 39926 569
rect 53004 8884 53060 8940
rect 44195 7983 44251 8039
rect 45013 7983 45069 8039
rect 44696 7648 44752 7704
rect 46182 7648 46238 7704
rect 44195 5778 44251 5834
rect 45013 5778 45069 5834
rect 45681 5778 45737 5834
rect 46499 5778 46555 5834
rect 44696 5443 44752 5499
rect 46182 5444 46238 5500
rect 44195 3573 44251 3629
rect 45013 3573 45069 3629
rect 45681 3574 45737 3630
rect 46499 3574 46555 3630
rect 44696 3238 44752 3294
rect 41344 1215 43112 1355
rect 52804 5661 52860 5717
rect 47794 3511 47994 4311
rect 49342 2853 49398 2909
rect 52184 3511 52484 4311
rect 49750 2853 49806 2909
rect 49756 2401 50356 2541
rect 50816 3175 52584 3315
rect 44195 1368 44251 1424
rect 45013 1368 45069 1424
rect 43429 1250 43485 1306
rect 40278 513 40334 569
rect 42712 231 43012 1031
rect 49756 2001 50356 2141
rect 46975 -169 47031 -49
rect 49342 513 49398 569
rect 53667 7983 53723 8039
rect 54485 7983 54541 8039
rect 54168 7648 54224 7704
rect 55654 7648 55710 7704
rect 53667 5778 53723 5834
rect 54485 5778 54541 5834
rect 55153 5778 55209 5834
rect 55971 5778 56027 5834
rect 54168 5443 54224 5499
rect 55654 5444 55710 5500
rect 53667 3573 53723 3629
rect 54485 3573 54541 3629
rect 55153 3574 55209 3630
rect 55971 3574 56027 3630
rect 54168 3238 54224 3294
rect 50816 1215 52584 1355
rect 53667 1368 53723 1424
rect 54485 1368 54541 1424
rect 52901 1250 52957 1306
rect 49750 513 49806 569
rect 52184 231 52484 1031
<< metal3 >>
rect 6796 9908 6882 9912
rect 6796 9852 6808 9908
rect 6864 9852 6882 9908
rect 6796 9840 6882 9852
rect 16268 9908 16354 9912
rect 16268 9852 16280 9908
rect 16336 9852 16354 9908
rect 16268 9840 16354 9852
rect 25740 9909 25826 9913
rect 25740 9853 25752 9909
rect 25808 9853 25826 9909
rect 25740 9841 25826 9853
rect 35212 9909 35298 9913
rect 35212 9853 35224 9909
rect 35280 9853 35298 9909
rect 35212 9841 35298 9853
rect 44684 9909 44770 9913
rect 44684 9853 44696 9909
rect 44752 9853 44770 9909
rect 44684 9841 44770 9853
rect 54156 9909 54242 9913
rect 54156 9853 54168 9909
rect 54224 9853 54242 9909
rect 54156 9841 54242 9853
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 6295 8038 6375 8050
rect 6295 7982 6307 8038
rect 6363 7982 6375 8038
rect 6295 7970 6375 7982
rect 7113 8038 7193 8050
rect 7113 7982 7125 8038
rect 7181 7982 7193 8038
rect 7113 7970 7193 7982
rect 15767 8038 15847 8050
rect 15767 7982 15779 8038
rect 15835 7982 15847 8038
rect 15767 7970 15847 7982
rect 16585 8038 16665 8050
rect 16585 7982 16597 8038
rect 16653 7982 16665 8038
rect 16585 7970 16665 7982
rect 25239 8039 25319 8051
rect 25239 7983 25251 8039
rect 25307 7983 25319 8039
rect 25239 7971 25319 7983
rect 26057 8039 26137 8051
rect 26057 7983 26069 8039
rect 26125 7983 26137 8039
rect 26057 7971 26137 7983
rect 34711 8039 34791 8051
rect 34711 7983 34723 8039
rect 34779 7983 34791 8039
rect 34711 7971 34791 7983
rect 35529 8039 35609 8051
rect 35529 7983 35541 8039
rect 35597 7983 35609 8039
rect 35529 7971 35609 7983
rect 44183 8039 44263 8051
rect 44183 7983 44195 8039
rect 44251 7983 44263 8039
rect 44183 7971 44263 7983
rect 45001 8039 45081 8051
rect 45001 7983 45013 8039
rect 45069 7983 45081 8039
rect 45001 7971 45081 7983
rect 53655 8039 53735 8051
rect 53655 7983 53667 8039
rect 53723 7983 53735 8039
rect 53655 7971 53735 7983
rect 54473 8039 54553 8051
rect 54473 7983 54485 8039
rect 54541 7983 54553 8039
rect 54473 7971 54553 7983
rect 6796 7703 6882 7707
rect 6796 7647 6808 7703
rect 6864 7647 6882 7703
rect 6796 7635 6882 7647
rect 8282 7703 8368 7707
rect 8282 7647 8294 7703
rect 8350 7647 8368 7703
rect 8282 7635 8368 7647
rect 16268 7703 16354 7707
rect 16268 7647 16280 7703
rect 16336 7647 16354 7703
rect 16268 7635 16354 7647
rect 17754 7703 17840 7707
rect 17754 7647 17766 7703
rect 17822 7647 17840 7703
rect 17754 7635 17840 7647
rect 25740 7704 25826 7708
rect 25740 7648 25752 7704
rect 25808 7648 25826 7704
rect 25740 7636 25826 7648
rect 27226 7704 27312 7708
rect 27226 7648 27238 7704
rect 27294 7648 27312 7704
rect 27226 7636 27312 7648
rect 35212 7704 35298 7708
rect 35212 7648 35224 7704
rect 35280 7648 35298 7704
rect 35212 7636 35298 7648
rect 36698 7704 36784 7708
rect 36698 7648 36710 7704
rect 36766 7648 36784 7704
rect 36698 7636 36784 7648
rect 44684 7704 44770 7708
rect 44684 7648 44696 7704
rect 44752 7648 44770 7704
rect 44684 7636 44770 7648
rect 46170 7704 46256 7708
rect 46170 7648 46182 7704
rect 46238 7648 46256 7704
rect 46170 7636 46256 7648
rect 54156 7704 54242 7708
rect 54156 7648 54168 7704
rect 54224 7648 54242 7704
rect 54156 7636 54242 7648
rect 55642 7704 55728 7708
rect 55642 7648 55654 7704
rect 55710 7648 55728 7704
rect 55642 7636 55728 7648
rect 6295 5833 6375 5845
rect 6295 5777 6307 5833
rect 6363 5777 6375 5833
rect 6295 5765 6375 5777
rect 7113 5833 7193 5845
rect 7113 5777 7125 5833
rect 7181 5777 7193 5833
rect 7113 5765 7193 5777
rect 7781 5833 7861 5845
rect 7781 5777 7793 5833
rect 7849 5777 7861 5833
rect 7781 5765 7861 5777
rect 8599 5833 8679 5845
rect 8599 5777 8611 5833
rect 8667 5777 8679 5833
rect 8599 5765 8679 5777
rect 15767 5833 15847 5845
rect 15767 5777 15779 5833
rect 15835 5777 15847 5833
rect 15767 5765 15847 5777
rect 16585 5833 16665 5845
rect 16585 5777 16597 5833
rect 16653 5777 16665 5833
rect 16585 5765 16665 5777
rect 17253 5833 17333 5845
rect 17253 5777 17265 5833
rect 17321 5777 17333 5833
rect 17253 5765 17333 5777
rect 18071 5833 18151 5845
rect 18071 5777 18083 5833
rect 18139 5777 18151 5833
rect 18071 5765 18151 5777
rect 25239 5834 25319 5846
rect 25239 5778 25251 5834
rect 25307 5778 25319 5834
rect 25239 5766 25319 5778
rect 26057 5834 26137 5846
rect 26057 5778 26069 5834
rect 26125 5778 26137 5834
rect 26057 5766 26137 5778
rect 26725 5834 26805 5846
rect 26725 5778 26737 5834
rect 26793 5778 26805 5834
rect 26725 5766 26805 5778
rect 27543 5834 27623 5846
rect 27543 5778 27555 5834
rect 27611 5778 27623 5834
rect 27543 5766 27623 5778
rect 34711 5834 34791 5846
rect 34711 5778 34723 5834
rect 34779 5778 34791 5834
rect 34711 5766 34791 5778
rect 35529 5834 35609 5846
rect 35529 5778 35541 5834
rect 35597 5778 35609 5834
rect 35529 5766 35609 5778
rect 36197 5834 36277 5846
rect 36197 5778 36209 5834
rect 36265 5778 36277 5834
rect 36197 5766 36277 5778
rect 37015 5834 37095 5846
rect 37015 5778 37027 5834
rect 37083 5778 37095 5834
rect 37015 5766 37095 5778
rect 44183 5834 44263 5846
rect 44183 5778 44195 5834
rect 44251 5778 44263 5834
rect 44183 5766 44263 5778
rect 45001 5834 45081 5846
rect 45001 5778 45013 5834
rect 45069 5778 45081 5834
rect 45001 5766 45081 5778
rect 45669 5834 45749 5846
rect 45669 5778 45681 5834
rect 45737 5778 45749 5834
rect 45669 5766 45749 5778
rect 46487 5834 46567 5846
rect 46487 5778 46499 5834
rect 46555 5778 46567 5834
rect 46487 5766 46567 5778
rect 53655 5834 53735 5846
rect 53655 5778 53667 5834
rect 53723 5778 53735 5834
rect 53655 5766 53735 5778
rect 54473 5834 54553 5846
rect 54473 5778 54485 5834
rect 54541 5778 54553 5834
rect 54473 5766 54553 5778
rect 55141 5834 55221 5846
rect 55141 5778 55153 5834
rect 55209 5778 55221 5834
rect 55141 5766 55221 5778
rect 55959 5834 56039 5846
rect 55959 5778 55971 5834
rect 56027 5778 56039 5834
rect 55959 5766 56039 5778
rect 5430 5716 5512 5728
rect 3058 5660 5444 5716
rect 5500 5709 5512 5716
rect 14902 5716 14984 5728
rect 14902 5709 14916 5716
rect 5500 5660 14916 5709
rect 14972 5709 14984 5716
rect 24374 5717 24456 5729
rect 24374 5709 24388 5717
rect 14972 5661 24388 5709
rect 24444 5709 24456 5717
rect 33846 5717 33928 5729
rect 33846 5709 33860 5717
rect 24444 5661 33860 5709
rect 33916 5709 33928 5717
rect 43318 5717 43400 5729
rect 43318 5709 43332 5717
rect 33916 5661 43332 5709
rect 43388 5709 43400 5717
rect 52790 5717 52872 5729
rect 52790 5709 52804 5717
rect 43388 5661 52804 5709
rect 52860 5661 52872 5717
rect 14972 5660 52872 5661
rect 3058 5655 52872 5660
rect 5430 5649 52872 5655
rect 5430 5648 52790 5649
rect 6796 5498 6882 5502
rect 6796 5442 6808 5498
rect 6864 5442 6882 5498
rect 6796 5430 6882 5442
rect 8282 5499 8368 5503
rect 8282 5443 8294 5499
rect 8350 5443 8368 5499
rect 8282 5431 8368 5443
rect 16268 5498 16354 5502
rect 16268 5442 16280 5498
rect 16336 5442 16354 5498
rect 16268 5430 16354 5442
rect 17754 5499 17840 5503
rect 17754 5443 17766 5499
rect 17822 5443 17840 5499
rect 17754 5431 17840 5443
rect 25740 5499 25826 5503
rect 25740 5443 25752 5499
rect 25808 5443 25826 5499
rect 25740 5431 25826 5443
rect 27226 5500 27312 5504
rect 27226 5444 27238 5500
rect 27294 5444 27312 5500
rect 27226 5432 27312 5444
rect 35212 5499 35298 5503
rect 35212 5443 35224 5499
rect 35280 5443 35298 5499
rect 35212 5431 35298 5443
rect 36698 5500 36784 5504
rect 36698 5444 36710 5500
rect 36766 5444 36784 5500
rect 36698 5432 36784 5444
rect 44684 5499 44770 5503
rect 44684 5443 44696 5499
rect 44752 5443 44770 5499
rect 44684 5431 44770 5443
rect 46170 5500 46256 5504
rect 46170 5444 46182 5500
rect 46238 5444 46256 5500
rect 46170 5432 46256 5444
rect 54156 5499 54242 5503
rect 54156 5443 54168 5499
rect 54224 5443 54242 5499
rect 54156 5431 54242 5443
rect 55642 5500 55728 5504
rect 55642 5444 55654 5500
rect 55710 5444 55728 5500
rect 55642 5432 55728 5444
rect 4814 4310 5134 4320
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 9896 4310 10116 4320
rect 6295 3628 6375 3640
rect 6295 3572 6307 3628
rect 6363 3572 6375 3628
rect 6295 3560 6375 3572
rect 7113 3628 7193 3640
rect 7113 3572 7125 3628
rect 7181 3572 7193 3628
rect 7113 3560 7193 3572
rect 7781 3629 7861 3641
rect 7781 3573 7793 3629
rect 7849 3573 7861 3629
rect 7781 3561 7861 3573
rect 8599 3629 8679 3641
rect 8599 3573 8611 3629
rect 8667 3573 8679 3629
rect 8599 3561 8679 3573
rect 4814 3500 5134 3510
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 9896 3500 10116 3510
rect 14286 4310 14606 4320
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 19368 4311 19588 4321
rect 15767 3628 15847 3640
rect 15767 3572 15779 3628
rect 15835 3572 15847 3628
rect 15767 3560 15847 3572
rect 16585 3628 16665 3640
rect 16585 3572 16597 3628
rect 16653 3572 16665 3628
rect 16585 3560 16665 3572
rect 17253 3629 17333 3641
rect 17253 3573 17265 3629
rect 17321 3573 17333 3629
rect 17253 3561 17333 3573
rect 18071 3629 18151 3641
rect 18071 3573 18083 3629
rect 18139 3573 18151 3629
rect 18071 3561 18151 3573
rect 14286 3500 14606 3510
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 19368 3501 19588 3511
rect 23758 4311 24078 4321
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 28840 4311 29060 4321
rect 25239 3629 25319 3641
rect 25239 3573 25251 3629
rect 25307 3573 25319 3629
rect 25239 3561 25319 3573
rect 26057 3629 26137 3641
rect 26057 3573 26069 3629
rect 26125 3573 26137 3629
rect 26057 3561 26137 3573
rect 26725 3630 26805 3642
rect 26725 3574 26737 3630
rect 26793 3574 26805 3630
rect 26725 3562 26805 3574
rect 27543 3630 27623 3642
rect 27543 3574 27555 3630
rect 27611 3574 27623 3630
rect 27543 3562 27623 3574
rect 23758 3501 24078 3511
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 28840 3501 29060 3511
rect 33230 4311 33550 4321
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 38312 4311 38532 4321
rect 34711 3629 34791 3641
rect 34711 3573 34723 3629
rect 34779 3573 34791 3629
rect 34711 3561 34791 3573
rect 35529 3629 35609 3641
rect 35529 3573 35541 3629
rect 35597 3573 35609 3629
rect 35529 3561 35609 3573
rect 36197 3630 36277 3642
rect 36197 3574 36209 3630
rect 36265 3574 36277 3630
rect 36197 3562 36277 3574
rect 37015 3630 37095 3642
rect 37015 3574 37027 3630
rect 37083 3574 37095 3630
rect 37015 3562 37095 3574
rect 33230 3501 33550 3511
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 38312 3501 38532 3511
rect 42702 4311 43022 4321
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 47784 4311 48004 4321
rect 44183 3629 44263 3641
rect 44183 3573 44195 3629
rect 44251 3573 44263 3629
rect 44183 3561 44263 3573
rect 45001 3629 45081 3641
rect 45001 3573 45013 3629
rect 45069 3573 45081 3629
rect 45001 3561 45081 3573
rect 45669 3630 45749 3642
rect 45669 3574 45681 3630
rect 45737 3574 45749 3630
rect 45669 3562 45749 3574
rect 46487 3630 46567 3642
rect 46487 3574 46499 3630
rect 46555 3574 46567 3630
rect 46487 3562 46567 3574
rect 42702 3501 43022 3511
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 47784 3501 48004 3511
rect 52174 4311 52494 4321
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 53655 3629 53735 3641
rect 53655 3573 53667 3629
rect 53723 3573 53735 3629
rect 53655 3561 53735 3573
rect 54473 3629 54553 3641
rect 54473 3573 54485 3629
rect 54541 3573 54553 3629
rect 54473 3561 54553 3573
rect 55141 3630 55221 3642
rect 55141 3574 55153 3630
rect 55209 3574 55221 3630
rect 55141 3562 55221 3574
rect 55959 3630 56039 3642
rect 55959 3574 55971 3630
rect 56027 3574 56039 3630
rect 55959 3562 56039 3574
rect 52174 3501 52494 3511
rect 940 3346 1020 3356
rect 940 3290 952 3346
rect 1008 3290 1020 3346
rect 940 2517 1020 3290
rect 3444 3314 5236 3326
rect 3444 3174 3456 3314
rect 5224 3174 5236 3314
rect 12916 3314 14708 3326
rect 6796 3293 6882 3297
rect 6796 3237 6808 3293
rect 6864 3237 6882 3293
rect 6796 3225 6882 3237
rect 1970 2908 2458 2918
rect 1970 2852 1982 2908
rect 2038 2852 2390 2908
rect 2446 2852 2458 2908
rect 1970 2842 2458 2852
rect 2384 2540 3008 2552
rect 940 2507 1256 2517
rect 940 2431 1166 2507
rect 1246 2431 1256 2507
rect 940 2421 1256 2431
rect 2384 2400 2396 2540
rect 2996 2400 3008 2540
rect 2384 2388 3008 2400
rect 3444 2152 5236 3174
rect 12916 3174 12928 3314
rect 14696 3174 14708 3314
rect 22388 3315 24180 3327
rect 16268 3293 16354 3297
rect 16268 3237 16280 3293
rect 16336 3237 16354 3293
rect 16268 3225 16354 3237
rect 11442 2908 11930 2918
rect 11442 2852 11454 2908
rect 11510 2852 11862 2908
rect 11918 2852 11930 2908
rect 11442 2842 11930 2852
rect 11856 2540 12480 2552
rect 11856 2400 11868 2540
rect 12468 2400 12480 2540
rect 11856 2388 12480 2400
rect 12916 2152 14708 3174
rect 22388 3175 22400 3315
rect 24168 3175 24180 3315
rect 31860 3315 33652 3327
rect 25740 3294 25826 3298
rect 25740 3238 25752 3294
rect 25808 3238 25826 3294
rect 25740 3226 25826 3238
rect 20914 2909 21402 2919
rect 20914 2853 20926 2909
rect 20982 2853 21334 2909
rect 21390 2853 21402 2909
rect 20914 2843 21402 2853
rect 21328 2541 21952 2553
rect 21328 2401 21340 2541
rect 21940 2401 21952 2541
rect 21328 2389 21952 2401
rect 22388 2153 24180 3175
rect 31860 3175 31872 3315
rect 33640 3175 33652 3315
rect 41332 3315 43124 3327
rect 35212 3294 35298 3298
rect 35212 3238 35224 3294
rect 35280 3238 35298 3294
rect 35212 3226 35298 3238
rect 30386 2909 30874 2919
rect 30386 2853 30398 2909
rect 30454 2853 30806 2909
rect 30862 2853 30874 2909
rect 30386 2843 30874 2853
rect 30800 2541 31424 2553
rect 30800 2401 30812 2541
rect 31412 2401 31424 2541
rect 30800 2389 31424 2401
rect 31860 2153 33652 3175
rect 41332 3175 41344 3315
rect 43112 3175 43124 3315
rect 50804 3315 52596 3327
rect 44684 3294 44770 3298
rect 44684 3238 44696 3294
rect 44752 3238 44770 3294
rect 44684 3226 44770 3238
rect 39858 2909 40346 2919
rect 39858 2853 39870 2909
rect 39926 2853 40278 2909
rect 40334 2853 40346 2909
rect 39858 2843 40346 2853
rect 40272 2541 40896 2553
rect 40272 2401 40284 2541
rect 40884 2401 40896 2541
rect 40272 2389 40896 2401
rect 41332 2153 43124 3175
rect 50804 3175 50816 3315
rect 52584 3175 52596 3315
rect 54156 3294 54242 3298
rect 54156 3238 54168 3294
rect 54224 3238 54242 3294
rect 54156 3226 54242 3238
rect 49330 2909 49818 2919
rect 49330 2853 49342 2909
rect 49398 2853 49750 2909
rect 49806 2853 49818 2909
rect 49330 2843 49818 2853
rect 49744 2541 50368 2553
rect 49744 2401 49756 2541
rect 50356 2401 50368 2541
rect 49744 2389 50368 2401
rect 50804 2153 52596 3175
rect 2384 2140 5236 2152
rect 2384 2000 2396 2140
rect 2996 2000 5236 2140
rect 2384 1988 5236 2000
rect 11856 2140 14708 2152
rect 11856 2000 11868 2140
rect 12468 2000 14708 2140
rect 11856 1988 14708 2000
rect 21328 2141 24180 2153
rect 21328 2001 21340 2141
rect 21940 2001 24180 2141
rect 21328 1989 24180 2001
rect 30800 2141 33652 2153
rect 30800 2001 30812 2141
rect 31412 2001 33652 2141
rect 30800 1989 33652 2001
rect 40272 2141 43124 2153
rect 40272 2001 40284 2141
rect 40884 2001 43124 2141
rect 40272 1989 43124 2001
rect 49744 2141 52596 2153
rect 49744 2001 49756 2141
rect 50356 2001 52596 2141
rect 49744 1989 52596 2001
rect 6295 1423 6375 1435
rect 6295 1367 6307 1423
rect 6363 1367 6375 1423
rect 3444 1354 5236 1366
rect 6295 1355 6375 1367
rect 7113 1423 7193 1435
rect 7113 1367 7125 1423
rect 7181 1367 7193 1423
rect 7113 1355 7193 1367
rect 15767 1423 15847 1435
rect 15767 1367 15779 1423
rect 15835 1367 15847 1423
rect 3444 1214 3456 1354
rect 5224 1214 5236 1354
rect 12916 1354 14708 1366
rect 15767 1355 15847 1367
rect 16585 1423 16665 1435
rect 16585 1367 16597 1423
rect 16653 1367 16665 1423
rect 25239 1424 25319 1436
rect 25239 1368 25251 1424
rect 25307 1368 25319 1424
rect 16585 1355 16665 1367
rect 22388 1355 24180 1367
rect 25239 1356 25319 1368
rect 26057 1424 26137 1436
rect 26057 1368 26069 1424
rect 26125 1368 26137 1424
rect 26057 1356 26137 1368
rect 34711 1424 34791 1436
rect 34711 1368 34723 1424
rect 34779 1368 34791 1424
rect 5529 1305 5615 1317
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 3444 1202 5236 1214
rect 12916 1214 12928 1354
rect 14696 1214 14708 1354
rect 15001 1305 15087 1317
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 12916 1202 14708 1214
rect 22388 1215 22400 1355
rect 24168 1215 24180 1355
rect 31860 1355 33652 1367
rect 34711 1356 34791 1368
rect 35529 1424 35609 1436
rect 35529 1368 35541 1424
rect 35597 1368 35609 1424
rect 35529 1356 35609 1368
rect 44183 1424 44263 1436
rect 44183 1368 44195 1424
rect 44251 1368 44263 1424
rect 24473 1306 24559 1318
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 22388 1203 24180 1215
rect 31860 1215 31872 1355
rect 33640 1215 33652 1355
rect 41332 1355 43124 1367
rect 44183 1356 44263 1368
rect 45001 1424 45081 1436
rect 45001 1368 45013 1424
rect 45069 1368 45081 1424
rect 45001 1356 45081 1368
rect 53655 1424 53735 1436
rect 53655 1368 53667 1424
rect 53723 1368 53735 1424
rect 33945 1306 34031 1318
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 31860 1203 33652 1215
rect 41332 1215 41344 1355
rect 43112 1215 43124 1355
rect 50804 1355 52596 1367
rect 53655 1356 53735 1368
rect 54473 1424 54553 1436
rect 54473 1368 54485 1424
rect 54541 1368 54553 1424
rect 54473 1356 54553 1368
rect 43417 1306 43503 1318
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 41332 1203 43124 1215
rect 50804 1215 50816 1355
rect 52584 1215 52596 1355
rect 52889 1306 52975 1318
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 50804 1203 52596 1215
rect 4814 1030 5134 1040
rect 1970 568 2458 578
rect 1970 512 1982 568
rect 2038 512 2390 568
rect 2446 512 2458 568
rect 1970 502 2458 512
rect 4814 230 4824 1030
rect 5124 230 5134 1030
rect 14286 1030 14606 1040
rect 11442 568 11930 578
rect 11442 512 11454 568
rect 11510 512 11862 568
rect 11918 512 11930 568
rect 11442 502 11930 512
rect 4814 220 5134 230
rect 14286 230 14296 1030
rect 14596 230 14606 1030
rect 23758 1031 24078 1041
rect 20914 569 21402 579
rect 20914 513 20926 569
rect 20982 513 21334 569
rect 21390 513 21402 569
rect 20914 503 21402 513
rect 14286 220 14606 230
rect 23758 231 23768 1031
rect 24068 231 24078 1031
rect 33230 1031 33550 1041
rect 30386 569 30874 579
rect 30386 513 30398 569
rect 30454 513 30806 569
rect 30862 513 30874 569
rect 30386 503 30874 513
rect 23758 221 24078 231
rect 33230 231 33240 1031
rect 33540 231 33550 1031
rect 42702 1031 43022 1041
rect 39858 569 40346 579
rect 39858 513 39870 569
rect 39926 513 40278 569
rect 40334 513 40346 569
rect 39858 503 40346 513
rect 33230 221 33550 231
rect 42702 231 42712 1031
rect 43012 231 43022 1031
rect 52174 1031 52494 1041
rect 49330 569 49818 579
rect 49330 513 49342 569
rect 49398 513 49750 569
rect 49806 513 49818 569
rect 49330 503 49818 513
rect 42702 221 43022 231
rect 52174 231 52184 1031
rect 52484 231 52494 1031
rect 52174 221 52494 231
rect 9077 -51 9087 -50
rect -689 -169 -441 -51
rect -451 -171 -441 -169
rect -385 -169 9087 -51
rect -385 -171 -375 -169
rect 9077 -170 9087 -169
rect 9143 -51 9153 -50
rect 18549 -51 18559 -50
rect 9143 -169 18559 -51
rect 9143 -170 9153 -169
rect 18549 -170 18559 -169
rect 18615 -51 18625 -50
rect 28021 -51 28031 -49
rect 18615 -169 28031 -51
rect 28087 -51 28097 -49
rect 37493 -51 37503 -49
rect 28087 -169 37503 -51
rect 37559 -51 37569 -49
rect 46965 -51 46975 -49
rect 37559 -169 46975 -51
rect 47031 -169 47041 -49
rect 18615 -170 18625 -169
<< via3 >>
rect 6808 9852 6864 9908
rect 16280 9852 16336 9908
rect 25752 9853 25808 9909
rect 35224 9853 35280 9909
rect 44696 9853 44752 9909
rect 54168 9853 54224 9909
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 24588 8884 24644 8940
rect 34060 8884 34116 8940
rect 43532 8884 43588 8940
rect 53004 8884 53060 8940
rect 6307 7982 6363 8038
rect 7125 7982 7181 8038
rect 15779 7982 15835 8038
rect 16597 7982 16653 8038
rect 25251 7983 25307 8039
rect 26069 7983 26125 8039
rect 34723 7983 34779 8039
rect 35541 7983 35597 8039
rect 44195 7983 44251 8039
rect 45013 7983 45069 8039
rect 53667 7983 53723 8039
rect 54485 7983 54541 8039
rect 6808 7647 6864 7703
rect 8294 7647 8350 7703
rect 16280 7647 16336 7703
rect 17766 7647 17822 7703
rect 25752 7648 25808 7704
rect 27238 7648 27294 7704
rect 35224 7648 35280 7704
rect 36710 7648 36766 7704
rect 44696 7648 44752 7704
rect 46182 7648 46238 7704
rect 54168 7648 54224 7704
rect 55654 7648 55710 7704
rect 6307 5777 6363 5833
rect 7125 5777 7181 5833
rect 7793 5777 7849 5833
rect 8611 5777 8667 5833
rect 15779 5777 15835 5833
rect 16597 5777 16653 5833
rect 17265 5777 17321 5833
rect 18083 5777 18139 5833
rect 25251 5778 25307 5834
rect 26069 5778 26125 5834
rect 26737 5778 26793 5834
rect 27555 5778 27611 5834
rect 34723 5778 34779 5834
rect 35541 5778 35597 5834
rect 36209 5778 36265 5834
rect 37027 5778 37083 5834
rect 44195 5778 44251 5834
rect 45013 5778 45069 5834
rect 45681 5778 45737 5834
rect 46499 5778 46555 5834
rect 53667 5778 53723 5834
rect 54485 5778 54541 5834
rect 55153 5778 55209 5834
rect 55971 5778 56027 5834
rect 6808 5442 6864 5498
rect 8294 5443 8350 5499
rect 16280 5442 16336 5498
rect 17766 5443 17822 5499
rect 25752 5443 25808 5499
rect 27238 5444 27294 5500
rect 35224 5443 35280 5499
rect 36710 5444 36766 5500
rect 44696 5443 44752 5499
rect 46182 5444 46238 5500
rect 54168 5443 54224 5499
rect 55654 5444 55710 5500
rect 4824 3510 5124 4310
rect 6307 3572 6363 3628
rect 7125 3572 7181 3628
rect 7793 3573 7849 3629
rect 8611 3573 8667 3629
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 15779 3572 15835 3628
rect 16597 3572 16653 3628
rect 17265 3573 17321 3629
rect 18083 3573 18139 3629
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 25251 3573 25307 3629
rect 26069 3573 26125 3629
rect 26737 3574 26793 3630
rect 27555 3574 27611 3630
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 34723 3573 34779 3629
rect 35541 3573 35597 3629
rect 36209 3574 36265 3630
rect 37027 3574 37083 3630
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 44195 3573 44251 3629
rect 45013 3573 45069 3629
rect 45681 3574 45737 3630
rect 46499 3574 46555 3630
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 53667 3573 53723 3629
rect 54485 3573 54541 3629
rect 55153 3574 55209 3630
rect 55971 3574 56027 3630
rect 6808 3237 6864 3293
rect 2396 2400 2996 2540
rect 16280 3237 16336 3293
rect 11868 2400 12468 2540
rect 25752 3238 25808 3294
rect 21340 2401 21940 2541
rect 35224 3238 35280 3294
rect 30812 2401 31412 2541
rect 44696 3238 44752 3294
rect 40284 2401 40884 2541
rect 54168 3238 54224 3294
rect 49756 2401 50356 2541
rect 6307 1367 6363 1423
rect 7125 1367 7181 1423
rect 15779 1367 15835 1423
rect 3456 1214 5224 1354
rect 16597 1367 16653 1423
rect 25251 1368 25307 1424
rect 26069 1368 26125 1424
rect 34723 1368 34779 1424
rect 5541 1249 5597 1305
rect 12928 1214 14696 1354
rect 15013 1249 15069 1305
rect 22400 1215 24168 1355
rect 35541 1368 35597 1424
rect 44195 1368 44251 1424
rect 24485 1250 24541 1306
rect 31872 1215 33640 1355
rect 45013 1368 45069 1424
rect 53667 1368 53723 1424
rect 33957 1250 34013 1306
rect 41344 1215 43112 1355
rect 54485 1368 54541 1424
rect 43429 1250 43485 1306
rect 50816 1215 52584 1355
rect 52901 1250 52957 1306
rect 4824 230 5124 1030
rect 14296 230 14596 1030
rect 23768 231 24068 1031
rect 33240 231 33540 1031
rect 42712 231 43012 1031
rect 52184 231 52484 1031
<< metal4 >>
rect 6796 9908 6882 9912
rect 6796 9852 6808 9908
rect 6864 9852 6882 9908
rect 6796 9840 6882 9852
rect 16268 9908 16354 9912
rect 16268 9852 16280 9908
rect 16336 9852 16354 9908
rect 16268 9840 16354 9852
rect 25740 9909 25826 9913
rect 25740 9853 25752 9909
rect 25808 9853 25826 9909
rect 25740 9841 25826 9853
rect 35212 9909 35298 9913
rect 35212 9853 35224 9909
rect 35280 9853 35298 9909
rect 35212 9841 35298 9853
rect 44684 9909 44770 9913
rect 44684 9853 44696 9909
rect 44752 9853 44770 9909
rect 44684 9841 44770 9853
rect 54156 9909 54242 9913
rect 54156 9853 54168 9909
rect 54224 9853 54242 9909
rect 54156 9841 54242 9853
rect 5630 8939 5718 8951
rect 5630 8883 5644 8939
rect 5700 8883 5718 8939
rect 5630 8871 5718 8883
rect 5782 8038 9082 9704
rect 15102 8939 15190 8951
rect 15102 8883 15116 8939
rect 15172 8883 15190 8939
rect 15102 8871 15190 8883
rect 5782 7982 6307 8038
rect 6363 7982 7125 8038
rect 7181 7982 9082 8038
rect 5782 7864 9082 7982
rect 5782 7499 6614 7864
rect 6796 7703 6882 7707
rect 6796 7647 6808 7703
rect 6864 7647 6882 7703
rect 6796 7635 6882 7647
rect 7064 7499 8100 7864
rect 8282 7703 8368 7707
rect 8282 7647 8294 7703
rect 8350 7647 8368 7703
rect 8282 7635 8368 7647
rect 8550 7499 9082 7864
rect 5782 5833 9082 7499
rect 5782 5777 6307 5833
rect 6363 5777 7125 5833
rect 7181 5777 7793 5833
rect 7849 5777 8611 5833
rect 8667 5777 9082 5833
rect 5782 5659 9082 5777
rect 5782 5294 6614 5659
rect 6796 5498 6882 5502
rect 6796 5442 6808 5498
rect 6864 5442 6882 5498
rect 6796 5430 6882 5442
rect 7064 5294 8100 5659
rect 8282 5499 8368 5503
rect 8282 5443 8294 5499
rect 8350 5443 8368 5499
rect 8282 5431 8368 5443
rect 8550 5294 9082 5659
rect 4814 4310 5134 4320
rect 4814 3510 4824 4310
rect 5124 3510 5134 4310
rect 4814 3500 5134 3510
rect 5782 3629 9082 5294
rect 15254 8038 18554 9704
rect 24574 8940 24662 8952
rect 24574 8884 24588 8940
rect 24644 8884 24662 8940
rect 24574 8872 24662 8884
rect 15254 7982 15779 8038
rect 15835 7982 16597 8038
rect 16653 7982 18554 8038
rect 15254 7864 18554 7982
rect 15254 7499 16086 7864
rect 16268 7703 16354 7707
rect 16268 7647 16280 7703
rect 16336 7647 16354 7703
rect 16268 7635 16354 7647
rect 16536 7499 17572 7864
rect 17754 7703 17840 7707
rect 17754 7647 17766 7703
rect 17822 7647 17840 7703
rect 17754 7635 17840 7647
rect 18022 7499 18554 7864
rect 15254 5833 18554 7499
rect 15254 5777 15779 5833
rect 15835 5777 16597 5833
rect 16653 5777 17265 5833
rect 17321 5777 18083 5833
rect 18139 5777 18554 5833
rect 15254 5659 18554 5777
rect 15254 5294 16086 5659
rect 16268 5498 16354 5502
rect 16268 5442 16280 5498
rect 16336 5442 16354 5498
rect 16268 5430 16354 5442
rect 16536 5294 17572 5659
rect 17754 5499 17840 5503
rect 17754 5443 17766 5499
rect 17822 5443 17840 5499
rect 17754 5431 17840 5443
rect 18022 5294 18554 5659
rect 5782 3628 7793 3629
rect 5782 3572 6307 3628
rect 6363 3572 7125 3628
rect 7181 3573 7793 3628
rect 7849 3573 8611 3629
rect 8667 3573 9082 3629
rect 7181 3572 9082 3573
rect 5782 3454 9082 3572
rect 9896 4310 10116 4320
rect 9896 3510 9906 4310
rect 10106 3510 10116 4310
rect 9896 3500 10116 3510
rect 14286 4310 14606 4320
rect 14286 3510 14296 4310
rect 14596 3510 14606 4310
rect 14286 3500 14606 3510
rect 15254 3629 18554 5294
rect 24726 8039 28026 9705
rect 34046 8940 34134 8952
rect 34046 8884 34060 8940
rect 34116 8884 34134 8940
rect 34046 8872 34134 8884
rect 24726 7983 25251 8039
rect 25307 7983 26069 8039
rect 26125 7983 28026 8039
rect 24726 7865 28026 7983
rect 24726 7500 25558 7865
rect 25740 7704 25826 7708
rect 25740 7648 25752 7704
rect 25808 7648 25826 7704
rect 25740 7636 25826 7648
rect 26008 7500 27044 7865
rect 27226 7704 27312 7708
rect 27226 7648 27238 7704
rect 27294 7648 27312 7704
rect 27226 7636 27312 7648
rect 27494 7500 28026 7865
rect 24726 5834 28026 7500
rect 24726 5778 25251 5834
rect 25307 5778 26069 5834
rect 26125 5778 26737 5834
rect 26793 5778 27555 5834
rect 27611 5778 28026 5834
rect 24726 5660 28026 5778
rect 24726 5295 25558 5660
rect 25740 5499 25826 5503
rect 25740 5443 25752 5499
rect 25808 5443 25826 5499
rect 25740 5431 25826 5443
rect 26008 5295 27044 5660
rect 27226 5500 27312 5504
rect 27226 5444 27238 5500
rect 27294 5444 27312 5500
rect 27226 5432 27312 5444
rect 27494 5295 28026 5660
rect 15254 3628 17265 3629
rect 15254 3572 15779 3628
rect 15835 3572 16597 3628
rect 16653 3573 17265 3628
rect 17321 3573 18083 3629
rect 18139 3573 18554 3629
rect 16653 3572 18554 3573
rect 5782 3089 6614 3454
rect 6796 3293 6882 3297
rect 6796 3237 6808 3293
rect 6864 3237 6882 3293
rect 6796 3225 6882 3237
rect 7064 3089 9082 3454
rect 2384 2540 5236 2552
rect 2384 2400 2396 2540
rect 2996 2400 5236 2540
rect 2384 2388 5236 2400
rect 3444 1354 5236 2388
rect 3444 1214 3456 1354
rect 5224 1214 5236 1354
rect 5782 1423 9082 3089
rect 15254 3454 18554 3572
rect 19368 4311 19588 4321
rect 19368 3511 19378 4311
rect 19578 3511 19588 4311
rect 19368 3501 19588 3511
rect 23758 4311 24078 4321
rect 23758 3511 23768 4311
rect 24068 3511 24078 4311
rect 23758 3501 24078 3511
rect 24726 3630 28026 5295
rect 34198 8039 37498 9705
rect 43518 8940 43606 8952
rect 43518 8884 43532 8940
rect 43588 8884 43606 8940
rect 43518 8872 43606 8884
rect 34198 7983 34723 8039
rect 34779 7983 35541 8039
rect 35597 7983 37498 8039
rect 34198 7865 37498 7983
rect 34198 7500 35030 7865
rect 35212 7704 35298 7708
rect 35212 7648 35224 7704
rect 35280 7648 35298 7704
rect 35212 7636 35298 7648
rect 35480 7500 36516 7865
rect 36698 7704 36784 7708
rect 36698 7648 36710 7704
rect 36766 7648 36784 7704
rect 36698 7636 36784 7648
rect 36966 7500 37498 7865
rect 34198 5834 37498 7500
rect 34198 5778 34723 5834
rect 34779 5778 35541 5834
rect 35597 5778 36209 5834
rect 36265 5778 37027 5834
rect 37083 5778 37498 5834
rect 34198 5660 37498 5778
rect 34198 5295 35030 5660
rect 35212 5499 35298 5503
rect 35212 5443 35224 5499
rect 35280 5443 35298 5499
rect 35212 5431 35298 5443
rect 35480 5295 36516 5660
rect 36698 5500 36784 5504
rect 36698 5444 36710 5500
rect 36766 5444 36784 5500
rect 36698 5432 36784 5444
rect 36966 5295 37498 5660
rect 24726 3629 26737 3630
rect 24726 3573 25251 3629
rect 25307 3573 26069 3629
rect 26125 3574 26737 3629
rect 26793 3574 27555 3630
rect 27611 3574 28026 3630
rect 26125 3573 28026 3574
rect 15254 3089 16086 3454
rect 16268 3293 16354 3297
rect 16268 3237 16280 3293
rect 16336 3237 16354 3293
rect 16268 3225 16354 3237
rect 16536 3089 18554 3454
rect 11856 2540 14708 2552
rect 11856 2400 11868 2540
rect 12468 2400 14708 2540
rect 11856 2388 14708 2400
rect 5782 1367 6307 1423
rect 6363 1367 7125 1423
rect 7181 1367 9082 1423
rect 5529 1305 5615 1317
rect 5529 1249 5541 1305
rect 5597 1249 5615 1305
rect 5529 1237 5615 1249
rect 5782 1237 9082 1367
rect 12916 1354 14708 2388
rect 3444 1202 5236 1214
rect 5782 1040 7078 1237
rect 12916 1214 12928 1354
rect 14696 1214 14708 1354
rect 15254 1423 18554 3089
rect 24726 3455 28026 3573
rect 28840 4311 29060 4321
rect 28840 3511 28850 4311
rect 29050 3511 29060 4311
rect 28840 3501 29060 3511
rect 33230 4311 33550 4321
rect 33230 3511 33240 4311
rect 33540 3511 33550 4311
rect 33230 3501 33550 3511
rect 34198 3630 37498 5295
rect 43670 8039 46970 9705
rect 52990 8940 53078 8952
rect 52990 8884 53004 8940
rect 53060 8884 53078 8940
rect 52990 8872 53078 8884
rect 43670 7983 44195 8039
rect 44251 7983 45013 8039
rect 45069 7983 46970 8039
rect 43670 7865 46970 7983
rect 43670 7500 44502 7865
rect 44684 7704 44770 7708
rect 44684 7648 44696 7704
rect 44752 7648 44770 7704
rect 44684 7636 44770 7648
rect 44952 7500 45988 7865
rect 46170 7704 46256 7708
rect 46170 7648 46182 7704
rect 46238 7648 46256 7704
rect 46170 7636 46256 7648
rect 46438 7500 46970 7865
rect 43670 5834 46970 7500
rect 43670 5778 44195 5834
rect 44251 5778 45013 5834
rect 45069 5778 45681 5834
rect 45737 5778 46499 5834
rect 46555 5778 46970 5834
rect 43670 5660 46970 5778
rect 43670 5295 44502 5660
rect 44684 5499 44770 5503
rect 44684 5443 44696 5499
rect 44752 5443 44770 5499
rect 44684 5431 44770 5443
rect 44952 5295 45988 5660
rect 46170 5500 46256 5504
rect 46170 5444 46182 5500
rect 46238 5444 46256 5500
rect 46170 5432 46256 5444
rect 46438 5295 46970 5660
rect 34198 3629 36209 3630
rect 34198 3573 34723 3629
rect 34779 3573 35541 3629
rect 35597 3574 36209 3629
rect 36265 3574 37027 3630
rect 37083 3574 37498 3630
rect 35597 3573 37498 3574
rect 24726 3090 25558 3455
rect 25740 3294 25826 3298
rect 25740 3238 25752 3294
rect 25808 3238 25826 3294
rect 25740 3226 25826 3238
rect 26008 3090 28026 3455
rect 21328 2541 24180 2553
rect 21328 2401 21340 2541
rect 21940 2401 24180 2541
rect 21328 2389 24180 2401
rect 15254 1367 15779 1423
rect 15835 1367 16597 1423
rect 16653 1367 18554 1423
rect 15001 1305 15087 1317
rect 15001 1249 15013 1305
rect 15069 1249 15087 1305
rect 15001 1237 15087 1249
rect 15254 1237 18554 1367
rect 22388 1355 24180 2389
rect 12916 1202 14708 1214
rect 15254 1040 16550 1237
rect 22388 1215 22400 1355
rect 24168 1215 24180 1355
rect 24726 1424 28026 3090
rect 34198 3455 37498 3573
rect 38312 4311 38532 4321
rect 38312 3511 38322 4311
rect 38522 3511 38532 4311
rect 38312 3501 38532 3511
rect 42702 4311 43022 4321
rect 42702 3511 42712 4311
rect 43012 3511 43022 4311
rect 42702 3501 43022 3511
rect 43670 3630 46970 5295
rect 53142 8039 56442 9705
rect 53142 7983 53667 8039
rect 53723 7983 54485 8039
rect 54541 7983 56442 8039
rect 53142 7865 56442 7983
rect 53142 7500 53974 7865
rect 54156 7704 54242 7708
rect 54156 7648 54168 7704
rect 54224 7648 54242 7704
rect 54156 7636 54242 7648
rect 54424 7500 55460 7865
rect 55642 7704 55728 7708
rect 55642 7648 55654 7704
rect 55710 7648 55728 7704
rect 55642 7636 55728 7648
rect 55910 7500 56442 7865
rect 53142 5834 56442 7500
rect 53142 5778 53667 5834
rect 53723 5778 54485 5834
rect 54541 5778 55153 5834
rect 55209 5778 55971 5834
rect 56027 5778 56442 5834
rect 53142 5660 56442 5778
rect 53142 5295 53974 5660
rect 54156 5499 54242 5503
rect 54156 5443 54168 5499
rect 54224 5443 54242 5499
rect 54156 5431 54242 5443
rect 54424 5295 55460 5660
rect 55642 5500 55728 5504
rect 55642 5444 55654 5500
rect 55710 5444 55728 5500
rect 55642 5432 55728 5444
rect 55910 5295 56442 5660
rect 43670 3629 45681 3630
rect 43670 3573 44195 3629
rect 44251 3573 45013 3629
rect 45069 3574 45681 3629
rect 45737 3574 46499 3630
rect 46555 3574 46970 3630
rect 45069 3573 46970 3574
rect 34198 3090 35030 3455
rect 35212 3294 35298 3298
rect 35212 3238 35224 3294
rect 35280 3238 35298 3294
rect 35212 3226 35298 3238
rect 35480 3090 37498 3455
rect 30800 2541 33652 2553
rect 30800 2401 30812 2541
rect 31412 2401 33652 2541
rect 30800 2389 33652 2401
rect 24726 1368 25251 1424
rect 25307 1368 26069 1424
rect 26125 1368 28026 1424
rect 24473 1306 24559 1318
rect 24473 1250 24485 1306
rect 24541 1250 24559 1306
rect 24473 1238 24559 1250
rect 24726 1238 28026 1368
rect 31860 1355 33652 2389
rect 22388 1203 24180 1215
rect 24726 1041 26022 1238
rect 31860 1215 31872 1355
rect 33640 1215 33652 1355
rect 34198 1424 37498 3090
rect 43670 3455 46970 3573
rect 47784 4311 48004 4321
rect 47784 3511 47794 4311
rect 47994 3511 48004 4311
rect 47784 3501 48004 3511
rect 52174 4311 52494 4321
rect 52174 3511 52184 4311
rect 52484 3511 52494 4311
rect 52174 3501 52494 3511
rect 53142 3630 56442 5295
rect 53142 3629 55153 3630
rect 53142 3573 53667 3629
rect 53723 3573 54485 3629
rect 54541 3574 55153 3629
rect 55209 3574 55971 3630
rect 56027 3574 56442 3630
rect 54541 3573 56442 3574
rect 43670 3090 44502 3455
rect 44684 3294 44770 3298
rect 44684 3238 44696 3294
rect 44752 3238 44770 3294
rect 44684 3226 44770 3238
rect 44952 3090 46970 3455
rect 40272 2541 43124 2553
rect 40272 2401 40284 2541
rect 40884 2401 43124 2541
rect 40272 2389 43124 2401
rect 34198 1368 34723 1424
rect 34779 1368 35541 1424
rect 35597 1368 37498 1424
rect 33945 1306 34031 1318
rect 33945 1250 33957 1306
rect 34013 1250 34031 1306
rect 33945 1238 34031 1250
rect 34198 1238 37498 1368
rect 41332 1355 43124 2389
rect 31860 1203 33652 1215
rect 34198 1041 35494 1238
rect 41332 1215 41344 1355
rect 43112 1215 43124 1355
rect 43670 1424 46970 3090
rect 53142 3455 56442 3573
rect 53142 3090 53974 3455
rect 54156 3294 54242 3298
rect 54156 3238 54168 3294
rect 54224 3238 54242 3294
rect 54156 3226 54242 3238
rect 54424 3090 56442 3455
rect 49744 2541 52596 2553
rect 49744 2401 49756 2541
rect 50356 2401 52596 2541
rect 49744 2389 52596 2401
rect 43670 1368 44195 1424
rect 44251 1368 45013 1424
rect 45069 1368 46970 1424
rect 43417 1306 43503 1318
rect 43417 1250 43429 1306
rect 43485 1250 43503 1306
rect 43417 1238 43503 1250
rect 43670 1238 46970 1368
rect 50804 1355 52596 2389
rect 41332 1203 43124 1215
rect 43670 1041 44966 1238
rect 50804 1215 50816 1355
rect 52584 1215 52596 1355
rect 53142 1424 56442 3090
rect 53142 1368 53667 1424
rect 53723 1368 54485 1424
rect 54541 1368 56442 1424
rect 52889 1306 52975 1318
rect 52889 1250 52901 1306
rect 52957 1250 52975 1306
rect 52889 1238 52975 1250
rect 53142 1238 56442 1368
rect 50804 1203 52596 1215
rect 53142 1041 54438 1238
rect 4814 1030 7078 1040
rect 4814 230 4824 1030
rect 5124 230 7078 1030
rect 4814 220 7078 230
rect 14286 1030 16550 1040
rect 14286 230 14296 1030
rect 14596 230 16550 1030
rect 14286 220 16550 230
rect 23758 1031 26022 1041
rect 23758 231 23768 1031
rect 24068 231 26022 1031
rect 23758 221 26022 231
rect 33230 1031 35494 1041
rect 33230 231 33240 1031
rect 33540 231 35494 1031
rect 33230 221 35494 231
rect 42702 1031 44966 1041
rect 42702 231 42712 1031
rect 43012 231 44966 1031
rect 42702 221 44966 231
rect 52174 1031 54438 1041
rect 52174 231 52184 1031
rect 52484 231 54438 1031
rect 52174 221 54438 231
<< via4 >>
rect 6808 9852 6864 9908
rect 16280 9852 16336 9908
rect 25752 9853 25808 9909
rect 35224 9853 35280 9909
rect 44696 9853 44752 9909
rect 54168 9853 54224 9909
rect 5644 8883 5700 8939
rect 15116 8883 15172 8939
rect 6808 7647 6864 7703
rect 8294 7647 8350 7703
rect 6808 5442 6864 5498
rect 8294 5443 8350 5499
rect 4824 3510 5124 4310
rect 24588 8884 24644 8940
rect 16280 7647 16336 7703
rect 17766 7647 17822 7703
rect 16280 5442 16336 5498
rect 17766 5443 17822 5499
rect 9906 3510 10106 4310
rect 14296 3510 14596 4310
rect 34060 8884 34116 8940
rect 25752 7648 25808 7704
rect 27238 7648 27294 7704
rect 25752 5443 25808 5499
rect 27238 5444 27294 5500
rect 6808 3237 6864 3293
rect 19378 3511 19578 4311
rect 23768 3511 24068 4311
rect 43532 8884 43588 8940
rect 35224 7648 35280 7704
rect 36710 7648 36766 7704
rect 35224 5443 35280 5499
rect 36710 5444 36766 5500
rect 16280 3237 16336 3293
rect 5541 1249 5597 1305
rect 28850 3511 29050 4311
rect 33240 3511 33540 4311
rect 53004 8884 53060 8940
rect 44696 7648 44752 7704
rect 46182 7648 46238 7704
rect 44696 5443 44752 5499
rect 46182 5444 46238 5500
rect 25752 3238 25808 3294
rect 15013 1249 15069 1305
rect 38322 3511 38522 4311
rect 42712 3511 43012 4311
rect 54168 7648 54224 7704
rect 55654 7648 55710 7704
rect 54168 5443 54224 5499
rect 55654 5444 55710 5500
rect 35224 3238 35280 3294
rect 24485 1250 24541 1306
rect 47794 3511 47994 4311
rect 52184 3511 52484 4311
rect 44696 3238 44752 3294
rect 33957 1250 34013 1306
rect 54168 3238 54224 3294
rect 43429 1250 43485 1306
rect 52901 1250 52957 1306
<< metal5 >>
rect 5782 9908 9082 10016
rect 5782 9852 6808 9908
rect 6864 9852 9082 9908
rect 5782 9031 9082 9852
rect 15254 9908 18554 10016
rect 15254 9852 16280 9908
rect 16336 9852 18554 9908
rect 15254 9031 18554 9852
rect 24726 9909 28026 10017
rect 24726 9853 25752 9909
rect 25808 9853 28026 9909
rect 24726 9032 28026 9853
rect 34198 9909 37498 10017
rect 34198 9853 35224 9909
rect 35280 9853 37498 9909
rect 34198 9032 37498 9853
rect 43670 9909 46970 10017
rect 43670 9853 44696 9909
rect 44752 9853 46970 9909
rect 43670 9032 46970 9853
rect 53142 9909 56442 10017
rect 53142 9853 54168 9909
rect 54224 9853 56442 9909
rect 53142 9032 56442 9853
rect 5630 8939 9082 9031
rect 5630 8883 5644 8939
rect 5700 8883 9082 8939
rect 5630 8871 9082 8883
rect 15102 8939 18554 9031
rect 15102 8883 15116 8939
rect 15172 8883 18554 8939
rect 15102 8871 18554 8883
rect 24574 8940 28026 9032
rect 24574 8884 24588 8940
rect 24644 8884 28026 8940
rect 24574 8872 28026 8884
rect 34046 8940 37498 9032
rect 34046 8884 34060 8940
rect 34116 8884 37498 8940
rect 34046 8872 37498 8884
rect 43518 8940 46970 9032
rect 43518 8884 43532 8940
rect 43588 8884 46970 8940
rect 43518 8872 46970 8884
rect 52990 8940 56442 9032
rect 52990 8884 53004 8940
rect 53060 8884 56442 8940
rect 52990 8872 56442 8884
rect 5782 7703 9082 8871
rect 5782 7647 6808 7703
rect 6864 7647 8294 7703
rect 8350 7647 9082 7703
rect 5782 5499 9082 7647
rect 5782 5498 8294 5499
rect 5782 5442 6808 5498
rect 6864 5443 8294 5498
rect 8350 5443 9082 5499
rect 6864 5442 9082 5443
rect 5782 4320 9082 5442
rect 15254 7703 18554 8871
rect 15254 7647 16280 7703
rect 16336 7647 17766 7703
rect 17822 7647 18554 7703
rect 15254 5499 18554 7647
rect 15254 5498 17766 5499
rect 15254 5442 16280 5498
rect 16336 5443 17766 5498
rect 17822 5443 18554 5499
rect 16336 5442 18554 5443
rect 15254 4321 18554 5442
rect 24726 7704 28026 8872
rect 24726 7648 25752 7704
rect 25808 7648 27238 7704
rect 27294 7648 28026 7704
rect 24726 5500 28026 7648
rect 24726 5499 27238 5500
rect 24726 5443 25752 5499
rect 25808 5444 27238 5499
rect 27294 5444 28026 5500
rect 25808 5443 28026 5444
rect 24726 4321 28026 5443
rect 34198 7704 37498 8872
rect 34198 7648 35224 7704
rect 35280 7648 36710 7704
rect 36766 7648 37498 7704
rect 34198 5500 37498 7648
rect 34198 5499 36710 5500
rect 34198 5443 35224 5499
rect 35280 5444 36710 5499
rect 36766 5444 37498 5500
rect 35280 5443 37498 5444
rect 34198 4321 37498 5443
rect 43670 7704 46970 8872
rect 43670 7648 44696 7704
rect 44752 7648 46182 7704
rect 46238 7648 46970 7704
rect 43670 5500 46970 7648
rect 43670 5499 46182 5500
rect 43670 5443 44696 5499
rect 44752 5444 46182 5499
rect 46238 5444 46970 5500
rect 44752 5443 46970 5444
rect 43670 4321 46970 5443
rect 53142 7704 56442 8872
rect 53142 7648 54168 7704
rect 54224 7648 55654 7704
rect 55710 7648 56442 7704
rect 53142 5500 56442 7648
rect 53142 5499 55654 5500
rect 53142 5443 54168 5499
rect 54224 5444 55654 5499
rect 55710 5444 56442 5500
rect 54224 5443 56442 5444
rect 53142 4321 56442 5443
rect 15254 4320 19588 4321
rect 4814 4310 10116 4320
rect 4814 3510 4824 4310
rect 5124 3510 9906 4310
rect 10106 3510 10116 4310
rect 4814 3500 10116 3510
rect 14286 4311 19588 4320
rect 14286 4310 19378 4311
rect 14286 3510 14296 4310
rect 14596 3511 19378 4310
rect 19578 3511 19588 4311
rect 14596 3510 19588 3511
rect 14286 3501 19588 3510
rect 23758 4311 29060 4321
rect 23758 3511 23768 4311
rect 24068 3511 28850 4311
rect 29050 3511 29060 4311
rect 23758 3501 29060 3511
rect 33230 4311 38532 4321
rect 33230 3511 33240 4311
rect 33540 3511 38322 4311
rect 38522 3511 38532 4311
rect 33230 3501 38532 3511
rect 42702 4311 48004 4321
rect 42702 3511 42712 4311
rect 43012 3511 47794 4311
rect 47994 3511 48004 4311
rect 42702 3501 48004 3511
rect 52174 4311 56442 4321
rect 52174 3511 52184 4311
rect 52484 3511 56442 4311
rect 52174 3501 56442 3511
rect 14286 3500 18554 3501
rect 5782 3293 9082 3500
rect 5782 3237 6808 3293
rect 6864 3237 9082 3293
rect 5782 1397 9082 3237
rect 15254 3293 18554 3500
rect 15254 3237 16280 3293
rect 16336 3237 18554 3293
rect 15254 1397 18554 3237
rect 24726 3294 28026 3501
rect 24726 3238 25752 3294
rect 25808 3238 28026 3294
rect 24726 1398 28026 3238
rect 34198 3294 37498 3501
rect 34198 3238 35224 3294
rect 35280 3238 37498 3294
rect 34198 1398 37498 3238
rect 43670 3294 46970 3501
rect 43670 3238 44696 3294
rect 44752 3238 46970 3294
rect 43670 1398 46970 3238
rect 53142 3294 56442 3501
rect 53142 3238 54168 3294
rect 54224 3238 56442 3294
rect 53142 1398 56442 3238
rect 5529 1305 9082 1397
rect 5529 1249 5541 1305
rect 5597 1249 9082 1305
rect 5529 1237 9082 1249
rect 15001 1305 18554 1397
rect 15001 1249 15013 1305
rect 15069 1249 18554 1305
rect 15001 1237 18554 1249
rect 24473 1306 28026 1398
rect 24473 1250 24485 1306
rect 24541 1250 28026 1306
rect 24473 1238 28026 1250
rect 33945 1306 37498 1398
rect 33945 1250 33957 1306
rect 34013 1250 37498 1306
rect 33945 1238 37498 1250
rect 43417 1306 46970 1398
rect 43417 1250 43429 1306
rect 43485 1250 46970 1306
rect 43417 1238 46970 1250
rect 52889 1306 56442 1398
rect 52889 1250 52901 1306
rect 52957 1250 56442 1306
rect 52889 1238 56442 1250
<< labels >>
rlabel metal3 -689 -113 -689 -113 7 load
port 0 w
rlabel metal2 39 -370 39 -370 5 B6
port 1 s
rlabel metal2 9511 -370 9511 -370 5 B5
port 2 s
rlabel metal2 18983 -370 18983 -370 5 B4
port 3 s
rlabel metal2 56875 9891 56875 9891 1 serial_out
port 4 n
rlabel metal1 230 4493 230 4493 7 avdd
port 5 w
rlabel metal2 28455 -369 28455 -369 5 B3
port 6 s
rlabel metal1 230 54 230 54 7 avss
port 7 w
rlabel metal2 37927 -369 37927 -369 5 B2
port 8 s
rlabel metal2 47398 -369 47398 -369 5 B1
port 9 s
rlabel metal3 3058 5685 3058 5685 7 clk
port 10 w
rlabel metal2 10 3317 10 3317 7 2inmux_0.Bit
rlabel metal2 10 3161 10 3161 7 2inmux_0.Load
rlabel metal1 565 4510 565 4510 1 2inmux_0.VDD
rlabel metal2 5384 2064 5384 2064 3 2inmux_0.OUT
rlabel metal1 534 30 534 30 5 2inmux_0.VSS
rlabel metal2 10 821 10 821 7 2inmux_0.In
rlabel metal2 9482 3317 9482 3317 7 2inmux_2.Bit
rlabel metal2 9482 3161 9482 3161 7 2inmux_2.Load
rlabel metal1 10037 4510 10037 4510 1 2inmux_2.VDD
rlabel metal2 14856 2064 14856 2064 3 2inmux_2.OUT
rlabel metal1 10006 30 10006 30 5 2inmux_2.VSS
rlabel metal2 9482 821 9482 821 7 2inmux_2.In
rlabel metal1 5644 8911 5644 8911 7 dffrs_0.setb
rlabel metal1 5644 5688 5644 5688 7 dffrs_0.clk
rlabel metal1 5644 2063 5644 2063 7 dffrs_0.d
rlabel metal1 5661 1276 5661 1276 7 dffrs_0.resetb
rlabel metal2 9112 6590 9112 6590 3 dffrs_0.Q
rlabel metal2 9112 4385 9112 4385 3 dffrs_0.Qb
rlabel metal5 7752 10016 7752 10016 1 dffrs_0.vdd
rlabel metal4 7711 1237 7711 1237 5 dffrs_0.vss
rlabel metal1 15116 8911 15116 8911 7 dffrs_1.setb
rlabel metal1 15116 5688 15116 5688 7 dffrs_1.clk
rlabel metal1 15116 2063 15116 2063 7 dffrs_1.d
rlabel metal1 15133 1276 15133 1276 7 dffrs_1.resetb
rlabel metal2 18584 6590 18584 6590 3 dffrs_1.Q
rlabel metal2 18584 4385 18584 4385 3 dffrs_1.Qb
rlabel metal5 17224 10016 17224 10016 1 dffrs_1.vdd
rlabel metal4 17183 1237 17183 1237 5 dffrs_1.vss
rlabel metal2 18954 3318 18954 3318 7 2inmux_3.Bit
rlabel metal2 18954 3162 18954 3162 7 2inmux_3.Load
rlabel metal1 19509 4511 19509 4511 1 2inmux_3.VDD
rlabel metal2 24328 2065 24328 2065 3 2inmux_3.OUT
rlabel metal1 19478 31 19478 31 5 2inmux_3.VSS
rlabel metal2 18954 822 18954 822 7 2inmux_3.In
rlabel metal1 24588 8912 24588 8912 7 dffrs_2.setb
rlabel metal1 24588 5689 24588 5689 7 dffrs_2.clk
rlabel metal1 24588 2064 24588 2064 7 dffrs_2.d
rlabel metal1 24605 1277 24605 1277 7 dffrs_2.resetb
rlabel metal2 28056 6591 28056 6591 3 dffrs_2.Q
rlabel metal2 28056 4386 28056 4386 3 dffrs_2.Qb
rlabel metal5 26696 10017 26696 10017 1 dffrs_2.vdd
rlabel metal4 26655 1238 26655 1238 5 dffrs_2.vss
rlabel metal2 28426 3318 28426 3318 7 2inmux_4.Bit
rlabel metal2 28426 3162 28426 3162 7 2inmux_4.Load
rlabel metal1 28981 4511 28981 4511 1 2inmux_4.VDD
rlabel metal2 33800 2065 33800 2065 3 2inmux_4.OUT
rlabel metal1 28950 31 28950 31 5 2inmux_4.VSS
rlabel metal2 28426 822 28426 822 7 2inmux_4.In
rlabel metal1 34060 8912 34060 8912 7 dffrs_3.setb
rlabel metal1 34060 5689 34060 5689 7 dffrs_3.clk
rlabel metal1 34060 2064 34060 2064 7 dffrs_3.d
rlabel metal1 34077 1277 34077 1277 7 dffrs_3.resetb
rlabel metal2 37528 6591 37528 6591 3 dffrs_3.Q
rlabel metal2 37528 4386 37528 4386 3 dffrs_3.Qb
rlabel metal5 36168 10017 36168 10017 1 dffrs_3.vdd
rlabel metal4 36127 1238 36127 1238 5 dffrs_3.vss
rlabel metal2 37898 3318 37898 3318 7 2inmux_5.Bit
rlabel metal2 37898 3162 37898 3162 7 2inmux_5.Load
rlabel metal1 38453 4511 38453 4511 1 2inmux_5.VDD
rlabel metal2 43272 2065 43272 2065 3 2inmux_5.OUT
rlabel metal1 38422 31 38422 31 5 2inmux_5.VSS
rlabel metal2 37898 822 37898 822 7 2inmux_5.In
rlabel metal2 47370 3318 47370 3318 7 2inmux_1.Bit
rlabel metal2 47370 3162 47370 3162 7 2inmux_1.Load
rlabel metal1 47925 4511 47925 4511 1 2inmux_1.VDD
rlabel metal2 52744 2065 52744 2065 3 2inmux_1.OUT
rlabel metal1 47894 31 47894 31 5 2inmux_1.VSS
rlabel metal2 47370 822 47370 822 7 2inmux_1.In
rlabel metal1 43532 8912 43532 8912 7 dffrs_4.setb
rlabel metal1 43532 5689 43532 5689 7 dffrs_4.clk
rlabel metal1 43532 2064 43532 2064 7 dffrs_4.d
rlabel metal1 43549 1277 43549 1277 7 dffrs_4.resetb
rlabel metal2 47000 6591 47000 6591 3 dffrs_4.Q
rlabel metal2 47000 4386 47000 4386 3 dffrs_4.Qb
rlabel metal5 45640 10017 45640 10017 1 dffrs_4.vdd
rlabel metal4 45599 1238 45599 1238 5 dffrs_4.vss
rlabel metal1 53004 8912 53004 8912 7 dffrs_5.setb
rlabel metal1 53004 5689 53004 5689 7 dffrs_5.clk
rlabel metal1 53004 2064 53004 2064 7 dffrs_5.d
rlabel metal1 53021 1277 53021 1277 7 dffrs_5.resetb
rlabel metal2 56472 6591 56472 6591 3 dffrs_5.Q
rlabel metal2 56472 4386 56472 4386 3 dffrs_5.Qb
rlabel metal5 55112 10017 55112 10017 1 dffrs_5.vdd
rlabel metal4 55071 1238 55071 1238 5 dffrs_5.vss
<< end >>
