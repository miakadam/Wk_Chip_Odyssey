magic
tech gf180mcuD
magscale 1 10
timestamp 1757859367
<< metal1 >>
rect 200 1346 640 1396
rect 80 1120 160 1130
rect 80 1030 100 1120
rect 80 1020 160 1030
rect 270 1020 350 1130
rect 450 1120 530 1130
rect 450 1030 469 1120
rect 529 1030 530 1120
rect 450 1020 530 1030
rect 640 430 730 440
rect 277 410 347 423
rect 277 320 290 410
rect 343 320 347 410
rect 640 340 660 430
rect 714 340 730 430
rect 640 320 730 340
rect 277 303 347 320
<< via1 >>
rect 100 1030 160 1120
rect 469 1030 529 1120
rect 290 320 343 410
rect 660 340 714 430
<< metal2 >>
rect -120 1120 980 1150
rect -120 1030 100 1120
rect 160 1030 469 1120
rect 529 1030 980 1120
rect -120 1000 980 1030
rect -60 430 1040 440
rect -60 410 660 430
rect -60 320 290 410
rect 343 340 660 410
rect 714 340 1040 430
rect 343 320 1040 340
rect -60 290 1040 320
use nfet_03v3_QDTW5R  XM1
timestamp 1757859367
transform 1 0 414 0 1 726
box -474 -786 474 786
<< end >>
