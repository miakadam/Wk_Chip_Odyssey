* NGSPICE file created from osu_sc_and2_1.ext - technology: gf180mcuD

.subckt osu_sc_and2_1 A B Y VDD VSS
X0 VSS B a_280_210# VSS nfet_03v3 ad=0.3825p pd=1.75u as=0.10625p ps=1.1u w=0.85u l=0.3u
X1 a_120_210# A VDD VDD pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 Y a_120_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.3825p ps=1.75u w=0.85u l=0.3u
X3 VDD B a_120_210# VDD pfet_03v3 ad=0.6375p pd=2.45u as=0.4675p ps=2.25u w=1.7u l=0.3u
X4 Y a_120_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.6375p ps=2.45u w=1.7u l=0.3u
X5 a_280_210# A a_120_210# VSS nfet_03v3 ad=0.10625p pd=1.1u as=0.425p ps=2.7u w=0.85u l=0.3u
.ends

