* NGSPICE file created from osu_sc_buf_4.ext - technology: gf180mcuD

.subckt osu_sc_buf_4 A Y VDD VSS
X0 Y.t5 a_100_200 VDD.t7 VDD.t6 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 Y.t1 a_100_200 VSS.t7 VSS.t6 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X2 VSS.t9 A.t0 a_100_200 VSS.t8 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X3 VSS.t5 a_100_200 Y.t0 VSS.t4 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 Y.t4 a_100_200 VDD.t5 VDD.t4 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 VDD.t9 A.t1 a_100_200 VDD.t8 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X6 VSS.t3 a_100_200 Y.t7 VSS.t2 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X7 VDD.t3 a_100_200 Y.t3 VDD.t2 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X8 Y.t6 a_100_200 VSS.t1 VSS.t0 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X9 VDD.t1 a_100_200 Y.t2 VDD.t0 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
R0 VDD.t2 VDD.t4 265.625
R1 VDD.t8 VDD.n9 242.189
R2 VDD.t6 VDD.n5 195.312
R3 VDD.n6 VDD.t6 179.689
R4 VDD.n10 VDD.t8 145.413
R5 VDD.n6 VDD.t2 85.938
R6 VDD.n5 VDD.t0 70.313
R7 VDD.n9 VDD.t4 23.438
R8 VDD.n5 VDD.n4 12.6005
R9 VDD.n7 VDD.n6 12.6005
R10 VDD.n9 VDD.n8 12.6005
R11 VDD.n4 VDD.t1 3.38176
R12 VDD.n1 VDD.n0 2.16583
R13 VDD.n3 VDD.n2 2.16583
R14 VDD.n0 VDD.t5 1.13285
R15 VDD.n0 VDD.t9 1.13285
R16 VDD.n2 VDD.t7 1.13285
R17 VDD.n2 VDD.t3 1.13285
R18 VDD.n8 VDD.n7 0.154786
R19 VDD.n4 VDD.n3 0.1355
R20 VDD.n10 VDD.n1 0.109786
R21 VDD.n8 VDD.n1 0.0455
R22 VDD.n7 VDD.n3 0.0197857
R23 VDD VDD.n10 0.00371429
R24 Y.n5 Y.n4 6.5435
R25 Y.n2 Y.n1 6.5435
R26 Y Y.n8 4.5005
R27 Y.n6 Y.n3 2.17483
R28 Y.n4 Y.t0 2.03874
R29 Y.n4 Y.t1 2.03874
R30 Y.n1 Y.t7 2.03874
R31 Y.n1 Y.t6 2.03874
R32 Y.n8 Y.n0 2.00383
R33 Y.n0 Y.t2 1.13285
R34 Y.n0 Y.t5 1.13285
R35 Y.n3 Y.t3 1.13285
R36 Y.n3 Y.t4 1.13285
R37 Y.n5 Y.n2 0.5105
R38 Y.n7 Y.n6 0.5105
R39 Y.n7 Y.n2 0.2165
R40 Y.n6 Y.n5 0.2165
R41 Y.n8 Y.n7 0.1175
R42 VSS.t4 VSS.t6 876.985
R43 VSS.t8 VSS.n9 799.604
R44 VSS.t0 VSS.n5 644.841
R45 VSS.n6 VSS.t0 593.255
R46 VSS.n10 VSS.t8 448.892
R47 VSS.n6 VSS.t4 283.731
R48 VSS.n5 VSS.t2 232.143
R49 VSS.n9 VSS.t6 77.3815
R50 VSS.n5 VSS.n4 10.4005
R51 VSS.n7 VSS.n6 10.4005
R52 VSS.n9 VSS.n8 10.4005
R53 VSS.n4 VSS.t3 8.70131
R54 VSS.n3 VSS.n2 6.5795
R55 VSS.n1 VSS.n0 6.5795
R56 VSS.n2 VSS.t1 2.03874
R57 VSS.n2 VSS.t5 2.03874
R58 VSS.n0 VSS.t7 2.03874
R59 VSS.n0 VSS.t9 2.03874
R60 VSS.n8 VSS.n7 0.154786
R61 VSS.n4 VSS.n3 0.1355
R62 VSS.n10 VSS.n1 0.109786
R63 VSS.n8 VSS.n1 0.0455
R64 VSS.n7 VSS.n3 0.0197857
R65 VSS VSS.n10 0.00371429
R66 A.n0 A.t1 45.6255
R67 A.n0 A.t0 20.6838
R68 A A.n0 12.5005
.ends

