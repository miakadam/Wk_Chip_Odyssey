* NGSPICE file created from osu_sc_inv_1.ext - technology: gf180mcuD

.subckt osu_sc_inv_1 A Y VDD VSS
X0 Y A VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 Y A VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
.ends

