magic
tech gf180mcuD
magscale 1 10
timestamp 1757578771
<< metal1 >>
rect 2097 -500 3063 -420
rect 2097 -629 2143 -500
rect 2312 -631 2388 -598
rect 2772 -631 2848 -598
rect 3017 -629 3063 -500
rect 2130 -897 2236 -723
rect 2402 -782 2482 -772
rect 2402 -838 2414 -782
rect 2470 -838 2482 -782
rect 2402 -848 2482 -838
rect 2678 -782 2758 -772
rect 2678 -838 2690 -782
rect 2746 -838 2758 -782
rect 2678 -848 2758 -838
rect 2924 -897 3030 -723
rect 2322 -1176 2378 -989
rect 2540 -1040 2610 -1038
rect 2782 -1040 2838 -989
rect 2540 -1096 2552 -1040
rect 2608 -1096 2838 -1040
rect 2540 -1098 2610 -1096
rect 2322 -1178 2620 -1176
rect 2322 -1234 2552 -1178
rect 2608 -1234 2620 -1178
rect 2322 -1236 2620 -1234
rect 2312 -1451 2388 -1418
rect 2772 -1451 2848 -1418
rect 2136 -1717 2242 -1543
rect 2402 -1602 2482 -1592
rect 2402 -1658 2414 -1602
rect 2470 -1658 2482 -1602
rect 2402 -1668 2482 -1658
rect 2678 -1602 2758 -1592
rect 2678 -1658 2690 -1602
rect 2746 -1658 2758 -1602
rect 2678 -1668 2758 -1658
rect 2915 -1717 3021 -1543
rect 2310 -1778 2390 -1768
rect 2097 -1940 2143 -1800
rect 2310 -1834 2322 -1778
rect 2378 -1834 2390 -1778
rect 2310 -1844 2390 -1834
rect 2770 -1778 2850 -1768
rect 2770 -1834 2782 -1778
rect 2838 -1834 2850 -1778
rect 2770 -1844 2850 -1834
rect 3017 -1940 3063 -1800
rect 2097 -2020 3063 -1940
<< via1 >>
rect 2414 -838 2470 -782
rect 2690 -838 2746 -782
rect 2552 -1096 2608 -1040
rect 2552 -1234 2608 -1178
rect 2414 -1658 2470 -1602
rect 2690 -1658 2746 -1602
rect 2322 -1834 2378 -1778
rect 2782 -1834 2838 -1778
<< metal2 >>
rect 2402 -782 2482 -772
rect 2402 -838 2414 -782
rect 2470 -838 2482 -782
rect 2402 -848 2482 -838
rect 2678 -782 2758 -772
rect 2678 -838 2690 -782
rect 2746 -838 2758 -782
rect 2678 -848 2758 -838
rect 2414 -1040 2470 -848
rect 2539 -1040 2619 -1028
rect 2414 -1096 2552 -1040
rect 2608 -1096 2619 -1040
rect 2414 -1288 2470 -1096
rect 2539 -1108 2619 -1096
rect 2540 -1178 2620 -1168
rect 2690 -1178 2746 -848
rect 2540 -1234 2552 -1178
rect 2608 -1234 2746 -1178
rect 2540 -1244 2620 -1234
rect 1870 -1344 2470 -1288
rect 2414 -1592 2470 -1344
rect 2690 -1288 2746 -1234
rect 2690 -1344 3290 -1288
rect 2690 -1592 2746 -1344
rect 2402 -1602 2482 -1592
rect 2402 -1658 2414 -1602
rect 2470 -1658 2482 -1602
rect 2402 -1668 2482 -1658
rect 2678 -1602 2758 -1592
rect 2678 -1658 2690 -1602
rect 2746 -1658 2758 -1602
rect 2678 -1668 2758 -1658
rect 2310 -1778 2390 -1768
rect 2310 -1834 2322 -1778
rect 2378 -1834 2390 -1778
rect 2310 -1844 2390 -1834
rect 2770 -1778 2850 -1768
rect 2770 -1834 2782 -1778
rect 2838 -1834 2850 -1778
rect 2770 -1844 2850 -1834
rect 2322 -2178 2378 -1844
rect 2782 -2178 2838 -1844
use nfet_03v3_EKTWUP  M2
timestamp 1757566850
transform 1 0 2810 0 1 -1630
box -290 -310 290 310
use pfet_03v3_L25D84  M3
timestamp 1757566850
transform 1 0 2350 0 1 -810
box -290 -310 290 310
use nfet_03v3_EKTWUP  nfet_03v3_EKTWUP_0
timestamp 1757566850
transform 1 0 2350 0 1 -1630
box -290 -310 290 310
use pfet_03v3_L25D84  pfet_03v3_L25D84_0
timestamp 1757566850
transform 1 0 2810 0 1 -810
box -290 -310 290 310
<< labels >>
rlabel metal1 2578 -420 2578 -420 1 VDD
port 0 n
rlabel metal2 1870 -1318 1870 -1318 7 Vout1
port 1 w
rlabel metal2 3290 -1318 3290 -1318 3 Vout2
port 2 e
rlabel metal2 2350 -2178 2350 -2178 5 Vin1
port 3 s
rlabel metal2 2811 -2178 2811 -2178 5 Vin2
port 4 s
rlabel metal1 2583 -2020 2583 -2020 5 VSS
port 5 s
<< end >>
