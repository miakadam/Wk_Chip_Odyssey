magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< nwell >>
rect -954 -13022 954 13022
<< pmos >>
rect -704 9812 -304 12812
rect -200 9812 200 12812
rect 304 9812 704 12812
rect -704 6580 -304 9580
rect -200 6580 200 9580
rect 304 6580 704 9580
rect -704 3348 -304 6348
rect -200 3348 200 6348
rect 304 3348 704 6348
rect -704 116 -304 3116
rect -200 116 200 3116
rect 304 116 704 3116
rect -704 -3116 -304 -116
rect -200 -3116 200 -116
rect 304 -3116 704 -116
rect -704 -6348 -304 -3348
rect -200 -6348 200 -3348
rect 304 -6348 704 -3348
rect -704 -9580 -304 -6580
rect -200 -9580 200 -6580
rect 304 -9580 704 -6580
rect -704 -12812 -304 -9812
rect -200 -12812 200 -9812
rect 304 -12812 704 -9812
<< pdiff >>
rect -792 12799 -704 12812
rect -792 9825 -779 12799
rect -733 9825 -704 12799
rect -792 9812 -704 9825
rect -304 12799 -200 12812
rect -304 9825 -275 12799
rect -229 9825 -200 12799
rect -304 9812 -200 9825
rect 200 12799 304 12812
rect 200 9825 229 12799
rect 275 9825 304 12799
rect 200 9812 304 9825
rect 704 12799 792 12812
rect 704 9825 733 12799
rect 779 9825 792 12799
rect 704 9812 792 9825
rect -792 9567 -704 9580
rect -792 6593 -779 9567
rect -733 6593 -704 9567
rect -792 6580 -704 6593
rect -304 9567 -200 9580
rect -304 6593 -275 9567
rect -229 6593 -200 9567
rect -304 6580 -200 6593
rect 200 9567 304 9580
rect 200 6593 229 9567
rect 275 6593 304 9567
rect 200 6580 304 6593
rect 704 9567 792 9580
rect 704 6593 733 9567
rect 779 6593 792 9567
rect 704 6580 792 6593
rect -792 6335 -704 6348
rect -792 3361 -779 6335
rect -733 3361 -704 6335
rect -792 3348 -704 3361
rect -304 6335 -200 6348
rect -304 3361 -275 6335
rect -229 3361 -200 6335
rect -304 3348 -200 3361
rect 200 6335 304 6348
rect 200 3361 229 6335
rect 275 3361 304 6335
rect 200 3348 304 3361
rect 704 6335 792 6348
rect 704 3361 733 6335
rect 779 3361 792 6335
rect 704 3348 792 3361
rect -792 3103 -704 3116
rect -792 129 -779 3103
rect -733 129 -704 3103
rect -792 116 -704 129
rect -304 3103 -200 3116
rect -304 129 -275 3103
rect -229 129 -200 3103
rect -304 116 -200 129
rect 200 3103 304 3116
rect 200 129 229 3103
rect 275 129 304 3103
rect 200 116 304 129
rect 704 3103 792 3116
rect 704 129 733 3103
rect 779 129 792 3103
rect 704 116 792 129
rect -792 -129 -704 -116
rect -792 -3103 -779 -129
rect -733 -3103 -704 -129
rect -792 -3116 -704 -3103
rect -304 -129 -200 -116
rect -304 -3103 -275 -129
rect -229 -3103 -200 -129
rect -304 -3116 -200 -3103
rect 200 -129 304 -116
rect 200 -3103 229 -129
rect 275 -3103 304 -129
rect 200 -3116 304 -3103
rect 704 -129 792 -116
rect 704 -3103 733 -129
rect 779 -3103 792 -129
rect 704 -3116 792 -3103
rect -792 -3361 -704 -3348
rect -792 -6335 -779 -3361
rect -733 -6335 -704 -3361
rect -792 -6348 -704 -6335
rect -304 -3361 -200 -3348
rect -304 -6335 -275 -3361
rect -229 -6335 -200 -3361
rect -304 -6348 -200 -6335
rect 200 -3361 304 -3348
rect 200 -6335 229 -3361
rect 275 -6335 304 -3361
rect 200 -6348 304 -6335
rect 704 -3361 792 -3348
rect 704 -6335 733 -3361
rect 779 -6335 792 -3361
rect 704 -6348 792 -6335
rect -792 -6593 -704 -6580
rect -792 -9567 -779 -6593
rect -733 -9567 -704 -6593
rect -792 -9580 -704 -9567
rect -304 -6593 -200 -6580
rect -304 -9567 -275 -6593
rect -229 -9567 -200 -6593
rect -304 -9580 -200 -9567
rect 200 -6593 304 -6580
rect 200 -9567 229 -6593
rect 275 -9567 304 -6593
rect 200 -9580 304 -9567
rect 704 -6593 792 -6580
rect 704 -9567 733 -6593
rect 779 -9567 792 -6593
rect 704 -9580 792 -9567
rect -792 -9825 -704 -9812
rect -792 -12799 -779 -9825
rect -733 -12799 -704 -9825
rect -792 -12812 -704 -12799
rect -304 -9825 -200 -9812
rect -304 -12799 -275 -9825
rect -229 -12799 -200 -9825
rect -304 -12812 -200 -12799
rect 200 -9825 304 -9812
rect 200 -12799 229 -9825
rect 275 -12799 304 -9825
rect 200 -12812 304 -12799
rect 704 -9825 792 -9812
rect 704 -12799 733 -9825
rect 779 -12799 792 -9825
rect 704 -12812 792 -12799
<< pdiffc >>
rect -779 9825 -733 12799
rect -275 9825 -229 12799
rect 229 9825 275 12799
rect 733 9825 779 12799
rect -779 6593 -733 9567
rect -275 6593 -229 9567
rect 229 6593 275 9567
rect 733 6593 779 9567
rect -779 3361 -733 6335
rect -275 3361 -229 6335
rect 229 3361 275 6335
rect 733 3361 779 6335
rect -779 129 -733 3103
rect -275 129 -229 3103
rect 229 129 275 3103
rect 733 129 779 3103
rect -779 -3103 -733 -129
rect -275 -3103 -229 -129
rect 229 -3103 275 -129
rect 733 -3103 779 -129
rect -779 -6335 -733 -3361
rect -275 -6335 -229 -3361
rect 229 -6335 275 -3361
rect 733 -6335 779 -3361
rect -779 -9567 -733 -6593
rect -275 -9567 -229 -6593
rect 229 -9567 275 -6593
rect 733 -9567 779 -6593
rect -779 -12799 -733 -9825
rect -275 -12799 -229 -9825
rect 229 -12799 275 -9825
rect 733 -12799 779 -9825
<< nsubdiff >>
rect -930 12926 930 12998
rect -930 12882 -858 12926
rect -930 -12882 -917 12882
rect -871 -12882 -858 12882
rect 858 12882 930 12926
rect -930 -12926 -858 -12882
rect 858 -12882 871 12882
rect 917 -12882 930 12882
rect 858 -12926 930 -12882
rect -930 -12998 930 -12926
<< nsubdiffcont >>
rect -917 -12882 -871 12882
rect 871 -12882 917 12882
<< polysilicon >>
rect -704 12891 -304 12904
rect -704 12845 -691 12891
rect -317 12845 -304 12891
rect -704 12812 -304 12845
rect -200 12891 200 12904
rect -200 12845 -187 12891
rect 187 12845 200 12891
rect -200 12812 200 12845
rect 304 12891 704 12904
rect 304 12845 317 12891
rect 691 12845 704 12891
rect 304 12812 704 12845
rect -704 9779 -304 9812
rect -704 9733 -691 9779
rect -317 9733 -304 9779
rect -704 9720 -304 9733
rect -200 9779 200 9812
rect -200 9733 -187 9779
rect 187 9733 200 9779
rect -200 9720 200 9733
rect 304 9779 704 9812
rect 304 9733 317 9779
rect 691 9733 704 9779
rect 304 9720 704 9733
rect -704 9659 -304 9672
rect -704 9613 -691 9659
rect -317 9613 -304 9659
rect -704 9580 -304 9613
rect -200 9659 200 9672
rect -200 9613 -187 9659
rect 187 9613 200 9659
rect -200 9580 200 9613
rect 304 9659 704 9672
rect 304 9613 317 9659
rect 691 9613 704 9659
rect 304 9580 704 9613
rect -704 6547 -304 6580
rect -704 6501 -691 6547
rect -317 6501 -304 6547
rect -704 6488 -304 6501
rect -200 6547 200 6580
rect -200 6501 -187 6547
rect 187 6501 200 6547
rect -200 6488 200 6501
rect 304 6547 704 6580
rect 304 6501 317 6547
rect 691 6501 704 6547
rect 304 6488 704 6501
rect -704 6427 -304 6440
rect -704 6381 -691 6427
rect -317 6381 -304 6427
rect -704 6348 -304 6381
rect -200 6427 200 6440
rect -200 6381 -187 6427
rect 187 6381 200 6427
rect -200 6348 200 6381
rect 304 6427 704 6440
rect 304 6381 317 6427
rect 691 6381 704 6427
rect 304 6348 704 6381
rect -704 3315 -304 3348
rect -704 3269 -691 3315
rect -317 3269 -304 3315
rect -704 3256 -304 3269
rect -200 3315 200 3348
rect -200 3269 -187 3315
rect 187 3269 200 3315
rect -200 3256 200 3269
rect 304 3315 704 3348
rect 304 3269 317 3315
rect 691 3269 704 3315
rect 304 3256 704 3269
rect -704 3195 -304 3208
rect -704 3149 -691 3195
rect -317 3149 -304 3195
rect -704 3116 -304 3149
rect -200 3195 200 3208
rect -200 3149 -187 3195
rect 187 3149 200 3195
rect -200 3116 200 3149
rect 304 3195 704 3208
rect 304 3149 317 3195
rect 691 3149 704 3195
rect 304 3116 704 3149
rect -704 83 -304 116
rect -704 37 -691 83
rect -317 37 -304 83
rect -704 24 -304 37
rect -200 83 200 116
rect -200 37 -187 83
rect 187 37 200 83
rect -200 24 200 37
rect 304 83 704 116
rect 304 37 317 83
rect 691 37 704 83
rect 304 24 704 37
rect -704 -37 -304 -24
rect -704 -83 -691 -37
rect -317 -83 -304 -37
rect -704 -116 -304 -83
rect -200 -37 200 -24
rect -200 -83 -187 -37
rect 187 -83 200 -37
rect -200 -116 200 -83
rect 304 -37 704 -24
rect 304 -83 317 -37
rect 691 -83 704 -37
rect 304 -116 704 -83
rect -704 -3149 -304 -3116
rect -704 -3195 -691 -3149
rect -317 -3195 -304 -3149
rect -704 -3208 -304 -3195
rect -200 -3149 200 -3116
rect -200 -3195 -187 -3149
rect 187 -3195 200 -3149
rect -200 -3208 200 -3195
rect 304 -3149 704 -3116
rect 304 -3195 317 -3149
rect 691 -3195 704 -3149
rect 304 -3208 704 -3195
rect -704 -3269 -304 -3256
rect -704 -3315 -691 -3269
rect -317 -3315 -304 -3269
rect -704 -3348 -304 -3315
rect -200 -3269 200 -3256
rect -200 -3315 -187 -3269
rect 187 -3315 200 -3269
rect -200 -3348 200 -3315
rect 304 -3269 704 -3256
rect 304 -3315 317 -3269
rect 691 -3315 704 -3269
rect 304 -3348 704 -3315
rect -704 -6381 -304 -6348
rect -704 -6427 -691 -6381
rect -317 -6427 -304 -6381
rect -704 -6440 -304 -6427
rect -200 -6381 200 -6348
rect -200 -6427 -187 -6381
rect 187 -6427 200 -6381
rect -200 -6440 200 -6427
rect 304 -6381 704 -6348
rect 304 -6427 317 -6381
rect 691 -6427 704 -6381
rect 304 -6440 704 -6427
rect -704 -6501 -304 -6488
rect -704 -6547 -691 -6501
rect -317 -6547 -304 -6501
rect -704 -6580 -304 -6547
rect -200 -6501 200 -6488
rect -200 -6547 -187 -6501
rect 187 -6547 200 -6501
rect -200 -6580 200 -6547
rect 304 -6501 704 -6488
rect 304 -6547 317 -6501
rect 691 -6547 704 -6501
rect 304 -6580 704 -6547
rect -704 -9613 -304 -9580
rect -704 -9659 -691 -9613
rect -317 -9659 -304 -9613
rect -704 -9672 -304 -9659
rect -200 -9613 200 -9580
rect -200 -9659 -187 -9613
rect 187 -9659 200 -9613
rect -200 -9672 200 -9659
rect 304 -9613 704 -9580
rect 304 -9659 317 -9613
rect 691 -9659 704 -9613
rect 304 -9672 704 -9659
rect -704 -9733 -304 -9720
rect -704 -9779 -691 -9733
rect -317 -9779 -304 -9733
rect -704 -9812 -304 -9779
rect -200 -9733 200 -9720
rect -200 -9779 -187 -9733
rect 187 -9779 200 -9733
rect -200 -9812 200 -9779
rect 304 -9733 704 -9720
rect 304 -9779 317 -9733
rect 691 -9779 704 -9733
rect 304 -9812 704 -9779
rect -704 -12845 -304 -12812
rect -704 -12891 -691 -12845
rect -317 -12891 -304 -12845
rect -704 -12904 -304 -12891
rect -200 -12845 200 -12812
rect -200 -12891 -187 -12845
rect 187 -12891 200 -12845
rect -200 -12904 200 -12891
rect 304 -12845 704 -12812
rect 304 -12891 317 -12845
rect 691 -12891 704 -12845
rect 304 -12904 704 -12891
<< polycontact >>
rect -691 12845 -317 12891
rect -187 12845 187 12891
rect 317 12845 691 12891
rect -691 9733 -317 9779
rect -187 9733 187 9779
rect 317 9733 691 9779
rect -691 9613 -317 9659
rect -187 9613 187 9659
rect 317 9613 691 9659
rect -691 6501 -317 6547
rect -187 6501 187 6547
rect 317 6501 691 6547
rect -691 6381 -317 6427
rect -187 6381 187 6427
rect 317 6381 691 6427
rect -691 3269 -317 3315
rect -187 3269 187 3315
rect 317 3269 691 3315
rect -691 3149 -317 3195
rect -187 3149 187 3195
rect 317 3149 691 3195
rect -691 37 -317 83
rect -187 37 187 83
rect 317 37 691 83
rect -691 -83 -317 -37
rect -187 -83 187 -37
rect 317 -83 691 -37
rect -691 -3195 -317 -3149
rect -187 -3195 187 -3149
rect 317 -3195 691 -3149
rect -691 -3315 -317 -3269
rect -187 -3315 187 -3269
rect 317 -3315 691 -3269
rect -691 -6427 -317 -6381
rect -187 -6427 187 -6381
rect 317 -6427 691 -6381
rect -691 -6547 -317 -6501
rect -187 -6547 187 -6501
rect 317 -6547 691 -6501
rect -691 -9659 -317 -9613
rect -187 -9659 187 -9613
rect 317 -9659 691 -9613
rect -691 -9779 -317 -9733
rect -187 -9779 187 -9733
rect 317 -9779 691 -9733
rect -691 -12891 -317 -12845
rect -187 -12891 187 -12845
rect 317 -12891 691 -12845
<< metal1 >>
rect -917 12939 917 12985
rect -917 12882 -871 12939
rect -702 12845 -691 12891
rect -317 12845 -306 12891
rect -198 12845 -187 12891
rect 187 12845 198 12891
rect 306 12845 317 12891
rect 691 12845 702 12891
rect 871 12882 917 12939
rect -779 12799 -733 12810
rect -779 9814 -733 9825
rect -275 12799 -229 12810
rect -275 9814 -229 9825
rect 229 12799 275 12810
rect 229 9814 275 9825
rect 733 12799 779 12810
rect 733 9814 779 9825
rect -702 9733 -691 9779
rect -317 9733 -306 9779
rect -198 9733 -187 9779
rect 187 9733 198 9779
rect 306 9733 317 9779
rect 691 9733 702 9779
rect -702 9613 -691 9659
rect -317 9613 -306 9659
rect -198 9613 -187 9659
rect 187 9613 198 9659
rect 306 9613 317 9659
rect 691 9613 702 9659
rect -779 9567 -733 9578
rect -779 6582 -733 6593
rect -275 9567 -229 9578
rect -275 6582 -229 6593
rect 229 9567 275 9578
rect 229 6582 275 6593
rect 733 9567 779 9578
rect 733 6582 779 6593
rect -702 6501 -691 6547
rect -317 6501 -306 6547
rect -198 6501 -187 6547
rect 187 6501 198 6547
rect 306 6501 317 6547
rect 691 6501 702 6547
rect -702 6381 -691 6427
rect -317 6381 -306 6427
rect -198 6381 -187 6427
rect 187 6381 198 6427
rect 306 6381 317 6427
rect 691 6381 702 6427
rect -779 6335 -733 6346
rect -779 3350 -733 3361
rect -275 6335 -229 6346
rect -275 3350 -229 3361
rect 229 6335 275 6346
rect 229 3350 275 3361
rect 733 6335 779 6346
rect 733 3350 779 3361
rect -702 3269 -691 3315
rect -317 3269 -306 3315
rect -198 3269 -187 3315
rect 187 3269 198 3315
rect 306 3269 317 3315
rect 691 3269 702 3315
rect -702 3149 -691 3195
rect -317 3149 -306 3195
rect -198 3149 -187 3195
rect 187 3149 198 3195
rect 306 3149 317 3195
rect 691 3149 702 3195
rect -779 3103 -733 3114
rect -779 118 -733 129
rect -275 3103 -229 3114
rect -275 118 -229 129
rect 229 3103 275 3114
rect 229 118 275 129
rect 733 3103 779 3114
rect 733 118 779 129
rect -702 37 -691 83
rect -317 37 -306 83
rect -198 37 -187 83
rect 187 37 198 83
rect 306 37 317 83
rect 691 37 702 83
rect -702 -83 -691 -37
rect -317 -83 -306 -37
rect -198 -83 -187 -37
rect 187 -83 198 -37
rect 306 -83 317 -37
rect 691 -83 702 -37
rect -779 -129 -733 -118
rect -779 -3114 -733 -3103
rect -275 -129 -229 -118
rect -275 -3114 -229 -3103
rect 229 -129 275 -118
rect 229 -3114 275 -3103
rect 733 -129 779 -118
rect 733 -3114 779 -3103
rect -702 -3195 -691 -3149
rect -317 -3195 -306 -3149
rect -198 -3195 -187 -3149
rect 187 -3195 198 -3149
rect 306 -3195 317 -3149
rect 691 -3195 702 -3149
rect -702 -3315 -691 -3269
rect -317 -3315 -306 -3269
rect -198 -3315 -187 -3269
rect 187 -3315 198 -3269
rect 306 -3315 317 -3269
rect 691 -3315 702 -3269
rect -779 -3361 -733 -3350
rect -779 -6346 -733 -6335
rect -275 -3361 -229 -3350
rect -275 -6346 -229 -6335
rect 229 -3361 275 -3350
rect 229 -6346 275 -6335
rect 733 -3361 779 -3350
rect 733 -6346 779 -6335
rect -702 -6427 -691 -6381
rect -317 -6427 -306 -6381
rect -198 -6427 -187 -6381
rect 187 -6427 198 -6381
rect 306 -6427 317 -6381
rect 691 -6427 702 -6381
rect -702 -6547 -691 -6501
rect -317 -6547 -306 -6501
rect -198 -6547 -187 -6501
rect 187 -6547 198 -6501
rect 306 -6547 317 -6501
rect 691 -6547 702 -6501
rect -779 -6593 -733 -6582
rect -779 -9578 -733 -9567
rect -275 -6593 -229 -6582
rect -275 -9578 -229 -9567
rect 229 -6593 275 -6582
rect 229 -9578 275 -9567
rect 733 -6593 779 -6582
rect 733 -9578 779 -9567
rect -702 -9659 -691 -9613
rect -317 -9659 -306 -9613
rect -198 -9659 -187 -9613
rect 187 -9659 198 -9613
rect 306 -9659 317 -9613
rect 691 -9659 702 -9613
rect -702 -9779 -691 -9733
rect -317 -9779 -306 -9733
rect -198 -9779 -187 -9733
rect 187 -9779 198 -9733
rect 306 -9779 317 -9733
rect 691 -9779 702 -9733
rect -779 -9825 -733 -9814
rect -779 -12810 -733 -12799
rect -275 -9825 -229 -9814
rect -275 -12810 -229 -12799
rect 229 -9825 275 -9814
rect 229 -12810 275 -12799
rect 733 -9825 779 -9814
rect 733 -12810 779 -12799
rect -917 -12939 -871 -12882
rect -702 -12891 -691 -12845
rect -317 -12891 -306 -12845
rect -198 -12891 -187 -12845
rect 187 -12891 198 -12845
rect 306 -12891 317 -12845
rect 691 -12891 702 -12845
rect 871 -12939 917 -12882
rect -917 -12985 917 -12939
<< properties >>
string FIXED_BBOX -894 -12962 894 12962
string gencell pfet_03v3
string library gf180mcu
string parameters w 15.0 l 2.0 m 8 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
