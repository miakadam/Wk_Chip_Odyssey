magic
tech gf180mcuD
magscale 1 10
timestamp 1758180527
<< nwell >>
rect 5065 2693 6205 3333
rect 6445 1255 7025 2427
rect 7415 2360 8455 2980
rect 8845 1255 9425 2427
rect 6217 -210 9653 -190
rect 4897 -790 5477 -210
rect 5757 -790 10113 -210
rect 10393 -790 10973 -210
rect 6217 -810 9653 -790
<< pwell >>
rect 7415 1540 8455 2160
rect 6445 455 7025 1227
rect 8845 455 9425 1227
rect 6079 -1966 9791 -1146
rect 9415 -2304 9495 -2182
rect 5717 -5100 10153 -2304
<< nmos >>
rect 5265 2273 5325 2443
rect 5435 2273 5495 2443
rect 5605 2273 5665 2443
rect 5775 2273 5835 2443
rect 5945 2273 6005 2443
rect 7665 1750 7745 1950
rect 8125 1750 8205 1950
rect 6695 617 6775 1017
rect 9095 617 9175 1017
rect 6329 -1756 6529 -1356
rect 6633 -1756 6833 -1356
rect 6937 -1756 7137 -1356
rect 7241 -1756 7441 -1356
rect 7545 -1756 7745 -1356
rect 8125 -1756 8325 -1356
rect 8429 -1756 8629 -1356
rect 8733 -1756 8933 -1356
rect 9037 -1756 9237 -1356
rect 9341 -1756 9541 -1356
rect 6163 -3141 6363 -2841
rect 6467 -3141 6667 -2841
rect 6771 -3141 6971 -2841
rect 7075 -3141 7275 -2841
rect 7379 -3141 7579 -2841
rect 7683 -3141 7883 -2841
rect 7987 -3141 8187 -2841
rect 8291 -3141 8491 -2841
rect 8595 -3141 8795 -2841
rect 8899 -3141 9099 -2841
rect 9203 -3141 9403 -2841
rect 9507 -3141 9707 -2841
rect 6163 -4104 6363 -3804
rect 6467 -4104 6667 -3804
rect 6771 -4104 6971 -3804
rect 7075 -4104 7275 -3804
rect 7379 -4104 7579 -3804
rect 7683 -4104 7883 -3804
rect 7987 -4104 8187 -3804
rect 8291 -4104 8491 -3804
rect 8595 -4104 8795 -3804
rect 8899 -4104 9099 -3804
rect 9203 -4104 9403 -3804
rect 9507 -4104 9707 -3804
rect 7711 -4890 7791 -4730
rect 7895 -4890 7975 -4730
rect 8079 -4890 8159 -4730
<< pmos >>
rect 5265 2783 5325 3123
rect 5435 2783 5495 3123
rect 5605 2783 5665 3123
rect 5775 2783 5835 3123
rect 5945 2783 6005 3123
rect 7665 2570 7745 2770
rect 8125 2570 8205 2770
rect 6695 1465 6775 2265
rect 9095 1465 9175 2265
rect 5147 -580 5227 -420
rect 6007 -580 6087 -420
rect 6467 -600 6667 -400
rect 6771 -600 6971 -400
rect 7075 -600 7275 -400
rect 7379 -600 7579 -400
rect 7683 -600 7883 -400
rect 7987 -600 8187 -400
rect 8291 -600 8491 -400
rect 8595 -600 8795 -400
rect 8899 -600 9099 -400
rect 9203 -600 9403 -400
rect 9783 -580 9863 -420
rect 10643 -580 10723 -420
<< ndiff >>
rect 5165 2381 5265 2443
rect 5165 2335 5187 2381
rect 5233 2335 5265 2381
rect 5165 2273 5265 2335
rect 5325 2381 5435 2443
rect 5325 2335 5357 2381
rect 5403 2335 5435 2381
rect 5325 2273 5435 2335
rect 5495 2381 5605 2443
rect 5495 2335 5527 2381
rect 5573 2335 5605 2381
rect 5495 2273 5605 2335
rect 5665 2381 5775 2443
rect 5665 2335 5697 2381
rect 5743 2335 5775 2381
rect 5665 2273 5775 2335
rect 5835 2381 5945 2443
rect 5835 2335 5867 2381
rect 5913 2335 5945 2381
rect 5835 2273 5945 2335
rect 6005 2381 6105 2443
rect 6005 2335 6037 2381
rect 6083 2335 6105 2381
rect 6005 2273 6105 2335
rect 7577 1937 7665 1950
rect 7577 1763 7590 1937
rect 7636 1763 7665 1937
rect 7577 1750 7665 1763
rect 7745 1937 7833 1950
rect 7745 1763 7774 1937
rect 7820 1763 7833 1937
rect 7745 1750 7833 1763
rect 8037 1937 8125 1950
rect 8037 1763 8050 1937
rect 8096 1763 8125 1937
rect 8037 1750 8125 1763
rect 8205 1937 8293 1950
rect 8205 1763 8234 1937
rect 8280 1763 8293 1937
rect 8205 1750 8293 1763
rect 6607 1004 6695 1017
rect 6607 630 6620 1004
rect 6666 630 6695 1004
rect 6607 617 6695 630
rect 6775 1004 6863 1017
rect 6775 630 6804 1004
rect 6850 630 6863 1004
rect 6775 617 6863 630
rect 9007 1004 9095 1017
rect 9007 630 9020 1004
rect 9066 630 9095 1004
rect 9007 617 9095 630
rect 9175 1004 9263 1017
rect 9175 630 9204 1004
rect 9250 630 9263 1004
rect 9175 617 9263 630
rect 6241 -1369 6329 -1356
rect 6241 -1743 6254 -1369
rect 6300 -1743 6329 -1369
rect 6241 -1756 6329 -1743
rect 6529 -1369 6633 -1356
rect 6529 -1743 6558 -1369
rect 6604 -1743 6633 -1369
rect 6529 -1756 6633 -1743
rect 6833 -1369 6937 -1356
rect 6833 -1743 6862 -1369
rect 6908 -1743 6937 -1369
rect 6833 -1756 6937 -1743
rect 7137 -1369 7241 -1356
rect 7137 -1743 7166 -1369
rect 7212 -1743 7241 -1369
rect 7137 -1756 7241 -1743
rect 7441 -1369 7545 -1356
rect 7441 -1743 7470 -1369
rect 7516 -1743 7545 -1369
rect 7441 -1756 7545 -1743
rect 7745 -1369 7833 -1356
rect 7745 -1743 7774 -1369
rect 7820 -1743 7833 -1369
rect 7745 -1756 7833 -1743
rect 8037 -1369 8125 -1356
rect 8037 -1743 8050 -1369
rect 8096 -1743 8125 -1369
rect 8037 -1756 8125 -1743
rect 8325 -1369 8429 -1356
rect 8325 -1743 8354 -1369
rect 8400 -1743 8429 -1369
rect 8325 -1756 8429 -1743
rect 8629 -1369 8733 -1356
rect 8629 -1743 8658 -1369
rect 8704 -1743 8733 -1369
rect 8629 -1756 8733 -1743
rect 8933 -1369 9037 -1356
rect 8933 -1743 8962 -1369
rect 9008 -1743 9037 -1369
rect 8933 -1756 9037 -1743
rect 9237 -1369 9341 -1356
rect 9237 -1743 9266 -1369
rect 9312 -1743 9341 -1369
rect 9237 -1756 9341 -1743
rect 9541 -1369 9629 -1356
rect 9541 -1743 9570 -1369
rect 9616 -1743 9629 -1369
rect 9541 -1756 9629 -1743
rect 6075 -2854 6163 -2841
rect 6075 -3128 6088 -2854
rect 6134 -3128 6163 -2854
rect 6075 -3141 6163 -3128
rect 6363 -2854 6467 -2841
rect 6363 -3128 6392 -2854
rect 6438 -3128 6467 -2854
rect 6363 -3141 6467 -3128
rect 6667 -2854 6771 -2841
rect 6667 -3128 6696 -2854
rect 6742 -3128 6771 -2854
rect 6667 -3141 6771 -3128
rect 6971 -2854 7075 -2841
rect 6971 -3128 7000 -2854
rect 7046 -3128 7075 -2854
rect 6971 -3141 7075 -3128
rect 7275 -2854 7379 -2841
rect 7275 -3128 7304 -2854
rect 7350 -3128 7379 -2854
rect 7275 -3141 7379 -3128
rect 7579 -2854 7683 -2841
rect 7579 -3128 7608 -2854
rect 7654 -3128 7683 -2854
rect 7579 -3141 7683 -3128
rect 7883 -2854 7987 -2841
rect 7883 -3128 7912 -2854
rect 7958 -3128 7987 -2854
rect 7883 -3141 7987 -3128
rect 8187 -2854 8291 -2841
rect 8187 -3128 8216 -2854
rect 8262 -3128 8291 -2854
rect 8187 -3141 8291 -3128
rect 8491 -2854 8595 -2841
rect 8491 -3128 8520 -2854
rect 8566 -3128 8595 -2854
rect 8491 -3141 8595 -3128
rect 8795 -2854 8899 -2841
rect 8795 -3128 8824 -2854
rect 8870 -3128 8899 -2854
rect 8795 -3141 8899 -3128
rect 9099 -2854 9203 -2841
rect 9099 -3128 9128 -2854
rect 9174 -3128 9203 -2854
rect 9099 -3141 9203 -3128
rect 9403 -2854 9507 -2841
rect 9403 -3128 9432 -2854
rect 9478 -3128 9507 -2854
rect 9403 -3141 9507 -3128
rect 9707 -2854 9795 -2841
rect 9707 -3128 9736 -2854
rect 9782 -3128 9795 -2854
rect 9707 -3141 9795 -3128
rect 6075 -3817 6163 -3804
rect 6075 -4091 6088 -3817
rect 6134 -4091 6163 -3817
rect 6075 -4104 6163 -4091
rect 6363 -3817 6467 -3804
rect 6363 -4091 6392 -3817
rect 6438 -4091 6467 -3817
rect 6363 -4104 6467 -4091
rect 6667 -3817 6771 -3804
rect 6667 -4091 6696 -3817
rect 6742 -4091 6771 -3817
rect 6667 -4104 6771 -4091
rect 6971 -3817 7075 -3804
rect 6971 -4091 7000 -3817
rect 7046 -4091 7075 -3817
rect 6971 -4104 7075 -4091
rect 7275 -3817 7379 -3804
rect 7275 -4091 7304 -3817
rect 7350 -4091 7379 -3817
rect 7275 -4104 7379 -4091
rect 7579 -3817 7683 -3804
rect 7579 -4091 7608 -3817
rect 7654 -4091 7683 -3817
rect 7579 -4104 7683 -4091
rect 7883 -3817 7987 -3804
rect 7883 -4091 7912 -3817
rect 7958 -4091 7987 -3817
rect 7883 -4104 7987 -4091
rect 8187 -3817 8291 -3804
rect 8187 -4091 8216 -3817
rect 8262 -4091 8291 -3817
rect 8187 -4104 8291 -4091
rect 8491 -3817 8595 -3804
rect 8491 -4091 8520 -3817
rect 8566 -4091 8595 -3817
rect 8491 -4104 8595 -4091
rect 8795 -3817 8899 -3804
rect 8795 -4091 8824 -3817
rect 8870 -4091 8899 -3817
rect 8795 -4104 8899 -4091
rect 9099 -3817 9203 -3804
rect 9099 -4091 9128 -3817
rect 9174 -4091 9203 -3817
rect 9099 -4104 9203 -4091
rect 9403 -3817 9507 -3804
rect 9403 -4091 9432 -3817
rect 9478 -4091 9507 -3817
rect 9403 -4104 9507 -4091
rect 9707 -3817 9795 -3804
rect 9707 -4091 9736 -3817
rect 9782 -4091 9795 -3817
rect 9707 -4104 9795 -4091
rect 7623 -4743 7711 -4730
rect 7623 -4877 7636 -4743
rect 7682 -4877 7711 -4743
rect 7623 -4890 7711 -4877
rect 7791 -4743 7895 -4730
rect 7791 -4877 7820 -4743
rect 7866 -4877 7895 -4743
rect 7791 -4890 7895 -4877
rect 7975 -4743 8079 -4730
rect 7975 -4877 8004 -4743
rect 8050 -4877 8079 -4743
rect 7975 -4890 8079 -4877
rect 8159 -4743 8247 -4730
rect 8159 -4877 8188 -4743
rect 8234 -4877 8247 -4743
rect 8159 -4890 8247 -4877
<< pdiff >>
rect 5165 3070 5265 3123
rect 5165 2836 5187 3070
rect 5233 2836 5265 3070
rect 5165 2783 5265 2836
rect 5325 3095 5435 3123
rect 5325 2861 5357 3095
rect 5403 2861 5435 3095
rect 5325 2783 5435 2861
rect 5495 3070 5605 3123
rect 5495 2836 5527 3070
rect 5573 2836 5605 3070
rect 5495 2783 5605 2836
rect 5665 3095 5775 3123
rect 5665 2861 5697 3095
rect 5743 2861 5775 3095
rect 5665 2783 5775 2861
rect 5835 3070 5945 3123
rect 5835 2836 5867 3070
rect 5913 2836 5945 3070
rect 5835 2783 5945 2836
rect 6005 3070 6105 3123
rect 6005 2836 6037 3070
rect 6083 2836 6105 3070
rect 6005 2783 6105 2836
rect 7577 2757 7665 2770
rect 7577 2583 7590 2757
rect 7636 2583 7665 2757
rect 7577 2570 7665 2583
rect 7745 2757 7833 2770
rect 7745 2583 7774 2757
rect 7820 2583 7833 2757
rect 7745 2570 7833 2583
rect 8037 2757 8125 2770
rect 8037 2583 8050 2757
rect 8096 2583 8125 2757
rect 8037 2570 8125 2583
rect 8205 2757 8293 2770
rect 8205 2583 8234 2757
rect 8280 2583 8293 2757
rect 8205 2570 8293 2583
rect 6607 2252 6695 2265
rect 6607 1478 6620 2252
rect 6666 1478 6695 2252
rect 6607 1465 6695 1478
rect 6775 2252 6863 2265
rect 6775 1478 6804 2252
rect 6850 1478 6863 2252
rect 6775 1465 6863 1478
rect 9007 2252 9095 2265
rect 9007 1478 9020 2252
rect 9066 1478 9095 2252
rect 9007 1465 9095 1478
rect 9175 2252 9263 2265
rect 9175 1478 9204 2252
rect 9250 1478 9263 2252
rect 9175 1465 9263 1478
rect 5059 -433 5147 -420
rect 5059 -567 5072 -433
rect 5118 -567 5147 -433
rect 5059 -580 5147 -567
rect 5227 -433 5315 -420
rect 5227 -567 5256 -433
rect 5302 -567 5315 -433
rect 5227 -580 5315 -567
rect 5919 -433 6007 -420
rect 5919 -567 5932 -433
rect 5978 -567 6007 -433
rect 5919 -580 6007 -567
rect 6087 -433 6175 -420
rect 6087 -567 6116 -433
rect 6162 -567 6175 -433
rect 6087 -580 6175 -567
rect 6379 -413 6467 -400
rect 6379 -587 6392 -413
rect 6438 -587 6467 -413
rect 6379 -600 6467 -587
rect 6667 -413 6771 -400
rect 6667 -587 6696 -413
rect 6742 -587 6771 -413
rect 6667 -600 6771 -587
rect 6971 -413 7075 -400
rect 6971 -587 7000 -413
rect 7046 -587 7075 -413
rect 6971 -600 7075 -587
rect 7275 -413 7379 -400
rect 7275 -587 7304 -413
rect 7350 -587 7379 -413
rect 7275 -600 7379 -587
rect 7579 -413 7683 -400
rect 7579 -587 7608 -413
rect 7654 -587 7683 -413
rect 7579 -600 7683 -587
rect 7883 -413 7987 -400
rect 7883 -587 7912 -413
rect 7958 -587 7987 -413
rect 7883 -600 7987 -587
rect 8187 -413 8291 -400
rect 8187 -587 8216 -413
rect 8262 -587 8291 -413
rect 8187 -600 8291 -587
rect 8491 -413 8595 -400
rect 8491 -587 8520 -413
rect 8566 -587 8595 -413
rect 8491 -600 8595 -587
rect 8795 -413 8899 -400
rect 8795 -587 8824 -413
rect 8870 -587 8899 -413
rect 8795 -600 8899 -587
rect 9099 -413 9203 -400
rect 9099 -587 9128 -413
rect 9174 -587 9203 -413
rect 9099 -600 9203 -587
rect 9403 -413 9491 -400
rect 9403 -587 9432 -413
rect 9478 -587 9491 -413
rect 9403 -600 9491 -587
rect 9695 -433 9783 -420
rect 9695 -567 9708 -433
rect 9754 -567 9783 -433
rect 9695 -580 9783 -567
rect 9863 -433 9951 -420
rect 9863 -567 9892 -433
rect 9938 -567 9951 -433
rect 9863 -580 9951 -567
rect 10555 -433 10643 -420
rect 10555 -567 10568 -433
rect 10614 -567 10643 -433
rect 10555 -580 10643 -567
rect 10723 -433 10811 -420
rect 10723 -567 10752 -433
rect 10798 -567 10811 -433
rect 10723 -580 10811 -567
<< ndiffc >>
rect 5187 2335 5233 2381
rect 5357 2335 5403 2381
rect 5527 2335 5573 2381
rect 5697 2335 5743 2381
rect 5867 2335 5913 2381
rect 6037 2335 6083 2381
rect 7590 1763 7636 1937
rect 7774 1763 7820 1937
rect 8050 1763 8096 1937
rect 8234 1763 8280 1937
rect 6620 630 6666 1004
rect 6804 630 6850 1004
rect 9020 630 9066 1004
rect 9204 630 9250 1004
rect 6254 -1743 6300 -1369
rect 6558 -1743 6604 -1369
rect 6862 -1743 6908 -1369
rect 7166 -1743 7212 -1369
rect 7470 -1743 7516 -1369
rect 7774 -1743 7820 -1369
rect 8050 -1743 8096 -1369
rect 8354 -1743 8400 -1369
rect 8658 -1743 8704 -1369
rect 8962 -1743 9008 -1369
rect 9266 -1743 9312 -1369
rect 9570 -1743 9616 -1369
rect 6088 -3128 6134 -2854
rect 6392 -3128 6438 -2854
rect 6696 -3128 6742 -2854
rect 7000 -3128 7046 -2854
rect 7304 -3128 7350 -2854
rect 7608 -3128 7654 -2854
rect 7912 -3128 7958 -2854
rect 8216 -3128 8262 -2854
rect 8520 -3128 8566 -2854
rect 8824 -3128 8870 -2854
rect 9128 -3128 9174 -2854
rect 9432 -3128 9478 -2854
rect 9736 -3128 9782 -2854
rect 6088 -4091 6134 -3817
rect 6392 -4091 6438 -3817
rect 6696 -4091 6742 -3817
rect 7000 -4091 7046 -3817
rect 7304 -4091 7350 -3817
rect 7608 -4091 7654 -3817
rect 7912 -4091 7958 -3817
rect 8216 -4091 8262 -3817
rect 8520 -4091 8566 -3817
rect 8824 -4091 8870 -3817
rect 9128 -4091 9174 -3817
rect 9432 -4091 9478 -3817
rect 9736 -4091 9782 -3817
rect 7636 -4877 7682 -4743
rect 7820 -4877 7866 -4743
rect 8004 -4877 8050 -4743
rect 8188 -4877 8234 -4743
<< pdiffc >>
rect 5187 2836 5233 3070
rect 5357 2861 5403 3095
rect 5527 2836 5573 3070
rect 5697 2861 5743 3095
rect 5867 2836 5913 3070
rect 6037 2836 6083 3070
rect 7590 2583 7636 2757
rect 7774 2583 7820 2757
rect 8050 2583 8096 2757
rect 8234 2583 8280 2757
rect 6620 1478 6666 2252
rect 6804 1478 6850 2252
rect 9020 1478 9066 2252
rect 9204 1478 9250 2252
rect 5072 -567 5118 -433
rect 5256 -567 5302 -433
rect 5932 -567 5978 -433
rect 6116 -567 6162 -433
rect 6392 -587 6438 -413
rect 6696 -587 6742 -413
rect 7000 -587 7046 -413
rect 7304 -587 7350 -413
rect 7608 -587 7654 -413
rect 7912 -587 7958 -413
rect 8216 -587 8262 -413
rect 8520 -587 8566 -413
rect 8824 -587 8870 -413
rect 9128 -587 9174 -413
rect 9432 -587 9478 -413
rect 9708 -567 9754 -433
rect 9892 -567 9938 -433
rect 10568 -567 10614 -433
rect 10752 -567 10798 -433
<< psubdiff >>
rect 5265 2181 5415 2203
rect 5265 2135 5317 2181
rect 5363 2135 5415 2181
rect 5265 2113 5415 2135
rect 5505 2181 5655 2203
rect 5505 2135 5557 2181
rect 5603 2135 5655 2181
rect 5505 2113 5655 2135
rect 5745 2181 5895 2203
rect 5745 2135 5797 2181
rect 5843 2135 5895 2181
rect 5745 2113 5895 2135
rect 5985 2181 6135 2203
rect 5985 2135 6037 2181
rect 6083 2135 6135 2181
rect 5985 2113 6135 2135
rect 7439 2064 8431 2136
rect 7439 2020 7511 2064
rect 7439 1680 7452 2020
rect 7498 1680 7511 2020
rect 7899 2020 7971 2064
rect 7439 1636 7511 1680
rect 7899 1680 7912 2020
rect 7958 1680 7971 2020
rect 8359 2020 8431 2064
rect 7899 1636 7971 1680
rect 8359 1680 8372 2020
rect 8418 1680 8431 2020
rect 8359 1636 8431 1680
rect 7439 1564 8431 1636
rect 6469 1131 7001 1203
rect 6469 551 6541 1131
rect 6929 551 7001 1131
rect 6469 538 7001 551
rect 6469 492 6585 538
rect 6885 492 7001 538
rect 6469 479 7001 492
rect 8869 1131 9401 1203
rect 8869 551 8941 1131
rect 9329 551 9401 1131
rect 8869 538 9401 551
rect 8869 492 8985 538
rect 9285 492 9401 538
rect 8869 479 9401 492
rect 6103 -1242 9767 -1170
rect 6103 -1286 6175 -1242
rect 6103 -1826 6116 -1286
rect 6162 -1826 6175 -1286
rect 7899 -1286 7971 -1242
rect 6103 -1870 6175 -1826
rect 7899 -1826 7912 -1286
rect 7958 -1826 7971 -1286
rect 9695 -1286 9767 -1242
rect 7899 -1870 7971 -1826
rect 9695 -1826 9708 -1286
rect 9754 -1826 9767 -1286
rect 9695 -1870 9767 -1826
rect 6103 -1942 9767 -1870
rect 5742 -2401 10128 -2329
rect 5742 -2500 5942 -2401
rect 5742 -3000 5792 -2500
rect 5892 -3000 5942 -2500
rect 9928 -2500 10128 -2401
rect 5742 -3945 5942 -3000
rect 9928 -3000 9978 -2500
rect 10078 -3000 10128 -2500
rect 5742 -4445 5792 -3945
rect 5892 -4445 5942 -3945
rect 9928 -3945 10128 -3000
rect 5742 -4544 5942 -4445
rect 9928 -4445 9978 -3945
rect 10078 -4445 10128 -3945
rect 9928 -4544 10128 -4445
rect 5742 -4616 10128 -4544
rect 7485 -4660 7557 -4616
rect 7485 -4960 7498 -4660
rect 7544 -4960 7557 -4660
rect 8313 -4660 8385 -4616
rect 7485 -5004 7557 -4960
rect 8313 -4960 8326 -4660
rect 8372 -4960 8385 -4660
rect 8313 -5004 8385 -4960
rect 7485 -5076 8385 -5004
<< nsubdiff >>
rect 5265 3261 5415 3283
rect 5265 3215 5317 3261
rect 5363 3215 5415 3261
rect 5265 3193 5415 3215
rect 5505 3261 5655 3283
rect 5505 3215 5557 3261
rect 5603 3215 5655 3261
rect 5505 3193 5655 3215
rect 5745 3261 5895 3283
rect 5745 3215 5797 3261
rect 5843 3215 5895 3261
rect 5745 3193 5895 3215
rect 5985 3261 6135 3283
rect 5985 3215 6037 3261
rect 6083 3215 6135 3261
rect 5985 3193 6135 3215
rect 7439 2884 8431 2956
rect 7439 2840 7511 2884
rect 7439 2500 7452 2840
rect 7498 2500 7511 2840
rect 7899 2840 7971 2884
rect 7439 2456 7511 2500
rect 7899 2500 7912 2840
rect 7958 2500 7971 2840
rect 8359 2840 8431 2884
rect 7899 2456 7971 2500
rect 8359 2500 8372 2840
rect 8418 2500 8431 2840
rect 8359 2456 8431 2500
rect 6469 2390 7001 2403
rect 6469 2344 6585 2390
rect 6885 2344 7001 2390
rect 7439 2384 8431 2456
rect 8869 2390 9401 2403
rect 6469 2331 7001 2344
rect 6469 1351 6541 2331
rect 6929 1351 7001 2331
rect 8869 2344 8985 2390
rect 9285 2344 9401 2390
rect 8869 2331 9401 2344
rect 6469 1279 7001 1351
rect 8869 1351 8941 2331
rect 9329 1351 9401 2331
rect 8869 1279 9401 1351
rect 6241 -234 9629 -214
rect 4921 -306 5453 -234
rect 4921 -350 4993 -306
rect 4921 -650 4934 -350
rect 4980 -650 4993 -350
rect 5381 -350 5453 -306
rect 4921 -694 4993 -650
rect 5381 -650 5394 -350
rect 5440 -650 5453 -350
rect 5381 -694 5453 -650
rect 4921 -766 5453 -694
rect 5781 -286 10089 -234
rect 5781 -306 6313 -286
rect 5781 -350 5853 -306
rect 5781 -650 5794 -350
rect 5840 -650 5853 -350
rect 6241 -330 6313 -306
rect 9557 -306 10089 -286
rect 5781 -694 5853 -650
rect 6241 -670 6254 -330
rect 6300 -670 6313 -330
rect 9557 -330 9629 -306
rect 6241 -694 6313 -670
rect 9557 -670 9570 -330
rect 9616 -670 9629 -330
rect 10017 -350 10089 -306
rect 5781 -714 6313 -694
rect 9557 -694 9629 -670
rect 10017 -650 10030 -350
rect 10076 -650 10089 -350
rect 10017 -694 10089 -650
rect 9557 -714 10089 -694
rect 5781 -766 10089 -714
rect 10417 -306 10949 -234
rect 10417 -350 10489 -306
rect 10417 -650 10430 -350
rect 10476 -650 10489 -350
rect 10877 -350 10949 -306
rect 10417 -694 10489 -650
rect 10877 -650 10890 -350
rect 10936 -650 10949 -350
rect 10877 -694 10949 -650
rect 10417 -766 10949 -694
rect 6241 -786 9629 -766
<< psubdiffcont >>
rect 5317 2135 5363 2181
rect 5557 2135 5603 2181
rect 5797 2135 5843 2181
rect 6037 2135 6083 2181
rect 7452 1680 7498 2020
rect 7912 1680 7958 2020
rect 8372 1680 8418 2020
rect 6585 492 6885 538
rect 8985 492 9285 538
rect 6116 -1826 6162 -1286
rect 7912 -1826 7958 -1286
rect 9708 -1826 9754 -1286
rect 5792 -3000 5892 -2500
rect 9978 -3000 10078 -2500
rect 5792 -4445 5892 -3945
rect 9978 -4445 10078 -3945
rect 7498 -4960 7544 -4660
rect 8326 -4960 8372 -4660
<< nsubdiffcont >>
rect 5317 3215 5363 3261
rect 5557 3215 5603 3261
rect 5797 3215 5843 3261
rect 6037 3215 6083 3261
rect 7452 2500 7498 2840
rect 7912 2500 7958 2840
rect 8372 2500 8418 2840
rect 6585 2344 6885 2390
rect 8985 2344 9285 2390
rect 4934 -650 4980 -350
rect 5394 -650 5440 -350
rect 5794 -650 5840 -350
rect 6254 -670 6300 -330
rect 9570 -670 9616 -330
rect 10030 -650 10076 -350
rect 10430 -650 10476 -350
rect 10890 -650 10936 -350
<< polysilicon >>
rect 5265 3123 5325 3173
rect 5435 3123 5495 3173
rect 5605 3123 5665 3173
rect 5775 3123 5835 3173
rect 5945 3123 6005 3173
rect 5265 2763 5325 2783
rect 5435 2763 5495 2783
rect 5605 2763 5665 2783
rect 5775 2763 5835 2783
rect 5265 2753 5835 2763
rect 5265 2726 5895 2753
rect 5265 2703 5822 2726
rect 5435 2523 5495 2703
rect 5775 2680 5822 2703
rect 5868 2680 5895 2726
rect 5775 2653 5895 2680
rect 5775 2523 5835 2653
rect 5945 2603 6005 2783
rect 5265 2463 5835 2523
rect 5885 2576 6005 2603
rect 5885 2530 5912 2576
rect 5958 2530 6005 2576
rect 5885 2503 6005 2530
rect 5265 2443 5325 2463
rect 5435 2443 5495 2463
rect 5605 2443 5665 2463
rect 5775 2443 5835 2463
rect 5945 2443 6005 2503
rect 7665 2849 7745 2862
rect 7665 2803 7678 2849
rect 7732 2803 7745 2849
rect 7665 2770 7745 2803
rect 7665 2537 7745 2570
rect 7665 2491 7678 2537
rect 7732 2491 7745 2537
rect 7665 2478 7745 2491
rect 8125 2849 8205 2862
rect 8125 2803 8138 2849
rect 8192 2803 8205 2849
rect 8125 2770 8205 2803
rect 8125 2537 8205 2570
rect 8125 2491 8138 2537
rect 8192 2491 8205 2537
rect 8125 2478 8205 2491
rect 5265 2223 5325 2273
rect 5435 2223 5495 2273
rect 5605 2223 5665 2273
rect 5775 2223 5835 2273
rect 5945 2223 6005 2273
rect 6695 2265 6775 2309
rect 6695 1432 6775 1465
rect 6695 1386 6708 1432
rect 6762 1386 6775 1432
rect 6695 1373 6775 1386
rect 7665 2029 7745 2042
rect 7665 1983 7678 2029
rect 7732 1983 7745 2029
rect 7665 1950 7745 1983
rect 7665 1717 7745 1750
rect 7665 1671 7678 1717
rect 7732 1671 7745 1717
rect 7665 1658 7745 1671
rect 8125 2029 8205 2042
rect 8125 1983 8138 2029
rect 8192 1983 8205 2029
rect 8125 1950 8205 1983
rect 8125 1717 8205 1750
rect 8125 1671 8138 1717
rect 8192 1671 8205 1717
rect 8125 1658 8205 1671
rect 9095 2265 9175 2309
rect 9095 1432 9175 1465
rect 9095 1386 9108 1432
rect 9162 1386 9175 1432
rect 9095 1373 9175 1386
rect 6695 1096 6775 1109
rect 6695 1050 6708 1096
rect 6762 1050 6775 1096
rect 6695 1017 6775 1050
rect 6695 573 6775 617
rect 9095 1096 9175 1109
rect 9095 1050 9108 1096
rect 9162 1050 9175 1096
rect 9095 1017 9175 1050
rect 9095 573 9175 617
rect 5147 -341 5227 -328
rect 5147 -387 5160 -341
rect 5214 -387 5227 -341
rect 5147 -420 5227 -387
rect 5147 -613 5227 -580
rect 5147 -659 5160 -613
rect 5214 -659 5227 -613
rect 5147 -672 5227 -659
rect 6007 -341 6087 -328
rect 6007 -387 6020 -341
rect 6074 -387 6087 -341
rect 6007 -420 6087 -387
rect 6007 -613 6087 -580
rect 6007 -659 6020 -613
rect 6074 -659 6087 -613
rect 6007 -672 6087 -659
rect 6467 -321 6667 -308
rect 6467 -367 6480 -321
rect 6654 -367 6667 -321
rect 6467 -400 6667 -367
rect 6771 -321 6971 -308
rect 6771 -367 6784 -321
rect 6958 -367 6971 -321
rect 6771 -400 6971 -367
rect 7075 -321 7275 -308
rect 7075 -367 7088 -321
rect 7262 -367 7275 -321
rect 7075 -400 7275 -367
rect 7379 -321 7579 -308
rect 7379 -367 7392 -321
rect 7566 -367 7579 -321
rect 7379 -400 7579 -367
rect 7683 -321 7883 -308
rect 7683 -367 7696 -321
rect 7870 -367 7883 -321
rect 7683 -400 7883 -367
rect 7987 -321 8187 -308
rect 7987 -367 8000 -321
rect 8174 -367 8187 -321
rect 7987 -400 8187 -367
rect 8291 -321 8491 -308
rect 8291 -367 8304 -321
rect 8478 -367 8491 -321
rect 8291 -400 8491 -367
rect 8595 -321 8795 -308
rect 8595 -367 8608 -321
rect 8782 -367 8795 -321
rect 8595 -400 8795 -367
rect 8899 -321 9099 -308
rect 8899 -367 8912 -321
rect 9086 -367 9099 -321
rect 8899 -400 9099 -367
rect 9203 -321 9403 -308
rect 9203 -367 9216 -321
rect 9390 -367 9403 -321
rect 9203 -400 9403 -367
rect 6467 -633 6667 -600
rect 6467 -679 6480 -633
rect 6654 -679 6667 -633
rect 6467 -692 6667 -679
rect 6771 -633 6971 -600
rect 6771 -679 6784 -633
rect 6958 -679 6971 -633
rect 6771 -692 6971 -679
rect 7075 -633 7275 -600
rect 7075 -679 7088 -633
rect 7262 -679 7275 -633
rect 7075 -692 7275 -679
rect 7379 -633 7579 -600
rect 7379 -679 7392 -633
rect 7566 -679 7579 -633
rect 7379 -692 7579 -679
rect 7683 -633 7883 -600
rect 7683 -679 7696 -633
rect 7870 -679 7883 -633
rect 7683 -692 7883 -679
rect 7987 -633 8187 -600
rect 7987 -679 8000 -633
rect 8174 -679 8187 -633
rect 7987 -692 8187 -679
rect 8291 -633 8491 -600
rect 8291 -679 8304 -633
rect 8478 -679 8491 -633
rect 8291 -692 8491 -679
rect 8595 -633 8795 -600
rect 8595 -679 8608 -633
rect 8782 -679 8795 -633
rect 8595 -692 8795 -679
rect 8899 -633 9099 -600
rect 8899 -679 8912 -633
rect 9086 -679 9099 -633
rect 8899 -692 9099 -679
rect 9203 -633 9403 -600
rect 9203 -679 9216 -633
rect 9390 -679 9403 -633
rect 9203 -692 9403 -679
rect 9783 -341 9863 -328
rect 9783 -387 9796 -341
rect 9850 -387 9863 -341
rect 9783 -420 9863 -387
rect 9783 -613 9863 -580
rect 9783 -659 9796 -613
rect 9850 -659 9863 -613
rect 9783 -672 9863 -659
rect 10643 -341 10723 -328
rect 10643 -387 10656 -341
rect 10710 -387 10723 -341
rect 10643 -420 10723 -387
rect 10643 -613 10723 -580
rect 10643 -659 10656 -613
rect 10710 -659 10723 -613
rect 10643 -672 10723 -659
rect 6329 -1277 6529 -1264
rect 6329 -1323 6342 -1277
rect 6516 -1323 6529 -1277
rect 6329 -1356 6529 -1323
rect 6633 -1277 6833 -1264
rect 6633 -1323 6646 -1277
rect 6820 -1323 6833 -1277
rect 6633 -1356 6833 -1323
rect 6937 -1277 7137 -1264
rect 6937 -1323 6950 -1277
rect 7124 -1323 7137 -1277
rect 6937 -1356 7137 -1323
rect 7241 -1277 7441 -1264
rect 7241 -1323 7254 -1277
rect 7428 -1323 7441 -1277
rect 7241 -1356 7441 -1323
rect 7545 -1277 7745 -1264
rect 7545 -1323 7558 -1277
rect 7732 -1323 7745 -1277
rect 7545 -1356 7745 -1323
rect 6329 -1789 6529 -1756
rect 6329 -1835 6342 -1789
rect 6516 -1835 6529 -1789
rect 6329 -1848 6529 -1835
rect 6633 -1789 6833 -1756
rect 6633 -1835 6646 -1789
rect 6820 -1835 6833 -1789
rect 6633 -1848 6833 -1835
rect 6937 -1789 7137 -1756
rect 6937 -1835 6950 -1789
rect 7124 -1835 7137 -1789
rect 6937 -1848 7137 -1835
rect 7241 -1789 7441 -1756
rect 7241 -1835 7254 -1789
rect 7428 -1835 7441 -1789
rect 7241 -1848 7441 -1835
rect 7545 -1789 7745 -1756
rect 7545 -1835 7558 -1789
rect 7732 -1835 7745 -1789
rect 7545 -1848 7745 -1835
rect 8125 -1277 8325 -1264
rect 8125 -1323 8138 -1277
rect 8312 -1323 8325 -1277
rect 8125 -1356 8325 -1323
rect 8429 -1277 8629 -1264
rect 8429 -1323 8442 -1277
rect 8616 -1323 8629 -1277
rect 8429 -1356 8629 -1323
rect 8733 -1277 8933 -1264
rect 8733 -1323 8746 -1277
rect 8920 -1323 8933 -1277
rect 8733 -1356 8933 -1323
rect 9037 -1277 9237 -1264
rect 9037 -1323 9050 -1277
rect 9224 -1323 9237 -1277
rect 9037 -1356 9237 -1323
rect 9341 -1277 9541 -1264
rect 9341 -1323 9354 -1277
rect 9528 -1323 9541 -1277
rect 9341 -1356 9541 -1323
rect 8125 -1789 8325 -1756
rect 8125 -1835 8138 -1789
rect 8312 -1835 8325 -1789
rect 8125 -1848 8325 -1835
rect 8429 -1789 8629 -1756
rect 8429 -1835 8442 -1789
rect 8616 -1835 8629 -1789
rect 8429 -1848 8629 -1835
rect 8733 -1789 8933 -1756
rect 8733 -1835 8746 -1789
rect 8920 -1835 8933 -1789
rect 8733 -1848 8933 -1835
rect 9037 -1789 9237 -1756
rect 9037 -1835 9050 -1789
rect 9224 -1835 9237 -1789
rect 9037 -1848 9237 -1835
rect 9341 -1789 9541 -1756
rect 9341 -1835 9354 -1789
rect 9528 -1835 9541 -1789
rect 9341 -1848 9541 -1835
rect 6163 -2762 6363 -2749
rect 6163 -2808 6176 -2762
rect 6350 -2808 6363 -2762
rect 6163 -2841 6363 -2808
rect 6467 -2762 6667 -2749
rect 6467 -2808 6480 -2762
rect 6654 -2808 6667 -2762
rect 6467 -2841 6667 -2808
rect 6771 -2762 6971 -2749
rect 6771 -2808 6784 -2762
rect 6958 -2808 6971 -2762
rect 6771 -2841 6971 -2808
rect 7075 -2762 7275 -2749
rect 7075 -2808 7088 -2762
rect 7262 -2808 7275 -2762
rect 7075 -2841 7275 -2808
rect 7379 -2762 7579 -2749
rect 7379 -2808 7392 -2762
rect 7566 -2808 7579 -2762
rect 7379 -2841 7579 -2808
rect 7683 -2762 7883 -2749
rect 7683 -2808 7696 -2762
rect 7870 -2808 7883 -2762
rect 7683 -2841 7883 -2808
rect 7987 -2762 8187 -2749
rect 7987 -2808 8000 -2762
rect 8174 -2808 8187 -2762
rect 7987 -2841 8187 -2808
rect 8291 -2762 8491 -2749
rect 8291 -2808 8304 -2762
rect 8478 -2808 8491 -2762
rect 8291 -2841 8491 -2808
rect 8595 -2762 8795 -2749
rect 8595 -2808 8608 -2762
rect 8782 -2808 8795 -2762
rect 8595 -2841 8795 -2808
rect 8899 -2762 9099 -2749
rect 8899 -2808 8912 -2762
rect 9086 -2808 9099 -2762
rect 8899 -2841 9099 -2808
rect 9203 -2762 9403 -2749
rect 9203 -2808 9216 -2762
rect 9390 -2808 9403 -2762
rect 9203 -2841 9403 -2808
rect 9507 -2762 9707 -2749
rect 9507 -2808 9520 -2762
rect 9694 -2808 9707 -2762
rect 9507 -2841 9707 -2808
rect 6163 -3174 6363 -3141
rect 6163 -3220 6176 -3174
rect 6350 -3220 6363 -3174
rect 6163 -3233 6363 -3220
rect 6467 -3174 6667 -3141
rect 6467 -3220 6480 -3174
rect 6654 -3220 6667 -3174
rect 6467 -3233 6667 -3220
rect 6771 -3174 6971 -3141
rect 6771 -3220 6784 -3174
rect 6958 -3220 6971 -3174
rect 6771 -3233 6971 -3220
rect 7075 -3174 7275 -3141
rect 7075 -3220 7088 -3174
rect 7262 -3220 7275 -3174
rect 7075 -3233 7275 -3220
rect 7379 -3174 7579 -3141
rect 7379 -3220 7392 -3174
rect 7566 -3220 7579 -3174
rect 7379 -3233 7579 -3220
rect 7683 -3174 7883 -3141
rect 7683 -3220 7696 -3174
rect 7870 -3220 7883 -3174
rect 7683 -3233 7883 -3220
rect 7987 -3174 8187 -3141
rect 7987 -3220 8000 -3174
rect 8174 -3220 8187 -3174
rect 7987 -3233 8187 -3220
rect 8291 -3174 8491 -3141
rect 8291 -3220 8304 -3174
rect 8478 -3220 8491 -3174
rect 8291 -3233 8491 -3220
rect 8595 -3174 8795 -3141
rect 8595 -3220 8608 -3174
rect 8782 -3220 8795 -3174
rect 8595 -3233 8795 -3220
rect 8899 -3174 9099 -3141
rect 8899 -3220 8912 -3174
rect 9086 -3220 9099 -3174
rect 8899 -3233 9099 -3220
rect 9203 -3174 9403 -3141
rect 9203 -3220 9216 -3174
rect 9390 -3220 9403 -3174
rect 9203 -3233 9403 -3220
rect 9507 -3174 9707 -3141
rect 9507 -3220 9520 -3174
rect 9694 -3220 9707 -3174
rect 9507 -3233 9707 -3220
rect 6825 -3235 6915 -3233
rect 6163 -3725 6363 -3712
rect 6163 -3771 6176 -3725
rect 6350 -3771 6363 -3725
rect 6163 -3804 6363 -3771
rect 6467 -3725 6667 -3712
rect 6467 -3771 6480 -3725
rect 6654 -3771 6667 -3725
rect 6467 -3804 6667 -3771
rect 6771 -3725 6971 -3712
rect 6771 -3771 6784 -3725
rect 6958 -3771 6971 -3725
rect 6771 -3804 6971 -3771
rect 7075 -3725 7275 -3712
rect 7075 -3771 7088 -3725
rect 7262 -3771 7275 -3725
rect 7075 -3804 7275 -3771
rect 7379 -3725 7579 -3712
rect 7379 -3771 7392 -3725
rect 7566 -3771 7579 -3725
rect 7379 -3804 7579 -3771
rect 7683 -3725 7883 -3712
rect 7683 -3771 7696 -3725
rect 7870 -3771 7883 -3725
rect 7683 -3804 7883 -3771
rect 7987 -3725 8187 -3712
rect 7987 -3771 8000 -3725
rect 8174 -3771 8187 -3725
rect 7987 -3804 8187 -3771
rect 8291 -3725 8491 -3712
rect 8291 -3771 8304 -3725
rect 8478 -3771 8491 -3725
rect 8291 -3804 8491 -3771
rect 8595 -3725 8795 -3712
rect 8595 -3771 8608 -3725
rect 8782 -3771 8795 -3725
rect 8595 -3804 8795 -3771
rect 8899 -3725 9099 -3712
rect 8899 -3771 8912 -3725
rect 9086 -3771 9099 -3725
rect 8899 -3804 9099 -3771
rect 9203 -3725 9403 -3712
rect 9203 -3771 9216 -3725
rect 9390 -3771 9403 -3725
rect 9203 -3804 9403 -3771
rect 9507 -3725 9707 -3712
rect 9507 -3771 9520 -3725
rect 9694 -3771 9707 -3725
rect 9507 -3804 9707 -3771
rect 6163 -4137 6363 -4104
rect 6163 -4183 6176 -4137
rect 6350 -4183 6363 -4137
rect 6163 -4196 6363 -4183
rect 6467 -4137 6667 -4104
rect 6467 -4183 6480 -4137
rect 6654 -4183 6667 -4137
rect 6467 -4196 6667 -4183
rect 6771 -4137 6971 -4104
rect 6771 -4183 6784 -4137
rect 6958 -4183 6971 -4137
rect 6771 -4196 6971 -4183
rect 7075 -4137 7275 -4104
rect 7075 -4183 7088 -4137
rect 7262 -4183 7275 -4137
rect 7075 -4196 7275 -4183
rect 7379 -4137 7579 -4104
rect 7379 -4183 7392 -4137
rect 7566 -4183 7579 -4137
rect 7379 -4196 7579 -4183
rect 7683 -4137 7883 -4104
rect 7683 -4183 7696 -4137
rect 7870 -4183 7883 -4137
rect 7683 -4196 7883 -4183
rect 7987 -4137 8187 -4104
rect 7987 -4183 8000 -4137
rect 8174 -4183 8187 -4137
rect 7987 -4196 8187 -4183
rect 8291 -4137 8491 -4104
rect 8291 -4183 8304 -4137
rect 8478 -4183 8491 -4137
rect 8291 -4196 8491 -4183
rect 8595 -4137 8795 -4104
rect 8595 -4183 8608 -4137
rect 8782 -4183 8795 -4137
rect 8595 -4196 8795 -4183
rect 8899 -4137 9099 -4104
rect 8899 -4183 8912 -4137
rect 9086 -4183 9099 -4137
rect 8899 -4196 9099 -4183
rect 9203 -4137 9403 -4104
rect 9203 -4183 9216 -4137
rect 9390 -4183 9403 -4137
rect 9203 -4196 9403 -4183
rect 9507 -4137 9707 -4104
rect 9507 -4183 9520 -4137
rect 9694 -4183 9707 -4137
rect 9507 -4196 9707 -4183
rect 7711 -4651 7791 -4638
rect 7711 -4697 7724 -4651
rect 7778 -4697 7791 -4651
rect 7711 -4730 7791 -4697
rect 7895 -4651 7975 -4638
rect 7895 -4697 7908 -4651
rect 7962 -4697 7975 -4651
rect 7895 -4730 7975 -4697
rect 8079 -4651 8159 -4638
rect 8079 -4697 8092 -4651
rect 8146 -4697 8159 -4651
rect 8079 -4730 8159 -4697
rect 7711 -4923 7791 -4890
rect 7711 -4969 7724 -4923
rect 7778 -4969 7791 -4923
rect 7711 -4982 7791 -4969
rect 7895 -4923 7975 -4890
rect 7895 -4969 7908 -4923
rect 7962 -4969 7975 -4923
rect 7895 -4982 7975 -4969
rect 8079 -4923 8159 -4890
rect 8079 -4969 8092 -4923
rect 8146 -4969 8159 -4923
rect 8079 -4982 8159 -4969
<< polycontact >>
rect 5822 2680 5868 2726
rect 5912 2530 5958 2576
rect 7678 2803 7732 2849
rect 7678 2491 7732 2537
rect 8138 2803 8192 2849
rect 8138 2491 8192 2537
rect 6708 1386 6762 1432
rect 7678 1983 7732 2029
rect 7678 1671 7732 1717
rect 8138 1983 8192 2029
rect 8138 1671 8192 1717
rect 9108 1386 9162 1432
rect 6708 1050 6762 1096
rect 9108 1050 9162 1096
rect 5160 -387 5214 -341
rect 5160 -659 5214 -613
rect 6020 -387 6074 -341
rect 6020 -659 6074 -613
rect 6480 -367 6654 -321
rect 6784 -367 6958 -321
rect 7088 -367 7262 -321
rect 7392 -367 7566 -321
rect 7696 -367 7870 -321
rect 8000 -367 8174 -321
rect 8304 -367 8478 -321
rect 8608 -367 8782 -321
rect 8912 -367 9086 -321
rect 9216 -367 9390 -321
rect 6480 -679 6654 -633
rect 6784 -679 6958 -633
rect 7088 -679 7262 -633
rect 7392 -679 7566 -633
rect 7696 -679 7870 -633
rect 8000 -679 8174 -633
rect 8304 -679 8478 -633
rect 8608 -679 8782 -633
rect 8912 -679 9086 -633
rect 9216 -679 9390 -633
rect 9796 -387 9850 -341
rect 9796 -659 9850 -613
rect 10656 -387 10710 -341
rect 10656 -659 10710 -613
rect 6342 -1323 6516 -1277
rect 6646 -1323 6820 -1277
rect 6950 -1323 7124 -1277
rect 7254 -1323 7428 -1277
rect 7558 -1323 7732 -1277
rect 6342 -1835 6516 -1789
rect 6646 -1835 6820 -1789
rect 6950 -1835 7124 -1789
rect 7254 -1835 7428 -1789
rect 7558 -1835 7732 -1789
rect 8138 -1323 8312 -1277
rect 8442 -1323 8616 -1277
rect 8746 -1323 8920 -1277
rect 9050 -1323 9224 -1277
rect 9354 -1323 9528 -1277
rect 8138 -1835 8312 -1789
rect 8442 -1835 8616 -1789
rect 8746 -1835 8920 -1789
rect 9050 -1835 9224 -1789
rect 9354 -1835 9528 -1789
rect 6176 -2808 6350 -2762
rect 6480 -2808 6654 -2762
rect 6784 -2808 6958 -2762
rect 7088 -2808 7262 -2762
rect 7392 -2808 7566 -2762
rect 7696 -2808 7870 -2762
rect 8000 -2808 8174 -2762
rect 8304 -2808 8478 -2762
rect 8608 -2808 8782 -2762
rect 8912 -2808 9086 -2762
rect 9216 -2808 9390 -2762
rect 9520 -2808 9694 -2762
rect 6176 -3220 6350 -3174
rect 6480 -3220 6654 -3174
rect 6784 -3220 6958 -3174
rect 7088 -3220 7262 -3174
rect 7392 -3220 7566 -3174
rect 7696 -3220 7870 -3174
rect 8000 -3220 8174 -3174
rect 8304 -3220 8478 -3174
rect 8608 -3220 8782 -3174
rect 8912 -3220 9086 -3174
rect 9216 -3220 9390 -3174
rect 9520 -3220 9694 -3174
rect 6176 -3771 6350 -3725
rect 6480 -3771 6654 -3725
rect 6784 -3771 6958 -3725
rect 7088 -3771 7262 -3725
rect 7392 -3771 7566 -3725
rect 7696 -3771 7870 -3725
rect 8000 -3771 8174 -3725
rect 8304 -3771 8478 -3725
rect 8608 -3771 8782 -3725
rect 8912 -3771 9086 -3725
rect 9216 -3771 9390 -3725
rect 9520 -3771 9694 -3725
rect 6176 -4183 6350 -4137
rect 6480 -4183 6654 -4137
rect 6784 -4183 6958 -4137
rect 7088 -4183 7262 -4137
rect 7392 -4183 7566 -4137
rect 7696 -4183 7870 -4137
rect 8000 -4183 8174 -4137
rect 8304 -4183 8478 -4137
rect 8608 -4183 8782 -4137
rect 8912 -4183 9086 -4137
rect 9216 -4183 9390 -4137
rect 9520 -4183 9694 -4137
rect 7724 -4697 7778 -4651
rect 7908 -4697 7962 -4651
rect 8092 -4697 8146 -4651
rect 7724 -4969 7778 -4923
rect 7908 -4969 7962 -4923
rect 8092 -4969 8146 -4923
<< metal1 >>
rect 3654 4000 11642 4380
rect 4011 1082 4089 4000
rect 5620 3333 5700 4000
rect 5065 3261 6205 3333
rect 5065 3215 5317 3261
rect 5363 3215 5557 3261
rect 5603 3215 5797 3261
rect 5843 3215 6037 3261
rect 6083 3215 6205 3261
rect 5065 3193 6205 3215
rect 5185 3070 5235 3193
rect 5185 2836 5187 3070
rect 5233 2836 5235 3070
rect 5355 3095 5405 3123
rect 5355 2861 5357 3095
rect 5403 2861 5405 3095
rect 5355 2843 5405 2861
rect 5525 3070 5575 3193
rect 5185 2783 5235 2836
rect 5325 2839 5425 2843
rect 5325 2787 5349 2839
rect 5401 2787 5425 2839
rect 5325 2783 5425 2787
rect 5525 2836 5527 3070
rect 5573 2836 5575 3070
rect 5525 2783 5575 2836
rect 5695 3095 5745 3123
rect 5695 2861 5697 3095
rect 5743 2861 5745 3095
rect 5355 2733 5405 2783
rect 5695 2733 5745 2861
rect 5865 3070 5915 3193
rect 5865 2836 5867 3070
rect 5913 2836 5915 3070
rect 5865 2783 5915 2836
rect 6035 3070 6085 3123
rect 6035 2836 6037 3070
rect 6083 2836 6085 3070
rect 6035 2733 6085 2836
rect 5355 2673 5745 2733
rect 5795 2726 6085 2733
rect 5795 2680 5822 2726
rect 5868 2680 6085 2726
rect 5795 2673 6085 2680
rect 5355 2553 5405 2673
rect 5695 2553 5745 2673
rect 5355 2493 5745 2553
rect 5885 2579 5985 2583
rect 5885 2527 5909 2579
rect 5961 2527 5985 2579
rect 5885 2523 5985 2527
rect 5185 2381 5235 2443
rect 5185 2335 5187 2381
rect 5233 2335 5235 2381
rect 5185 2203 5235 2335
rect 5355 2381 5405 2493
rect 5355 2335 5357 2381
rect 5403 2335 5405 2381
rect 5355 2273 5405 2335
rect 5525 2381 5575 2443
rect 5525 2335 5527 2381
rect 5573 2335 5575 2381
rect 5525 2203 5575 2335
rect 5695 2381 5745 2493
rect 5695 2335 5697 2381
rect 5743 2335 5745 2381
rect 5695 2273 5745 2335
rect 5865 2381 5915 2443
rect 5865 2335 5867 2381
rect 5913 2335 5915 2381
rect 5865 2203 5915 2335
rect 6035 2381 6085 2673
rect 6700 2390 6780 4000
rect 7880 3060 7960 4000
rect 7452 2980 8418 3060
rect 7452 2840 7498 2980
rect 7667 2849 7743 2882
rect 7667 2803 7678 2849
rect 7732 2803 7743 2849
rect 7912 2840 7958 2851
rect 7590 2757 7636 2768
rect 7498 2583 7590 2757
rect 7774 2757 7820 2768
rect 7757 2698 7774 2708
rect 7820 2698 7837 2708
rect 7757 2642 7769 2698
rect 7825 2642 7837 2698
rect 7757 2632 7774 2642
rect 7590 2572 7636 2583
rect 7820 2632 7837 2642
rect 7774 2572 7820 2583
rect 7452 2489 7498 2500
rect 7667 2491 7678 2537
rect 7732 2491 7743 2537
rect 8127 2849 8203 2882
rect 8127 2803 8138 2849
rect 8192 2803 8203 2849
rect 8372 2840 8418 2980
rect 8050 2757 8096 2768
rect 8033 2698 8050 2708
rect 8234 2757 8280 2768
rect 8096 2698 8113 2708
rect 8033 2642 8045 2698
rect 8101 2642 8113 2698
rect 8033 2632 8050 2642
rect 8096 2632 8113 2642
rect 8050 2572 8096 2583
rect 8280 2583 8372 2757
rect 8234 2572 8280 2583
rect 6574 2389 6585 2390
rect 6035 2335 6037 2381
rect 6083 2335 6085 2381
rect 6503 2344 6585 2389
rect 6885 2389 6896 2390
rect 6885 2344 6953 2389
rect 6503 2337 6953 2344
rect 6035 2273 6085 2335
rect 6511 2329 6953 2337
rect 6611 2252 6671 2329
rect 7677 2304 7733 2491
rect 7912 2489 7958 2500
rect 8127 2491 8138 2537
rect 8192 2491 8203 2537
rect 7895 2440 7965 2442
rect 8137 2440 8193 2491
rect 8372 2489 8418 2500
rect 7895 2384 7907 2440
rect 7963 2384 8193 2440
rect 9100 2390 9180 4000
rect 8974 2389 8985 2390
rect 7895 2382 7965 2384
rect 8917 2344 8985 2389
rect 9285 2389 9296 2390
rect 9285 2344 9367 2389
rect 8917 2337 9367 2344
rect 8917 2329 9359 2337
rect 7677 2302 7975 2304
rect 5065 2181 6205 2203
rect 5065 2135 5317 2181
rect 5363 2135 5557 2181
rect 5603 2135 5797 2181
rect 5843 2135 6037 2181
rect 6083 2135 6205 2181
rect 5065 2063 6205 2135
rect 6611 2105 6620 2252
rect 6666 2105 6671 2252
rect 6804 2261 6850 2263
rect 6804 2252 6887 2261
rect 6620 1467 6666 1478
rect 6850 1478 6887 2252
rect 7677 2246 7907 2302
rect 7963 2246 7975 2302
rect 9020 2261 9066 2263
rect 7677 2244 7975 2246
rect 8983 2252 9066 2261
rect 6804 1467 6887 1478
rect 6697 1405 6708 1432
rect 6695 1386 6708 1405
rect 6762 1405 6773 1432
rect 6762 1386 6775 1405
rect 5565 1279 5659 1291
rect 6695 1279 6775 1386
rect 5565 1203 5577 1279
rect 5657 1203 6775 1279
rect 5565 1201 5659 1203
rect 6695 1096 6775 1203
rect 6695 1085 6708 1096
rect 4010 881 4090 1082
rect 6697 1050 6708 1085
rect 6762 1085 6775 1096
rect 6823 1349 6887 1467
rect 7452 2020 7498 2031
rect 7667 2029 7743 2062
rect 7667 1983 7678 2029
rect 7732 1983 7743 2029
rect 7912 2020 7958 2031
rect 7590 1937 7636 1948
rect 7498 1763 7590 1937
rect 7774 1937 7820 1948
rect 7757 1878 7774 1888
rect 7820 1878 7837 1888
rect 7757 1822 7769 1878
rect 7825 1822 7837 1878
rect 7757 1812 7774 1822
rect 7590 1752 7636 1763
rect 7820 1812 7837 1822
rect 7774 1752 7820 1763
rect 7667 1712 7678 1717
rect 7452 1540 7498 1680
rect 7665 1702 7678 1712
rect 7732 1712 7743 1717
rect 7732 1702 7745 1712
rect 7665 1646 7677 1702
rect 7733 1646 7745 1702
rect 8127 2029 8203 2062
rect 8127 1983 8138 2029
rect 8192 1983 8203 2029
rect 8372 2020 8418 2031
rect 8050 1937 8096 1948
rect 8033 1878 8050 1888
rect 8234 1937 8280 1948
rect 8096 1878 8113 1888
rect 8033 1822 8045 1878
rect 8101 1822 8113 1878
rect 8033 1812 8050 1822
rect 8096 1812 8113 1822
rect 8050 1752 8096 1763
rect 8280 1763 8372 1937
rect 8234 1752 8280 1763
rect 8127 1712 8138 1717
rect 7912 1669 7958 1680
rect 8125 1702 8138 1712
rect 8192 1712 8203 1717
rect 8192 1702 8205 1712
rect 7665 1636 7745 1646
rect 8125 1646 8137 1702
rect 8193 1646 8205 1702
rect 8125 1636 8205 1646
rect 8372 1540 8418 1680
rect 7452 1460 8418 1540
rect 8983 1478 9020 2252
rect 9199 2252 9259 2329
rect 9199 2105 9204 2252
rect 8983 1467 9066 1478
rect 9250 2105 9259 2252
rect 9204 1467 9250 1478
rect 6823 1279 6891 1349
rect 7675 1279 7747 1281
rect 6823 1203 7677 1279
rect 7733 1203 7747 1279
rect 6762 1050 6773 1085
rect 6823 1015 6891 1203
rect 7675 1191 7747 1203
rect 6620 1004 6666 1015
rect 3993 864 4106 881
rect 3993 786 4010 864
rect 4090 786 4106 864
rect 3993 775 4106 786
rect 6619 630 6620 713
rect 6804 1004 6891 1015
rect 6666 630 6667 713
rect 6619 546 6667 630
rect 6850 633 6891 1004
rect 6804 619 6850 630
rect 4869 543 7471 546
rect 7891 543 7957 1460
rect 8983 1349 9047 1467
rect 9097 1405 9108 1432
rect 8123 1279 8195 1281
rect 8979 1279 9047 1349
rect 8123 1203 8137 1279
rect 8193 1203 9047 1279
rect 8123 1191 8195 1203
rect 8979 1015 9047 1203
rect 9095 1386 9108 1405
rect 9162 1405 9173 1432
rect 9162 1386 9175 1405
rect 9095 1279 9175 1386
rect 10201 1279 10305 1291
rect 9095 1203 10213 1279
rect 10293 1203 10305 1279
rect 9095 1096 9175 1203
rect 10201 1201 10305 1203
rect 10421 1100 10499 4000
rect 9095 1085 9108 1096
rect 9097 1050 9108 1085
rect 9162 1085 9175 1096
rect 9162 1050 9173 1085
rect 8979 1004 9066 1015
rect 8979 633 9020 1004
rect 9204 1004 9250 1015
rect 9020 619 9066 630
rect 9203 630 9204 713
rect 10420 930 10500 1100
rect 10400 750 10520 930
rect 9250 630 9251 713
rect 10400 690 10420 750
rect 10500 690 10520 750
rect 9203 546 9251 630
rect 11305 552 11463 567
rect 11305 546 11332 552
rect 9182 545 11332 546
rect 8965 543 11332 545
rect 4396 538 11332 543
rect 4396 492 6585 538
rect 6885 492 8985 538
rect 9285 492 11332 538
rect 4396 483 11332 492
rect 4396 454 4599 483
rect 4869 481 11332 483
rect 4396 365 4454 454
rect 4545 365 4599 454
rect 11305 445 11332 481
rect 11441 445 11463 552
rect 11305 434 11463 445
rect 4396 336 4599 365
rect 4705 335 4809 349
rect 11061 335 11165 347
rect 4705 259 4717 335
rect 4797 259 11073 335
rect 11153 259 11165 335
rect 4705 249 4809 259
rect 4934 -350 4980 -339
rect 5149 -341 5225 259
rect 5149 -387 5160 -341
rect 5214 -387 5225 -341
rect 5394 -350 5440 -339
rect 5072 -431 5118 -422
rect 5256 -431 5302 -422
rect 4980 -433 5135 -431
rect 4980 -567 5067 -433
rect 5123 -567 5135 -433
rect 4980 -569 5135 -567
rect 5239 -433 5319 -431
rect 5239 -567 5251 -433
rect 5307 -567 5319 -433
rect 5239 -569 5319 -567
rect 5377 -433 5394 -431
rect 5794 -350 5840 -339
rect 5440 -433 5457 -431
rect 5377 -567 5389 -433
rect 5445 -567 5457 -433
rect 5377 -569 5394 -567
rect 5072 -578 5118 -569
rect 5256 -578 5302 -569
rect 4934 -661 4980 -650
rect 5149 -659 5160 -613
rect 5214 -659 5225 -613
rect 5149 -689 5225 -659
rect 5440 -569 5457 -567
rect 5394 -661 5440 -650
rect 6009 -341 6085 259
rect 6009 -387 6020 -341
rect 6074 -387 6085 -341
rect 6254 -330 6300 -319
rect 6773 -321 7273 -265
rect 5932 -431 5978 -422
rect 6116 -431 6162 -422
rect 5840 -433 5995 -431
rect 5840 -567 5927 -433
rect 5983 -567 5995 -433
rect 5840 -569 5995 -567
rect 6099 -433 6179 -431
rect 6099 -567 6111 -433
rect 6167 -567 6179 -433
rect 6099 -569 6179 -567
rect 6237 -433 6254 -431
rect 6469 -367 6480 -321
rect 6654 -367 6665 -321
rect 6773 -367 6784 -321
rect 6958 -367 6969 -321
rect 7077 -367 7088 -321
rect 7262 -367 7273 -321
rect 7381 -321 7881 -265
rect 7381 -367 7392 -321
rect 7566 -367 7577 -321
rect 7685 -367 7696 -321
rect 7870 -367 7881 -321
rect 7989 -321 8489 -265
rect 7989 -367 8000 -321
rect 8174 -367 8185 -321
rect 8293 -367 8304 -321
rect 8478 -367 8489 -321
rect 8597 -321 9097 -265
rect 8597 -367 8608 -321
rect 8782 -367 8793 -321
rect 8901 -367 8912 -321
rect 9086 -367 9097 -321
rect 9205 -367 9216 -321
rect 9390 -367 9401 -321
rect 9570 -330 9616 -319
rect 6392 -413 6438 -402
rect 6300 -433 6317 -431
rect 6237 -567 6249 -433
rect 6305 -567 6317 -433
rect 6237 -569 6254 -567
rect 5932 -578 5978 -569
rect 6116 -578 6162 -569
rect 5794 -661 5840 -650
rect 6009 -659 6020 -613
rect 6074 -659 6085 -613
rect 6009 -689 6085 -659
rect 6300 -569 6317 -567
rect 6696 -413 6742 -402
rect 6679 -420 6696 -418
rect 7000 -413 7046 -402
rect 6742 -420 6759 -418
rect 6679 -564 6691 -420
rect 6747 -564 6759 -420
rect 6679 -566 6696 -564
rect 6392 -598 6438 -587
rect 6742 -566 6759 -564
rect 6983 -521 7000 -511
rect 7304 -413 7350 -402
rect 7287 -420 7304 -418
rect 7608 -413 7654 -402
rect 7350 -420 7367 -418
rect 7046 -521 7063 -511
rect 6983 -577 6995 -521
rect 7051 -577 7063 -521
rect 7287 -564 7299 -420
rect 7355 -564 7367 -420
rect 7287 -566 7304 -564
rect 6983 -587 7000 -577
rect 7046 -587 7063 -577
rect 7350 -566 7367 -564
rect 7591 -521 7608 -511
rect 7912 -413 7958 -402
rect 7895 -420 7912 -418
rect 8216 -413 8262 -402
rect 7958 -420 7975 -418
rect 7654 -521 7671 -511
rect 7591 -577 7603 -521
rect 7659 -577 7671 -521
rect 7895 -564 7907 -420
rect 7963 -564 7975 -420
rect 7895 -566 7912 -564
rect 7591 -587 7608 -577
rect 7654 -587 7671 -577
rect 7958 -566 7975 -564
rect 8199 -521 8216 -511
rect 8520 -413 8566 -402
rect 8503 -420 8520 -418
rect 8824 -413 8870 -402
rect 8566 -420 8583 -418
rect 8262 -521 8279 -511
rect 8199 -577 8211 -521
rect 8267 -577 8279 -521
rect 8503 -564 8515 -420
rect 8571 -564 8583 -420
rect 8503 -566 8520 -564
rect 8199 -587 8216 -577
rect 8262 -587 8279 -577
rect 8566 -566 8583 -564
rect 8807 -521 8824 -511
rect 9128 -413 9174 -402
rect 9111 -420 9128 -418
rect 9432 -413 9478 -402
rect 9174 -420 9191 -418
rect 8870 -521 8887 -511
rect 8807 -577 8819 -521
rect 8875 -577 8887 -521
rect 9111 -564 9123 -420
rect 9179 -564 9191 -420
rect 9111 -566 9128 -564
rect 8807 -587 8824 -577
rect 8870 -587 8887 -577
rect 9174 -566 9191 -564
rect 6696 -598 6742 -587
rect 7000 -598 7046 -587
rect 7304 -598 7350 -587
rect 7608 -598 7654 -587
rect 7912 -598 7958 -587
rect 8216 -598 8262 -587
rect 8520 -598 8566 -587
rect 8824 -598 8870 -587
rect 9128 -598 9174 -587
rect 9553 -433 9570 -431
rect 9785 -341 9861 259
rect 9785 -387 9796 -341
rect 9850 -387 9861 -341
rect 10030 -350 10076 -339
rect 9708 -431 9754 -422
rect 9892 -431 9938 -422
rect 9616 -433 9633 -431
rect 9553 -567 9565 -433
rect 9621 -567 9633 -433
rect 9553 -569 9570 -567
rect 9432 -598 9478 -587
rect 7786 -628 7866 -618
rect 7786 -633 7798 -628
rect 7854 -633 7866 -628
rect 8004 -628 8084 -618
rect 8004 -633 8016 -628
rect 8072 -633 8084 -628
rect 6254 -681 6300 -670
rect 6469 -679 6480 -633
rect 6654 -679 6665 -633
rect 6773 -679 6784 -633
rect 6958 -644 6969 -633
rect 7077 -644 7088 -633
rect 6958 -679 7088 -644
rect 7262 -679 7273 -633
rect 7381 -679 7392 -633
rect 7566 -679 7577 -633
rect 7685 -679 7696 -633
rect 7870 -679 7881 -633
rect 7989 -679 8000 -633
rect 8174 -679 8185 -633
rect 8293 -679 8304 -633
rect 8478 -679 8489 -633
rect 8597 -679 8608 -633
rect 8782 -644 8793 -633
rect 8901 -644 8912 -633
rect 8782 -679 8912 -644
rect 9086 -679 9097 -633
rect 9205 -679 9216 -633
rect 9390 -679 9401 -633
rect 9616 -569 9633 -567
rect 9691 -433 9771 -431
rect 9691 -567 9703 -433
rect 9759 -567 9771 -433
rect 9691 -569 9771 -567
rect 9875 -433 10030 -431
rect 9875 -567 9887 -433
rect 9943 -567 10030 -433
rect 9875 -569 10030 -567
rect 9708 -578 9754 -569
rect 9892 -578 9938 -569
rect 6833 -690 7273 -679
rect 7786 -684 7798 -679
rect 7854 -684 7866 -679
rect 5565 -936 5669 -924
rect 6087 -936 6191 -926
rect 6833 -936 6937 -690
rect 7786 -694 7866 -684
rect 8004 -684 8016 -679
rect 8072 -684 8084 -679
rect 8004 -694 8084 -684
rect 8597 -690 9037 -679
rect 9570 -681 9616 -670
rect 9785 -659 9796 -613
rect 9850 -659 9861 -613
rect 9785 -689 9861 -659
rect 10430 -350 10476 -339
rect 10413 -433 10430 -431
rect 10645 -341 10721 259
rect 11061 247 11165 259
rect 10645 -387 10656 -341
rect 10710 -387 10721 -341
rect 10890 -350 10936 -339
rect 10568 -431 10614 -422
rect 10752 -431 10798 -422
rect 10476 -433 10493 -431
rect 10413 -567 10425 -433
rect 10481 -567 10493 -433
rect 10413 -569 10430 -567
rect 10030 -661 10076 -650
rect 10476 -569 10493 -567
rect 10551 -433 10631 -431
rect 10551 -567 10563 -433
rect 10619 -567 10631 -433
rect 10551 -569 10631 -567
rect 10735 -433 10890 -431
rect 10735 -567 10747 -433
rect 10803 -567 10890 -433
rect 10735 -569 10890 -567
rect 10568 -578 10614 -569
rect 10752 -578 10798 -569
rect 10430 -661 10476 -650
rect 10645 -659 10656 -613
rect 10710 -659 10721 -613
rect 10645 -689 10721 -659
rect 10890 -661 10936 -650
rect 7441 -936 7681 -928
rect 5565 -1020 5577 -936
rect 5657 -1020 6099 -936
rect 6179 -938 7681 -936
rect 6179 -1018 6845 -938
rect 6925 -1018 7453 -938
rect 7533 -1018 7591 -938
rect 7671 -1018 7681 -938
rect 6179 -1020 7681 -1018
rect 5565 -1030 5669 -1020
rect 6087 -1030 6191 -1020
rect 6833 -1032 6937 -1020
rect 7441 -1032 7681 -1020
rect 8187 -936 8429 -928
rect 8933 -936 9037 -690
rect 9679 -936 9783 -926
rect 10201 -936 10305 -926
rect 8187 -938 9691 -936
rect 8187 -1018 8199 -938
rect 8279 -1018 8337 -938
rect 8417 -1018 8945 -938
rect 9025 -1018 9691 -938
rect 8187 -1020 9691 -1018
rect 9771 -1020 10213 -936
rect 10293 -1020 10305 -936
rect 8187 -1032 8429 -1020
rect 8933 -1031 9037 -1020
rect 9679 -1030 9783 -1020
rect 10201 -1030 10305 -1020
rect 6635 -1232 7439 -1217
rect 6116 -1286 6162 -1275
rect 6635 -1277 7254 -1232
rect 7334 -1277 7439 -1232
rect 8431 -1232 9235 -1217
rect 6099 -1682 6116 -1672
rect 6331 -1323 6342 -1277
rect 6516 -1323 6527 -1277
rect 6635 -1323 6646 -1277
rect 6820 -1323 6831 -1277
rect 6939 -1323 6950 -1277
rect 7124 -1323 7135 -1277
rect 7243 -1323 7254 -1277
rect 7428 -1323 7439 -1277
rect 7547 -1323 7558 -1277
rect 7732 -1323 7743 -1277
rect 7912 -1286 7958 -1275
rect 8431 -1277 8536 -1232
rect 8616 -1277 9235 -1232
rect 6254 -1369 6300 -1358
rect 6162 -1682 6179 -1672
rect 6099 -1826 6111 -1682
rect 6167 -1826 6179 -1682
rect 6558 -1369 6604 -1358
rect 6541 -1592 6558 -1590
rect 6862 -1369 6908 -1358
rect 6845 -1376 6862 -1374
rect 7166 -1369 7212 -1358
rect 6908 -1376 6925 -1374
rect 6845 -1520 6857 -1376
rect 6913 -1520 6925 -1376
rect 6845 -1522 6862 -1520
rect 6604 -1592 6621 -1590
rect 6541 -1736 6553 -1592
rect 6609 -1736 6621 -1592
rect 6541 -1738 6558 -1736
rect 6254 -1754 6300 -1743
rect 6604 -1738 6621 -1736
rect 6558 -1754 6604 -1743
rect 6908 -1522 6925 -1520
rect 7149 -1592 7166 -1590
rect 7470 -1369 7516 -1358
rect 7453 -1376 7470 -1374
rect 7774 -1369 7820 -1358
rect 7516 -1376 7533 -1374
rect 7453 -1520 7465 -1376
rect 7521 -1520 7533 -1376
rect 7453 -1522 7470 -1520
rect 7212 -1592 7229 -1590
rect 7149 -1736 7161 -1592
rect 7217 -1736 7229 -1592
rect 7149 -1738 7166 -1736
rect 6862 -1754 6908 -1743
rect 7212 -1738 7229 -1736
rect 7166 -1754 7212 -1743
rect 7516 -1522 7533 -1520
rect 7470 -1754 7516 -1743
rect 7774 -1754 7820 -1743
rect 6099 -1837 6179 -1826
rect 6331 -1835 6342 -1789
rect 6516 -1835 6527 -1789
rect 6635 -1835 6646 -1789
rect 6820 -1835 6831 -1789
rect 6939 -1835 6950 -1789
rect 7124 -1835 7135 -1789
rect 7243 -1835 7254 -1789
rect 7428 -1835 7439 -1789
rect 7547 -1835 7558 -1789
rect 7732 -1835 7743 -1789
rect 8127 -1323 8138 -1277
rect 8312 -1323 8323 -1277
rect 8431 -1323 8442 -1277
rect 8616 -1323 8627 -1277
rect 8735 -1323 8746 -1277
rect 8920 -1323 8931 -1277
rect 9039 -1323 9050 -1277
rect 9224 -1323 9235 -1277
rect 9343 -1323 9354 -1277
rect 9528 -1323 9539 -1277
rect 9708 -1286 9754 -1275
rect 8050 -1369 8096 -1358
rect 8354 -1369 8400 -1358
rect 8337 -1376 8354 -1374
rect 8658 -1369 8704 -1358
rect 8400 -1376 8417 -1374
rect 8337 -1520 8349 -1376
rect 8405 -1520 8417 -1376
rect 8337 -1522 8354 -1520
rect 8050 -1754 8096 -1743
rect 8400 -1522 8417 -1520
rect 8641 -1592 8658 -1590
rect 8962 -1369 9008 -1358
rect 8945 -1376 8962 -1374
rect 9266 -1369 9312 -1358
rect 9008 -1376 9025 -1374
rect 8945 -1520 8957 -1376
rect 9013 -1520 9025 -1376
rect 8945 -1522 8962 -1520
rect 8704 -1592 8721 -1590
rect 8641 -1736 8653 -1592
rect 8709 -1736 8721 -1592
rect 8641 -1738 8658 -1736
rect 8354 -1754 8400 -1743
rect 8704 -1738 8721 -1736
rect 8658 -1754 8704 -1743
rect 9008 -1522 9025 -1520
rect 9249 -1592 9266 -1590
rect 9570 -1369 9616 -1358
rect 9312 -1592 9329 -1590
rect 9249 -1736 9261 -1592
rect 9317 -1736 9329 -1592
rect 9249 -1738 9266 -1736
rect 8962 -1754 9008 -1743
rect 9312 -1738 9329 -1736
rect 9266 -1754 9312 -1743
rect 9570 -1754 9616 -1743
rect 9691 -1682 9708 -1672
rect 9754 -1682 9771 -1672
rect 7912 -1837 7958 -1826
rect 8127 -1835 8138 -1789
rect 8312 -1835 8323 -1789
rect 8431 -1835 8442 -1789
rect 8616 -1835 8627 -1789
rect 8735 -1835 8746 -1789
rect 8920 -1835 8931 -1789
rect 9039 -1835 9050 -1789
rect 9224 -1835 9235 -1789
rect 9343 -1835 9354 -1789
rect 9528 -1835 9539 -1789
rect 9691 -1826 9703 -1682
rect 9759 -1826 9771 -1682
rect 9691 -1837 9771 -1826
rect 5227 -2102 5331 -2092
rect 6363 -2102 6467 -2090
rect 6529 -2102 6633 -2090
rect 7137 -2102 7241 -2090
rect 5227 -2182 5239 -2102
rect 5319 -2182 6375 -2102
rect 6455 -2182 6541 -2102
rect 6621 -2182 7149 -2102
rect 7229 -2182 7241 -2102
rect 5227 -2192 5331 -2182
rect 6363 -2194 6467 -2182
rect 6529 -2194 6633 -2182
rect 7137 -2194 7241 -2182
rect 8629 -2102 8733 -2090
rect 9237 -2102 9341 -2090
rect 9403 -2102 9507 -2090
rect 10539 -2102 10643 -2092
rect 8629 -2182 8641 -2102
rect 8721 -2182 9249 -2102
rect 9329 -2182 9415 -2102
rect 9495 -2182 10551 -2102
rect 10631 -2182 10643 -2102
rect 8629 -2194 8733 -2182
rect 9237 -2194 9341 -2182
rect 9403 -2194 9507 -2182
rect 10539 -2192 10643 -2182
rect 5781 -2500 5903 -2489
rect 5781 -3000 5792 -2500
rect 5892 -3000 5903 -2500
rect 9967 -2500 10089 -2489
rect 6165 -2808 6176 -2762
rect 6350 -2808 6361 -2762
rect 6469 -2808 6480 -2762
rect 6654 -2808 6665 -2762
rect 6773 -2808 6784 -2762
rect 6958 -2808 6969 -2762
rect 7077 -2808 7088 -2762
rect 7262 -2808 7273 -2762
rect 7381 -2808 7392 -2762
rect 7566 -2808 7577 -2762
rect 7685 -2808 7696 -2762
rect 7870 -2808 7881 -2762
rect 7989 -2808 8000 -2762
rect 8174 -2808 8185 -2762
rect 8293 -2808 8304 -2762
rect 8478 -2808 8489 -2762
rect 8597 -2808 8608 -2762
rect 8782 -2808 8793 -2762
rect 8901 -2808 8912 -2762
rect 9086 -2808 9097 -2762
rect 9205 -2808 9216 -2762
rect 9390 -2808 9401 -2762
rect 9509 -2808 9520 -2762
rect 9694 -2808 9705 -2762
rect 5781 -3011 5903 -3000
rect 6088 -2854 6134 -2843
rect 6392 -2854 6438 -2843
rect 6375 -2910 6392 -2900
rect 6696 -2854 6742 -2843
rect 6438 -2910 6455 -2900
rect 6375 -3071 6387 -2910
rect 6443 -3071 6455 -2910
rect 6375 -3081 6392 -3071
rect 6088 -3139 6134 -3128
rect 6438 -3081 6455 -3071
rect 6679 -2958 6696 -2948
rect 7000 -2854 7046 -2843
rect 6983 -2874 7000 -2864
rect 7304 -2854 7350 -2843
rect 7046 -2874 7063 -2864
rect 6742 -2958 6759 -2948
rect 6392 -3139 6438 -3128
rect 6679 -3119 6691 -2958
rect 6747 -3119 6759 -2958
rect 6983 -3091 6995 -2874
rect 7051 -3091 7063 -2874
rect 6983 -3099 7000 -3091
rect 6679 -3128 6696 -3119
rect 6742 -3128 6759 -3119
rect 6679 -3129 6759 -3128
rect 7046 -3099 7063 -3091
rect 7287 -2958 7304 -2948
rect 7608 -2854 7654 -2843
rect 7591 -2874 7608 -2864
rect 7912 -2854 7958 -2843
rect 7654 -2874 7671 -2864
rect 7591 -2930 7603 -2874
rect 7659 -2930 7671 -2874
rect 7591 -2940 7608 -2930
rect 7350 -2958 7367 -2948
rect 6696 -3139 6742 -3129
rect 7000 -3139 7046 -3128
rect 7287 -3119 7299 -2958
rect 7355 -3119 7367 -2958
rect 7287 -3128 7304 -3119
rect 7350 -3128 7367 -3119
rect 7287 -3129 7367 -3128
rect 7654 -2940 7671 -2930
rect 7304 -3139 7350 -3129
rect 7608 -3139 7654 -3128
rect 7895 -2958 7912 -2948
rect 8216 -2854 8262 -2843
rect 8199 -2874 8216 -2864
rect 8520 -2854 8566 -2843
rect 8262 -2874 8279 -2864
rect 8199 -2930 8211 -2874
rect 8267 -2930 8279 -2874
rect 8199 -2940 8216 -2930
rect 7958 -2958 7975 -2948
rect 7895 -3119 7907 -2958
rect 7963 -3119 7975 -2958
rect 7895 -3128 7912 -3119
rect 7958 -3128 7975 -3119
rect 7895 -3129 7975 -3128
rect 8262 -2940 8279 -2930
rect 7912 -3139 7958 -3129
rect 8216 -3139 8262 -3128
rect 8503 -2958 8520 -2948
rect 8824 -2854 8870 -2843
rect 8807 -2874 8824 -2864
rect 9128 -2854 9174 -2843
rect 8870 -2874 8887 -2864
rect 8566 -2958 8583 -2948
rect 8503 -3119 8515 -2958
rect 8571 -3119 8583 -2958
rect 8503 -3128 8520 -3119
rect 8566 -3128 8583 -3119
rect 8503 -3129 8583 -3128
rect 8807 -3119 8819 -2874
rect 8875 -3119 8887 -2874
rect 8807 -3128 8824 -3119
rect 8870 -3128 8887 -3119
rect 8807 -3129 8887 -3128
rect 9111 -2958 9128 -2948
rect 9432 -2854 9478 -2843
rect 9415 -2910 9432 -2900
rect 9736 -2854 9782 -2843
rect 9478 -2910 9495 -2900
rect 9174 -2958 9191 -2948
rect 9111 -3119 9123 -2958
rect 9179 -3119 9191 -2958
rect 9415 -3071 9427 -2910
rect 9483 -3071 9495 -2910
rect 9415 -3081 9432 -3071
rect 9111 -3128 9128 -3119
rect 9174 -3128 9191 -3119
rect 9111 -3129 9191 -3128
rect 9478 -3081 9495 -3071
rect 8520 -3139 8566 -3129
rect 8824 -3139 8870 -3129
rect 9128 -3139 9174 -3129
rect 9432 -3139 9478 -3128
rect 9967 -3000 9978 -2500
rect 10078 -3000 10089 -2500
rect 9967 -3011 10089 -3000
rect 9736 -3139 9782 -3128
rect 6820 -3174 6835 -3165
rect 6905 -3174 6920 -3165
rect 7125 -3174 7140 -3165
rect 7210 -3174 7225 -3165
rect 8035 -3174 8050 -3165
rect 8120 -3174 8135 -3165
rect 8340 -3174 8355 -3165
rect 8425 -3174 8440 -3165
rect 9255 -3174 9270 -3165
rect 9340 -3174 9355 -3165
rect 6165 -3220 6176 -3174
rect 6350 -3220 6361 -3174
rect 6469 -3220 6480 -3174
rect 6654 -3220 6665 -3174
rect 6773 -3220 6784 -3174
rect 6958 -3220 6969 -3174
rect 7077 -3220 7088 -3174
rect 7262 -3220 7273 -3174
rect 7381 -3220 7392 -3174
rect 7566 -3220 7577 -3174
rect 7685 -3220 7696 -3174
rect 7870 -3220 7881 -3174
rect 7989 -3220 8000 -3174
rect 8174 -3220 8185 -3174
rect 8293 -3220 8304 -3174
rect 8478 -3220 8489 -3174
rect 8597 -3220 8608 -3174
rect 8782 -3220 8793 -3174
rect 8901 -3220 8912 -3174
rect 9086 -3220 9097 -3174
rect 9205 -3220 9216 -3174
rect 9390 -3220 9401 -3174
rect 9509 -3220 9520 -3174
rect 9694 -3220 9705 -3174
rect 6470 -3275 6665 -3220
rect 6775 -3225 6835 -3220
rect 6905 -3225 6960 -3220
rect 7125 -3225 7140 -3220
rect 7210 -3225 7225 -3220
rect 7380 -3275 7575 -3220
rect 7685 -3275 7880 -3220
rect 8035 -3225 8050 -3220
rect 8120 -3225 8135 -3220
rect 8340 -3225 8355 -3220
rect 8425 -3225 8440 -3220
rect 8600 -3275 8795 -3220
rect 8900 -3275 9095 -3220
rect 9255 -3225 9270 -3220
rect 9340 -3225 9355 -3220
rect 3581 -3290 10065 -3275
rect 3581 -3323 9585 -3290
rect 3581 -3350 6842 -3323
rect 6830 -3379 6842 -3350
rect 6898 -3350 8057 -3323
rect 6898 -3379 6910 -3350
rect 6830 -3389 6910 -3379
rect 8045 -3379 8057 -3350
rect 8113 -3350 9585 -3323
rect 9645 -3350 10065 -3290
rect 8113 -3379 8125 -3350
rect 8045 -3389 8125 -3379
rect 7135 -3571 7215 -3561
rect 7135 -3600 7147 -3571
rect 3581 -3627 7147 -3600
rect 7203 -3600 7215 -3571
rect 8350 -3571 8430 -3561
rect 8350 -3600 8362 -3571
rect 7203 -3627 8362 -3600
rect 8418 -3600 8430 -3571
rect 8418 -3627 9845 -3600
rect 3581 -3660 9845 -3627
rect 9905 -3660 10065 -3600
rect 3581 -3675 10065 -3660
rect 6470 -3725 6665 -3675
rect 7380 -3725 7575 -3675
rect 7685 -3725 7880 -3675
rect 8595 -3725 8790 -3675
rect 8900 -3725 9095 -3675
rect 6165 -3771 6176 -3725
rect 6350 -3771 6361 -3725
rect 6469 -3771 6480 -3725
rect 6654 -3771 6665 -3725
rect 6773 -3771 6784 -3725
rect 6958 -3771 6969 -3725
rect 7077 -3771 7088 -3725
rect 7262 -3771 7273 -3725
rect 7381 -3771 7392 -3725
rect 7566 -3771 7577 -3725
rect 7685 -3771 7696 -3725
rect 7870 -3771 7881 -3725
rect 7989 -3771 8000 -3725
rect 8174 -3771 8185 -3725
rect 8293 -3771 8304 -3725
rect 8478 -3771 8489 -3725
rect 8597 -3771 8608 -3725
rect 8782 -3771 8793 -3725
rect 8901 -3771 8912 -3725
rect 9086 -3771 9097 -3725
rect 9205 -3771 9216 -3725
rect 9390 -3771 9401 -3725
rect 9509 -3771 9520 -3725
rect 9694 -3771 9705 -3725
rect 6820 -3785 6835 -3771
rect 6905 -3785 6920 -3771
rect 7125 -3785 7140 -3771
rect 7210 -3785 7225 -3771
rect 8035 -3785 8050 -3771
rect 8120 -3785 8135 -3771
rect 8340 -3785 8355 -3771
rect 8425 -3785 8440 -3771
rect 9255 -3785 9270 -3771
rect 9340 -3785 9355 -3771
rect 6088 -3817 6134 -3806
rect 5781 -3945 5903 -3934
rect 5781 -4445 5792 -3945
rect 5892 -4445 5903 -3945
rect 6392 -3817 6438 -3806
rect 6375 -4018 6392 -4008
rect 6696 -3817 6742 -3806
rect 6679 -3829 6696 -3819
rect 7000 -3817 7046 -3806
rect 6742 -3829 6759 -3819
rect 6679 -3990 6691 -3829
rect 6747 -3990 6759 -3829
rect 6679 -4000 6696 -3990
rect 6438 -4018 6455 -4008
rect 6375 -4074 6387 -4018
rect 6443 -4074 6455 -4018
rect 6375 -4084 6392 -4074
rect 6088 -4102 6134 -4091
rect 6438 -4084 6455 -4074
rect 6392 -4102 6438 -4091
rect 6742 -4000 6759 -3990
rect 6983 -3863 7000 -3853
rect 7304 -3817 7350 -3806
rect 7287 -3829 7304 -3819
rect 7608 -3817 7654 -3806
rect 7350 -3829 7367 -3819
rect 7046 -3863 7063 -3853
rect 6983 -4074 6995 -3863
rect 7051 -4074 7063 -3863
rect 7287 -3990 7299 -3829
rect 7355 -3990 7367 -3829
rect 7287 -4000 7304 -3990
rect 6983 -4084 7000 -4074
rect 6696 -4102 6742 -4091
rect 7046 -4084 7063 -4074
rect 7000 -4102 7046 -4091
rect 7350 -4000 7367 -3990
rect 7591 -3829 7608 -3819
rect 7912 -3817 7958 -3806
rect 7654 -3829 7671 -3819
rect 7591 -4074 7603 -3829
rect 7659 -4074 7671 -3829
rect 7895 -3829 7912 -3819
rect 8216 -3817 8262 -3806
rect 7958 -3829 7975 -3819
rect 7895 -3990 7907 -3829
rect 7963 -3990 7975 -3829
rect 7895 -4000 7912 -3990
rect 7591 -4084 7608 -4074
rect 7304 -4102 7350 -4091
rect 7654 -4084 7671 -4074
rect 7608 -4102 7654 -4091
rect 7958 -4000 7975 -3990
rect 8199 -3863 8216 -3853
rect 8520 -3817 8566 -3806
rect 8503 -3829 8520 -3819
rect 8824 -3817 8870 -3806
rect 8566 -3829 8583 -3819
rect 8262 -3863 8279 -3853
rect 8199 -4074 8211 -3863
rect 8267 -4074 8279 -3863
rect 8503 -3990 8515 -3829
rect 8571 -3990 8583 -3829
rect 8503 -4000 8520 -3990
rect 8199 -4084 8216 -4074
rect 7912 -4102 7958 -4091
rect 8262 -4084 8279 -4074
rect 8216 -4102 8262 -4091
rect 8566 -4000 8583 -3990
rect 8807 -3829 8824 -3819
rect 9128 -3817 9174 -3806
rect 8870 -3829 8887 -3819
rect 8807 -4074 8819 -3829
rect 8875 -4074 8887 -3829
rect 8807 -4084 8824 -4074
rect 8520 -4102 8566 -4091
rect 8870 -4084 8887 -4074
rect 9111 -3829 9128 -3819
rect 9432 -3817 9478 -3806
rect 9174 -3829 9191 -3819
rect 9111 -4074 9123 -3829
rect 9179 -4074 9191 -3829
rect 9111 -4084 9128 -4074
rect 8824 -4102 8870 -4091
rect 9174 -4084 9191 -4074
rect 9415 -4017 9432 -4007
rect 9736 -3817 9782 -3806
rect 9478 -4017 9495 -4007
rect 9415 -4074 9427 -4017
rect 9483 -4074 9495 -4017
rect 9415 -4084 9432 -4074
rect 9128 -4102 9174 -4091
rect 9478 -4084 9495 -4074
rect 9432 -4102 9478 -4091
rect 9736 -4102 9782 -4091
rect 9967 -3945 10089 -3934
rect 6165 -4183 6176 -4137
rect 6350 -4183 6361 -4137
rect 6469 -4183 6480 -4137
rect 6654 -4183 6665 -4137
rect 6773 -4183 6784 -4137
rect 6958 -4183 6969 -4137
rect 7077 -4183 7088 -4137
rect 7262 -4183 7273 -4137
rect 7381 -4183 7392 -4137
rect 7566 -4183 7577 -4137
rect 7685 -4183 7696 -4137
rect 7870 -4183 7881 -4137
rect 7989 -4183 8000 -4137
rect 8174 -4183 8185 -4137
rect 8293 -4183 8304 -4137
rect 8478 -4183 8489 -4137
rect 8597 -4183 8608 -4137
rect 8782 -4183 8793 -4137
rect 8901 -4183 8912 -4137
rect 9086 -4183 9097 -4137
rect 9205 -4183 9216 -4137
rect 9390 -4183 9401 -4137
rect 9509 -4183 9520 -4137
rect 9694 -4183 9705 -4137
rect 9967 -4241 9978 -3945
rect 9953 -4257 9978 -4241
rect 10078 -4241 10089 -3945
rect 9953 -4394 9967 -4257
rect 5781 -4456 5903 -4445
rect 9952 -4467 9967 -4394
rect 10078 -4405 10094 -4241
rect 10078 -4445 10089 -4405
rect 10072 -4467 10089 -4445
rect 9952 -4485 10089 -4467
rect 7498 -4660 7544 -4649
rect 7481 -4749 7498 -4747
rect 7713 -4651 7789 -4621
rect 7713 -4697 7724 -4651
rect 7778 -4697 7789 -4651
rect 7897 -4651 7973 -4621
rect 7897 -4697 7908 -4651
rect 7962 -4697 7973 -4651
rect 8081 -4651 8157 -4621
rect 8081 -4697 8092 -4651
rect 8146 -4697 8157 -4651
rect 8326 -4660 8372 -4649
rect 7636 -4743 7682 -4732
rect 7544 -4749 7561 -4747
rect 7481 -4871 7493 -4749
rect 7549 -4871 7561 -4749
rect 7481 -4873 7498 -4871
rect 7544 -4873 7561 -4871
rect 7820 -4743 7866 -4732
rect 7803 -4749 7820 -4747
rect 8004 -4743 8050 -4732
rect 7866 -4749 7883 -4747
rect 7803 -4871 7815 -4749
rect 7871 -4871 7883 -4749
rect 7803 -4873 7820 -4871
rect 7636 -4888 7682 -4877
rect 7866 -4873 7883 -4871
rect 7987 -4749 8004 -4747
rect 8188 -4743 8234 -4732
rect 8050 -4749 8067 -4747
rect 7987 -4871 7999 -4749
rect 8055 -4871 8067 -4749
rect 7987 -4873 8004 -4871
rect 7820 -4888 7866 -4877
rect 8050 -4873 8067 -4871
rect 8004 -4888 8050 -4877
rect 8188 -4888 8234 -4877
rect 7498 -4971 7544 -4960
rect 7713 -4969 7724 -4923
rect 7778 -4969 7789 -4923
rect 7713 -4999 7789 -4969
rect 7897 -4969 7908 -4923
rect 7962 -4969 7973 -4923
rect 4705 -5100 4809 -5090
rect 7897 -5100 7973 -4969
rect 8081 -4969 8092 -4923
rect 8146 -4969 8157 -4923
rect 8081 -4999 8157 -4969
rect 8326 -4971 8372 -4960
rect 11061 -5100 11165 -5090
rect 3570 -5180 4717 -5100
rect 4797 -5180 11073 -5100
rect 11153 -5180 11165 -5100
rect 4705 -5190 4809 -5180
rect 11061 -5190 11165 -5180
rect 3562 -5472 11642 -5418
rect 3562 -5473 9964 -5472
rect 3562 -5540 5457 -5473
rect 3562 -5627 4456 -5540
rect 4541 -5560 5457 -5540
rect 5546 -5478 9964 -5473
rect 5546 -5560 6013 -5478
rect 4541 -5627 6013 -5560
rect 3562 -5689 6013 -5627
rect 6368 -5675 9964 -5478
rect 10078 -5526 11642 -5472
rect 10078 -5628 10442 -5526
rect 10546 -5548 11642 -5526
rect 10546 -5628 11332 -5548
rect 10078 -5655 11332 -5628
rect 11441 -5655 11642 -5548
rect 10078 -5675 11642 -5655
rect 6368 -5689 11642 -5675
rect 3562 -5798 11642 -5689
<< via1 >>
rect 5349 2787 5401 2839
rect 5909 2576 5961 2579
rect 5909 2530 5912 2576
rect 5912 2530 5958 2576
rect 5958 2530 5961 2576
rect 5909 2527 5961 2530
rect 7769 2642 7774 2698
rect 7774 2642 7820 2698
rect 7820 2642 7825 2698
rect 8045 2642 8050 2698
rect 8050 2642 8096 2698
rect 8096 2642 8101 2698
rect 7907 2384 7963 2440
rect 7907 2246 7963 2302
rect 5577 1203 5657 1279
rect 7769 1822 7774 1878
rect 7774 1822 7820 1878
rect 7820 1822 7825 1878
rect 7677 1671 7678 1702
rect 7678 1671 7732 1702
rect 7732 1671 7733 1702
rect 7677 1646 7733 1671
rect 8045 1822 8050 1878
rect 8050 1822 8096 1878
rect 8096 1822 8101 1878
rect 8137 1671 8138 1702
rect 8138 1671 8192 1702
rect 8192 1671 8193 1702
rect 8137 1646 8193 1671
rect 7677 1203 7733 1279
rect 4010 786 4090 864
rect 8137 1203 8193 1279
rect 10213 1203 10293 1279
rect 10420 690 10500 750
rect 4454 365 4545 454
rect 11332 445 11441 552
rect 4717 259 4797 335
rect 11073 259 11153 335
rect 5067 -567 5072 -433
rect 5072 -567 5118 -433
rect 5118 -567 5123 -433
rect 5251 -567 5256 -433
rect 5256 -567 5302 -433
rect 5302 -567 5307 -433
rect 5389 -567 5394 -433
rect 5394 -567 5440 -433
rect 5440 -567 5445 -433
rect 5927 -567 5932 -433
rect 5932 -567 5978 -433
rect 5978 -567 5983 -433
rect 6111 -567 6116 -433
rect 6116 -567 6162 -433
rect 6162 -567 6167 -433
rect 6249 -567 6254 -433
rect 6254 -567 6300 -433
rect 6300 -567 6305 -433
rect 6691 -564 6696 -420
rect 6696 -564 6742 -420
rect 6742 -564 6747 -420
rect 6995 -577 7000 -521
rect 7000 -577 7046 -521
rect 7046 -577 7051 -521
rect 7299 -564 7304 -420
rect 7304 -564 7350 -420
rect 7350 -564 7355 -420
rect 7603 -577 7608 -521
rect 7608 -577 7654 -521
rect 7654 -577 7659 -521
rect 7907 -564 7912 -420
rect 7912 -564 7958 -420
rect 7958 -564 7963 -420
rect 8211 -577 8216 -521
rect 8216 -577 8262 -521
rect 8262 -577 8267 -521
rect 8515 -564 8520 -420
rect 8520 -564 8566 -420
rect 8566 -564 8571 -420
rect 8819 -577 8824 -521
rect 8824 -577 8870 -521
rect 8870 -577 8875 -521
rect 9123 -564 9128 -420
rect 9128 -564 9174 -420
rect 9174 -564 9179 -420
rect 9565 -567 9570 -433
rect 9570 -567 9616 -433
rect 9616 -567 9621 -433
rect 7798 -633 7854 -628
rect 8016 -633 8072 -628
rect 7798 -679 7854 -633
rect 8016 -679 8072 -633
rect 9703 -567 9708 -433
rect 9708 -567 9754 -433
rect 9754 -567 9759 -433
rect 9887 -567 9892 -433
rect 9892 -567 9938 -433
rect 9938 -567 9943 -433
rect 7798 -684 7854 -679
rect 8016 -684 8072 -679
rect 10425 -567 10430 -433
rect 10430 -567 10476 -433
rect 10476 -567 10481 -433
rect 10563 -567 10568 -433
rect 10568 -567 10614 -433
rect 10614 -567 10619 -433
rect 10747 -567 10752 -433
rect 10752 -567 10798 -433
rect 10798 -567 10803 -433
rect 5577 -1020 5657 -936
rect 6099 -1020 6179 -936
rect 6845 -1018 6925 -938
rect 7453 -1018 7533 -938
rect 7591 -1018 7671 -938
rect 8199 -1018 8279 -938
rect 8337 -1018 8417 -938
rect 8945 -1018 9025 -938
rect 9691 -1020 9771 -936
rect 10213 -1020 10293 -936
rect 7254 -1277 7334 -1232
rect 7254 -1312 7334 -1277
rect 8536 -1277 8616 -1232
rect 6111 -1826 6116 -1682
rect 6116 -1826 6162 -1682
rect 6162 -1826 6167 -1682
rect 6857 -1520 6862 -1376
rect 6862 -1520 6908 -1376
rect 6908 -1520 6913 -1376
rect 6553 -1736 6558 -1592
rect 6558 -1736 6604 -1592
rect 6604 -1736 6609 -1592
rect 7465 -1520 7470 -1376
rect 7470 -1520 7516 -1376
rect 7516 -1520 7521 -1376
rect 7161 -1736 7166 -1592
rect 7166 -1736 7212 -1592
rect 7212 -1736 7217 -1592
rect 8536 -1312 8616 -1277
rect 8349 -1520 8354 -1376
rect 8354 -1520 8400 -1376
rect 8400 -1520 8405 -1376
rect 8957 -1520 8962 -1376
rect 8962 -1520 9008 -1376
rect 9008 -1520 9013 -1376
rect 8653 -1736 8658 -1592
rect 8658 -1736 8704 -1592
rect 8704 -1736 8709 -1592
rect 9261 -1736 9266 -1592
rect 9266 -1736 9312 -1592
rect 9312 -1736 9317 -1592
rect 9703 -1826 9708 -1682
rect 9708 -1826 9754 -1682
rect 9754 -1826 9759 -1682
rect 5239 -2182 5319 -2102
rect 6375 -2182 6455 -2102
rect 6541 -2182 6621 -2102
rect 7149 -2182 7229 -2102
rect 8641 -2182 8721 -2102
rect 9249 -2182 9329 -2102
rect 9415 -2182 9495 -2102
rect 10551 -2182 10631 -2102
rect 5792 -2661 5892 -2500
rect 6387 -3071 6392 -2910
rect 6392 -3071 6438 -2910
rect 6438 -3071 6443 -2910
rect 6691 -3119 6696 -2958
rect 6696 -3119 6742 -2958
rect 6742 -3119 6747 -2958
rect 6995 -3091 7000 -2874
rect 7000 -3091 7046 -2874
rect 7046 -3091 7051 -2874
rect 7603 -2930 7608 -2874
rect 7608 -2930 7654 -2874
rect 7654 -2930 7659 -2874
rect 7299 -3119 7304 -2958
rect 7304 -3119 7350 -2958
rect 7350 -3119 7355 -2958
rect 8211 -2930 8216 -2874
rect 8216 -2930 8262 -2874
rect 8262 -2930 8267 -2874
rect 7907 -3119 7912 -2958
rect 7912 -3119 7958 -2958
rect 7958 -3119 7963 -2958
rect 8515 -3119 8520 -2958
rect 8520 -3119 8566 -2958
rect 8566 -3119 8571 -2958
rect 8819 -3119 8824 -2874
rect 8824 -3119 8870 -2874
rect 8870 -3119 8875 -2874
rect 9123 -3119 9128 -2958
rect 9128 -3119 9174 -2958
rect 9174 -3119 9179 -2958
rect 9427 -3071 9432 -2910
rect 9432 -3071 9478 -2910
rect 9478 -3071 9483 -2910
rect 9978 -2661 10078 -2500
rect 6835 -3174 6905 -3165
rect 7140 -3174 7210 -3165
rect 8050 -3174 8120 -3165
rect 8355 -3174 8425 -3165
rect 9270 -3174 9340 -3165
rect 6835 -3220 6905 -3174
rect 7140 -3220 7210 -3174
rect 8050 -3220 8120 -3174
rect 8355 -3220 8425 -3174
rect 9270 -3220 9340 -3174
rect 6835 -3225 6905 -3220
rect 7140 -3225 7210 -3220
rect 8050 -3225 8120 -3220
rect 8355 -3225 8425 -3220
rect 9270 -3225 9340 -3220
rect 6842 -3379 6898 -3323
rect 8057 -3379 8113 -3323
rect 9585 -3350 9645 -3290
rect 7147 -3627 7203 -3571
rect 8362 -3627 8418 -3571
rect 9845 -3660 9905 -3600
rect 6835 -3771 6905 -3725
rect 7140 -3771 7210 -3725
rect 8050 -3771 8120 -3725
rect 8355 -3771 8425 -3725
rect 9270 -3771 9340 -3725
rect 6835 -3785 6905 -3771
rect 7140 -3785 7210 -3771
rect 8050 -3785 8120 -3771
rect 8355 -3785 8425 -3771
rect 9270 -3785 9340 -3771
rect 5792 -4445 5892 -4284
rect 6691 -3990 6696 -3829
rect 6696 -3990 6742 -3829
rect 6742 -3990 6747 -3829
rect 6387 -4074 6392 -4018
rect 6392 -4074 6438 -4018
rect 6438 -4074 6443 -4018
rect 6995 -4074 7000 -3863
rect 7000 -4074 7046 -3863
rect 7046 -4074 7051 -3863
rect 7299 -3990 7304 -3829
rect 7304 -3990 7350 -3829
rect 7350 -3990 7355 -3829
rect 7603 -4074 7608 -3829
rect 7608 -4074 7654 -3829
rect 7654 -4074 7659 -3829
rect 7907 -3990 7912 -3829
rect 7912 -3990 7958 -3829
rect 7958 -3990 7963 -3829
rect 8211 -4074 8216 -3863
rect 8216 -4074 8262 -3863
rect 8262 -4074 8267 -3863
rect 8515 -3990 8520 -3829
rect 8520 -3990 8566 -3829
rect 8566 -3990 8571 -3829
rect 8819 -4074 8824 -3829
rect 8824 -4074 8870 -3829
rect 8870 -4074 8875 -3829
rect 9123 -4074 9128 -3829
rect 9128 -4074 9174 -3829
rect 9174 -4074 9179 -3829
rect 9427 -4074 9432 -4017
rect 9432 -4074 9478 -4017
rect 9478 -4074 9483 -4017
rect 9967 -4445 9978 -4257
rect 9978 -4445 10072 -4257
rect 9967 -4467 10072 -4445
rect 7493 -4871 7498 -4749
rect 7498 -4871 7544 -4749
rect 7544 -4871 7549 -4749
rect 7815 -4871 7820 -4749
rect 7820 -4871 7866 -4749
rect 7866 -4871 7871 -4749
rect 7999 -4871 8004 -4749
rect 8004 -4871 8050 -4749
rect 8050 -4871 8055 -4749
rect 4717 -5180 4797 -5100
rect 11073 -5180 11153 -5100
rect 4456 -5627 4541 -5540
rect 5457 -5560 5546 -5473
rect 6013 -5689 6368 -5478
rect 9964 -5675 10078 -5472
rect 10442 -5628 10546 -5526
rect 11332 -5655 11441 -5548
<< metal2 >>
rect 5325 2843 5425 2853
rect 3730 2839 5425 2843
rect 3730 2787 5349 2839
rect 5401 2787 5425 2839
rect 3730 2783 5425 2787
rect 5325 2773 5425 2783
rect 7757 2698 7837 2708
rect 7757 2642 7769 2698
rect 7825 2642 7837 2698
rect 7757 2632 7837 2642
rect 8033 2698 8113 2708
rect 8033 2642 8045 2698
rect 8101 2642 8113 2698
rect 8033 2632 8113 2642
rect 5895 2583 5975 2593
rect 5885 2579 5985 2583
rect 5885 2527 5909 2579
rect 5961 2527 7276 2579
rect 5885 2523 7276 2527
rect 5895 2513 5975 2523
rect 7220 2192 7276 2523
rect 7769 2440 7825 2632
rect 7894 2440 7974 2452
rect 7769 2384 7907 2440
rect 7963 2384 7974 2440
rect 7769 2192 7825 2384
rect 7894 2372 7974 2384
rect 7895 2302 7975 2312
rect 8045 2302 8101 2632
rect 7895 2246 7907 2302
rect 7963 2246 8101 2302
rect 7895 2236 7975 2246
rect 7220 2136 7825 2192
rect 7769 1888 7825 2136
rect 8045 2192 8101 2246
rect 8045 2136 8645 2192
rect 8045 1888 8101 2136
rect 7757 1878 7837 1888
rect 7757 1822 7769 1878
rect 7825 1822 7837 1878
rect 7757 1812 7837 1822
rect 8033 1878 8113 1888
rect 8033 1822 8045 1878
rect 8101 1822 8113 1878
rect 8033 1812 8113 1822
rect 7665 1702 7745 1712
rect 7665 1646 7677 1702
rect 7733 1646 7745 1702
rect 7665 1636 7745 1646
rect 8125 1702 8205 1712
rect 8125 1646 8137 1702
rect 8193 1646 8205 1702
rect 8125 1636 8205 1646
rect 5565 1279 5659 1291
rect 7677 1281 7733 1636
rect 8137 1281 8193 1636
rect 5565 1203 5577 1279
rect 5657 1203 5659 1279
rect 5565 1201 5659 1203
rect 7675 1279 7747 1281
rect 7675 1203 7677 1279
rect 7733 1203 7747 1279
rect 3993 864 4106 881
rect 3993 786 4010 864
rect 4090 786 4106 864
rect 3993 775 4106 786
rect 4010 320 4090 775
rect 4446 454 4555 467
rect 4446 365 4454 454
rect 4545 365 4555 454
rect 4446 358 4555 365
rect 4000 300 4100 320
rect 4000 220 4010 300
rect 4090 220 4100 300
rect 4000 210 4100 220
rect 4454 -1018 4545 358
rect 4705 335 4809 349
rect 4705 259 4717 335
rect 4797 259 4809 335
rect 4705 249 4809 259
rect 4456 -5518 4543 -1018
rect 4717 -5090 4797 249
rect 5045 26 5145 36
rect 5045 -54 5055 26
rect 5135 -54 5145 26
rect 5045 -64 5145 -54
rect 5367 26 5467 36
rect 5367 -54 5377 26
rect 5457 -54 5467 26
rect 5367 -64 5467 -54
rect 5055 -433 5135 -64
rect 5251 -431 5307 -423
rect 5055 -567 5067 -433
rect 5123 -567 5135 -433
rect 5055 -569 5135 -567
rect 5239 -433 5319 -431
rect 5239 -567 5251 -433
rect 5307 -567 5319 -433
rect 5067 -577 5123 -569
rect 5239 -2092 5319 -567
rect 5377 -433 5457 -64
rect 5377 -567 5389 -433
rect 5445 -567 5457 -433
rect 5377 -569 5457 -567
rect 5389 -577 5445 -569
rect 5577 -924 5657 1201
rect 7675 1191 7747 1203
rect 8123 1279 8195 1281
rect 8123 1203 8137 1279
rect 8193 1203 8195 1279
rect 8123 1191 8195 1203
rect 10201 1279 10305 1291
rect 10201 1203 10213 1279
rect 10293 1203 10305 1279
rect 10201 1201 10305 1203
rect 5905 26 6005 36
rect 5905 -54 5915 26
rect 5995 -54 6005 26
rect 5905 -64 6005 -54
rect 6227 26 6327 36
rect 6227 -54 6237 26
rect 6317 -54 6327 26
rect 6227 -64 6327 -54
rect 6669 26 6769 36
rect 6669 -54 6679 26
rect 6759 -54 6769 26
rect 6669 -64 6769 -54
rect 7277 26 7377 36
rect 7277 -54 7287 26
rect 7367 -54 7377 26
rect 7277 -64 7377 -54
rect 7885 26 7985 36
rect 7885 -54 7895 26
rect 7975 -54 7985 26
rect 7885 -64 7985 -54
rect 8493 26 8593 36
rect 8493 -54 8503 26
rect 8583 -54 8593 26
rect 8493 -64 8593 -54
rect 9101 26 9201 36
rect 9101 -54 9111 26
rect 9191 -54 9201 26
rect 9101 -64 9201 -54
rect 9543 26 9643 36
rect 9543 -54 9553 26
rect 9633 -54 9643 26
rect 9543 -64 9643 -54
rect 9865 26 9965 36
rect 9865 -54 9875 26
rect 9955 -54 9965 26
rect 9865 -64 9965 -54
rect 5915 -433 5995 -64
rect 6111 -431 6167 -423
rect 5915 -567 5927 -433
rect 5983 -567 5995 -433
rect 5915 -569 5995 -567
rect 6099 -433 6179 -431
rect 6099 -567 6111 -433
rect 6167 -567 6179 -433
rect 5927 -577 5983 -569
rect 5565 -936 5669 -924
rect 6099 -926 6179 -567
rect 6237 -433 6317 -64
rect 6237 -567 6249 -433
rect 6305 -567 6317 -433
rect 6679 -420 6759 -64
rect 6679 -564 6691 -420
rect 6747 -564 6759 -420
rect 7287 -420 7367 -64
rect 6679 -566 6759 -564
rect 6983 -521 7063 -511
rect 6237 -569 6317 -567
rect 6249 -577 6305 -569
rect 6691 -574 6747 -566
rect 6983 -577 6995 -521
rect 7051 -577 7063 -521
rect 7287 -564 7299 -420
rect 7355 -564 7367 -420
rect 7895 -420 7975 -64
rect 7287 -566 7367 -564
rect 7591 -521 7671 -511
rect 7299 -574 7355 -566
rect 6983 -587 7063 -577
rect 7591 -577 7603 -521
rect 7659 -577 7671 -521
rect 7895 -564 7907 -420
rect 7963 -564 7975 -420
rect 8503 -420 8583 -64
rect 7895 -566 7975 -564
rect 8199 -521 8279 -511
rect 7907 -574 7963 -566
rect 5565 -1020 5577 -936
rect 5657 -1020 5669 -936
rect 5565 -1030 5669 -1020
rect 6087 -936 6191 -926
rect 7591 -928 7671 -577
rect 8199 -577 8211 -521
rect 8267 -577 8279 -521
rect 8503 -564 8515 -420
rect 8571 -564 8583 -420
rect 9111 -420 9191 -64
rect 8503 -566 8583 -564
rect 8807 -521 8887 -511
rect 8515 -574 8571 -566
rect 7786 -628 7866 -618
rect 7786 -684 7798 -628
rect 7854 -684 7866 -628
rect 7786 -758 7866 -684
rect 8004 -628 8084 -618
rect 8004 -684 8016 -628
rect 8072 -684 8084 -628
rect 7776 -768 7876 -758
rect 7776 -848 7786 -768
rect 7866 -848 7876 -768
rect 7776 -858 7876 -848
rect 8004 -928 8084 -684
rect 8199 -758 8279 -577
rect 8807 -577 8819 -521
rect 8875 -577 8887 -521
rect 9111 -564 9123 -420
rect 9179 -564 9191 -420
rect 9111 -566 9191 -564
rect 9553 -433 9633 -64
rect 9703 -431 9759 -423
rect 9123 -574 9179 -566
rect 9553 -567 9565 -433
rect 9621 -567 9633 -433
rect 9553 -569 9633 -567
rect 9691 -433 9771 -431
rect 9691 -567 9703 -433
rect 9759 -567 9771 -433
rect 9565 -577 9621 -569
rect 8807 -587 8887 -577
rect 8189 -768 8289 -758
rect 8189 -848 8199 -768
rect 8279 -848 8289 -768
rect 8189 -858 8289 -848
rect 8199 -928 8279 -858
rect 9691 -926 9771 -567
rect 9875 -433 9955 -64
rect 9875 -567 9887 -433
rect 9943 -567 9955 -433
rect 9875 -569 9955 -567
rect 9887 -577 9943 -569
rect 10213 -926 10293 1201
rect 10400 790 10520 810
rect 10400 690 10420 790
rect 10500 690 10520 790
rect 10400 670 10520 690
rect 11305 552 11463 567
rect 11305 445 11332 552
rect 11441 445 11463 552
rect 11305 434 11463 445
rect 11061 335 11165 347
rect 11061 259 11073 335
rect 11153 259 11165 335
rect 11061 247 11165 259
rect 10403 26 10503 36
rect 10403 -54 10413 26
rect 10493 -54 10503 26
rect 10403 -64 10503 -54
rect 10725 26 10825 36
rect 10725 -54 10735 26
rect 10815 -54 10825 26
rect 10725 -64 10825 -54
rect 10413 -433 10493 -64
rect 10563 -431 10619 -423
rect 10413 -567 10425 -433
rect 10481 -567 10493 -433
rect 10413 -569 10493 -567
rect 10551 -433 10631 -431
rect 10551 -567 10563 -433
rect 10619 -567 10631 -433
rect 10425 -577 10481 -569
rect 6087 -1020 6099 -936
rect 6179 -1020 6191 -936
rect 6087 -1030 6191 -1020
rect 6833 -938 6937 -928
rect 6833 -1018 6845 -938
rect 6925 -1018 6937 -938
rect 6833 -1032 6937 -1018
rect 7441 -938 7681 -928
rect 7994 -938 8094 -928
rect 7441 -1018 7453 -938
rect 7533 -1018 7591 -938
rect 7671 -1018 8004 -938
rect 8084 -1018 8094 -938
rect 7441 -1032 7681 -1018
rect 7994 -1028 8094 -1018
rect 8187 -938 8429 -928
rect 8187 -1018 8199 -938
rect 8279 -1018 8337 -938
rect 8417 -1018 8429 -938
rect 8187 -1032 8429 -1018
rect 8933 -938 9037 -927
rect 8933 -1018 8945 -938
rect 9025 -1018 9037 -938
rect 8933 -1031 9037 -1018
rect 9679 -936 9783 -926
rect 9679 -1020 9691 -936
rect 9771 -1020 9783 -936
rect 9679 -1030 9783 -1020
rect 10201 -936 10305 -926
rect 10201 -1020 10213 -936
rect 10293 -1020 10305 -936
rect 10201 -1030 10305 -1020
rect 6845 -1376 6925 -1032
rect 7244 -1232 7344 -1222
rect 7244 -1312 7254 -1232
rect 7334 -1312 7344 -1232
rect 7244 -1322 7344 -1312
rect 6845 -1520 6857 -1376
rect 6913 -1520 6925 -1376
rect 6845 -1522 6925 -1520
rect 7453 -1376 7533 -1032
rect 7453 -1520 7465 -1376
rect 7521 -1520 7533 -1376
rect 7453 -1522 7533 -1520
rect 8337 -1376 8417 -1032
rect 8526 -1232 8626 -1222
rect 8526 -1312 8536 -1232
rect 8616 -1312 8626 -1232
rect 8526 -1322 8626 -1312
rect 8337 -1520 8349 -1376
rect 8405 -1520 8417 -1376
rect 8337 -1522 8417 -1520
rect 8945 -1376 9025 -1031
rect 8945 -1520 8957 -1376
rect 9013 -1520 9025 -1376
rect 8945 -1522 9025 -1520
rect 6857 -1530 6913 -1522
rect 7465 -1530 7521 -1522
rect 8349 -1530 8405 -1522
rect 8957 -1530 9013 -1522
rect 6553 -1590 6609 -1582
rect 7161 -1590 7217 -1582
rect 8653 -1590 8709 -1582
rect 9261 -1590 9317 -1582
rect 6541 -1592 6621 -1590
rect 6099 -1682 6179 -1672
rect 5790 -1826 6111 -1682
rect 6167 -1826 6179 -1682
rect 5227 -2102 5331 -2092
rect 5227 -2182 5239 -2102
rect 5319 -2182 5331 -2102
rect 5227 -2192 5331 -2182
rect 5790 -2362 5894 -1826
rect 6099 -1837 6179 -1826
rect 6541 -1736 6553 -1592
rect 6609 -1736 6621 -1592
rect 6541 -2090 6621 -1736
rect 7149 -1592 7229 -1590
rect 7149 -1736 7161 -1592
rect 7217 -1736 7229 -1592
rect 7149 -2090 7229 -1736
rect 8641 -1592 8721 -1590
rect 8641 -1736 8653 -1592
rect 8709 -1736 8721 -1592
rect 8641 -2090 8721 -1736
rect 9249 -1592 9329 -1590
rect 9249 -1736 9261 -1592
rect 9317 -1736 9329 -1592
rect 9249 -2090 9329 -1736
rect 9691 -1682 9771 -1672
rect 9691 -1826 9703 -1682
rect 9759 -1826 10080 -1682
rect 9691 -1837 9771 -1826
rect 6363 -2102 6467 -2090
rect 6363 -2182 6375 -2102
rect 6455 -2182 6467 -2102
rect 6363 -2194 6467 -2182
rect 6529 -2102 6633 -2090
rect 6529 -2182 6541 -2102
rect 6621 -2182 6633 -2102
rect 6529 -2194 6633 -2182
rect 7137 -2102 7241 -2090
rect 7137 -2182 7149 -2102
rect 7229 -2182 7241 -2102
rect 7137 -2194 7241 -2182
rect 8629 -2102 8733 -2090
rect 8629 -2182 8641 -2102
rect 8721 -2182 8733 -2102
rect 8629 -2194 8733 -2182
rect 9237 -2102 9341 -2090
rect 9237 -2182 9249 -2102
rect 9329 -2182 9341 -2102
rect 9237 -2194 9341 -2182
rect 9403 -2102 9507 -2090
rect 9403 -2182 9415 -2102
rect 9495 -2182 9507 -2102
rect 9403 -2194 9507 -2182
rect 5449 -2466 5894 -2362
rect 4705 -5100 4809 -5090
rect 4705 -5180 4717 -5100
rect 4797 -5180 4809 -5100
rect 4705 -5190 4809 -5180
rect 5457 -5220 5546 -2466
rect 5790 -2500 5894 -2466
rect 5790 -2661 5792 -2500
rect 5892 -2661 5894 -2500
rect 5790 -2673 5894 -2661
rect 6375 -2910 6455 -2194
rect 9415 -2672 9495 -2194
rect 6375 -3071 6387 -2910
rect 6443 -3071 6455 -2910
rect 6983 -2728 9495 -2672
rect 9976 -2353 10080 -1826
rect 10551 -2092 10631 -567
rect 10735 -433 10815 -64
rect 10735 -567 10747 -433
rect 10803 -567 10815 -433
rect 10735 -569 10815 -567
rect 10747 -577 10803 -569
rect 10539 -2102 10643 -2092
rect 10539 -2182 10551 -2102
rect 10631 -2182 10643 -2102
rect 10539 -2192 10643 -2182
rect 9976 -2457 10546 -2353
rect 9976 -2500 10080 -2457
rect 9976 -2661 9978 -2500
rect 10078 -2661 10080 -2500
rect 9976 -2673 10080 -2661
rect 6983 -2874 7063 -2728
rect 6375 -3081 6455 -3071
rect 6679 -2958 6759 -2948
rect 6679 -3119 6691 -2958
rect 6747 -3119 6759 -2958
rect 6983 -3091 6995 -2874
rect 7051 -3091 7063 -2874
rect 7591 -2874 7671 -2864
rect 7591 -2930 7603 -2874
rect 7659 -2930 7671 -2874
rect 7591 -2940 7671 -2930
rect 8199 -2874 8279 -2728
rect 8199 -2930 8211 -2874
rect 8267 -2930 8279 -2874
rect 8199 -2940 8279 -2930
rect 8807 -2874 8887 -2864
rect 6983 -3099 7063 -3091
rect 7287 -2958 7367 -2948
rect 6679 -3449 6759 -3119
rect 7287 -3119 7299 -2958
rect 7355 -3119 7367 -2958
rect 6820 -3165 7225 -3155
rect 6820 -3225 6835 -3165
rect 6905 -3225 7140 -3165
rect 7210 -3225 7225 -3165
rect 6820 -3235 7225 -3225
rect 6830 -3323 6910 -3313
rect 6830 -3379 6842 -3323
rect 6898 -3379 6910 -3323
rect 6830 -3389 6910 -3379
rect 7287 -3449 7367 -3119
rect 7895 -2958 7975 -2948
rect 7895 -3119 7907 -2958
rect 7963 -3119 7975 -2958
rect 7895 -3449 7975 -3119
rect 8503 -2958 8583 -2948
rect 8503 -3119 8515 -2958
rect 8571 -3119 8583 -2958
rect 8035 -3165 8440 -3155
rect 8035 -3225 8050 -3165
rect 8120 -3225 8355 -3165
rect 8425 -3225 8440 -3165
rect 8035 -3235 8440 -3225
rect 8045 -3323 8125 -3313
rect 8045 -3379 8057 -3323
rect 8113 -3379 8125 -3323
rect 8045 -3389 8125 -3379
rect 8503 -3449 8583 -3119
rect 8807 -3119 8819 -2874
rect 8875 -3119 8887 -2874
rect 9415 -2910 9495 -2728
rect 8807 -3129 8887 -3119
rect 9111 -2958 9191 -2948
rect 9111 -3119 9123 -2958
rect 9179 -3119 9191 -2958
rect 9415 -3071 9427 -2910
rect 9483 -3071 9495 -2910
rect 9415 -3081 9495 -3071
rect 9111 -3449 9191 -3119
rect 9255 -3165 9355 -3155
rect 9549 -3165 9775 -3164
rect 9255 -3225 9270 -3165
rect 9340 -3224 9775 -3165
rect 9340 -3225 9514 -3224
rect 9255 -3235 9355 -3225
rect 9570 -3290 9655 -3280
rect 9570 -3350 9585 -3290
rect 9645 -3350 9655 -3290
rect 9570 -3365 9655 -3350
rect 6679 -3505 9191 -3449
rect 6679 -3829 6759 -3505
rect 7135 -3571 7215 -3561
rect 7135 -3627 7147 -3571
rect 7203 -3627 7215 -3571
rect 7135 -3637 7215 -3627
rect 6820 -3725 7225 -3715
rect 6820 -3785 6835 -3725
rect 6905 -3785 7140 -3725
rect 7210 -3785 7225 -3725
rect 6820 -3795 7225 -3785
rect 6679 -3990 6691 -3829
rect 6747 -3990 6759 -3829
rect 7287 -3829 7367 -3505
rect 6375 -4018 6455 -4008
rect 6375 -4074 6387 -4018
rect 6443 -4074 6455 -4018
rect 6375 -4084 6455 -4074
rect 5790 -4284 5894 -4272
rect 5790 -4445 5792 -4284
rect 5892 -4445 5894 -4284
rect 6679 -4336 6759 -3990
rect 6983 -3863 7063 -3853
rect 6983 -4074 6995 -3863
rect 7051 -4074 7063 -3863
rect 7287 -3990 7299 -3829
rect 7355 -3990 7367 -3829
rect 7287 -4000 7367 -3990
rect 7591 -3829 7671 -3819
rect 6983 -4220 7063 -4074
rect 7591 -4074 7603 -3829
rect 7659 -4074 7671 -3829
rect 7895 -3829 7975 -3505
rect 8350 -3571 8430 -3561
rect 8350 -3627 8362 -3571
rect 8418 -3627 8430 -3571
rect 8350 -3637 8430 -3627
rect 8035 -3725 8440 -3715
rect 8035 -3785 8050 -3725
rect 8120 -3785 8355 -3725
rect 8425 -3785 8440 -3725
rect 8035 -3795 8440 -3785
rect 7895 -3990 7907 -3829
rect 7963 -3990 7975 -3829
rect 8503 -3829 8583 -3505
rect 7895 -4000 7975 -3990
rect 8199 -3863 8279 -3853
rect 7591 -4084 7671 -4074
rect 8199 -4074 8211 -3863
rect 8267 -4074 8279 -3863
rect 8503 -3990 8515 -3829
rect 8571 -3990 8583 -3829
rect 8503 -4000 8583 -3990
rect 8807 -3829 8887 -3819
rect 8199 -4220 8279 -4074
rect 8807 -4074 8819 -3829
rect 8875 -4074 8887 -3829
rect 8807 -4084 8887 -4074
rect 9111 -3829 9191 -3505
rect 9585 -3505 9645 -3365
rect 9715 -3385 9775 -3224
rect 9715 -3445 9905 -3385
rect 9585 -3565 9775 -3505
rect 9255 -3725 9355 -3715
rect 9715 -3725 9775 -3565
rect 9845 -3590 9905 -3445
rect 9835 -3600 9915 -3590
rect 9835 -3660 9845 -3600
rect 9905 -3660 9915 -3600
rect 9835 -3670 9915 -3660
rect 9255 -3785 9270 -3725
rect 9340 -3785 9775 -3725
rect 9255 -3795 9355 -3785
rect 9111 -4074 9123 -3829
rect 9179 -4074 9191 -3829
rect 9111 -4084 9191 -4074
rect 9415 -4017 9495 -4007
rect 9415 -4074 9427 -4017
rect 9483 -4074 9495 -4017
rect 9415 -4220 9495 -4074
rect 6983 -4276 9495 -4220
rect 9953 -4257 10094 -4241
rect 6679 -4347 9201 -4336
rect 6679 -4403 9111 -4347
rect 9191 -4403 9201 -4347
rect 9953 -4394 9967 -4257
rect 6679 -4413 9201 -4403
rect 5790 -4747 5894 -4445
rect 5790 -4749 7883 -4747
rect 5790 -4871 7493 -4749
rect 7549 -4871 7815 -4749
rect 7871 -4871 7883 -4749
rect 5790 -4873 7883 -4871
rect 7987 -4749 8067 -4413
rect 9952 -4467 9967 -4394
rect 10072 -4405 10094 -4257
rect 10072 -4467 10089 -4405
rect 9952 -4485 10089 -4467
rect 7987 -4871 7999 -4749
rect 8055 -4871 8067 -4749
rect 7987 -4873 8067 -4871
rect 5431 -5473 5583 -5220
rect 6018 -5469 6368 -4873
rect 9970 -5408 10069 -4485
rect 9970 -5453 10087 -5408
rect 9960 -5464 10087 -5453
rect 4432 -5540 4567 -5518
rect 4432 -5627 4456 -5540
rect 4541 -5627 4567 -5540
rect 5431 -5560 5457 -5473
rect 5546 -5560 5583 -5473
rect 5431 -5593 5583 -5560
rect 5999 -5478 6389 -5469
rect 4432 -5642 4567 -5627
rect 5999 -5689 6013 -5478
rect 6368 -5689 6389 -5478
rect 5999 -5710 6389 -5689
rect 9960 -5472 10086 -5464
rect 9960 -5675 9964 -5472
rect 10078 -5675 10086 -5472
rect 10442 -5516 10546 -2457
rect 11073 -5090 11153 247
rect 11061 -5100 11165 -5090
rect 11061 -5180 11073 -5100
rect 11153 -5180 11165 -5100
rect 11061 -5190 11165 -5180
rect 10431 -5526 10559 -5516
rect 10431 -5628 10442 -5526
rect 10546 -5628 10559 -5526
rect 11332 -5536 11441 434
rect 10431 -5662 10559 -5628
rect 11322 -5548 11450 -5536
rect 11322 -5655 11332 -5548
rect 11441 -5655 11450 -5548
rect 9960 -5694 10086 -5675
rect 11322 -5677 11450 -5655
<< via2 >>
rect 4010 220 4090 300
rect 5055 -54 5135 26
rect 5377 -54 5457 26
rect 5915 -54 5995 26
rect 6237 -54 6317 26
rect 6679 -54 6759 26
rect 7287 -54 7367 26
rect 7895 -54 7975 26
rect 8503 -54 8583 26
rect 9111 -54 9191 26
rect 9553 -54 9633 26
rect 9875 -54 9955 26
rect 6995 -577 7051 -521
rect 7603 -577 7659 -521
rect 7786 -848 7866 -768
rect 8819 -577 8875 -521
rect 8199 -848 8279 -768
rect 10420 750 10500 790
rect 10420 710 10500 750
rect 10413 -54 10493 26
rect 10735 -54 10815 26
rect 8004 -1018 8084 -938
rect 7254 -1312 7334 -1232
rect 8536 -1312 8616 -1232
rect 6387 -3071 6443 -2910
rect 6995 -3091 7051 -3035
rect 7603 -2930 7659 -2874
rect 7147 -3223 7203 -3167
rect 6842 -3379 6898 -3323
rect 8362 -3223 8418 -3167
rect 8057 -3379 8113 -3323
rect 8819 -3119 8875 -2874
rect 9427 -3071 9483 -2910
rect 7147 -3627 7203 -3571
rect 6842 -3783 6898 -3727
rect 6387 -4074 6443 -4018
rect 6995 -3919 7051 -3863
rect 7603 -4074 7659 -3829
rect 8362 -3627 8418 -3571
rect 8057 -3783 8113 -3727
rect 8211 -3919 8267 -3863
rect 8819 -4074 8875 -3829
rect 9123 -4074 9179 -3829
rect 9111 -4403 9191 -4347
<< metal3 >>
rect 10400 790 10520 810
rect 10400 710 10420 790
rect 10500 710 10520 790
rect 10400 690 10520 710
rect 4000 300 4100 320
rect 4000 220 4010 300
rect 4090 220 4100 300
rect 4000 210 4100 220
rect 4010 26 4090 210
rect 5045 26 5145 36
rect 5367 26 5467 36
rect 5905 26 6005 36
rect 6227 26 6327 36
rect 6669 26 6769 36
rect 7885 26 7985 146
rect 10420 36 10500 690
rect 8493 26 8593 36
rect 9101 26 9201 36
rect 9543 26 9643 36
rect 9865 26 9965 36
rect 10403 26 10503 36
rect 10725 26 10825 36
rect 4010 -54 5055 26
rect 5135 -54 5377 26
rect 5457 -54 5915 26
rect 5995 -54 6237 26
rect 6317 -54 6679 26
rect 6759 -54 7287 26
rect 7367 -54 7895 26
rect 7975 -54 8503 26
rect 8583 -54 9111 26
rect 9191 -54 9553 26
rect 9633 -54 9875 26
rect 9955 -54 10413 26
rect 10493 -54 10735 26
rect 10815 -54 10825 26
rect 5045 -64 5145 -54
rect 5367 -64 5467 -54
rect 5905 -64 6005 -54
rect 6227 -64 6327 -54
rect 6669 -64 6769 -54
rect 7277 -64 7377 -54
rect 7885 -64 7985 -54
rect 8493 -64 8593 -54
rect 9101 -64 9201 -54
rect 9543 -64 9643 -54
rect 9865 -64 9965 -54
rect 10403 -64 10503 -54
rect 10725 -64 10825 -54
rect 6983 -521 7063 -511
rect 6983 -577 6995 -521
rect 7051 -577 7063 -521
rect 6983 -587 7063 -577
rect 7591 -521 7671 -511
rect 8807 -521 8887 -511
rect 7591 -577 7603 -521
rect 7659 -577 8819 -521
rect 8875 -577 8887 -521
rect 7591 -587 7671 -577
rect 8807 -587 8887 -577
rect 6995 -768 7051 -587
rect 7776 -768 7876 -758
rect 8189 -768 8289 -758
rect 6995 -848 7786 -768
rect 7866 -848 8199 -768
rect 8279 -848 8289 -768
rect 7244 -1232 7344 -848
rect 7776 -858 7876 -848
rect 8189 -858 8289 -848
rect 7994 -938 8094 -928
rect 7994 -1018 8004 -938
rect 8084 -1018 8094 -938
rect 7994 -1066 8094 -1018
rect 7994 -1146 8616 -1066
rect 8536 -1222 8616 -1146
rect 7244 -1312 7254 -1232
rect 7334 -1312 7344 -1232
rect 7244 -1322 7344 -1312
rect 8526 -1232 8626 -1222
rect 8526 -1312 8536 -1232
rect 8616 -1312 8626 -1232
rect 8526 -1322 8626 -1312
rect 6375 -2874 8887 -2864
rect 6375 -2910 7603 -2874
rect 6375 -3071 6387 -2910
rect 6443 -2930 7603 -2910
rect 7659 -2930 8819 -2874
rect 6443 -2940 8819 -2930
rect 6443 -3071 6455 -2940
rect 6375 -3081 6455 -3071
rect 6983 -3035 7063 -3025
rect 6382 -3505 6447 -3081
rect 6983 -3091 6995 -3035
rect 7051 -3091 7063 -3035
rect 6830 -3323 6910 -3313
rect 6830 -3379 6842 -3323
rect 6898 -3379 6910 -3323
rect 6830 -3389 6910 -3379
rect 6983 -3389 7063 -3091
rect 8807 -3119 8819 -2940
rect 8875 -3119 8887 -2874
rect 9415 -2910 9495 -2900
rect 9415 -3071 9427 -2910
rect 9483 -3071 9495 -2910
rect 9415 -3081 9495 -3071
rect 7125 -3167 7225 -3155
rect 7125 -3223 7147 -3167
rect 7203 -3223 7225 -3167
rect 7125 -3235 7225 -3223
rect 8340 -3167 8440 -3155
rect 8340 -3223 8362 -3167
rect 8418 -3223 8440 -3167
rect 8340 -3235 8440 -3223
rect 8045 -3323 8125 -3313
rect 8045 -3379 8057 -3323
rect 8113 -3379 8125 -3323
rect 8045 -3389 8125 -3379
rect 8807 -3389 8887 -3119
rect 6983 -3449 7671 -3389
rect 6382 -3565 7063 -3505
rect 6820 -3727 6920 -3715
rect 6820 -3783 6842 -3727
rect 6898 -3783 6920 -3727
rect 6820 -3795 6920 -3783
rect 6983 -3863 7063 -3565
rect 7135 -3571 7215 -3561
rect 7135 -3627 7147 -3571
rect 7203 -3627 7215 -3571
rect 7135 -3637 7215 -3627
rect 6983 -3919 6995 -3863
rect 7051 -3919 7063 -3863
rect 6983 -3929 7063 -3919
rect 7591 -3829 7671 -3449
rect 8199 -3449 8887 -3389
rect 8035 -3727 8135 -3715
rect 8035 -3783 8057 -3727
rect 8113 -3783 8135 -3727
rect 8035 -3795 8135 -3783
rect 7591 -4008 7603 -3829
rect 6375 -4018 7603 -4008
rect 6375 -4074 6387 -4018
rect 6443 -4074 7603 -4018
rect 7659 -4008 7671 -3829
rect 8199 -3863 8279 -3449
rect 9422 -3505 9487 -3081
rect 8350 -3571 8430 -3561
rect 8350 -3627 8362 -3571
rect 8418 -3627 8430 -3571
rect 8350 -3637 8430 -3627
rect 8807 -3565 9487 -3505
rect 8199 -3919 8211 -3863
rect 8267 -3919 8279 -3863
rect 8199 -3929 8279 -3919
rect 8807 -3829 8887 -3565
rect 8807 -4008 8819 -3829
rect 7659 -4074 8819 -4008
rect 8875 -4074 8887 -3829
rect 6375 -4084 8887 -4074
rect 9111 -3829 9191 -3819
rect 9111 -4074 9123 -3829
rect 9179 -4074 9191 -3829
rect 9111 -4336 9191 -4074
rect 9101 -4347 9201 -4336
rect 9101 -4403 9111 -4347
rect 9191 -4403 9201 -4347
rect 9101 -4413 9201 -4403
<< via3 >>
rect 6842 -3379 6898 -3323
rect 7147 -3223 7203 -3167
rect 8362 -3223 8418 -3167
rect 8057 -3379 8113 -3323
rect 6842 -3783 6898 -3727
rect 7147 -3627 7203 -3571
rect 8057 -3783 8113 -3727
rect 8362 -3627 8418 -3571
<< metal4 >>
rect 7125 -3167 7225 -3155
rect 7125 -3223 7147 -3167
rect 7203 -3223 7225 -3167
rect 7125 -3235 7225 -3223
rect 8340 -3167 8440 -3155
rect 8340 -3223 8362 -3167
rect 8418 -3223 8440 -3167
rect 8340 -3235 8440 -3223
rect 6830 -3323 6910 -3313
rect 6830 -3379 6842 -3323
rect 6898 -3379 6910 -3323
rect 6830 -3389 6910 -3379
rect 6842 -3715 6898 -3389
rect 7147 -3561 7203 -3235
rect 8045 -3323 8125 -3313
rect 8045 -3379 8057 -3323
rect 8113 -3379 8125 -3323
rect 8045 -3389 8125 -3379
rect 7135 -3571 7215 -3561
rect 7135 -3627 7147 -3571
rect 7203 -3627 7215 -3571
rect 7135 -3637 7215 -3627
rect 8057 -3715 8113 -3389
rect 8362 -3561 8418 -3235
rect 8350 -3571 8430 -3561
rect 8350 -3627 8362 -3571
rect 8418 -3627 8430 -3571
rect 8350 -3637 8430 -3627
rect 6820 -3727 6920 -3715
rect 6820 -3783 6842 -3727
rect 6898 -3783 6920 -3727
rect 6820 -3795 6920 -3783
rect 8035 -3727 8135 -3715
rect 8035 -3783 8057 -3727
rect 8113 -3783 8135 -3727
rect 8035 -3795 8135 -3783
<< labels >>
rlabel metal2 7297 -4817 7297 -4817 7 lvsclean_SAlatch_0.VSS
rlabel metal3 7934 146 7934 146 1 lvsclean_SAlatch_0.VDD
rlabel metal2 5618 180 5618 180 1 lvsclean_SAlatch_0.Vout1
rlabel metal2 10254 180 10254 180 1 lvsclean_SAlatch_0.Vout2
rlabel metal1 7933 335 7933 335 1 lvsclean_SAlatch_0.Clk
rlabel metal1 10065 -3636 10065 -3636 3 lvsclean_SAlatch_0.Vin2
rlabel metal1 10065 -3315 10065 -3315 3 lvsclean_SAlatch_0.Vin1
rlabel metal1 6159 -2102 6159 -2102 1 lvsclean_SAlatch_0.Vp
rlabel metal1 9758 -2102 9758 -2102 1 lvsclean_SAlatch_0.Vq
rlabel metal1 9367 2357 9367 2357 3 x5.avdd
rlabel metal1 9363 501 9363 501 3 x5.avss
rlabel metal1 9163 1229 9163 1229 3 x5.in
rlabel metal1 9011 1233 9011 1233 3 x5.out
rlabel metal2 5935 2553 5935 2553 6 x4.A
rlabel metal2 5375 2813 5375 2813 6 x4.Y
rlabel metal1 6065 3233 6065 3233 6 x4.VDD
rlabel metal1 6065 2153 6065 2153 6 x4.VSS
rlabel metal1 6503 2357 6503 2357 7 x3.avdd
rlabel metal1 6507 501 6507 501 7 x3.avss
rlabel metal1 6707 1229 6707 1229 7 x3.in
rlabel metal1 6859 1233 6859 1233 7 x3.out
rlabel metal1 7933 3060 7933 3060 1 x2.VDD
rlabel metal2 7225 2162 7225 2162 7 x2.Vout1
rlabel metal2 8645 2162 8645 2162 3 x2.Vout2
rlabel metal2 7705 1302 7705 1302 5 x2.Vin1
rlabel metal2 8166 1302 8166 1302 5 x2.Vin2
rlabel metal1 7938 1460 7938 1460 5 x2.VSS
rlabel metal1 3562 -5618 3562 -5618 7 VSS
port 2 w
rlabel metal1 3570 -5140 3570 -5140 7 CLK
port 4 w
rlabel metal1 3581 -3637 3581 -3637 7 Vin2
port 8 w
rlabel metal1 3581 -3315 3581 -3315 7 Vin1
port 6 w
rlabel metal2 3730 2815 3730 2815 7 Vout
port 10 w
rlabel metal1 3654 4186 3654 4186 7 VDD
port 1 w
<< end >>
