* NGSPICE file created from osu_sc_or2_1.ext - technology: gf180mcuD

.subckt osu_sc_or2_1 A B Y VDD VSS
X0 a_90_720# A VSS VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X1 VDD B a_250_720# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.2125p ps=1.95u w=1.7u l=0.3u
X2 VSS B a_90_720# VSS nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 Y a_90_720# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 a_250_720# A a_90_720# VDD pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
X5 Y a_90_720# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.595p ps=2.4u w=1.7u l=0.3u
.ends

