* NGSPICE file created from no_offsetLatch.ext - technology: (null)

.subckt no_offsetLatch Clk Vin1 Vin2 VDD VSS Vout1 Vout2
X0 VDD.t27 Clk.t0 Vq VDD.t26 pfet_03v3
**devattr s=14080,496 d=14080,496
X1 Vq Vin2.t0 a_15720_n2324.t10 VSS.t2 nfet_03v3
**devattr s=15600,404 d=15600,404
X2 Vout1.t3 Vout2.t9 VDD.t19 VDD.t18 pfet_03v3
**devattr s=10400,304 d=10400,304
X3 VDD.t17 a_15520_1088 a_15432_1180 VDD.t16 pfet_03v3
**devattr s=17600,576 d=10400,304
X4 a_18456_1180 a_18256_1088 VDD.t5 VDD.t4 pfet_03v3
**devattr s=10400,304 d=17600,576
X5 Vp.t3 a_15382_n68 a_15294_24 VSS.t14 nfet_03v3
**devattr s=35200,976 d=20800,504
X6 Vq Vin2.t1 a_15720_n2324.t9 VSS.t13 nfet_03v3
**devattr s=15600,404 d=15600,404
X7 a_15720_n2324.t11 Vin1.t0 Vp.t2 VSS.t6 nfet_03v3
**devattr s=15600,404 d=15600,404
X8 Vp.t7 a_15216_n1453 a_15128_n1361 VSS.t15 nfet_03v3
**devattr s=26400,776 d=15600,404
X9 Vout1.t6 Vout2.t10 Vp.t6 VSS.t16 nfet_03v3
**devattr s=20800,504 d=20800,504
X10 Vout1.t5 Vout2.t11 Vp.t5 VSS.t17 nfet_03v3
**devattr s=20800,504 d=20800,504
X11 Vp.t1 Vin1.t1 a_15720_n2324.t0 VSS.t2 nfet_03v3
**devattr s=15600,404 d=15600,404
X12 Vq Vout1.t9 Vout2.t0 VSS.t1 nfet_03v3
**devattr s=20800,504 d=20800,504
X13 a_15720_n2324.t18 Vin1.t2 Vp.t14 VSS.t10 nfet_03v3
**devattr s=15600,404 d=15600,404
X14 Vout1.t8 Clk.t1 VDD.t25 VDD.t24 pfet_03v3
**devattr s=14080,496 d=14080,496
X15 a_16798_24 a_16598_n68 Vout1.t7 VSS.t18 nfet_03v3
**devattr s=20800,504 d=35200,976
X16 Vq Vout1.t10 Vout2.t6 VSS.t22 nfet_03v3
**devattr s=20800,504 d=20800,504
X17 Vout2.t5 Vout1.t11 VDD.t15 VDD.t14 pfet_03v3
**devattr s=10400,304 d=10400,304
X18 a_18594_24 a_18394_n68 Vq VSS.t21 nfet_03v3
**devattr s=20800,504 d=35200,976
X19 Vout2.t7 Vout1.t12 Vq VSS.t23 nfet_03v3
**devattr s=20800,504 d=20800,504
X20 Vp.t12 Vin1.t3 a_15720_n2324.t16 VSS.t13 nfet_03v3
**devattr s=15600,404 d=15600,404
X21 VDD.t23 Clk.t2 Vout2.t8 VDD.t22 pfet_03v3
**devattr s=14080,496 d=14080,496
X22 Vq Vin2.t2 a_15720_n2324.t8 VSS.t12 nfet_03v3
**devattr s=15600,404 d=15600,404
X23 Vq a_15216_n2416 a_15128_n2324 VSS.t15 nfet_03v3
**devattr s=26400,776 d=15600,404
X24 a_17212_n3110 a_17132_n3202 a_15720_n2324.t19 VSS.t24 nfet_03v3
**devattr s=8320,264 d=14080,496
X25 Vout1.t2 Vout2.t12 VDD.t1 VDD.t0 pfet_03v3
**devattr s=10400,304 d=10400,304
X26 a_15720_n2324.t7 Vin2.t3 Vq VSS.t11 nfet_03v3
**devattr s=15600,404 d=15600,404
X27 a_18760_n1361 a_18560_n1453 Vq VSS.t0 nfet_03v3
**devattr s=15600,404 d=26400,776
X28 a_15720_n2324.t6 Vin2.t4 Vq VSS.t10 nfet_03v3
**devattr s=15600,404 d=15600,404
X29 a_15720_n2324.t13 Vin1.t4 Vp.t9 VSS.t9 nfet_03v3
**devattr s=15600,404 d=15600,404
X30 Vp.t8 Vin1.t5 a_15720_n2324.t12 VSS.t8 nfet_03v3
**devattr s=15600,404 d=15600,404
X31 Vout2.t3 Vout1.t13 VDD.t11 VDD.t10 pfet_03v3
**devattr s=10400,304 d=10400,304
X32 VDD.t3 Vout2.t13 Vout1.t1 VDD.t2 pfet_03v3
**devattr s=10400,304 d=10400,304
X33 VSS.t4 a_16764_n3202 a_16676_n3110 VSS.t3 nfet_03v3
**devattr s=14080,496 d=8320,264
X34 a_15720_n2324.t17 Vin1.t6 Vp.t13 VSS.t11 nfet_03v3
**devattr s=15600,404 d=15600,404
X35 Vp.t10 Vin1.t7 a_15720_n2324.t14 VSS.t12 nfet_03v3
**devattr s=15600,404 d=15600,404
X36 Vp.t16 Clk.t3 VDD.t21 VDD.t20 pfet_03v3
**devattr s=14080,496 d=14080,496
X37 Vout2.t4 a_17178_n68 a_17090_24 VSS.t19 nfet_03v3
**devattr s=35200,976 d=20800,504
X38 a_18760_n2324 a_18560_n2416 Vp.t0 VSS.t0 nfet_03v3
**devattr s=15600,404 d=26400,776
X39 a_15720_n2324.t21 Clk.t4 VSS.t26 VSS.t25 nfet_03v3
**devattr s=8320,264 d=8320,264
X40 VDD.t13 Vout2.t14 Vout1.t0 VDD.t12 pfet_03v3
**devattr s=10400,304 d=10400,304
X41 a_15720_n2324.t5 Vin2.t5 Vq VSS.t9 nfet_03v3
**devattr s=15600,404 d=15600,404
X42 Vq Vin2.t6 a_15720_n2324.t4 VSS.t8 nfet_03v3
**devattr s=15600,404 d=15600,404
X43 Vp.t15 Vin1.t8 a_15720_n2324.t20 VSS.t7 nfet_03v3
**devattr s=15600,404 d=15600,404
X44 a_15720_n2324.t15 Vin1.t9 Vp.t11 VSS.t5 nfet_03v3
**devattr s=15600,404 d=15600,404
X45 VDD.t7 Vout1.t14 Vout2.t1 VDD.t6 pfet_03v3
**devattr s=10400,304 d=10400,304
X46 Vp.t4 Vout2.t15 Vout1.t4 VSS.t20 nfet_03v3
**devattr s=20800,504 d=20800,504
X47 Vq Vin2.t7 a_15720_n2324.t3 VSS.t7 nfet_03v3
**devattr s=15600,404 d=15600,404
X48 VDD.t9 Vout1.t15 Vout2.t2 VDD.t8 pfet_03v3
**devattr s=10400,304 d=10400,304
X49 a_15720_n2324.t2 Vin2.t8 Vq VSS.t6 nfet_03v3
**devattr s=15600,404 d=15600,404
X50 a_15720_n2324.t1 Vin2.t9 Vq VSS.t5 nfet_03v3
**devattr s=15600,404 d=15600,404
R0 Clk.n3 Clk.t3 21.1483
R1 Clk.n4 Clk.t1 21.1483
R2 Clk.n0 Clk.t2 21.1483
R3 Clk.n1 Clk.t0 21.1483
R4 Clk.n2 Clk.t4 20.5929
R5 Clk.n2 Clk.n1 19.1491
R6 Clk.n3 Clk.n2 19.1064
R7 Clk Clk.n0 2.23866
R8 Clk Clk.n4 2.23392
R9 Clk.n1 Clk.n0 1.01892
R10 Clk.n4 Clk.n3 1.01892
R11 VDD.t2 VDD.t4 490.324
R12 VDD.t18 VDD.t2 490.324
R13 VDD.t6 VDD.t18 490.324
R14 VDD.t10 VDD.t6 490.324
R15 VDD.t12 VDD.t10 490.324
R16 VDD.t0 VDD.t12 490.324
R17 VDD.t8 VDD.t0 490.324
R18 VDD.t14 VDD.t8 490.324
R19 VDD.t16 VDD.t14 490.324
R20 VDD.t4 VDD.n16 467.743
R21 VDD.n19 VDD.t16 467.743
R22 VDD.n9 VDD.t22 398.652
R23 VDD.t24 VDD.n18 398.652
R24 VDD.n16 VDD.t22 389.878
R25 VDD.n19 VDD.t24 389.878
R26 VDD.n7 VDD.n5 287.351
R27 VDD.n6 VDD.n4 287.351
R28 VDD.n2 VDD.t20 200.351
R29 VDD.n8 VDD.t26 200.351
R30 VDD.n18 VDD.n5 54.0755
R31 VDD.n18 VDD.n4 54.0755
R32 VDD.n9 VDD.n6 54.0755
R33 VDD.n9 VDD.n7 54.0755
R34 VDD.n20 VDD.n4 20.1255
R35 VDD.n20 VDD.n5 20.1255
R36 VDD.n15 VDD.n6 20.1255
R37 VDD.n15 VDD.n7 20.1255
R38 VDD.n27 VDD.n26 12.136
R39 VDD.n1 VDD.n0 12.136
R40 VDD.n13 VDD.n12 12.136
R41 VDD.n23 VDD.n22 12.136
R42 VDD.n25 VDD.n24 12.136
R43 VDD.n15 VDD.n14 11.111
R44 VDD.n21 VDD.n20 11.111
R45 VDD.n2 VDD.t21 10.8009
R46 VDD.n8 VDD.t27 10.8009
R47 VDD.n17 VDD.n3 9.536
R48 VDD.n11 VDD.n10 9.536
R49 VDD.n17 VDD.t25 7.4755
R50 VDD.n10 VDD.t23 7.4755
R51 VDD.n3 VDD.n2 5.4855
R52 VDD.n11 VDD.n8 5.4855
R53 VDD.n18 VDD.n17 2.1905
R54 VDD.n10 VDD.n9 2.1905
R55 VDD.n26 VDD.t11 1.8205
R56 VDD.n26 VDD.t13 1.8205
R57 VDD.n0 VDD.t19 1.8205
R58 VDD.n0 VDD.t7 1.8205
R59 VDD.n12 VDD.t5 1.8205
R60 VDD.n12 VDD.t3 1.8205
R61 VDD.n22 VDD.t15 1.8205
R62 VDD.n22 VDD.t17 1.8205
R63 VDD.n24 VDD.t1 1.8205
R64 VDD.n24 VDD.t9 1.8205
R65 VDD.n20 VDD.n19 1.5755
R66 VDD.n16 VDD.n15 1.5755
R67 VDD.n25 VDD.n23 0.667
R68 VDD.n13 VDD.n1 0.662
R69 VDD.n27 VDD.n25 0.622
R70 VDD.n27 VDD.n1 0.617
R71 VDD.n23 VDD.n21 0.47525
R72 VDD.n14 VDD.n13 0.47525
R73 VDD.n21 VDD.n3 0.34025
R74 VDD.n14 VDD.n11 0.34025
R75 VDD VDD.n27 0.1445
R76 Vin2.n5 Vin2.n4 23.1032
R77 Vin2.n1 Vin2.n0 23.1032
R78 Vin2.n8 Vin2.t1 21.8636
R79 Vin2.n4 Vin2.t2 16.3656
R80 Vin2.n0 Vin2.t0 16.3641
R81 Vin2.n4 Vin2.t8 16.021
R82 Vin2.n0 Vin2.t3 16.0195
R83 Vin2.n1 Vin2.t5 12.1667
R84 Vin2.n7 Vin2.t9 11.5195
R85 Vin2.n6 Vin2.t6 11.5195
R86 Vin2.n3 Vin2.t4 11.5195
R87 Vin2.n2 Vin2.t7 11.5195
R88 Vin2.n2 Vin2.n1 2.53166
R89 Vin2.n7 Vin2.n6 2.48408
R90 Vin2.n6 Vin2.n5 1.40666
R91 Vin2.n8 Vin2.n7 0.987026
R92 Vin2.n5 Vin2.n3 0.647132
R93 Vin2.n3 Vin2.n2 0.234605
R94 Vin2 Vin2.n8 0.2285
R95 a_15720_n2324.n16 a_15720_n2324.n15 11.2899
R96 a_15720_n2324.n16 a_15720_n2324.n14 8.49339
R97 a_15720_n2324.n1 a_15720_n2324.n0 4.89725
R98 a_15720_n2324.n12 a_15720_n2324.n11 4.89725
R99 a_15720_n2324.n4 a_15720_n2324.n2 4.89725
R100 a_15720_n2324.n7 a_15720_n2324.n5 4.89725
R101 a_15720_n2324.n10 a_15720_n2324.n8 4.89725
R102 a_15720_n2324.n4 a_15720_n2324.n3 4.88712
R103 a_15720_n2324.n7 a_15720_n2324.n6 4.88712
R104 a_15720_n2324.n10 a_15720_n2324.n9 4.88712
R105 a_15720_n2324.n18 a_15720_n2324.n17 4.4
R106 a_15720_n2324.n14 a_15720_n2324.n13 4.35275
R107 a_15720_n2324.n15 a_15720_n2324.t19 2.048
R108 a_15720_n2324.n15 a_15720_n2324.t21 2.048
R109 a_15720_n2324.n17 a_15720_n2324.n16 1.95895
R110 a_15720_n2324.n0 a_15720_n2324.t10 1.0925
R111 a_15720_n2324.n0 a_15720_n2324.t13 1.0925
R112 a_15720_n2324.n11 a_15720_n2324.t9 1.0925
R113 a_15720_n2324.n11 a_15720_n2324.t15 1.0925
R114 a_15720_n2324.n13 a_15720_n2324.t16 1.0925
R115 a_15720_n2324.n13 a_15720_n2324.t1 1.0925
R116 a_15720_n2324.n2 a_15720_n2324.t20 1.0925
R117 a_15720_n2324.n2 a_15720_n2324.t7 1.0925
R118 a_15720_n2324.n3 a_15720_n2324.t3 1.0925
R119 a_15720_n2324.n3 a_15720_n2324.t17 1.0925
R120 a_15720_n2324.n5 a_15720_n2324.t8 1.0925
R121 a_15720_n2324.n5 a_15720_n2324.t18 1.0925
R122 a_15720_n2324.n6 a_15720_n2324.t14 1.0925
R123 a_15720_n2324.n6 a_15720_n2324.t6 1.0925
R124 a_15720_n2324.n8 a_15720_n2324.t12 1.0925
R125 a_15720_n2324.n8 a_15720_n2324.t2 1.0925
R126 a_15720_n2324.n9 a_15720_n2324.t4 1.0925
R127 a_15720_n2324.n9 a_15720_n2324.t11 1.0925
R128 a_15720_n2324.t0 a_15720_n2324.n18 1.0925
R129 a_15720_n2324.n18 a_15720_n2324.t5 1.0925
R130 a_15720_n2324.n4 a_15720_n2324.n1 0.849071
R131 a_15720_n2324.n7 a_15720_n2324.n4 0.849071
R132 a_15720_n2324.n10 a_15720_n2324.n7 0.849071
R133 a_15720_n2324.n12 a_15720_n2324.n10 0.849071
R134 a_15720_n2324.n14 a_15720_n2324.n12 0.534875
R135 a_15720_n2324.n17 a_15720_n2324.n1 0.487625
R136 VSS.n9 VSS.n3 85644.1
R137 VSS.n19 VSS.n4 414.478
R138 VSS.n11 VSS.n9 220.377
R139 VSS.n17 VSS.n3 220.377
R140 VSS.n10 VSS.n5 205.139
R141 VSS.n18 VSS.n5 205.139
R142 VSS.n18 VSS.n6 205.139
R143 VSS.n10 VSS.n6 205.139
R144 VSS.n8 VSS.n7 167.988
R145 VSS.n21 VSS.n2 166.989
R146 VSS.t21 VSS.t0 123.174
R147 VSS.t1 VSS.t13 123.174
R148 VSS.t23 VSS.t5 123.174
R149 VSS.t22 VSS.t8 123.174
R150 VSS.t11 VSS.t17 123.174
R151 VSS.t2 VSS.t20 123.174
R152 VSS.t9 VSS.t16 123.174
R153 VSS.t15 VSS.t14 123.174
R154 VSS.n15 VSS.n14 118.222
R155 VSS.t12 VSS.t25 112.785
R156 VSS.t25 VSS.t10 112.785
R157 VSS.t13 VSS.t21 102.397
R158 VSS.t5 VSS.t1 102.397
R159 VSS.t8 VSS.t23 102.397
R160 VSS.t6 VSS.t22 102.397
R161 VSS.t17 VSS.t7 102.397
R162 VSS.t20 VSS.t11 102.397
R163 VSS.t16 VSS.t2 102.397
R164 VSS.t14 VSS.t9 102.397
R165 VSS.t0 VSS.n11 92.0096
R166 VSS.n13 VSS.t19 92.0096
R167 VSS.n16 VSS.t18 92.0096
R168 VSS.n17 VSS.t15 92.0096
R169 VSS.n7 VSS.n2 80.5005
R170 VSS.t19 VSS.t24 78.6535
R171 VSS.t3 VSS.t18 78.6535
R172 VSS.n13 VSS.t6 31.1649
R173 VSS.t7 VSS.n16 31.1649
R174 VSS.n12 VSS.n5 30.5283
R175 VSS.n12 VSS.n6 30.5283
R176 VSS.t24 VSS.t12 23.7448
R177 VSS.t10 VSS.t3 23.7448
R178 VSS.n15 VSS.n2 18.8616
R179 VSS.n14 VSS.n7 18.8616
R180 VSS.n1 VSS.n0 11.0305
R181 VSS.n10 VSS.n4 9.94004
R182 VSS.n19 VSS.n18 9.94004
R183 VSS.n15 VSS.n1 6.23383
R184 VSS VSS.n21 4.78577
R185 VSS.n0 VSS.t26 2.048
R186 VSS.n0 VSS.t4 2.048
R187 VSS.n16 VSS.n15 1.73383
R188 VSS.n14 VSS.n13 1.73383
R189 VSS.n8 VSS.n4 0.999917
R190 VSS.n20 VSS.n19 0.999917
R191 VSS.n21 VSS.n20 0.999917
R192 VSS.n11 VSS.n10 0.867167
R193 VSS.t25 VSS.n12 0.867167
R194 VSS.n18 VSS.n17 0.867167
R195 VSS VSS.n1 0.1605
R196 VSS.n9 VSS.n8 0.0215413
R197 VSS.n20 VSS.n3 0.0215413
R198 Vout2.t14 Vout2.t12 19.735
R199 Vout2.n5 Vout2.t14 18.9075
R200 Vout2.n12 Vout2.t8 16.9998
R201 Vout2.n2 Vout2.t10 13.6729
R202 Vout2.n3 Vout2.t11 13.3844
R203 Vout2.n2 Vout2.t15 13.3445
R204 Vout2.n4 Vout2.n1 12.247
R205 Vout2.n11 Vout2.n10 11.2403
R206 Vout2.n4 Vout2.n3 9.4181
R207 Vout2.n6 Vout2.n0 7.4449
R208 Vout2.n8 Vout2.n7 6.75194
R209 Vout2 Vout2.n12 6.32761
R210 Vout2.n9 Vout2.t9 5.04666
R211 Vout2.n6 Vout2.n5 4.94262
R212 Vout2.n9 Vout2.t13 4.84137
R213 Vout2.n11 Vout2.n8 2.836
R214 Vout2.n11 Vout2.n9 2.75432
R215 Vout2.n1 Vout2.t2 1.8205
R216 Vout2.n1 Vout2.t5 1.8205
R217 Vout2.n0 Vout2.t1 1.8205
R218 Vout2.n0 Vout2.t3 1.8205
R219 Vout2.n7 Vout2.t6 0.8195
R220 Vout2.n7 Vout2.t4 0.8195
R221 Vout2.n10 Vout2.t0 0.8195
R222 Vout2.n10 Vout2.t7 0.8195
R223 Vout2.n12 Vout2.n11 0.733357
R224 Vout2.n5 Vout2.n4 0.5315
R225 Vout2.n3 Vout2.n2 0.289009
R226 Vout2.n8 Vout2.n6 0.184462
R227 Vout1.t13 Vout1.t14 19.735
R228 Vout1.n2 Vout1.n0 18.0852
R229 Vout1.n12 Vout1.t8 16.9998
R230 Vout1.n5 Vout1.t13 14.5537
R231 Vout1.n5 Vout1.n4 14.2885
R232 Vout1.n3 Vout1.t9 13.6729
R233 Vout1.n4 Vout1.t10 13.3844
R234 Vout1.n3 Vout1.t12 13.3445
R235 Vout1.n11 Vout1.n10 11.24
R236 Vout1.n2 Vout1.n1 7.16477
R237 Vout1.n8 Vout1.n7 6.75194
R238 Vout1 Vout1.n12 6.32624
R239 Vout1.n9 Vout1.t15 5.04666
R240 Vout1.n9 Vout1.t11 4.84137
R241 Vout1.n11 Vout1.n8 2.836
R242 Vout1.n11 Vout1.n9 2.75432
R243 Vout1.n1 Vout1.t0 1.8205
R244 Vout1.n1 Vout1.t2 1.8205
R245 Vout1.n0 Vout1.t1 1.8205
R246 Vout1.n0 Vout1.t3 1.8205
R247 Vout1.n7 Vout1.t7 0.8195
R248 Vout1.n7 Vout1.t5 0.8195
R249 Vout1.n10 Vout1.t4 0.8195
R250 Vout1.n10 Vout1.t6 0.8195
R251 Vout1.n12 Vout1.n11 0.733357
R252 Vout1.n6 Vout1.n5 0.440894
R253 Vout1.n6 Vout1.n2 0.426875
R254 Vout1.n4 Vout1.n3 0.289009
R255 Vout1.n8 Vout1.n6 0.0607115
R256 Vp.n5 Vp.t16 19.5626
R257 Vp.n4 Vp.n2 11.9065
R258 Vp.n4 Vp.n3 11.2495
R259 Vp.n10 Vp.n9 11.243
R260 Vp.n16 Vp.n15 8.80104
R261 Vp.n12 Vp.n11 6.60725
R262 Vp.n8 Vp.n1 6.52262
R263 Vp.n14 Vp.n12 6.386
R264 Vp.n7 Vp.n5 5.44213
R265 Vp.n14 Vp.n13 4.36738
R266 Vp.n1 Vp.n0 4.36738
R267 Vp.n7 Vp.n6 4.3505
R268 Vp.n8 Vp.n7 2.2505
R269 Vp.n15 Vp.n1 2.14009
R270 Vp.n12 Vp.n10 1.50001
R271 Vp.n10 Vp.n8 1.49326
R272 Vp.n13 Vp.t2 1.0925
R273 Vp.n13 Vp.t10 1.0925
R274 Vp.n11 Vp.t11 1.0925
R275 Vp.n11 Vp.t8 1.0925
R276 Vp.n9 Vp.t14 1.0925
R277 Vp.n9 Vp.t15 1.0925
R278 Vp.n6 Vp.t9 1.0925
R279 Vp.n6 Vp.t7 1.0925
R280 Vp.n0 Vp.t13 1.0925
R281 Vp.n0 Vp.t1 1.0925
R282 Vp.t0 Vp.n16 1.0925
R283 Vp.n16 Vp.t12 1.0925
R284 Vp.n3 Vp.t6 0.8195
R285 Vp.n3 Vp.t3 0.8195
R286 Vp.n2 Vp.t5 0.8195
R287 Vp.n2 Vp.t4 0.8195
R288 Vp.n15 Vp.n14 0.314375
R289 Vp.n5 Vp.n4 0.16025
R290 Vin1.n5 Vin1.n4 23.1032
R291 Vin1.n1 Vin1.n0 23.1032
R292 Vin1.n8 Vin1.t3 21.8564
R293 Vin1.n4 Vin1.t0 16.3641
R294 Vin1.n0 Vin1.t6 16.3626
R295 Vin1.n4 Vin1.t7 16.0225
R296 Vin1.n0 Vin1.t1 16.021
R297 Vin1.n1 Vin1.t4 11.7992
R298 Vin1.n7 Vin1.t9 11.5195
R299 Vin1.n6 Vin1.t5 11.5195
R300 Vin1.n3 Vin1.t2 11.5195
R301 Vin1.n2 Vin1.t8 11.5195
R302 Vin1.n7 Vin1.n6 4.00673
R303 Vin1.n2 Vin1.n1 3.16619
R304 Vin1.n8 Vin1.n7 0.673591
R305 Vin1.n6 Vin1.n5 0.650658
R306 Vin1 Vin1.n8 0.5405
R307 Vin1.n5 Vin1.n3 0.279681
R308 Vin1.n3 Vin1.n2 0.231705
.ends

