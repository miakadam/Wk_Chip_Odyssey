magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 541 -23 587
rect 23 541 34 552
rect -103 430 -57 506
rect 57 430 103 506
rect -34 349 -23 395
rect -34 229 -23 275
rect 23 229 34 240
rect -103 118 -57 194
rect 57 118 103 194
rect -34 37 -23 83
rect -34 -83 -23 -37
rect 23 -83 34 -72
rect -103 -194 -57 -118
rect 57 -194 103 -118
rect -34 -275 -23 -229
rect -34 -395 -23 -349
rect 23 -395 34 -384
rect -103 -506 -57 -430
rect 57 -506 103 -430
rect -34 -587 -23 -541
<< nwell >>
rect -278 -718 278 718
<< pmos >>
rect -28 428 28 508
rect -28 116 28 196
rect -28 -196 28 -116
rect -28 -508 28 -428
<< pdiff >>
rect -116 495 -28 508
rect -116 441 -103 495
rect -57 441 -28 495
rect -116 428 -28 441
rect 28 495 116 508
rect 28 441 57 495
rect 103 441 116 495
rect 28 428 116 441
rect -116 183 -28 196
rect -116 129 -103 183
rect -57 129 -28 183
rect -116 116 -28 129
rect 28 183 116 196
rect 28 129 57 183
rect 103 129 116 183
rect 28 116 116 129
rect -116 -129 -28 -116
rect -116 -183 -103 -129
rect -57 -183 -28 -129
rect -116 -196 -28 -183
rect 28 -129 116 -116
rect 28 -183 57 -129
rect 103 -183 116 -129
rect 28 -196 116 -183
rect -116 -441 -28 -428
rect -116 -495 -103 -441
rect -57 -495 -28 -441
rect -116 -508 -28 -495
rect 28 -441 116 -428
rect 28 -495 57 -441
rect 103 -495 116 -441
rect 28 -508 116 -495
<< pdiffc >>
rect -103 441 -57 495
rect 57 441 103 495
rect -103 129 -57 183
rect 57 129 103 183
rect -103 -183 -57 -129
rect 57 -183 103 -129
rect -103 -495 -57 -441
rect 57 -495 103 -441
<< nsubdiff >>
rect -254 622 254 694
rect -254 578 -182 622
rect -254 -578 -241 578
rect -195 -578 -182 578
rect 182 578 254 622
rect -254 -622 -182 -578
rect 182 -578 195 578
rect 241 -578 254 578
rect 182 -622 254 -578
rect -254 -694 254 -622
<< nsubdiffcont >>
rect -241 -578 -195 578
rect 195 -578 241 578
<< polysilicon >>
rect -36 587 36 600
rect -36 541 -23 587
rect 23 541 36 587
rect -36 528 36 541
rect -28 508 28 528
rect -28 408 28 428
rect -36 395 36 408
rect -36 349 -23 395
rect 23 349 36 395
rect -36 336 36 349
rect -36 275 36 288
rect -36 229 -23 275
rect 23 229 36 275
rect -36 216 36 229
rect -28 196 28 216
rect -28 96 28 116
rect -36 83 36 96
rect -36 37 -23 83
rect 23 37 36 83
rect -36 24 36 37
rect -36 -37 36 -24
rect -36 -83 -23 -37
rect 23 -83 36 -37
rect -36 -96 36 -83
rect -28 -116 28 -96
rect -28 -216 28 -196
rect -36 -229 36 -216
rect -36 -275 -23 -229
rect 23 -275 36 -229
rect -36 -288 36 -275
rect -36 -349 36 -336
rect -36 -395 -23 -349
rect 23 -395 36 -349
rect -36 -408 36 -395
rect -28 -428 28 -408
rect -28 -528 28 -508
rect -36 -541 36 -528
rect -36 -587 -23 -541
rect 23 -587 36 -541
rect -36 -600 36 -587
<< polycontact >>
rect -23 541 23 587
rect -23 349 23 395
rect -23 229 23 275
rect -23 37 23 83
rect -23 -83 23 -37
rect -23 -275 23 -229
rect -23 -395 23 -349
rect -23 -587 23 -541
<< metal1 >>
rect -241 635 241 681
rect -241 578 -195 635
rect -34 541 -23 587
rect 23 541 34 587
rect 195 578 241 635
rect -103 495 -57 506
rect -103 430 -57 441
rect 57 495 103 506
rect 57 430 103 441
rect -34 349 -23 395
rect 23 349 34 395
rect -34 229 -23 275
rect 23 229 34 275
rect -103 183 -57 194
rect -103 118 -57 129
rect 57 183 103 194
rect 57 118 103 129
rect -34 37 -23 83
rect 23 37 34 83
rect -34 -83 -23 -37
rect 23 -83 34 -37
rect -103 -129 -57 -118
rect -103 -194 -57 -183
rect 57 -129 103 -118
rect 57 -194 103 -183
rect -34 -275 -23 -229
rect 23 -275 34 -229
rect -34 -395 -23 -349
rect 23 -395 34 -349
rect -103 -441 -57 -430
rect -103 -506 -57 -495
rect 57 -441 103 -430
rect 57 -506 103 -495
rect -241 -635 -195 -578
rect -34 -587 -23 -541
rect 23 -587 34 -541
rect 195 -635 241 -578
rect -241 -681 241 -635
<< properties >>
string FIXED_BBOX -218 -658 218 658
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.4 l 0.28 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
