* NGSPICE file created from diffpairtest.ext - technology: gf180mcuD

.subckt nfet_03v3_RPTYYZ a_708_n150# a_n708_n242# a_404_n150# a_n404_n242# a_n796_n150#
+ a_100_n150# a_n100_n242# a_n508_n150# a_n204_n150# a_2580_n1506# a_508_n242# a_204_n242#
X0 a_n204_n150# a_n404_n242# a_n508_n150# a_2580_n1506# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X1 a_n508_n150# a_n708_n242# a_n796_n150# a_2580_n1506# nfet_03v3 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=1u
X2 a_404_n150# a_204_n242# a_100_n150# a_2580_n1506# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X3 a_100_n150# a_n100_n242# a_n204_n150# a_2580_n1506# nfet_03v3 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=1u
X4 a_708_n150# a_508_n242# a_404_n150# a_2580_n1506# nfet_03v3 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=1u
.ends

.subckt diffpairtest Vin1 VSS Vd1 Vd2 Vin2
XXM9 VSS Vin1 Vd1 m1_10425_2575# Vd1 VSS m1_10425_2575# VSS Vd2 VSS Vin1 Vin1 nfet_03v3_RPTYYZ
XXM20 VSS Vin2 Vd2 a_10430_3135# Vd2 VSS a_10430_3135# VSS Vd1 VSS Vin2 Vin2 nfet_03v3_RPTYYZ
Xnfet_03v3_RPTYYZ_0 Vd1 m1_11640_3135# VSS m1_11640_3135# VSS Vd2 Vin2 Vd1 VSS VSS
+ Vin1 Vin2 nfet_03v3_RPTYYZ
XXM10 Vd2 m1_11640_2575# VSS m1_11640_2575# VSS Vd1 Vin1 Vd2 VSS VSS Vin2 Vin1 nfet_03v3_RPTYYZ
.ends

