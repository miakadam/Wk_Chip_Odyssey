magic
tech gf180mcuD
magscale 1 10
timestamp 1757548363
<< error_s >>
rect 5586 -435 5592 -389
rect 5594 -464 5638 -435
rect 5463 -664 5526 -654
rect 5400 -1020 5417 -1018
rect 5542 -1314 5630 -1272
rect 5710 -1314 5798 -1272
rect 5391 -1560 5418 -1346
rect 5570 -1372 5770 -1328
rect 5476 -1380 5838 -1372
rect 5476 -1400 5604 -1380
rect 5610 -1400 5838 -1380
rect 5630 -1406 5710 -1400
rect 5584 -1448 5704 -1428
rect 5544 -1458 5744 -1448
rect 5460 -1500 5828 -1458
rect 5378 -1704 5386 -1672
rect 4988 -1864 5026 -1835
rect 5378 -2500 5934 -1704
rect 5380 -2524 5934 -2500
<< metal1 >>
rect 5208 232 5658 284
rect 5216 224 5658 232
rect 5316 0 5376 224
rect 5400 -1020 5480 -700
rect 5528 -756 5592 156
rect 5528 -1252 5596 -756
rect 5324 -1560 5372 -1392
rect 5532 -1472 5596 -1252
rect 5280 -1564 5610 -1560
rect 5208 -1624 5658 -1564
use nfet_03v3_Q7US5R  XM3
timestamp 1757548363
transform 1 0 5440 0 1 -1264
box -60 -1260 520 200
use pfet_03v3_YXHA8C  XM4
timestamp 1757548363
transform 1 0 5440 0 1 -264
box -60 -1260 520 200
use nfet_03v3_Q7US5R  XXM3
timestamp 1757548363
transform 1 0 4834 0 1 -1264
box -60 -1260 520 200
use pfet_03v3_YXHA8C  XXM4
timestamp 1757548363
transform 1 0 5414 0 1 -1264
box -60 -1260 520 200
<< labels >>
rlabel metal1 5208 252 5208 252 7 avdd
port 0 w
rlabel metal1 5212 -1604 5212 -1604 7 avss
port 1 w
rlabel metal1 5412 -876 5412 -876 7 in
port 2 w
rlabel metal1 5564 -872 5564 -872 7 out
port 3 w
<< end >>
