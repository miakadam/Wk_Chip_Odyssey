* NGSPICE file created from v2comp_SAR_final.ext - technology: (null)

.subckt comp_SAR_final Vdd Vss Clk Vin1 Vin2 Comp_out Reset SAR_in Clk_piso Load Piso_out
X0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t0 Clk.t0 Vdd.t19 Vdd.t18 pfet_03v3
**devattr s=14080,496 d=14080,496
X1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t38 nfet_03v3
**devattr s=20800,504 d=20800,504
X2 a_n9429_n3007.t18 Vin1.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t11 Vss.t39 nfet_03v3
**devattr s=15600,404 d=15600,404
X3 Vdd.t11 a_n10831_3320 Comp_out.t7 Vdd.t10 pfet_03v3
**devattr s=18700,450 d=18700,450
X4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t4 Vss.t23 nfet_03v3
**devattr s=20800,504 d=20800,504
X5 a_n9429_n3007.t21 Vin2.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t29 nfet_03v3
**devattr s=15600,404 d=15600,404
X6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t1 a_n9429_n3007.t2 Vss.t24 nfet_03v3
**devattr s=15600,404 d=15600,404
X7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq a_n9933_n3099 a_n10021_n3007 Vss.t3 nfet_03v3
**devattr s=26400,776 d=15600,404
X8 Vdd.t45 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t7 Vdd.t44 pfet_03v3
**devattr s=10400,304 d=10400,304
X9 a_n9429_n3007.t3 Vin2.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t25 nfet_03v3
**devattr s=15600,404 d=15600,404
X10 a_n8351_n659 a_n8551_n751 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t1 Vss.t14 nfet_03v3
**devattr s=20800,504 d=35200,976
X11 a_n9429_n3007.t7 Vin2.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t39 nfet_03v3
**devattr s=15600,404 d=15600,404
X12 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t41 Vdd.t40 pfet_03v3
**devattr s=17600,576 d=17600,576
X13 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x3.out Vss.t33 Vss.t32 nfet_03v3
**devattr s=17600,576 d=17600,576
X14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t2 Vss.t37 nfet_03v3
**devattr s=20800,504 d=20800,504
X15 Comp_out.t3 a_n10831_3320 Vss.t11 Vss.t10 nfet_03v3
**devattr s=17000,540 d=9350,280
X16 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t12 Vss.t36 Vss.t35 nfet_03v3
**devattr s=35200,976 d=35200,976
X17 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t10 Vdd.t39 Vdd.t38 pfet_03v3
**devattr s=10400,304 d=10400,304
X18 Vdd.t33 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t5 Vdd.t32 pfet_03v3
**devattr s=10400,304 d=10400,304
X19 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t9 Vin1.t1 a_n9429_n3007.t17 Vss.t24 nfet_03v3
**devattr s=15600,404 d=15600,404
X20 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t12 Vdd.t29 Vdd.t28 pfet_03v3
**devattr s=10400,304 d=10400,304
X21 Vdd.t17 Clk.t1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vdd.t16 pfet_03v3
**devattr s=14080,496 d=14080,496
X22 a_n6389_n2044 a_n6589_n2136 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t41 nfet_03v3
**devattr s=15600,404 d=26400,776
X23 a_n10831_3320 comparator_no_offsetcal_0.x4.A Vss.t16 Vss.t15 nfet_03v3
**devattr s=9350,280 d=17000,540
X24 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t10 Vin1.t2 a_n9429_n3007.t16 Vss.t26 nfet_03v3
**devattr s=15600,404 d=15600,404
X25 a_n9429_n3007.t15 Vin1.t3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t7 Vss.t25 nfet_03v3
**devattr s=15600,404 d=15600,404
X26 Vdd.t15 Clk.t2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t0 Vdd.t14 pfet_03v3
**devattr s=14080,496 d=14080,496
X27 Vss.t22 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t13 comparator_no_offsetcal_0.x5.out Vss.t21 nfet_03v3
**devattr s=35200,976 d=35200,976
X28 Vdd.t3 a_n9629_405 a_n9717_497 Vdd.t2 pfet_03v3
**devattr s=17600,576 d=10400,304
X29 Comp_out.t6 a_n10831_3320 Vdd.t9 Vdd.t8 pfet_03v3
**devattr s=34000,880 d=18700,450
X30 Comp_out.t2 a_n10831_3320 Vss.t9 Vss.t8 nfet_03v3
**devattr s=9350,280 d=9350,280
X31 Vdd.t21 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t2 Vdd.t20 pfet_03v3
**devattr s=10400,304 d=10400,304
X32 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t13 Vss.t20 nfet_03v3
**devattr s=20800,504 d=20800,504
X33 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t1 Vss.t34 nfet_03v3
**devattr s=20800,504 d=20800,504
X34 a_n6389_n3007 a_n6589_n3099 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t12 Vss.t41 nfet_03v3
**devattr s=15600,404 d=26400,776
X35 a_n10831_3320 comparator_no_offsetcal_0.x4.A Vdd.t25 Vdd.t24 pfet_03v3
**devattr s=18700,450 d=34000,880
X36 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t6 Vss.t19 nfet_03v3
**devattr s=20800,504 d=20800,504
X37 a_n9429_n3007.t8 Vin2.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t42 nfet_03v3
**devattr s=15600,404 d=15600,404
X38 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t5 a_n9429_n3007.t19 Vss.t17 nfet_03v3
**devattr s=15600,404 d=15600,404
X39 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t6 a_n9429_n3007.t20 Vss.t18 nfet_03v3
**devattr s=15600,404 d=15600,404
X40 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t7 a_n9429_n3007.t4 Vss.t26 nfet_03v3
**devattr s=15600,404 d=15600,404
X41 Vss.t44 a_n8385_n3885 a_n8473_n3793 Vss.t43 nfet_03v3
**devattr s=14080,496 d=8320,264
X42 Comp_out.t5 a_n10831_3320 Vdd.t7 Vdd.t6 pfet_03v3
**devattr s=18700,450 d=18700,450
X43 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t14 Vdd.t43 Vdd.t42 pfet_03v3
**devattr s=10400,304 d=10400,304
X44 a_n9429_n3007.t14 Vin1.t4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t8 Vss.t27 nfet_03v3
**devattr s=15600,404 d=15600,404
X45 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t14 Vin1.t5 a_n9429_n3007.t13 Vss.t28 nfet_03v3
**devattr s=15600,404 d=15600,404
X46 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t0 Clk.t3 Vdd.t13 Vdd.t12 pfet_03v3
**devattr s=14080,496 d=14080,496
X47 comparator_no_offsetcal_0.x3.out comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t15 Vdd.t35 Vdd.t34 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X48 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t16 Vdd.t37 Vdd.t36 pfet_03v3
**devattr s=10400,304 d=10400,304
X49 a_n6693_497 a_n6893_405 Vdd.t1 Vdd.t0 pfet_03v3
**devattr s=10400,304 d=17600,576
X50 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t8 a_n7971_n751 a_n8059_n659 Vss.t40 nfet_03v3
**devattr s=35200,976 d=20800,504
X51 a_n9429_n3007.t12 Vin1.t6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t15 Vss.t42 nfet_03v3
**devattr s=15600,404 d=15600,404
X52 Vss.t7 a_n10831_3320 Comp_out.t1 Vss.t6 nfet_03v3
**devattr s=9350,280 d=9350,280
X53 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t1 Vin1.t7 a_n9429_n3007.t11 Vss.t17 nfet_03v3
**devattr s=15600,404 d=15600,404
X54 Vdd.t31 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t17 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t4 Vdd.t30 pfet_03v3
**devattr s=10400,304 d=10400,304
X55 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t5 a_n9767_n751 a_n9855_n659 Vss.t30 nfet_03v3
**devattr s=35200,976 d=20800,504
X56 a_n9429_n3007.t5 Vin2.t8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t27 nfet_03v3
**devattr s=15600,404 d=15600,404
X57 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t2 Vin1.t8 a_n9429_n3007.t10 Vss.t18 nfet_03v3
**devattr s=15600,404 d=15600,404
X58 a_n9429_n3007.t1 Clk.t4 Vss.t13 Vss.t12 nfet_03v3
**devattr s=8320,264 d=8320,264
X59 Vdd.t27 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t17 comparator_no_offsetcal_0.x5.out Vdd.t26 pfet_03v3
**devattr s=70400,1776 d=70400,1776
X60 a_n9429_n3007.t9 Vin1.t9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t4 Vss.t29 nfet_03v3
**devattr s=15600,404 d=15600,404
X61 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vin2.t9 a_n9429_n3007.t6 Vss.t28 nfet_03v3
**devattr s=15600,404 d=15600,404
X62 Vss.t5 a_n10831_3320 Comp_out.t0 Vss.t4 nfet_03v3
**devattr s=9350,280 d=9350,280
X63 Vdd.t23 comparator_no_offsetcal_0.x4.A comparator_no_offsetcal_0.x2.Vout2 Vdd.t22 pfet_03v3
**devattr s=17600,576 d=17600,576
X64 a_n6555_n659 a_n6755_n751 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vq Vss.t31 nfet_03v3
**devattr s=20800,504 d=35200,976
X65 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t16 a_n9933_n2136 a_n10021_n2044 Vss.t3 nfet_03v3
**devattr s=26400,776 d=15600,404
X66 Vss.t1 comparator_no_offsetcal_0.x5.out comparator_no_offsetcal_0.x2.Vout2 Vss.t0 nfet_03v3
**devattr s=17600,576 d=17600,576
X67 Vdd.t5 a_n10831_3320 Comp_out.t4 Vdd.t4 pfet_03v3
**devattr s=18700,450 d=18700,450
X68 a_n7937_n3793 a_n8017_n3885 a_n9429_n3007.t0 Vss.t2 nfet_03v3
**devattr s=8320,264 d=14080,496
R0 Clk.n4 Clk.t0 21.1483
R1 Clk.n3 Clk.t3 21.1483
R2 Clk.n2 Clk.t2 21.1483
R3 Clk.n1 Clk.t1 21.1483
R4 Clk.n0 Clk.t4 20.5929
R5 Clk.n1 Clk.n0 19.1491
R6 Clk.n5 Clk.n4 15.5861
R7 comparator_no_offsetcal_0.CLK Clk 5.90242
R8 Clk.n3 Clk.n2 4.47208
R9 Clk.n5 Clk.n0 3.56405
R10 comparator_no_offsetcal_0.CLK Clk.n5 1.32418
R11 Clk.n2 Clk.n1 1.01892
R12 Clk.n4 Clk.n3 1.01892
R13 Vdd.n14 Vdd.t34 869.717
R14 Vdd.n24 Vdd.t26 869.717
R15 Vdd.t0 Vdd.t32 490.324
R16 Vdd.t32 Vdd.t28 490.324
R17 Vdd.t28 Vdd.t44 490.324
R18 Vdd.t44 Vdd.t36 490.324
R19 Vdd.t36 Vdd.t20 490.324
R20 Vdd.t20 Vdd.t38 490.324
R21 Vdd.t38 Vdd.t30 490.324
R22 Vdd.t30 Vdd.t42 490.324
R23 Vdd.t42 Vdd.t2 490.324
R24 Vdd.n51 Vdd.t0 467.743
R25 Vdd.t2 Vdd.n49 467.743
R26 Vdd.n44 Vdd.t12 398.652
R27 Vdd.n52 Vdd.t14 398.652
R28 Vdd.n49 Vdd.t12 389.878
R29 Vdd.t14 Vdd.n51 389.878
R30 Vdd.t22 Vdd.n18 372.543
R31 Vdd.n21 Vdd.t40 372.543
R32 Vdd.n20 Vdd.t22 370.969
R33 Vdd.t40 Vdd.n20 370.969
R34 Vdd.n29 Vdd.n27 287.351
R35 Vdd.n30 Vdd.n28 287.351
R36 Vdd.t6 Vdd.t4 265.625
R37 Vdd.n7 Vdd.t24 242.189
R38 Vdd.t10 Vdd.n9 195.312
R39 Vdd.n42 Vdd.t18 190.464
R40 Vdd.n55 Vdd.t16 190.464
R41 Vdd.n10 Vdd.t10 179.689
R42 Vdd.t24 Vdd.n6 145.413
R43 Vdd.n10 Vdd.t6 85.938
R44 Vdd.n9 Vdd.t8 70.313
R45 Vdd.n18 Vdd.n16 58.9755
R46 Vdd.n21 Vdd.n16 58.9755
R47 Vdd.n21 Vdd.n17 58.9755
R48 Vdd.n18 Vdd.n17 58.9755
R49 Vdd.n44 Vdd.n29 54.0755
R50 Vdd.n52 Vdd.n27 54.0755
R51 Vdd.n52 Vdd.n28 54.0755
R52 Vdd.n44 Vdd.n30 54.0755
R53 Vdd.n43 Vdd.n42 29.3622
R54 Vdd.n56 Vdd.n55 29.3622
R55 Vdd.t4 Vdd.n7 23.438
R56 Vdd.n50 Vdd.n27 20.1255
R57 Vdd.n50 Vdd.n28 20.1255
R58 Vdd.n48 Vdd.n29 20.1255
R59 Vdd.n48 Vdd.n30 20.1255
R60 Vdd.n42 Vdd.n41 19.9167
R61 Vdd.n55 Vdd.n25 19.9167
R62 Vdd.n19 Vdd.n16 18.7255
R63 Vdd.n19 Vdd.n17 18.7255
R64 Vdd.n63 Vdd.n0 14.6602
R65 Vdd.n58 Vdd.n57 13.4987
R66 Vdd.n7 Vdd.n1 12.6005
R67 Vdd.n11 Vdd.n10 12.6005
R68 Vdd.n9 Vdd.n8 12.6005
R69 Vdd.n32 Vdd.n31 12.136
R70 Vdd.n34 Vdd.n33 12.136
R71 Vdd.n36 Vdd.n35 12.136
R72 Vdd.n38 Vdd.n37 12.136
R73 Vdd.n40 Vdd.n39 12.136
R74 Vdd.n48 Vdd.n47 11.111
R75 Vdd.n50 Vdd.n26 11.111
R76 Vdd.n57 Vdd.n25 9.86945
R77 Vdd.n54 Vdd.n53 9.536
R78 Vdd.n46 Vdd.n45 9.536
R79 Vdd.n41 Vdd.n0 9.536
R80 Vdd.n53 Vdd.t15 7.4755
R81 Vdd.n45 Vdd.t13 7.4755
R82 Vdd.n41 Vdd.t19 7.4755
R83 Vdd.n25 Vdd.t17 7.4755
R84 Vdd.n58 Vdd 5.27311
R85 Vdd.n22 Vdd.t41 4.4205
R86 Vdd.n15 Vdd.t23 4.4205
R87 Vdd.n8 Vdd.t9 3.38176
R88 Vdd.n53 Vdd.n52 2.1905
R89 Vdd.n45 Vdd.n44 2.1905
R90 Vdd.n3 Vdd.n2 2.16583
R91 Vdd.n5 Vdd.n4 2.16583
R92 Vdd.n24 Vdd.t27 1.99236
R93 Vdd.n13 Vdd.t35 1.91107
R94 Vdd.n61 Vdd.n14 1.83762
R95 Vdd.n59 Vdd.n24 1.83762
R96 Vdd.n31 Vdd.t1 1.8205
R97 Vdd.n31 Vdd.t33 1.8205
R98 Vdd.n33 Vdd.t29 1.8205
R99 Vdd.n33 Vdd.t45 1.8205
R100 Vdd.n35 Vdd.t37 1.8205
R101 Vdd.n35 Vdd.t21 1.8205
R102 Vdd.n37 Vdd.t39 1.8205
R103 Vdd.n37 Vdd.t31 1.8205
R104 Vdd.n39 Vdd.t43 1.8205
R105 Vdd.n39 Vdd.t3 1.8205
R106 Vdd.n20 Vdd.n19 1.5755
R107 Vdd.n22 Vdd.n21 1.5755
R108 Vdd.n18 Vdd.n15 1.5755
R109 Vdd.n51 Vdd.n50 1.5755
R110 Vdd.n49 Vdd.n48 1.5755
R111 Vdd.n2 Vdd.t7 1.13285
R112 Vdd.n2 Vdd.t11 1.13285
R113 Vdd.n4 Vdd.t25 1.13285
R114 Vdd.n4 Vdd.t5 1.13285
R115 Vdd.n60 Vdd.n23 1.058
R116 Vdd.n23 Vdd.n15 1.01373
R117 Vdd.n23 Vdd.n22 0.979984
R118 Vdd.n62 Vdd.n12 0.750875
R119 Vdd.n40 Vdd.n38 0.667
R120 Vdd.n34 Vdd.n32 0.662
R121 Vdd.n38 Vdd.n36 0.643429
R122 Vdd.n36 Vdd.n34 0.638429
R123 Vdd.n46 Vdd.n43 0.58325
R124 Vdd.n56 Vdd.n54 0.58325
R125 Vdd.n47 Vdd.n40 0.47525
R126 Vdd.n32 Vdd.n26 0.47525
R127 Vdd.n63 Vdd.n62 0.381816
R128 Vdd.n43 Vdd.n0 0.34025
R129 Vdd.n47 Vdd.n46 0.34025
R130 Vdd.n54 Vdd.n26 0.34025
R131 Vdd.n59 Vdd.n58 0.313132
R132 Vdd.n60 Vdd.n59 0.289447
R133 Vdd.n61 Vdd.n60 0.279974
R134 Vdd.n62 Vdd.n61 0.256289
R135 Vdd.n13 comparator_no_offsetcal_0.x3.avdd 0.207699
R136 Vdd.n8 Vdd.n3 0.1355
R137 Vdd.n6 Vdd.n5 0.109786
R138 Vdd.n12 Vdd.n1 0.103357
R139 Vdd.n14 Vdd.n13 0.0965492
R140 comparator_no_offsetcal_0.VDD Vdd.n63 0.0942895
R141 Vdd.n12 Vdd.n11 0.0519286
R142 Vdd.n5 Vdd.n1 0.0455
R143 Vdd.n11 Vdd.n3 0.0197857
R144 Vdd.n57 Vdd.n56 0.0068
R145 Vdd.n6 comparator_no_offsetcal_0.x4.VDD 0.00371429
R146 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 19.5626
R147 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 11.9065
R148 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 11.2495
R149 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 11.243
R150 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 8.80104
R151 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 6.60725
R152 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 6.52262
R153 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 6.386
R154 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 5.44213
R155 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 4.36738
R156 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 4.36738
R157 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 4.3505
R158 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n15 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 2.2505
R159 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 2.14009
R160 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 1.50001
R161 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n4 1.49326
R162 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t8 1.0925
R163 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t16 1.0925
R164 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t15 1.0925
R165 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t9 1.0925
R166 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t12 1.0925
R167 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t2 1.0925
R168 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t7 1.0925
R169 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t1 1.0925
R170 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t11 1.0925
R171 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t14 1.0925
R172 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t4 1.0925
R173 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t10 1.0925
R174 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t6 0.8195
R175 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t5 0.8195
R176 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t13 0.8195
R177 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.t3 0.8195
R178 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n9 0.314375
R179 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vp.n2 0.16025
R180 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t15 49.7997
R181 comparator_no_offsetcal_0.x3.in comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t12 31.5367
R182 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t16 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t10 19.735
R183 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 18.0852
R184 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t0 16.9998
R185 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t16 14.5537
R186 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 14.2885
R187 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t13 13.6729
R188 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t11 13.3844
R189 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t9 13.3445
R190 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 11.24
R191 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 7.16477
R192 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 6.95627
R193 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 6.75194
R194 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 6.32624
R195 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t17 5.04666
R196 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t14 4.84137
R197 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 2.836
R198 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n10 2.75432
R199 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t2 1.8205
R200 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t7 1.8205
R201 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t5 1.8205
R202 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t3 1.8205
R203 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t1 0.8195
R204 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t8 0.8195
R205 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t4 0.8195
R206 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.t6 0.8195
R207 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n12 0.733357
R208 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n6 0.440894
R209 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n3 0.426875
R210 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n4 0.289009
R211 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n7 0.0607115
R212 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout1.n0 comparator_no_offsetcal_0.x3.in 0.014
R213 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t17 49.7997
R214 comparator_no_offsetcal_0.x5.in comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t13 31.5367
R215 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t14 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t10 19.735
R216 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t14 18.9075
R217 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t0 16.9998
R218 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t16 13.6729
R219 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t15 13.3844
R220 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t9 13.3445
R221 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 12.247
R222 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 11.2403
R223 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 9.4181
R224 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 7.4449
R225 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 6.95074
R226 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 6.75194
R227 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 6.32761
R228 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t12 5.04666
R229 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 4.94262
R230 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t11 4.84137
R231 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 2.836
R232 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n10 2.75432
R233 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t4 1.8205
R234 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n2 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t6 1.8205
R235 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t7 1.8205
R236 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n1 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t5 1.8205
R237 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t2 0.8195
R238 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n8 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t8 0.8195
R239 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t1 0.8195
R240 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n11 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.t3 0.8195
R241 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n13 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n12 0.733357
R242 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n6 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n5 0.5315
R243 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n4 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n3 0.289009
R244 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n9 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n7 0.184462
R245 comparator_no_offsetcal_0.lvsclean_SAlatch_0.Vout2.n0 comparator_no_offsetcal_0.x5.in 0.014
R246 Vss.n36 Vss.n35 259245
R247 Vss.n59 Vss.n58 148254
R248 Vss.n34 Vss.n33 59530.8
R249 Vss.n63 Vss.n4 25794.4
R250 Vss.n59 Vss.n4 23334.9
R251 Vss.n35 Vss.n34 18659
R252 Vss.n63 Vss.t15 10202.1
R253 Vss.n64 Vss.n63 5567.73
R254 Vss.n35 Vss.n19 2358.54
R255 Vss.n65 Vss.t35 1596.98
R256 Vss.n36 Vss.t21 1596.98
R257 Vss.t10 Vss.n59 1095.73
R258 Vss.n34 Vss.n4 924.742
R259 Vss.n65 Vss.n2 478.125
R260 Vss.n56 Vss.n15 414.478
R261 Vss.n33 Vss.n32 325
R262 Vss.n64 Vss.n3 325
R263 Vss.n32 Vss.t0 293.137
R264 Vss.n24 Vss.t0 293.137
R265 Vss.n24 Vss.t32 293.137
R266 Vss.t32 Vss.n3 293.137
R267 Vss.n36 Vss.n33 248.53
R268 Vss.n65 Vss.n64 248.53
R269 Vss.n52 Vss.n16 205.139
R270 Vss.n54 Vss.n16 205.139
R271 Vss.n54 Vss.n53 205.139
R272 Vss.n53 Vss.n52 205.139
R273 Vss.n58 Vss.n13 193.476
R274 Vss.n51 Vss.n19 192.703
R275 Vss.t6 Vss.t8 191.642
R276 Vss.t15 Vss.n62 174.732
R277 Vss.n42 Vss.n20 166.989
R278 Vss.n21 Vss.n14 166.989
R279 Vss.t4 Vss.n60 140.913
R280 Vss.n61 Vss.t4 129.641
R281 Vss.n49 Vss.n48 118.222
R282 Vss.t41 Vss.t31 108.138
R283 Vss.t18 Vss.t34 108.138
R284 Vss.t39 Vss.t38 108.138
R285 Vss.t28 Vss.t37 108.138
R286 Vss.t20 Vss.t42 108.138
R287 Vss.t23 Vss.t24 108.138
R288 Vss.t19 Vss.t27 108.138
R289 Vss.t30 Vss.t3 108.138
R290 Vss.t15 Vss.n2 105.561
R291 Vss.t12 Vss.t17 99.0183
R292 Vss.t29 Vss.t12 99.0183
R293 Vss.n66 Vss.n65 98.7258
R294 Vss.n37 Vss.n36 98.7258
R295 Vss.t31 Vss.t18 89.8983
R296 Vss.t34 Vss.t39 89.8983
R297 Vss.t38 Vss.t28 89.8983
R298 Vss.t37 Vss.t25 89.8983
R299 Vss.t26 Vss.t20 89.8983
R300 Vss.t42 Vss.t23 89.8983
R301 Vss.t24 Vss.t19 89.8983
R302 Vss.t27 Vss.t30 89.8983
R303 Vss.n50 Vss.t40 80.7782
R304 Vss.n47 Vss.t14 80.7782
R305 Vss.t3 Vss.n13 80.7782
R306 Vss.n21 Vss.n20 80.5005
R307 Vss.t2 Vss.t40 69.0524
R308 Vss.t14 Vss.t43 69.0524
R309 Vss.n51 Vss.t41 65.5624
R310 Vss.n31 Vss.n23 65.5283
R311 Vss.n27 Vss.n23 65.5283
R312 Vss.n27 Vss.n26 65.5283
R313 Vss.n31 Vss.n26 65.5283
R314 Vss.t8 Vss.n61 62.0024
R315 Vss.n60 Vss.t10 50.7294
R316 Vss.n17 Vss.n16 30.5283
R317 Vss.n53 Vss.n17 30.5283
R318 Vss.t25 Vss.n50 27.3607
R319 Vss.n47 Vss.t26 27.3607
R320 Vss.t17 Vss.t2 20.8464
R321 Vss.t43 Vss.t29 20.8464
R322 Vss.n25 Vss.n23 20.8061
R323 Vss.n26 Vss.n25 20.8061
R324 Vss.n48 Vss.n21 18.8616
R325 Vss.n49 Vss.n20 18.8616
R326 Vss.n68 comparator_no_offsetcal_0.x3.avss 17.8218
R327 Vss.n62 Vss.t6 16.9105
R328 Vss.n39 comparator_no_offsetcal_0.x5.avss 16.7565
R329 Vss.n61 Vss.n9 14.6641
R330 Vss.n60 Vss.n12 14.1923
R331 Vss.n62 Vss.n8 11.9681
R332 Vss.n46 Vss.n22 11.0305
R333 Vss.n6 Vss.n2 10.4005
R334 Vss.n39 Vss 9.06952
R335 Vss.n12 Vss.t11 8.70131
R336 Vss.n55 Vss.n0 7.7564
R337 Vss.n40 Vss.n18 7.59387
R338 Vss.n43 Vss.n42 6.65104
R339 Vss.n7 Vss.n5 6.5795
R340 Vss.n11 Vss.n10 6.5795
R341 Vss.n55 Vss.n54 6.33584
R342 Vss.n52 Vss.n18 6.32806
R343 Vss.n48 Vss.n46 6.23383
R344 Vss.n30 Vss.t1 4.7885
R345 Vss.n28 Vss.t33 4.7885
R346 Vss.n45 Vss.n14 3.8722
R347 Vss.n18 Vss.n15 3.52248
R348 Vss.n56 Vss.n55 3.51469
R349 Vss.n67 Vss.t36 2.9111
R350 Vss.n38 Vss.t22 2.9111
R351 Vss.n22 Vss.t13 2.048
R352 Vss.n22 Vss.t44 2.048
R353 Vss.n5 Vss.t16 2.03874
R354 Vss.n5 Vss.t7 2.03874
R355 Vss.n10 Vss.t9 2.03874
R356 Vss.n10 Vss.t5 2.03874
R357 Vss.n48 Vss.n47 1.73383
R358 Vss.n50 Vss.n49 1.73383
R359 Vss.n37 Vss.n1 1.70279
R360 Vss.n66 Vss.n1 1.62925
R361 Vss.n31 Vss.n30 1.3005
R362 Vss.n32 Vss.n31 1.3005
R363 Vss.n25 Vss.n24 1.3005
R364 Vss.n28 Vss.n27 1.3005
R365 Vss.n27 Vss.n3 1.3005
R366 Vss.n29 Vss.n1 1.29323
R367 Vss.n30 Vss.n29 1.00923
R368 Vss.n41 Vss.n15 0.999917
R369 Vss.n42 Vss.n41 0.999917
R370 Vss.n57 Vss.n56 0.999917
R371 Vss.n57 Vss.n14 0.999917
R372 Vss.n29 Vss.n28 0.984484
R373 Vss.n45 Vss.n44 0.949529
R374 Vss.n44 Vss.n43 0.907842
R375 Vss.n52 Vss.n51 0.867167
R376 Vss.t12 Vss.n17 0.867167
R377 Vss.n54 Vss.n13 0.867167
R378 comparator_no_offsetcal_0.lvsclean_SAlatch_0.VSS Vss.n45 0.664071
R379 Vss.n68 Vss.n0 0.238053
R380 comparator_no_offsetcal_0.VSS Vss.n68 0.222184
R381 Vss.n40 Vss.n39 0.211763
R382 comparator_no_offsetcal_0.x3.avss Vss.n67 0.188808
R383 comparator_no_offsetcal_0.x5.avss Vss.n38 0.188808
R384 Vss.n44 Vss.n0 0.163684
R385 Vss.n46 comparator_no_offsetcal_0.lvsclean_SAlatch_0.VSS 0.1605
R386 Vss.n9 Vss.n8 0.154786
R387 Vss.n12 Vss.n11 0.1355
R388 Vss.n38 Vss.n37 0.128901
R389 Vss.n67 Vss.n66 0.127885
R390 Vss.n43 Vss.n40 0.112526
R391 Vss.n7 Vss.n6 0.109786
R392 Vss.n8 Vss.n7 0.0455
R393 Vss.n41 Vss.n19 0.0215413
R394 Vss.n58 Vss.n57 0.0215413
R395 Vss.n11 Vss.n9 0.0197857
R396 Vss.n6 comparator_no_offsetcal_0.x4.VSS 0.00371429
R397 Vin1.n7 Vin1.n6 23.1032
R398 Vin1.n3 Vin1.n2 23.1032
R399 Vin1.n0 Vin1.t8 22.5295
R400 Vin1.n2 Vin1.t3 16.3641
R401 Vin1.n6 Vin1.t6 16.3626
R402 Vin1.n2 Vin1.t7 16.0225
R403 Vin1.n6 Vin1.t1 16.021
R404 Vin1.n8 Vin1.t4 11.5195
R405 Vin1.n5 Vin1.t2 11.5195
R406 Vin1.n4 Vin1.t9 11.5195
R407 Vin1.n1 Vin1.t5 11.5195
R408 Vin1.n0 Vin1.t0 11.5195
R409 comparator_no_offsetcal_0.Vin1 Vin1 6.1115
R410 Vin1.n1 Vin1.n0 4.00673
R411 comparator_no_offsetcal_0.Vin1 Vin1.n8 3.5169
R412 Vin1.n7 Vin1.n5 3.16619
R413 Vin1.n3 Vin1.n1 0.650658
R414 Vin1.n8 Vin1.n7 0.280193
R415 Vin1.n4 Vin1.n3 0.279681
R416 Vin1.n5 Vin1.n4 0.231705
R417 a_n9429_n3007.n18 a_n9429_n3007.n17 11.2899
R418 a_n9429_n3007.n17 a_n9429_n3007.n16 8.49339
R419 a_n9429_n3007.n10 a_n9429_n3007.n9 4.89725
R420 a_n9429_n3007.n14 a_n9429_n3007.n2 4.89725
R421 a_n9429_n3007.n13 a_n9429_n3007.n3 4.89725
R422 a_n9429_n3007.n12 a_n9429_n3007.n5 4.89725
R423 a_n9429_n3007.n11 a_n9429_n3007.n7 4.89725
R424 a_n9429_n3007.n13 a_n9429_n3007.n4 4.88712
R425 a_n9429_n3007.n12 a_n9429_n3007.n6 4.88712
R426 a_n9429_n3007.n11 a_n9429_n3007.n8 4.88712
R427 a_n9429_n3007.n1 a_n9429_n3007.n0 4.4
R428 a_n9429_n3007.n16 a_n9429_n3007.n15 4.35275
R429 a_n9429_n3007.t0 a_n9429_n3007.n18 2.048
R430 a_n9429_n3007.n18 a_n9429_n3007.t1 2.048
R431 a_n9429_n3007.n17 a_n9429_n3007.n1 1.95895
R432 a_n9429_n3007.n9 a_n9429_n3007.t2 1.0925
R433 a_n9429_n3007.n9 a_n9429_n3007.t14 1.0925
R434 a_n9429_n3007.n0 a_n9429_n3007.t17 1.0925
R435 a_n9429_n3007.n0 a_n9429_n3007.t5 1.0925
R436 a_n9429_n3007.n2 a_n9429_n3007.t20 1.0925
R437 a_n9429_n3007.n2 a_n9429_n3007.t18 1.0925
R438 a_n9429_n3007.n15 a_n9429_n3007.t10 1.0925
R439 a_n9429_n3007.n15 a_n9429_n3007.t7 1.0925
R440 a_n9429_n3007.n3 a_n9429_n3007.t13 1.0925
R441 a_n9429_n3007.n3 a_n9429_n3007.t3 1.0925
R442 a_n9429_n3007.n4 a_n9429_n3007.t6 1.0925
R443 a_n9429_n3007.n4 a_n9429_n3007.t15 1.0925
R444 a_n9429_n3007.n5 a_n9429_n3007.t19 1.0925
R445 a_n9429_n3007.n5 a_n9429_n3007.t9 1.0925
R446 a_n9429_n3007.n6 a_n9429_n3007.t11 1.0925
R447 a_n9429_n3007.n6 a_n9429_n3007.t21 1.0925
R448 a_n9429_n3007.n7 a_n9429_n3007.t16 1.0925
R449 a_n9429_n3007.n7 a_n9429_n3007.t8 1.0925
R450 a_n9429_n3007.n8 a_n9429_n3007.t4 1.0925
R451 a_n9429_n3007.n8 a_n9429_n3007.t12 1.0925
R452 a_n9429_n3007.n14 a_n9429_n3007.n13 0.849071
R453 a_n9429_n3007.n13 a_n9429_n3007.n12 0.849071
R454 a_n9429_n3007.n12 a_n9429_n3007.n11 0.849071
R455 a_n9429_n3007.n11 a_n9429_n3007.n10 0.849071
R456 a_n9429_n3007.n16 a_n9429_n3007.n14 0.534875
R457 a_n9429_n3007.n10 a_n9429_n3007.n1 0.487625
R458 Comp_out.n9 Comp_out 11.2807
R459 Comp_out.n5 Comp_out.n4 6.5435
R460 Comp_out.n2 Comp_out.n1 6.5435
R461 comparator_no_offsetcal_0.x4.Y Comp_out.n8 4.5005
R462 Comp_out.n9 comparator_no_offsetcal_0.x4.Y 2.3842
R463 Comp_out.n6 Comp_out.n3 2.17483
R464 Comp_out.n4 Comp_out.t1 2.03874
R465 Comp_out.n4 Comp_out.t2 2.03874
R466 Comp_out.n1 Comp_out.t0 2.03874
R467 Comp_out.n1 Comp_out.t3 2.03874
R468 Comp_out.n8 Comp_out.n0 2.00383
R469 Comp_out.n0 Comp_out.t7 1.13285
R470 Comp_out.n0 Comp_out.t6 1.13285
R471 Comp_out.n3 Comp_out.t4 1.13285
R472 Comp_out.n3 Comp_out.t5 1.13285
R473 Comp_out.n5 Comp_out.n2 0.5105
R474 Comp_out.n7 Comp_out.n6 0.5105
R475 Comp_out.n7 Comp_out.n2 0.2165
R476 Comp_out.n6 Comp_out.n5 0.2165
R477 Comp_out.n8 Comp_out.n7 0.1175
R478 comparator_no_offsetcal_0.Vout Comp_out.n9 0.0311818
R479 Vin2.n7 Vin2.n6 23.1032
R480 Vin2.n3 Vin2.n2 23.1032
R481 Vin2.n0 Vin2.t6 22.8502
R482 Vin2.n2 Vin2.t5 16.3656
R483 Vin2.n6 Vin2.t1 16.3641
R484 Vin2.n2 Vin2.t2 16.021
R485 Vin2.n6 Vin2.t4 16.0195
R486 Vin2.n8 Vin2.t8 11.5195
R487 Vin2.n5 Vin2.t7 11.5195
R488 Vin2.n4 Vin2.t0 11.5195
R489 Vin2.n1 Vin2.t9 11.5195
R490 Vin2.n0 Vin2.t3 11.5195
R491 comparator_no_offsetcal_0.Vin2 Vin2 6.1091
R492 comparator_no_offsetcal_0.Vin2 Vin2.n8 3.51835
R493 Vin2.n7 Vin2.n5 2.53166
R494 Vin2.n1 Vin2.n0 2.48408
R495 Vin2.n3 Vin2.n1 1.40666
R496 Vin2.n8 Vin2.n7 0.647658
R497 Vin2.n4 Vin2.n3 0.647132
R498 Vin2.n5 Vin2.n4 0.234605
R499 SARlogic_0.reset Reset 0.18425
R500 SARlogic_0.comp_in SAR_in 0.1775
.ends

