magic
tech gf180mcuD
magscale 1 10
timestamp 1758004169
<< nwell >>
rect 106 1180 2074 2200
<< pwell >>
rect 1726 1091 1812 1171
rect 106 460 706 1080
rect 790 990 1390 1080
rect 790 732 1436 990
rect 790 460 1390 732
rect 1474 460 2074 1080
<< nmos >>
rect 356 670 456 870
rect 1040 670 1140 870
rect 1724 670 1824 870
<< pmos >>
rect 356 1390 456 1990
rect 560 1390 660 1990
rect 1040 1390 1140 1990
rect 1244 1390 1344 1990
rect 1724 1390 1824 1990
<< ndiff >>
rect 268 857 356 870
rect 268 683 281 857
rect 327 683 356 857
rect 268 670 356 683
rect 456 857 544 870
rect 456 683 485 857
rect 531 683 544 857
rect 456 670 544 683
rect 952 857 1040 870
rect 952 683 965 857
rect 1011 683 1040 857
rect 952 670 1040 683
rect 1140 857 1228 870
rect 1140 683 1169 857
rect 1215 683 1228 857
rect 1140 670 1228 683
rect 1636 857 1724 870
rect 1636 683 1649 857
rect 1695 683 1724 857
rect 1636 670 1724 683
rect 1824 857 1912 870
rect 1824 683 1853 857
rect 1899 683 1912 857
rect 1824 670 1912 683
<< pdiff >>
rect 268 1977 356 1990
rect 268 1403 281 1977
rect 327 1403 356 1977
rect 268 1390 356 1403
rect 456 1977 560 1990
rect 456 1403 485 1977
rect 531 1403 560 1977
rect 456 1390 560 1403
rect 660 1977 748 1990
rect 660 1403 689 1977
rect 735 1403 748 1977
rect 660 1390 748 1403
rect 952 1977 1040 1990
rect 952 1403 965 1977
rect 1011 1403 1040 1977
rect 952 1390 1040 1403
rect 1140 1977 1244 1990
rect 1140 1403 1169 1977
rect 1215 1403 1244 1977
rect 1140 1390 1244 1403
rect 1344 1977 1432 1990
rect 1344 1403 1373 1977
rect 1419 1403 1432 1977
rect 1344 1390 1432 1403
rect 1636 1977 1724 1990
rect 1636 1403 1649 1977
rect 1695 1403 1724 1977
rect 1636 1390 1724 1403
rect 1824 1977 1912 1990
rect 1824 1403 1853 1977
rect 1899 1403 1912 1977
rect 1824 1390 1912 1403
<< ndiffc >>
rect 281 683 327 857
rect 485 683 531 857
rect 965 683 1011 857
rect 1169 683 1215 857
rect 1649 683 1695 857
rect 1853 683 1899 857
<< pdiffc >>
rect 281 1403 327 1977
rect 485 1403 531 1977
rect 689 1403 735 1977
rect 965 1403 1011 1977
rect 1169 1403 1215 1977
rect 1373 1403 1419 1977
rect 1649 1403 1695 1977
rect 1853 1403 1899 1977
<< psubdiff >>
rect 130 984 682 1056
rect 130 940 202 984
rect 130 600 143 940
rect 189 600 202 940
rect 610 940 682 984
rect 130 556 202 600
rect 610 600 623 940
rect 669 600 682 940
rect 610 556 682 600
rect 130 484 682 556
rect 814 984 1366 1056
rect 814 940 886 984
rect 814 600 827 940
rect 873 600 886 940
rect 1294 940 1366 984
rect 814 556 886 600
rect 1294 600 1307 940
rect 1353 600 1366 940
rect 1294 556 1366 600
rect 814 484 1366 556
rect 1498 984 2050 1056
rect 1498 940 1570 984
rect 1498 600 1511 940
rect 1557 600 1570 940
rect 1978 940 2050 984
rect 1498 556 1570 600
rect 1978 600 1991 940
rect 2037 600 2050 940
rect 1978 556 2050 600
rect 1498 484 2050 556
<< nsubdiff >>
rect 130 2104 2050 2176
rect 130 2060 202 2104
rect 130 1320 143 2060
rect 189 1320 202 2060
rect 814 2060 886 2104
rect 130 1276 202 1320
rect 814 1320 827 2060
rect 873 1320 886 2060
rect 1498 2060 1570 2104
rect 814 1276 886 1320
rect 1498 1320 1511 2060
rect 1557 1320 1570 2060
rect 1978 2060 2050 2104
rect 1498 1276 1570 1320
rect 1978 1320 1991 2060
rect 2037 1320 2050 2060
rect 1978 1276 2050 1320
rect 130 1204 2050 1276
<< psubdiffcont >>
rect 143 600 189 940
rect 623 600 669 940
rect 827 600 873 940
rect 1307 600 1353 940
rect 1511 600 1557 940
rect 1991 600 2037 940
<< nsubdiffcont >>
rect 143 1320 189 2060
rect 827 1320 873 2060
rect 1511 1320 1557 2060
rect 1991 1320 2037 2060
<< polysilicon >>
rect 356 2069 456 2082
rect 356 2023 369 2069
rect 443 2023 456 2069
rect 356 1990 456 2023
rect 560 2069 660 2082
rect 560 2023 573 2069
rect 647 2023 660 2069
rect 560 1990 660 2023
rect 356 1357 456 1390
rect 356 1311 369 1357
rect 443 1311 456 1357
rect 356 1298 456 1311
rect 560 1357 660 1390
rect 560 1311 573 1357
rect 647 1311 660 1357
rect 560 1298 660 1311
rect 1040 2069 1140 2082
rect 1040 2023 1053 2069
rect 1127 2023 1140 2069
rect 1040 1990 1140 2023
rect 1244 2069 1344 2082
rect 1244 2023 1257 2069
rect 1331 2023 1344 2069
rect 1244 1990 1344 2023
rect 1040 1357 1140 1390
rect 1040 1311 1053 1357
rect 1127 1311 1140 1357
rect 1040 1298 1140 1311
rect 1244 1357 1344 1390
rect 1244 1311 1257 1357
rect 1331 1311 1344 1357
rect 1244 1298 1344 1311
rect 1724 2069 1824 2082
rect 1724 2023 1737 2069
rect 1811 2023 1824 2069
rect 1724 1990 1824 2023
rect 1724 1357 1824 1390
rect 1724 1311 1737 1357
rect 1811 1311 1824 1357
rect 1724 1298 1824 1311
rect 356 949 456 962
rect 356 903 369 949
rect 443 903 456 949
rect 356 870 456 903
rect 356 637 456 670
rect 356 591 369 637
rect 443 591 456 637
rect 356 578 456 591
rect 1040 949 1140 962
rect 1040 903 1053 949
rect 1127 903 1140 949
rect 1040 870 1140 903
rect 1040 637 1140 670
rect 1040 591 1053 637
rect 1127 591 1140 637
rect 1040 578 1140 591
rect 1724 949 1824 962
rect 1724 903 1737 949
rect 1811 903 1824 949
rect 1724 870 1824 903
rect 1724 637 1824 670
rect 1724 591 1737 637
rect 1811 591 1824 637
rect 1724 578 1824 591
<< polycontact >>
rect 369 2023 443 2069
rect 573 2023 647 2069
rect 369 1311 443 1357
rect 573 1311 647 1357
rect 1053 2023 1127 2069
rect 1257 2023 1331 2069
rect 1053 1311 1127 1357
rect 1257 1311 1331 1357
rect 1737 2023 1811 2069
rect 1737 1311 1811 1357
rect 369 903 443 949
rect 369 591 443 637
rect 1053 903 1127 949
rect 1053 591 1127 637
rect 1737 903 1811 949
rect 1737 591 1811 637
<< metal1 >>
rect 106 2200 2074 2403
rect 143 2060 189 2200
rect 358 2069 454 2100
rect 358 2023 369 2069
rect 443 2023 454 2069
rect 562 2069 658 2100
rect 562 2023 573 2069
rect 647 2023 658 2069
rect 827 2060 873 2200
rect 189 1977 327 1988
rect 485 1977 531 1988
rect 689 1977 827 1988
rect 189 1403 281 1977
rect 468 1737 480 1977
rect 536 1737 548 1977
rect 189 1392 327 1403
rect 485 1392 531 1403
rect 735 1403 827 1977
rect 689 1392 827 1403
rect 143 1309 189 1320
rect 358 1311 369 1357
rect 443 1337 454 1357
rect 562 1337 573 1357
rect 443 1311 573 1337
rect 647 1311 658 1357
rect 358 1284 658 1311
rect 1042 2069 1138 2100
rect 1042 2023 1053 2069
rect 1127 2023 1138 2069
rect 1246 2069 1342 2100
rect 1246 2023 1257 2069
rect 1331 2023 1342 2069
rect 1511 2060 1557 2200
rect 965 1977 1011 1988
rect 1169 1977 1215 1988
rect 1373 1977 1419 1988
rect 1152 1737 1164 1977
rect 1220 1737 1232 1977
rect 948 1403 960 1643
rect 1016 1403 1028 1643
rect 1356 1403 1368 1643
rect 1424 1403 1436 1643
rect 965 1392 1011 1403
rect 1169 1392 1215 1403
rect 1373 1392 1419 1403
rect 827 1309 873 1320
rect 1042 1311 1053 1357
rect 1127 1337 1138 1357
rect 1246 1337 1257 1357
rect 1127 1311 1257 1337
rect 1331 1311 1342 1357
rect 1042 1284 1342 1311
rect 1726 2069 1822 2100
rect 1726 2023 1737 2069
rect 1811 2023 1822 2069
rect 1991 2060 2037 2200
rect 1557 1977 1695 1988
rect 1557 1403 1649 1977
rect 1853 1977 1899 1988
rect 1836 1693 1853 1703
rect 1899 1693 1916 1703
rect 1836 1453 1848 1693
rect 1904 1453 1916 1693
rect 1836 1443 1853 1453
rect 1557 1392 1695 1403
rect 1899 1443 1916 1453
rect 1853 1392 1899 1403
rect 1511 1309 1557 1320
rect 1726 1311 1737 1357
rect 1811 1311 1822 1357
rect 358 1236 454 1284
rect 358 1180 378 1236
rect 434 1180 454 1236
rect 143 940 189 951
rect 358 949 454 1180
rect 1042 1080 1138 1284
rect 1726 1170 1822 1311
rect 1991 1309 2037 1320
rect 1658 1158 1822 1170
rect 1658 1102 1670 1158
rect 1726 1102 1822 1158
rect 1658 1090 1822 1102
rect 1042 1024 1062 1080
rect 1118 1024 1138 1080
rect 358 903 369 949
rect 443 903 454 949
rect 623 940 873 951
rect 281 857 327 868
rect 264 798 281 808
rect 485 857 623 868
rect 327 798 344 808
rect 264 742 276 798
rect 332 742 344 798
rect 264 732 281 742
rect 327 732 344 742
rect 281 672 327 683
rect 531 683 623 857
rect 485 672 623 683
rect 143 460 189 600
rect 358 591 369 637
rect 443 591 454 637
rect 358 560 454 591
rect 669 600 827 940
rect 1042 949 1138 1024
rect 1042 903 1053 949
rect 1127 903 1138 949
rect 1307 940 1353 951
rect 873 857 1011 868
rect 873 683 965 857
rect 1169 857 1215 868
rect 1152 798 1169 808
rect 1215 798 1232 808
rect 1152 742 1164 798
rect 1220 742 1232 798
rect 1152 732 1169 742
rect 873 672 1011 683
rect 1215 732 1232 742
rect 1169 672 1215 683
rect 623 589 873 600
rect 1042 591 1053 637
rect 1127 591 1138 637
rect 669 460 827 589
rect 1042 560 1138 591
rect 1307 460 1353 600
rect 1511 940 1557 951
rect 1726 949 1822 1090
rect 1726 903 1737 949
rect 1811 903 1822 949
rect 1991 940 2037 951
rect 1557 857 1695 868
rect 1557 683 1649 857
rect 1853 857 1899 868
rect 1836 798 1853 808
rect 1899 798 1916 808
rect 1836 742 1848 798
rect 1904 742 1916 798
rect 1836 732 1853 742
rect 1557 672 1695 683
rect 1899 732 1916 742
rect 1853 672 1899 683
rect 1511 460 1557 600
rect 1726 591 1737 637
rect 1811 591 1822 637
rect 1726 560 1822 591
rect 1991 460 2037 600
rect 106 257 2074 460
<< via1 >>
rect 480 1737 485 1977
rect 485 1737 531 1977
rect 531 1737 536 1977
rect 1164 1737 1169 1977
rect 1169 1737 1215 1977
rect 1215 1737 1220 1977
rect 960 1403 965 1643
rect 965 1403 1011 1643
rect 1011 1403 1016 1643
rect 1368 1403 1373 1643
rect 1373 1403 1419 1643
rect 1419 1403 1424 1643
rect 1848 1453 1853 1693
rect 1853 1453 1899 1693
rect 1899 1453 1904 1693
rect 378 1180 434 1236
rect 1670 1102 1726 1158
rect 1062 1024 1118 1080
rect 276 742 281 798
rect 281 742 327 798
rect 327 742 332 798
rect 1164 742 1169 798
rect 1169 742 1215 798
rect 1215 742 1220 798
rect 1848 742 1853 798
rect 1853 742 1899 798
rect 1899 742 1904 798
<< metal2 >>
rect 468 1977 1232 1987
rect 468 1737 480 1977
rect 536 1737 1164 1977
rect 1220 1737 1232 1977
rect 468 1727 1232 1737
rect 1836 1693 1916 1703
rect 948 1643 1436 1653
rect 948 1403 960 1643
rect 1016 1403 1368 1643
rect 1424 1403 1436 1643
rect 948 1393 1436 1403
rect 358 1236 454 1248
rect 46 1180 378 1236
rect 434 1180 454 1236
rect 358 1168 454 1180
rect 1356 1158 1436 1393
rect 1836 1453 1848 1693
rect 1904 1453 1916 1693
rect 1658 1158 1728 1170
rect 1356 1102 1670 1158
rect 1726 1102 1728 1158
rect 1042 1080 1138 1090
rect 46 1024 1062 1080
rect 1118 1024 1138 1080
rect 1042 1014 1138 1024
rect 1356 808 1436 1102
rect 1658 1090 1728 1102
rect 1836 1158 1916 1453
rect 1836 1102 2078 1158
rect 264 798 1436 808
rect 264 742 276 798
rect 332 742 1164 798
rect 1220 742 1436 798
rect 264 732 1436 742
rect 1836 798 1916 1102
rect 1836 742 1848 798
rect 1904 742 1916 798
rect 1836 732 1916 742
<< labels >>
rlabel metal1 1083 2403 1083 2403 1 VDD
port 0 n
rlabel metal1 1098 257 1098 257 5 VSS
port 1 s
rlabel metal2 2078 1130 2078 1130 3 OUT
port 2 e
rlabel metal2 46 1207 46 1207 7 A
port 3 w
rlabel metal2 46 1052 46 1052 7 B
port 4 w
<< end >>
