magic
tech gf180mcuD
magscale 1 10
timestamp 1755269543
<< error_p >>
rect 11144 9933 11155 9979
rect 11201 9933 11212 9944
rect -656 9813 -645 9859
rect -599 9813 -588 9824
rect 13424 9823 13435 9869
rect 21874 9843 21885 9889
rect 21931 9843 21942 9854
rect 13481 9823 13492 9834
rect 10374 9763 10385 9809
rect 10431 9763 10442 9774
rect 1624 9703 1635 9749
rect 1681 9703 1692 9714
rect 11904 9713 11915 9759
rect 11961 9713 11972 9724
rect 14114 9723 14125 9769
rect 14171 9723 14182 9734
rect -1426 9643 -1415 9689
rect 12664 9673 12675 9719
rect 14884 9693 14895 9739
rect 24154 9733 24165 9779
rect 24211 9733 24222 9744
rect 14941 9693 14952 9704
rect 12721 9673 12732 9684
rect 21104 9673 21115 9719
rect 21161 9673 21172 9684
rect -1369 9643 -1358 9654
rect 104 9593 115 9639
rect 161 9593 172 9604
rect 2314 9603 2325 9649
rect 2371 9603 2382 9614
rect 864 9553 875 9599
rect 3084 9573 3095 9619
rect 15614 9613 15625 9659
rect 15671 9613 15682 9624
rect 22634 9623 22645 9669
rect 22691 9623 22702 9634
rect 24844 9633 24855 9679
rect 24901 9633 24912 9644
rect 3141 9573 3152 9584
rect 921 9553 932 9564
rect 16414 9543 16425 9589
rect 23394 9583 23405 9629
rect 25614 9603 25625 9649
rect 25671 9603 25682 9614
rect 23451 9583 23462 9594
rect 16471 9543 16482 9554
rect 3814 9493 3825 9539
rect 10328 9532 10351 9543
rect 10465 9532 10488 9543
rect 26344 9523 26355 9569
rect 26401 9523 26412 9534
rect 3871 9493 3882 9504
rect 11098 9502 11121 9513
rect 11235 9502 11258 9513
rect 4614 9423 4625 9469
rect 10374 9451 10385 9497
rect 11858 9482 11881 9493
rect 11995 9482 12018 9493
rect 4671 9423 4682 9434
rect -1472 9412 -1449 9423
rect -1335 9412 -1312 9423
rect 11144 9421 11155 9467
rect 27144 9453 27155 9499
rect 32174 9493 32185 9539
rect 32231 9493 32242 9504
rect 42824 9493 42835 9539
rect 42881 9493 42892 9504
rect 27201 9453 27212 9464
rect 11904 9401 11915 9447
rect 12618 9442 12641 9453
rect 12755 9442 12778 9453
rect 21058 9442 21081 9453
rect 21195 9442 21218 9453
rect 21828 9412 21851 9423
rect 21965 9412 21988 9423
rect -702 9382 -679 9393
rect -565 9382 -542 9393
rect -1426 9331 -1415 9377
rect 58 9362 81 9373
rect 195 9362 218 9373
rect 12664 9361 12675 9407
rect 13378 9392 13401 9403
rect 13515 9392 13538 9403
rect 21104 9361 21115 9407
rect 22588 9392 22611 9403
rect 22725 9392 22748 9403
rect 34454 9383 34465 9429
rect 34511 9383 34522 9394
rect 45104 9383 45115 9429
rect 45161 9383 45172 9394
rect -656 9301 -645 9347
rect 104 9281 115 9327
rect 818 9322 841 9333
rect 955 9322 978 9333
rect 13424 9311 13435 9357
rect 21874 9331 21885 9377
rect 22634 9311 22645 9357
rect 23348 9352 23371 9363
rect 23485 9352 23508 9363
rect 31404 9323 31415 9369
rect 31461 9323 31472 9334
rect 14068 9292 14091 9303
rect 14205 9292 14228 9303
rect 864 9241 875 9287
rect 1578 9272 1601 9283
rect 1715 9272 1738 9283
rect 14838 9262 14861 9273
rect 14975 9262 14998 9273
rect 23394 9271 23405 9317
rect 24108 9302 24131 9313
rect 24245 9302 24268 9313
rect 32934 9273 32945 9319
rect 32991 9273 33002 9284
rect 35144 9283 35155 9329
rect 42054 9323 42065 9369
rect 42111 9323 42122 9334
rect 35201 9283 35212 9294
rect 1624 9191 1635 9237
rect 14114 9211 14125 9257
rect 2268 9172 2291 9183
rect 2405 9172 2428 9183
rect 14884 9181 14895 9227
rect 24154 9221 24165 9267
rect 33694 9233 33705 9279
rect 35914 9253 35925 9299
rect 43584 9273 43595 9319
rect 43641 9273 43652 9284
rect 45794 9283 45805 9329
rect 45851 9283 45862 9294
rect 35971 9253 35982 9264
rect 33751 9233 33762 9244
rect 44344 9233 44355 9279
rect 46564 9253 46575 9299
rect 46621 9253 46632 9264
rect 44401 9233 44412 9244
rect 24798 9202 24821 9213
rect 24935 9202 24958 9213
rect 15570 9182 15591 9193
rect 15705 9182 15728 9193
rect 25568 9172 25591 9183
rect 25705 9172 25728 9183
rect 36644 9173 36655 9219
rect 36701 9173 36712 9184
rect 47294 9173 47305 9219
rect 47351 9173 47362 9184
rect 3038 9142 3061 9153
rect 3175 9142 3198 9153
rect 2314 9091 2325 9137
rect 3084 9061 3095 9107
rect 15614 9101 15625 9147
rect 16368 9112 16391 9123
rect 16505 9112 16528 9123
rect 24844 9121 24855 9167
rect 25614 9091 25625 9137
rect 37444 9103 37455 9149
rect 37501 9103 37512 9114
rect 48094 9103 48105 9149
rect 48151 9103 48162 9114
rect 26300 9092 26321 9103
rect 26435 9092 26458 9103
rect 31358 9092 31381 9103
rect 31495 9092 31518 9103
rect 42008 9092 42031 9103
rect 42145 9092 42168 9103
rect 3770 9062 3791 9073
rect 3905 9062 3928 9073
rect 16414 9031 16425 9077
rect 32128 9062 32151 9073
rect 32265 9062 32288 9073
rect 42778 9062 42801 9073
rect 42915 9062 42938 9073
rect 3814 8981 3825 9027
rect 26344 9011 26355 9057
rect 27098 9022 27121 9033
rect 27235 9022 27258 9033
rect 31404 9011 31415 9057
rect 32888 9042 32911 9053
rect 33025 9042 33048 9053
rect 4568 8992 4591 9003
rect 4705 8992 4728 9003
rect 4614 8911 4625 8957
rect 27144 8941 27155 8987
rect 32174 8981 32185 9027
rect 32934 8961 32945 9007
rect 33648 9002 33671 9013
rect 33785 9002 33808 9013
rect 42054 9011 42065 9057
rect 43538 9042 43561 9053
rect 43675 9042 43698 9053
rect 42824 8981 42835 9027
rect 33694 8921 33705 8967
rect 34408 8952 34431 8963
rect 34545 8952 34568 8963
rect 43584 8961 43595 9007
rect 44298 9002 44321 9013
rect 44435 9002 44458 9013
rect 44344 8921 44355 8967
rect 45058 8952 45081 8963
rect 45195 8952 45218 8963
rect 34454 8871 34465 8917
rect 45104 8871 45115 8917
rect 35098 8852 35121 8863
rect 35235 8852 35258 8863
rect 45748 8852 45771 8863
rect 45885 8852 45908 8863
rect 35868 8822 35891 8833
rect 36005 8822 36028 8833
rect 46518 8822 46541 8833
rect 46655 8822 46678 8833
rect 35144 8771 35155 8817
rect 35914 8741 35925 8787
rect 45794 8771 45805 8817
rect 36600 8742 36621 8753
rect 36735 8742 36758 8753
rect 46564 8741 46575 8787
rect 47250 8742 47271 8753
rect 47385 8742 47408 8753
rect 10364 8633 10375 8679
rect 36644 8661 36655 8707
rect 37398 8672 37421 8683
rect 37535 8672 37558 8683
rect 47294 8661 47305 8707
rect 48048 8672 48071 8683
rect 48185 8672 48208 8683
rect 10421 8633 10432 8644
rect 11154 8613 11165 8659
rect 11211 8613 11222 8624
rect 37444 8591 37455 8637
rect 48094 8591 48105 8637
rect -1436 8513 -1425 8559
rect 21094 8543 21105 8589
rect 21151 8543 21162 8554
rect -1379 8513 -1368 8524
rect -646 8493 -635 8539
rect -589 8493 -578 8504
rect 11984 8463 11995 8509
rect 12684 8493 12695 8539
rect 21884 8523 21895 8569
rect 21941 8523 21952 8534
rect 12741 8493 12752 8504
rect 12041 8463 12052 8474
rect 13424 8453 13435 8499
rect 13481 8453 13492 8464
rect 184 8343 195 8389
rect 884 8373 895 8419
rect 941 8373 952 8384
rect 241 8343 252 8354
rect 1624 8333 1635 8379
rect 22714 8373 22725 8419
rect 23414 8403 23425 8449
rect 23471 8403 23482 8414
rect 22771 8373 22782 8384
rect 24154 8363 24165 8409
rect 24211 8363 24222 8374
rect 1681 8333 1692 8344
rect 12638 8262 12661 8273
rect 12775 8262 12798 8273
rect 11938 8232 11961 8243
rect 12075 8232 12098 8243
rect 10318 8202 10341 8213
rect 10455 8202 10478 8213
rect 11108 8182 11131 8193
rect 11245 8182 11268 8193
rect 838 8142 861 8153
rect 975 8142 998 8153
rect 138 8112 161 8123
rect 275 8112 298 8123
rect 10364 8121 10375 8167
rect 11984 8151 11995 8197
rect 12684 8181 12695 8227
rect 14154 8183 14165 8229
rect 14211 8183 14222 8194
rect 14834 8163 14845 8209
rect 15634 8183 15645 8229
rect 15691 8183 15702 8194
rect 31394 8193 31405 8239
rect 31451 8193 31462 8204
rect 14891 8163 14902 8174
rect 23368 8172 23391 8183
rect 23505 8172 23528 8183
rect 32184 8173 32195 8219
rect 42044 8193 42055 8239
rect 42101 8193 42112 8204
rect 32241 8173 32252 8184
rect 42834 8173 42845 8219
rect 42891 8173 42902 8184
rect -1482 8082 -1459 8093
rect -1345 8082 -1322 8093
rect -692 8062 -669 8073
rect -555 8062 -532 8073
rect -1436 8001 -1425 8047
rect 184 8031 195 8077
rect 884 8061 895 8107
rect 2354 8063 2365 8109
rect 2411 8063 2422 8074
rect 3034 8043 3045 8089
rect 3834 8063 3845 8109
rect 11154 8101 11165 8147
rect 16374 8123 16385 8169
rect 22668 8142 22691 8153
rect 22805 8142 22828 8153
rect 16431 8123 16442 8134
rect 21048 8112 21071 8123
rect 21185 8112 21208 8123
rect 21838 8092 21861 8103
rect 21975 8092 21998 8103
rect 3891 8063 3902 8074
rect 3091 8043 3102 8054
rect -646 7981 -635 8027
rect 4574 8003 4585 8049
rect 13378 8022 13401 8033
rect 13515 8022 13538 8033
rect 21094 8031 21105 8077
rect 22714 8061 22725 8107
rect 23414 8091 23425 8137
rect 24884 8093 24895 8139
rect 24941 8093 24952 8104
rect 25564 8073 25575 8119
rect 26364 8093 26375 8139
rect 26421 8093 26432 8104
rect 25621 8073 25632 8084
rect 4631 8003 4642 8014
rect 21884 8011 21895 8057
rect 27104 8033 27115 8079
rect 27161 8033 27172 8044
rect 33014 8023 33025 8069
rect 33714 8053 33725 8099
rect 33771 8053 33782 8064
rect 33071 8023 33082 8034
rect 34454 8013 34465 8059
rect 34511 8013 34522 8024
rect 43664 8023 43675 8069
rect 44364 8053 44375 8099
rect 44421 8053 44432 8064
rect 43721 8023 43732 8034
rect 45104 8013 45115 8059
rect 45161 8013 45172 8024
rect 13424 7941 13435 7987
rect 14108 7952 14131 7963
rect 14245 7952 14268 7963
rect 15588 7952 15611 7963
rect 15725 7952 15748 7963
rect 14788 7932 14811 7943
rect 14925 7932 14948 7943
rect 24108 7932 24131 7943
rect 24245 7932 24268 7943
rect 1578 7902 1601 7913
rect 1715 7902 1738 7913
rect 14154 7871 14165 7917
rect 1624 7821 1635 7867
rect 14834 7851 14845 7897
rect 15634 7871 15645 7917
rect 16328 7892 16351 7903
rect 16465 7892 16488 7903
rect 2308 7832 2331 7843
rect 2445 7832 2468 7843
rect 3788 7832 3811 7843
rect 3925 7832 3948 7843
rect 2988 7812 3011 7823
rect 3125 7812 3148 7823
rect 16374 7811 16385 7857
rect 24154 7851 24165 7897
rect 24838 7862 24861 7873
rect 24975 7862 24998 7873
rect 26318 7862 26341 7873
rect 26455 7862 26478 7873
rect 25518 7842 25541 7853
rect 25655 7842 25678 7853
rect 2354 7751 2365 7797
rect 3034 7731 3045 7777
rect 3834 7751 3845 7797
rect 4528 7772 4551 7783
rect 4665 7772 4688 7783
rect 24884 7781 24895 7827
rect 25564 7761 25575 7807
rect 26364 7781 26375 7827
rect 33668 7822 33691 7833
rect 33805 7822 33828 7833
rect 44318 7822 44341 7833
rect 44455 7822 44478 7833
rect 27058 7802 27081 7813
rect 27195 7802 27218 7813
rect 32968 7792 32991 7803
rect 33105 7792 33128 7803
rect 43618 7792 43641 7803
rect 43755 7792 43778 7803
rect 4574 7691 4585 7737
rect 27104 7721 27115 7767
rect 31348 7762 31371 7773
rect 31485 7762 31508 7773
rect 32138 7742 32161 7753
rect 32275 7742 32298 7753
rect 31394 7681 31405 7727
rect 33014 7711 33025 7757
rect 33714 7741 33725 7787
rect 35184 7743 35195 7789
rect 35241 7743 35252 7754
rect 35864 7723 35875 7769
rect 36664 7743 36675 7789
rect 41998 7762 42021 7773
rect 42135 7762 42158 7773
rect 36721 7743 36732 7754
rect 42788 7742 42811 7753
rect 42925 7742 42948 7753
rect 35921 7723 35932 7734
rect 32184 7661 32195 7707
rect 37404 7683 37415 7729
rect 37461 7683 37472 7694
rect 42044 7681 42055 7727
rect 43664 7711 43675 7757
rect 44364 7741 44375 7787
rect 45834 7743 45845 7789
rect 45891 7743 45902 7754
rect 46514 7723 46525 7769
rect 47314 7743 47325 7789
rect 47371 7743 47382 7754
rect 46571 7723 46582 7734
rect 42834 7661 42845 7707
rect 48054 7683 48065 7729
rect 48111 7683 48122 7694
rect 34408 7582 34431 7593
rect 34545 7582 34568 7593
rect 45058 7582 45081 7593
rect 45195 7582 45218 7593
rect 34454 7501 34465 7547
rect 35138 7512 35161 7523
rect 35275 7512 35298 7523
rect 36618 7512 36641 7523
rect 36755 7512 36778 7523
rect 35818 7492 35841 7503
rect 35955 7492 35978 7503
rect 45104 7501 45115 7547
rect 45788 7512 45811 7523
rect 45925 7512 45948 7523
rect 47268 7512 47291 7523
rect 47405 7512 47428 7523
rect 46468 7492 46491 7503
rect 46605 7492 46628 7503
rect 35184 7431 35195 7477
rect 35864 7411 35875 7457
rect 36664 7431 36675 7477
rect 37358 7452 37381 7463
rect 37495 7452 37518 7463
rect 45834 7431 45845 7477
rect 37404 7371 37415 7417
rect 46514 7411 46525 7457
rect 47314 7431 47325 7477
rect 48008 7452 48031 7463
rect 48145 7452 48168 7463
rect 48054 7371 48065 7417
rect 21094 4523 21105 4569
rect 21151 4523 21162 4534
rect 23374 4413 23385 4459
rect 23431 4413 23442 4424
rect 10624 4353 10635 4399
rect 10681 4353 10692 4364
rect 20324 4353 20335 4399
rect 20381 4353 20392 4364
rect 21854 4303 21865 4349
rect 21911 4303 21922 4314
rect 24064 4313 24075 4359
rect 24121 4313 24132 4324
rect 12904 4243 12915 4289
rect 22614 4263 22625 4309
rect 24834 4283 24845 4329
rect 24891 4283 24902 4294
rect 22671 4263 22682 4274
rect 12961 4243 12972 4254
rect -286 4173 -275 4219
rect -229 4173 -218 4184
rect 9854 4183 9865 4229
rect 25564 4203 25575 4249
rect 25621 4203 25632 4214
rect 9911 4183 9922 4194
rect 11384 4133 11395 4179
rect 11441 4133 11452 4144
rect 13594 4143 13605 4189
rect 13651 4143 13662 4154
rect 1994 4063 2005 4109
rect 12144 4093 12155 4139
rect 14364 4113 14375 4159
rect 26364 4133 26375 4179
rect 31914 4173 31925 4219
rect 31971 4173 31982 4184
rect 26421 4133 26432 4144
rect 14421 4113 14432 4124
rect 20278 4122 20301 4133
rect 20415 4122 20438 4133
rect 12201 4093 12212 4104
rect 21048 4092 21071 4103
rect 21185 4092 21208 4103
rect 2051 4063 2062 4074
rect -1056 4003 -1045 4049
rect 15094 4033 15105 4079
rect 15151 4033 15162 4044
rect 20324 4041 20335 4087
rect 21808 4072 21831 4083
rect 21945 4072 21968 4083
rect 34194 4063 34205 4109
rect 42294 4083 42305 4129
rect 42351 4083 42362 4094
rect 34251 4063 34262 4074
rect -999 4003 -988 4014
rect 21094 4011 21105 4057
rect 474 3953 485 3999
rect 531 3953 542 3964
rect 2684 3963 2695 4009
rect 2741 3963 2752 3974
rect 1234 3913 1245 3959
rect 3454 3933 3465 3979
rect 15894 3963 15905 4009
rect 21854 3991 21865 4037
rect 22568 4032 22591 4043
rect 22705 4032 22728 4043
rect 31144 4003 31155 4049
rect 31201 4003 31212 4014
rect 15951 3963 15962 3974
rect 9808 3952 9831 3963
rect 9945 3952 9968 3963
rect 22614 3951 22625 3997
rect 23328 3982 23351 3993
rect 23465 3982 23488 3993
rect 32674 3953 32685 3999
rect 32731 3953 32742 3964
rect 34884 3963 34895 4009
rect 34941 3963 34952 3974
rect 3511 3933 3522 3944
rect 1291 3913 1302 3924
rect 10578 3922 10601 3933
rect 10715 3922 10738 3933
rect 4184 3853 4195 3899
rect 9854 3871 9865 3917
rect 11338 3902 11361 3913
rect 11475 3902 11498 3913
rect 23374 3901 23385 3947
rect 33434 3913 33445 3959
rect 35654 3933 35665 3979
rect 44574 3973 44585 4019
rect 44631 3973 44642 3984
rect 35711 3933 35722 3944
rect 33491 3913 33502 3924
rect 41524 3913 41535 3959
rect 41581 3913 41592 3924
rect 4241 3853 4252 3864
rect 10624 3841 10635 3887
rect 24018 3882 24041 3893
rect 24155 3882 24178 3893
rect 4984 3783 4995 3829
rect 11384 3821 11395 3867
rect 12098 3862 12121 3873
rect 12235 3862 12258 3873
rect 24788 3852 24811 3863
rect 24925 3852 24948 3863
rect 36384 3853 36395 3899
rect 36441 3853 36452 3864
rect 43054 3863 43065 3909
rect 43111 3863 43122 3874
rect 45264 3873 45275 3919
rect 45321 3873 45332 3884
rect 5041 3783 5052 3794
rect -1102 3772 -1079 3783
rect -965 3772 -942 3783
rect 12144 3781 12155 3827
rect 12858 3812 12881 3823
rect 12995 3812 13018 3823
rect 24064 3801 24075 3847
rect -332 3742 -309 3753
rect -195 3742 -172 3753
rect -1056 3691 -1045 3737
rect 428 3722 451 3733
rect 565 3722 588 3733
rect 12904 3731 12915 3777
rect 24834 3771 24845 3817
rect 37184 3783 37195 3829
rect 43814 3823 43825 3869
rect 46034 3843 46045 3889
rect 46091 3843 46102 3854
rect 43871 3823 43882 3834
rect 37241 3783 37252 3794
rect 25520 3772 25541 3783
rect 25655 3772 25678 3783
rect 31098 3772 31121 3783
rect 31235 3772 31258 3783
rect 46764 3763 46775 3809
rect 46821 3763 46832 3774
rect 31868 3742 31891 3753
rect 32005 3742 32028 3753
rect 13548 3712 13571 3723
rect 13685 3712 13708 3723
rect -286 3661 -275 3707
rect 474 3641 485 3687
rect 1188 3682 1211 3693
rect 1325 3682 1348 3693
rect 14318 3682 14341 3693
rect 14455 3682 14478 3693
rect 25564 3691 25575 3737
rect 26318 3702 26341 3713
rect 26455 3702 26478 3713
rect 31144 3691 31155 3737
rect 32628 3722 32651 3733
rect 32765 3722 32788 3733
rect 1234 3601 1245 3647
rect 1948 3632 1971 3643
rect 2085 3632 2108 3643
rect 13594 3631 13605 3677
rect 14364 3601 14375 3647
rect 26364 3621 26375 3667
rect 31914 3661 31925 3707
rect 47564 3693 47575 3739
rect 47621 3693 47632 3704
rect 32674 3641 32685 3687
rect 33388 3682 33411 3693
rect 33525 3682 33548 3693
rect 41478 3682 41501 3693
rect 41615 3682 41638 3693
rect 42248 3652 42271 3663
rect 42385 3652 42408 3663
rect 15050 3602 15071 3613
rect 15185 3602 15208 3613
rect 33434 3601 33445 3647
rect 34148 3632 34171 3643
rect 34285 3632 34308 3643
rect 41524 3601 41535 3647
rect 43008 3632 43031 3643
rect 43145 3632 43168 3643
rect 1994 3551 2005 3597
rect 2638 3532 2661 3543
rect 2775 3532 2798 3543
rect 15094 3521 15105 3567
rect 34194 3551 34205 3597
rect 42294 3571 42305 3617
rect 43054 3551 43065 3597
rect 43768 3592 43791 3603
rect 43905 3592 43928 3603
rect 15848 3532 15871 3543
rect 15985 3532 16008 3543
rect 34838 3532 34861 3543
rect 34975 3532 34998 3543
rect 3408 3502 3431 3513
rect 3545 3502 3568 3513
rect 35608 3502 35631 3513
rect 35745 3502 35768 3513
rect 43814 3511 43825 3557
rect 44528 3542 44551 3553
rect 44665 3542 44688 3553
rect 2684 3451 2695 3497
rect 3454 3421 3465 3467
rect 15894 3451 15905 3497
rect 34884 3451 34895 3497
rect 4140 3422 4161 3433
rect 4275 3422 4298 3433
rect 35654 3421 35665 3467
rect 44574 3461 44585 3507
rect 45218 3442 45241 3453
rect 45355 3442 45378 3453
rect 36340 3422 36361 3433
rect 36475 3422 36498 3433
rect 45988 3412 46011 3423
rect 46125 3412 46148 3423
rect 4184 3341 4195 3387
rect 4938 3352 4961 3363
rect 5075 3352 5098 3363
rect 36384 3341 36395 3387
rect 37138 3352 37161 3363
rect 37275 3352 37298 3363
rect 45264 3361 45275 3407
rect 46034 3331 46045 3377
rect 46720 3332 46741 3343
rect 46855 3332 46878 3343
rect 4984 3271 4995 3317
rect 37184 3271 37195 3317
rect 20314 3223 20325 3269
rect 46764 3251 46775 3297
rect 47518 3262 47541 3273
rect 47655 3262 47678 3273
rect 20371 3223 20382 3234
rect 21104 3203 21115 3249
rect 21161 3203 21172 3214
rect 47564 3181 47575 3227
rect 9844 3053 9855 3099
rect 9901 3053 9912 3064
rect 10634 3033 10645 3079
rect 21934 3053 21945 3099
rect 22634 3083 22645 3129
rect 22691 3083 22702 3094
rect 21991 3053 22002 3064
rect 10691 3033 10702 3044
rect 23374 3043 23385 3089
rect 23431 3043 23442 3054
rect -1066 2873 -1055 2919
rect -1009 2873 -998 2884
rect -276 2853 -265 2899
rect 11464 2883 11475 2929
rect 12164 2913 12175 2959
rect 12221 2913 12232 2924
rect 11521 2883 11532 2894
rect 12904 2873 12915 2919
rect 12961 2873 12972 2884
rect 31134 2873 31145 2919
rect 31191 2873 31202 2884
rect -219 2853 -208 2864
rect 22588 2852 22611 2863
rect 22725 2852 22748 2863
rect 31924 2853 31935 2899
rect 31981 2853 31992 2864
rect 21888 2822 21911 2833
rect 22025 2822 22048 2833
rect 20268 2792 20291 2803
rect 20405 2792 20428 2803
rect 554 2703 565 2749
rect 1254 2733 1265 2779
rect 21058 2772 21081 2783
rect 21195 2772 21218 2783
rect 1311 2733 1322 2744
rect 611 2703 622 2714
rect 1994 2693 2005 2739
rect 20314 2711 20325 2757
rect 21934 2741 21945 2787
rect 22634 2771 22645 2817
rect 24104 2773 24115 2819
rect 24161 2773 24172 2784
rect 24784 2753 24795 2799
rect 25584 2773 25595 2819
rect 25641 2773 25652 2784
rect 41514 2783 41525 2829
rect 41571 2783 41582 2794
rect 24841 2753 24852 2764
rect 2051 2693 2062 2704
rect 12118 2682 12141 2693
rect 12255 2682 12278 2693
rect 21104 2691 21115 2737
rect 26324 2713 26335 2759
rect 26381 2713 26392 2724
rect 32754 2703 32765 2749
rect 33454 2733 33465 2779
rect 42304 2763 42315 2809
rect 42361 2763 42372 2774
rect 33511 2733 33522 2744
rect 32811 2703 32822 2714
rect 34194 2693 34205 2739
rect 34251 2693 34262 2704
rect 11418 2652 11441 2663
rect 11555 2652 11578 2663
rect 9798 2622 9821 2633
rect 9935 2622 9958 2633
rect 10588 2602 10611 2613
rect 10725 2602 10748 2613
rect 9844 2541 9855 2587
rect 11464 2571 11475 2617
rect 12164 2601 12175 2647
rect 13634 2603 13645 2649
rect 13691 2603 13702 2614
rect 14314 2583 14325 2629
rect 15114 2603 15125 2649
rect 15171 2603 15182 2614
rect 23328 2612 23351 2623
rect 23465 2612 23488 2623
rect 43134 2613 43145 2659
rect 43834 2643 43845 2689
rect 43891 2643 43902 2654
rect 43191 2613 43202 2624
rect 44574 2603 44585 2649
rect 44631 2603 44642 2614
rect 14371 2583 14382 2594
rect 10634 2521 10645 2567
rect 15854 2543 15865 2589
rect 15911 2543 15922 2554
rect 23374 2531 23385 2577
rect 24058 2542 24081 2553
rect 24195 2542 24218 2553
rect 25538 2542 25561 2553
rect 25675 2542 25698 2553
rect 24738 2522 24761 2533
rect 24875 2522 24898 2533
rect 1208 2502 1231 2513
rect 1345 2502 1368 2513
rect 508 2472 531 2483
rect 645 2472 668 2483
rect -1112 2442 -1089 2453
rect -975 2442 -952 2453
rect -322 2422 -299 2433
rect -185 2422 -162 2433
rect -1066 2361 -1055 2407
rect 554 2391 565 2437
rect 1254 2421 1265 2467
rect 2724 2423 2735 2469
rect 2781 2423 2792 2434
rect 3404 2403 3415 2449
rect 4204 2423 4215 2469
rect 24104 2461 24115 2507
rect 12858 2442 12881 2453
rect 12995 2442 13018 2453
rect 24784 2441 24795 2487
rect 25584 2461 25595 2507
rect 33408 2502 33431 2513
rect 33545 2502 33568 2513
rect 26278 2482 26301 2493
rect 26415 2482 26438 2493
rect 32708 2472 32731 2483
rect 32845 2472 32868 2483
rect 4261 2423 4272 2434
rect 3461 2403 3472 2414
rect -276 2341 -265 2387
rect 4944 2363 4955 2409
rect 5001 2363 5012 2374
rect 12904 2361 12915 2407
rect 26324 2401 26335 2447
rect 31088 2442 31111 2453
rect 31225 2442 31248 2453
rect 31878 2422 31901 2433
rect 32015 2422 32038 2433
rect 13588 2372 13611 2383
rect 13725 2372 13748 2383
rect 15068 2372 15091 2383
rect 15205 2372 15228 2383
rect 14268 2352 14291 2363
rect 14405 2352 14428 2363
rect 31134 2361 31145 2407
rect 32754 2391 32765 2437
rect 33454 2421 33465 2467
rect 34924 2423 34935 2469
rect 34981 2423 34992 2434
rect 35604 2403 35615 2449
rect 36404 2423 36415 2469
rect 36461 2423 36472 2434
rect 35661 2403 35672 2414
rect 43788 2412 43811 2423
rect 43925 2412 43948 2423
rect 31924 2341 31935 2387
rect 37144 2363 37155 2409
rect 43088 2382 43111 2393
rect 43225 2382 43248 2393
rect 37201 2363 37212 2374
rect 41468 2352 41491 2363
rect 41605 2352 41628 2363
rect 13634 2291 13645 2337
rect 1948 2262 1971 2273
rect 2085 2262 2108 2273
rect 14314 2271 14325 2317
rect 15114 2291 15125 2337
rect 42258 2332 42281 2343
rect 42395 2332 42418 2343
rect 15808 2312 15831 2323
rect 15945 2312 15968 2323
rect 15854 2231 15865 2277
rect 34148 2262 34171 2273
rect 34285 2262 34308 2273
rect 41514 2271 41525 2317
rect 43134 2301 43145 2347
rect 43834 2331 43845 2377
rect 45304 2333 45315 2379
rect 45361 2333 45372 2344
rect 45984 2313 45995 2359
rect 46784 2333 46795 2379
rect 46841 2333 46852 2344
rect 46041 2313 46052 2324
rect 42304 2251 42315 2297
rect 47524 2273 47535 2319
rect 47581 2273 47592 2284
rect 1994 2181 2005 2227
rect 2678 2192 2701 2203
rect 2815 2192 2838 2203
rect 4158 2192 4181 2203
rect 4295 2192 4318 2203
rect 3358 2172 3381 2183
rect 3495 2172 3518 2183
rect 34194 2181 34205 2227
rect 34878 2192 34901 2203
rect 35015 2192 35038 2203
rect 36358 2192 36381 2203
rect 36495 2192 36518 2203
rect 35558 2172 35581 2183
rect 35695 2172 35718 2183
rect 44528 2172 44551 2183
rect 44665 2172 44688 2183
rect 2724 2111 2735 2157
rect 3404 2091 3415 2137
rect 4204 2111 4215 2157
rect 4898 2132 4921 2143
rect 5035 2132 5058 2143
rect 34924 2111 34935 2157
rect 4944 2051 4955 2097
rect 35604 2091 35615 2137
rect 36404 2111 36415 2157
rect 37098 2132 37121 2143
rect 37235 2132 37258 2143
rect 37144 2051 37155 2097
rect 44574 2091 44585 2137
rect 45258 2102 45281 2113
rect 45395 2102 45418 2113
rect 46738 2102 46761 2113
rect 46875 2102 46898 2113
rect 45938 2082 45961 2093
rect 46075 2082 46098 2093
rect 45304 2021 45315 2067
rect 45984 2001 45995 2047
rect 46784 2021 46795 2067
rect 47478 2042 47501 2053
rect 47615 2042 47638 2053
rect 47524 1961 47535 2007
rect 32354 -1237 32365 -1191
rect 32411 -1237 32422 -1226
rect 34634 -1347 34645 -1301
rect 42564 -1327 42575 -1281
rect 42621 -1327 42632 -1316
rect 34691 -1347 34702 -1336
rect 31584 -1407 31595 -1361
rect 31641 -1407 31652 -1396
rect 33114 -1457 33125 -1411
rect 33171 -1457 33182 -1446
rect 35324 -1447 35335 -1401
rect 35381 -1447 35392 -1436
rect 33874 -1497 33885 -1451
rect 36094 -1477 36105 -1431
rect 44844 -1437 44855 -1391
rect 44901 -1437 44912 -1426
rect 36151 -1477 36162 -1466
rect 33931 -1497 33942 -1486
rect 41794 -1497 41805 -1451
rect 41851 -1497 41862 -1486
rect 36824 -1557 36835 -1511
rect 36881 -1557 36892 -1546
rect 43324 -1547 43335 -1501
rect 43381 -1547 43392 -1536
rect 45534 -1537 45545 -1491
rect 45591 -1537 45602 -1526
rect 37624 -1627 37635 -1581
rect 44084 -1587 44095 -1541
rect 46304 -1567 46315 -1521
rect 46361 -1567 46372 -1556
rect 44141 -1587 44152 -1576
rect 37681 -1627 37692 -1616
rect 154 -1677 165 -1631
rect 31538 -1638 31561 -1627
rect 31675 -1638 31698 -1627
rect 47034 -1647 47045 -1601
rect 47091 -1647 47102 -1636
rect 211 -1677 222 -1666
rect 32308 -1668 32331 -1657
rect 32445 -1668 32468 -1657
rect 31584 -1719 31595 -1673
rect 33068 -1688 33091 -1677
rect 33205 -1688 33228 -1677
rect 2434 -1787 2445 -1741
rect 32354 -1749 32365 -1703
rect 47834 -1717 47845 -1671
rect 47891 -1717 47902 -1706
rect 33114 -1769 33125 -1723
rect 33828 -1728 33851 -1717
rect 33965 -1728 33988 -1717
rect 41748 -1728 41771 -1717
rect 41885 -1728 41908 -1717
rect 42518 -1758 42541 -1747
rect 42655 -1758 42678 -1747
rect 2491 -1787 2502 -1776
rect -616 -1847 -605 -1801
rect -559 -1847 -548 -1836
rect 914 -1897 925 -1851
rect 971 -1897 982 -1886
rect 3124 -1887 3135 -1841
rect 21794 -1847 21805 -1801
rect 33874 -1809 33885 -1763
rect 34588 -1778 34611 -1767
rect 34725 -1778 34748 -1767
rect 41794 -1809 41805 -1763
rect 43278 -1778 43301 -1767
rect 43415 -1778 43438 -1767
rect 21851 -1847 21862 -1836
rect 34634 -1859 34645 -1813
rect 42564 -1839 42575 -1793
rect 43324 -1859 43335 -1813
rect 44038 -1818 44061 -1807
rect 44175 -1818 44198 -1807
rect 3181 -1887 3192 -1876
rect 1674 -1937 1685 -1891
rect 3894 -1917 3905 -1871
rect 35278 -1878 35301 -1867
rect 35415 -1878 35438 -1867
rect 3951 -1917 3962 -1906
rect 36048 -1908 36071 -1897
rect 36185 -1908 36208 -1897
rect 44084 -1899 44095 -1853
rect 44798 -1868 44821 -1857
rect 44935 -1868 44958 -1857
rect 1731 -1937 1742 -1926
rect 4624 -1997 4635 -1951
rect 24074 -1957 24085 -1911
rect 24131 -1957 24142 -1946
rect 35324 -1959 35335 -1913
rect 4681 -1997 4692 -1986
rect 21024 -2017 21035 -1971
rect 36094 -1989 36105 -1943
rect 44844 -1949 44855 -1903
rect 45488 -1968 45511 -1957
rect 45625 -1968 45648 -1957
rect 36780 -1988 36801 -1977
rect 36915 -1988 36938 -1977
rect 46258 -1998 46281 -1987
rect 46395 -1998 46418 -1987
rect 21081 -2017 21092 -2006
rect 5424 -2067 5435 -2021
rect 5481 -2067 5492 -2056
rect -662 -2078 -639 -2067
rect -525 -2078 -502 -2067
rect 108 -2108 131 -2097
rect 245 -2108 268 -2097
rect 10794 -2107 10805 -2061
rect 22554 -2067 22565 -2021
rect 22611 -2067 22622 -2056
rect 24764 -2057 24775 -2011
rect 24821 -2057 24832 -2046
rect 10851 -2107 10862 -2096
rect 23314 -2107 23325 -2061
rect 25534 -2087 25545 -2041
rect 36824 -2069 36835 -2023
rect 37578 -2058 37601 -2047
rect 37715 -2058 37738 -2047
rect 45534 -2049 45545 -2003
rect 25591 -2087 25602 -2076
rect 46304 -2079 46315 -2033
rect 46990 -2078 47011 -2067
rect 47125 -2078 47148 -2067
rect 23371 -2107 23382 -2096
rect -616 -2159 -605 -2113
rect 868 -2128 891 -2117
rect 1005 -2128 1028 -2117
rect 154 -2189 165 -2143
rect 914 -2209 925 -2163
rect 1628 -2168 1651 -2157
rect 1765 -2168 1788 -2157
rect 26264 -2167 26275 -2121
rect 37624 -2139 37635 -2093
rect 26321 -2167 26332 -2156
rect 47034 -2159 47045 -2113
rect 47788 -2148 47811 -2137
rect 47925 -2148 47948 -2137
rect 1674 -2249 1685 -2203
rect 2388 -2218 2411 -2207
rect 2525 -2218 2548 -2207
rect 13074 -2217 13085 -2171
rect 13131 -2217 13142 -2206
rect 2434 -2299 2445 -2253
rect 10024 -2277 10035 -2231
rect 27064 -2237 27075 -2191
rect 27121 -2237 27132 -2226
rect 47834 -2229 47845 -2183
rect 20978 -2248 21001 -2237
rect 21115 -2248 21138 -2237
rect 10081 -2277 10092 -2266
rect 3078 -2318 3101 -2307
rect 3215 -2318 3238 -2307
rect 11554 -2327 11565 -2281
rect 11611 -2327 11622 -2316
rect 13764 -2317 13775 -2271
rect 21748 -2278 21771 -2267
rect 21885 -2278 21908 -2267
rect 13821 -2317 13832 -2306
rect 3848 -2348 3871 -2337
rect 3985 -2348 4008 -2337
rect 3124 -2399 3135 -2353
rect 12314 -2367 12325 -2321
rect 14534 -2347 14545 -2301
rect 21024 -2329 21035 -2283
rect 22508 -2298 22531 -2287
rect 22645 -2298 22668 -2287
rect 14591 -2347 14602 -2336
rect 12371 -2367 12382 -2356
rect 21794 -2359 21805 -2313
rect 22554 -2379 22565 -2333
rect 23268 -2338 23291 -2327
rect 23405 -2338 23428 -2327
rect 3894 -2429 3905 -2383
rect 4580 -2428 4601 -2417
rect 4715 -2428 4738 -2417
rect 15264 -2427 15275 -2381
rect 15321 -2427 15332 -2416
rect 23314 -2419 23325 -2373
rect 24028 -2388 24051 -2377
rect 24165 -2388 24188 -2377
rect 4624 -2509 4635 -2463
rect 5378 -2498 5401 -2487
rect 5515 -2498 5538 -2487
rect 16064 -2497 16075 -2451
rect 24074 -2469 24085 -2423
rect 16121 -2497 16132 -2486
rect 24718 -2488 24741 -2477
rect 24855 -2488 24878 -2477
rect 9978 -2508 10001 -2497
rect 10115 -2508 10138 -2497
rect 25488 -2518 25511 -2507
rect 25625 -2518 25648 -2507
rect 5424 -2579 5435 -2533
rect 10748 -2538 10771 -2527
rect 10885 -2538 10908 -2527
rect 10024 -2589 10035 -2543
rect 11508 -2558 11531 -2547
rect 11645 -2558 11668 -2547
rect 24764 -2569 24775 -2523
rect 31574 -2537 31585 -2491
rect 31631 -2537 31642 -2526
rect 10794 -2619 10805 -2573
rect 11554 -2639 11565 -2593
rect 12268 -2598 12291 -2587
rect 12405 -2598 12428 -2587
rect 25534 -2599 25545 -2553
rect 32364 -2557 32375 -2511
rect 32421 -2557 32432 -2546
rect 26220 -2598 26241 -2587
rect 26355 -2598 26378 -2587
rect 41784 -2627 41795 -2581
rect 41841 -2627 41852 -2616
rect 12314 -2679 12325 -2633
rect 13028 -2648 13051 -2637
rect 13165 -2648 13188 -2637
rect 26264 -2679 26275 -2633
rect 27018 -2668 27041 -2657
rect 27155 -2668 27178 -2657
rect 13074 -2729 13085 -2683
rect 13718 -2748 13741 -2737
rect 13855 -2748 13878 -2737
rect 27064 -2749 27075 -2703
rect 33194 -2707 33205 -2661
rect 33894 -2677 33905 -2631
rect 42574 -2647 42585 -2601
rect 42631 -2647 42642 -2636
rect 33951 -2677 33962 -2666
rect 33251 -2707 33262 -2696
rect 34634 -2717 34645 -2671
rect 34691 -2717 34702 -2706
rect 14488 -2778 14511 -2767
rect 14625 -2778 14648 -2767
rect 13764 -2829 13775 -2783
rect 43404 -2797 43415 -2751
rect 44104 -2767 44115 -2721
rect 44161 -2767 44172 -2756
rect 43461 -2797 43472 -2786
rect 44844 -2807 44855 -2761
rect 44901 -2807 44912 -2796
rect 14534 -2859 14545 -2813
rect 15220 -2858 15241 -2847
rect 15355 -2858 15378 -2847
rect -626 -2977 -615 -2931
rect 15264 -2939 15275 -2893
rect 33848 -2908 33871 -2897
rect 33985 -2908 34008 -2897
rect 16018 -2928 16041 -2917
rect 16155 -2928 16178 -2917
rect 33148 -2938 33171 -2927
rect 33285 -2938 33308 -2927
rect -569 -2977 -558 -2966
rect 164 -2997 175 -2951
rect 221 -2997 232 -2986
rect 16064 -3009 16075 -2963
rect 31528 -2968 31551 -2957
rect 31665 -2968 31688 -2957
rect 32318 -2988 32341 -2977
rect 32455 -2988 32478 -2977
rect 31574 -3049 31585 -3003
rect 33194 -3019 33205 -2973
rect 33894 -2989 33905 -2943
rect 35364 -2987 35375 -2941
rect 35421 -2987 35432 -2976
rect 36044 -3007 36055 -2961
rect 36844 -2987 36855 -2941
rect 36901 -2987 36912 -2976
rect 36101 -3007 36112 -2996
rect 44058 -2998 44081 -2987
rect 44195 -2998 44218 -2987
rect 32364 -3069 32375 -3023
rect 37584 -3047 37595 -3001
rect 43358 -3028 43381 -3017
rect 43495 -3028 43518 -3017
rect 37641 -3047 37652 -3036
rect 41738 -3058 41761 -3047
rect 41875 -3058 41898 -3047
rect 994 -3147 1005 -3101
rect 1694 -3117 1705 -3071
rect 42528 -3078 42551 -3067
rect 42665 -3078 42688 -3067
rect 1751 -3117 1762 -3106
rect 1051 -3147 1062 -3136
rect 2434 -3157 2445 -3111
rect 2491 -3157 2502 -3146
rect 21014 -3147 21025 -3101
rect 21071 -3147 21082 -3136
rect 21804 -3167 21815 -3121
rect 34588 -3148 34611 -3137
rect 34725 -3148 34748 -3137
rect 41784 -3139 41795 -3093
rect 43404 -3109 43415 -3063
rect 44104 -3079 44115 -3033
rect 45574 -3077 45585 -3031
rect 45631 -3077 45642 -3066
rect 46254 -3097 46265 -3051
rect 47054 -3077 47065 -3031
rect 47111 -3077 47122 -3066
rect 46311 -3097 46322 -3086
rect 21861 -3167 21872 -3156
rect 42574 -3159 42585 -3113
rect 47794 -3137 47805 -3091
rect 47851 -3137 47862 -3126
rect 34634 -3229 34645 -3183
rect 35318 -3218 35341 -3207
rect 35455 -3218 35478 -3207
rect 36798 -3218 36821 -3207
rect 36935 -3218 36958 -3207
rect 35998 -3238 36021 -3227
rect 36135 -3238 36158 -3227
rect 44798 -3238 44821 -3227
rect 44935 -3238 44958 -3227
rect 22634 -3317 22645 -3271
rect 23334 -3287 23345 -3241
rect 23391 -3287 23402 -3276
rect 22691 -3317 22702 -3306
rect 24074 -3327 24085 -3281
rect 35364 -3299 35375 -3253
rect 24131 -3327 24142 -3316
rect 36044 -3319 36055 -3273
rect 36844 -3299 36855 -3253
rect 37538 -3278 37561 -3267
rect 37675 -3278 37698 -3267
rect 1648 -3348 1671 -3337
rect 1785 -3348 1808 -3337
rect 37584 -3359 37595 -3313
rect 44844 -3319 44855 -3273
rect 45528 -3308 45551 -3297
rect 45665 -3308 45688 -3297
rect 47008 -3308 47031 -3297
rect 47145 -3308 47168 -3297
rect 46208 -3328 46231 -3317
rect 46345 -3328 46368 -3317
rect 948 -3378 971 -3367
rect 1085 -3378 1108 -3367
rect -672 -3408 -649 -3397
rect -535 -3408 -512 -3397
rect 118 -3428 141 -3417
rect 255 -3428 278 -3417
rect -626 -3489 -615 -3443
rect 994 -3459 1005 -3413
rect 1694 -3429 1705 -3383
rect 3164 -3427 3175 -3381
rect 3221 -3427 3232 -3416
rect 3844 -3447 3855 -3401
rect 4644 -3427 4655 -3381
rect 10014 -3407 10025 -3361
rect 10071 -3407 10082 -3396
rect 4701 -3427 4712 -3416
rect 10804 -3427 10815 -3381
rect 45574 -3389 45585 -3343
rect 46254 -3409 46265 -3363
rect 47054 -3389 47065 -3343
rect 47748 -3368 47771 -3357
rect 47885 -3368 47908 -3357
rect 10861 -3427 10872 -3416
rect 3901 -3447 3912 -3436
rect 164 -3509 175 -3463
rect 5384 -3487 5395 -3441
rect 47794 -3449 47805 -3403
rect 5441 -3487 5452 -3476
rect 11634 -3577 11645 -3531
rect 12334 -3547 12345 -3501
rect 23288 -3518 23311 -3507
rect 23425 -3518 23448 -3507
rect 12391 -3547 12402 -3536
rect 11691 -3577 11702 -3566
rect 2388 -3588 2411 -3577
rect 2525 -3588 2548 -3577
rect 13074 -3587 13085 -3541
rect 22588 -3548 22611 -3537
rect 22725 -3548 22748 -3537
rect 13131 -3587 13142 -3576
rect 20968 -3578 20991 -3567
rect 21105 -3578 21128 -3567
rect 21758 -3598 21781 -3587
rect 21895 -3598 21918 -3587
rect 2434 -3669 2445 -3623
rect 3118 -3658 3141 -3647
rect 3255 -3658 3278 -3647
rect 4598 -3658 4621 -3647
rect 4735 -3658 4758 -3647
rect 21014 -3659 21025 -3613
rect 22634 -3629 22645 -3583
rect 23334 -3599 23345 -3553
rect 24804 -3597 24815 -3551
rect 24861 -3597 24872 -3586
rect 25484 -3617 25495 -3571
rect 26284 -3597 26295 -3551
rect 26341 -3597 26352 -3586
rect 25541 -3617 25552 -3606
rect 3798 -3678 3821 -3667
rect 3935 -3678 3958 -3667
rect 21804 -3679 21815 -3633
rect 27024 -3657 27035 -3611
rect 27081 -3657 27092 -3646
rect 3164 -3739 3175 -3693
rect 3844 -3759 3855 -3713
rect 4644 -3739 4655 -3693
rect 5338 -3718 5361 -3707
rect 5475 -3718 5498 -3707
rect 5384 -3799 5395 -3753
rect 24028 -3758 24051 -3747
rect 24165 -3758 24188 -3747
rect 12288 -3778 12311 -3767
rect 12425 -3778 12448 -3767
rect 11588 -3808 11611 -3797
rect 11725 -3808 11748 -3797
rect 9968 -3838 9991 -3827
rect 10105 -3838 10128 -3827
rect 10758 -3858 10781 -3847
rect 10895 -3858 10918 -3847
rect 10014 -3919 10025 -3873
rect 11634 -3889 11645 -3843
rect 12334 -3859 12345 -3813
rect 13804 -3857 13815 -3811
rect 13861 -3857 13872 -3846
rect 14484 -3877 14495 -3831
rect 15284 -3857 15295 -3811
rect 24074 -3839 24085 -3793
rect 24758 -3828 24781 -3817
rect 24895 -3828 24918 -3817
rect 26238 -3828 26261 -3817
rect 26375 -3828 26398 -3817
rect 15341 -3857 15352 -3846
rect 25438 -3848 25461 -3837
rect 25575 -3848 25598 -3837
rect 14541 -3877 14552 -3866
rect 10804 -3939 10815 -3893
rect 16024 -3917 16035 -3871
rect 16081 -3917 16092 -3906
rect 24804 -3909 24815 -3863
rect 25484 -3929 25495 -3883
rect 26284 -3909 26295 -3863
rect 26978 -3888 27001 -3877
rect 27115 -3888 27138 -3877
rect 27024 -3969 27035 -3923
rect 13028 -4018 13051 -4007
rect 13165 -4018 13188 -4007
rect 13074 -4099 13085 -4053
rect 13758 -4088 13781 -4077
rect 13895 -4088 13918 -4077
rect 15238 -4088 15261 -4077
rect 15375 -4088 15398 -4077
rect 14438 -4108 14461 -4097
rect 14575 -4108 14598 -4097
rect 13804 -4169 13815 -4123
rect 14484 -4189 14495 -4143
rect 15284 -4169 15295 -4123
rect 15978 -4148 16001 -4137
rect 16115 -4148 16138 -4137
rect 16024 -4229 16035 -4183
use tspc_flip_flop  x1
timestamp 1755256602
transform 1 0 -1610 0 1 12060
box -70 -4500 6536 -1390
use tspc_flip_flop  x2
timestamp 1755256602
transform 1 0 -1240 0 1 6420
box -70 -4500 6536 -1390
use tspc_flip_flop  x3
timestamp 1755256602
transform 1 0 -800 0 1 570
box -70 -4500 6536 -1390
use tspc_flip_flop  x4
timestamp 1755256602
transform 1 0 10190 0 1 12180
box -70 -4500 6536 -1390
use tspc_flip_flop  x5
timestamp 1755256602
transform 1 0 9670 0 1 6600
box -70 -4500 6536 -1390
use tspc_flip_flop  x6
timestamp 1755256602
transform 1 0 9840 0 1 140
box -70 -4500 6536 -1390
use tspc_flip_flop  x7
timestamp 1755256602
transform 1 0 20920 0 1 12090
box -70 -4500 6536 -1390
use tspc_flip_flop  x8
timestamp 1755256602
transform 1 0 20140 0 1 6770
box -70 -4500 6536 -1390
use tspc_flip_flop  x9
timestamp 1755256602
transform 1 0 20840 0 1 400
box -70 -4500 6536 -1390
use tspc_flip_flop  x10
timestamp 1755256602
transform 1 0 31220 0 1 11740
box -70 -4500 6536 -1390
use tspc_flip_flop  x11
timestamp 1755256602
transform 1 0 30960 0 1 6420
box -70 -4500 6536 -1390
use tspc_flip_flop  x12
timestamp 1755256602
transform 1 0 31400 0 1 1010
box -70 -4500 6536 -1390
use tspc_flip_flop  x13
timestamp 1755256602
transform 1 0 41870 0 1 11740
box -70 -4500 6536 -1390
use tspc_flip_flop  x14
timestamp 1755256602
transform 1 0 41340 0 1 6330
box -70 -4500 6536 -1390
use tspc_flip_flop  x15
timestamp 1755256602
transform 1 0 41610 0 1 920
box -70 -4500 6536 -1390
<< end >>
