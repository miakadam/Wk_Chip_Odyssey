* NGSPICE file created from or2.ext - technology: (null)

.subckt or2 VDD VSS OUT A B
X0 OUT.t0 a_268_670 VSS.t3 VSS.t2 nfet_03v3
**devattr s=17600,576 d=17600,576
X1 OUT.t1 a_268_670 VDD.t3 VDD.t2 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X2 a_456_1390 A.t0 VDD.t7 VDD.t6 pfet_03v3
**devattr s=52800,1376 d=31200,704
X3 a_456_1390 B.t0 a_268_670 VDD.t0 pfet_03v3
**devattr s=52800,1376 d=31200,704
X4 a_268_670 B.t1 a_456_1390 VDD.t1 pfet_03v3
**devattr s=31200,704 d=52800,1376
X5 VSS.t5 A.t1 a_268_670 VSS.t4 nfet_03v3
**devattr s=17600,576 d=17600,576
X6 VDD.t5 A.t2 a_456_1390 VDD.t4 pfet_03v3
**devattr s=31200,704 d=52800,1376
X7 a_268_670 B.t2 VSS.t1 VSS.t0 nfet_03v3
**devattr s=17600,576 d=17600,576
R0 VSS.n16 VSS.n15 916555
R1 VSS.n15 VSS.t2 845.071
R2 VSS.n10 VSS.t2 845.071
R3 VSS.n9 VSS.t0 845.071
R4 VSS.n6 VSS.t0 845.071
R5 VSS.n5 VSS.t4 845.071
R6 VSS.n16 VSS.t4 845.071
R7 VSS.n10 VSS.n9 718.311
R8 VSS.n6 VSS.n5 718.311
R9 VSS.n8 VSS.n7 44.1404
R10 VSS.n17 VSS.n3 44.1404
R11 VSS.n14 VSS.n11 44.1394
R12 VSS.n2 VSS.t5 4.84702
R13 VSS.n4 VSS.t1 4.84702
R14 VSS.n12 VSS.t3 4.7885
R15 VSS.n18 VSS.n17 2.16505
R16 VSS.n14 VSS.n13 2.11983
R17 VSS.n8 VSS.n0 1.90702
R18 VSS.n15 VSS.n14 1.3005
R19 VSS.n12 VSS.n11 1.3005
R20 VSS.n11 VSS.n10 1.3005
R21 VSS.n9 VSS.n8 1.3005
R22 VSS.n7 VSS.n4 1.3005
R23 VSS.n7 VSS.n6 1.3005
R24 VSS.n3 VSS.n2 1.3005
R25 VSS.n5 VSS.n3 1.3005
R26 VSS.n17 VSS.n16 1.3005
R27 VSS.n13 VSS.n12 0.463217
R28 VSS VSS.n18 0.155672
R29 VSS VSS.n0 0.103357
R30 VSS.n13 VSS.n0 0.0909434
R31 VSS.n18 VSS.n1 0.073981
R32 VSS.n4 VSS.n1 0.0258591
R33 VSS.n2 VSS.n1 0.0258591
R34 OUT.n0 OUT.t0 9.6935
R35 OUT.n0 OUT.t1 4.35383
R36 OUT OUT.n0 0.260857
R37 VDD.n5 VDD.t2 236.083
R38 VDD.n12 VDD.t6 236.083
R39 VDD.n9 VDD.t2 235.294
R40 VDD.t1 VDD.n9 235.294
R41 VDD.n11 VDD.t0 235.294
R42 VDD.t4 VDD.n11 235.294
R43 VDD.t0 VDD.t1 200
R44 VDD.t6 VDD.t4 200
R45 VDD.n12 VDD.n2 96.0755
R46 VDD.n12 VDD.n3 96.0755
R47 VDD.n5 VDD.n4 78.2255
R48 VDD.n6 VDD.n5 78.2255
R49 VDD.n4 VDD.n2 59.8505
R50 VDD.n6 VDD.n3 59.8505
R51 VDD.n10 VDD.n2 36.2255
R52 VDD.n10 VDD.n3 36.2255
R53 VDD.n8 VDD.n4 36.2255
R54 VDD.n8 VDD.n6 36.2255
R55 VDD.n5 VDD.n0 1.99863
R56 VDD.n13 VDD.t7 1.47383
R57 VDD.n1 VDD.t5 1.47383
R58 VDD.n7 VDD.t3 1.47383
R59 VDD.n14 VDD.n13 0.864295
R60 VDD.n10 VDD.n1 0.788
R61 VDD.n11 VDD.n10 0.788
R62 VDD.n8 VDD.n7 0.788
R63 VDD.n9 VDD.n8 0.788
R64 VDD.n13 VDD.n12 0.788
R65 VDD.n14 VDD.n1 0.561043
R66 VDD.n7 VDD.n0 0.561043
R67 VDD VDD.n0 0.200451
R68 VDD VDD.n14 0.1038
R69 A.n0 A.t2 34.2311
R70 A.n0 A.t0 34.011
R71 A.n1 A.t1 19.6529
R72 A A.n1 5.05593
R73 A.n1 A.n0 0.096125
R74 B.n0 B.t1 34.2311
R75 B.n0 B.t0 34.011
R76 B.n1 B.t2 19.5066
R77 B B.n1 6.15806
R78 B.n1 B.n0 0.242375
.ends

