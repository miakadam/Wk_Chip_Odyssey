magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -2718 -29110 2718 29110
<< nmos >>
rect -2468 26900 -2068 28900
rect -1964 26900 -1564 28900
rect -1460 26900 -1060 28900
rect -956 26900 -556 28900
rect -452 26900 -52 28900
rect 52 26900 452 28900
rect 556 26900 956 28900
rect 1060 26900 1460 28900
rect 1564 26900 1964 28900
rect 2068 26900 2468 28900
rect -2468 24668 -2068 26668
rect -1964 24668 -1564 26668
rect -1460 24668 -1060 26668
rect -956 24668 -556 26668
rect -452 24668 -52 26668
rect 52 24668 452 26668
rect 556 24668 956 26668
rect 1060 24668 1460 26668
rect 1564 24668 1964 26668
rect 2068 24668 2468 26668
rect -2468 22436 -2068 24436
rect -1964 22436 -1564 24436
rect -1460 22436 -1060 24436
rect -956 22436 -556 24436
rect -452 22436 -52 24436
rect 52 22436 452 24436
rect 556 22436 956 24436
rect 1060 22436 1460 24436
rect 1564 22436 1964 24436
rect 2068 22436 2468 24436
rect -2468 20204 -2068 22204
rect -1964 20204 -1564 22204
rect -1460 20204 -1060 22204
rect -956 20204 -556 22204
rect -452 20204 -52 22204
rect 52 20204 452 22204
rect 556 20204 956 22204
rect 1060 20204 1460 22204
rect 1564 20204 1964 22204
rect 2068 20204 2468 22204
rect -2468 17972 -2068 19972
rect -1964 17972 -1564 19972
rect -1460 17972 -1060 19972
rect -956 17972 -556 19972
rect -452 17972 -52 19972
rect 52 17972 452 19972
rect 556 17972 956 19972
rect 1060 17972 1460 19972
rect 1564 17972 1964 19972
rect 2068 17972 2468 19972
rect -2468 15740 -2068 17740
rect -1964 15740 -1564 17740
rect -1460 15740 -1060 17740
rect -956 15740 -556 17740
rect -452 15740 -52 17740
rect 52 15740 452 17740
rect 556 15740 956 17740
rect 1060 15740 1460 17740
rect 1564 15740 1964 17740
rect 2068 15740 2468 17740
rect -2468 13508 -2068 15508
rect -1964 13508 -1564 15508
rect -1460 13508 -1060 15508
rect -956 13508 -556 15508
rect -452 13508 -52 15508
rect 52 13508 452 15508
rect 556 13508 956 15508
rect 1060 13508 1460 15508
rect 1564 13508 1964 15508
rect 2068 13508 2468 15508
rect -2468 11276 -2068 13276
rect -1964 11276 -1564 13276
rect -1460 11276 -1060 13276
rect -956 11276 -556 13276
rect -452 11276 -52 13276
rect 52 11276 452 13276
rect 556 11276 956 13276
rect 1060 11276 1460 13276
rect 1564 11276 1964 13276
rect 2068 11276 2468 13276
rect -2468 9044 -2068 11044
rect -1964 9044 -1564 11044
rect -1460 9044 -1060 11044
rect -956 9044 -556 11044
rect -452 9044 -52 11044
rect 52 9044 452 11044
rect 556 9044 956 11044
rect 1060 9044 1460 11044
rect 1564 9044 1964 11044
rect 2068 9044 2468 11044
rect -2468 6812 -2068 8812
rect -1964 6812 -1564 8812
rect -1460 6812 -1060 8812
rect -956 6812 -556 8812
rect -452 6812 -52 8812
rect 52 6812 452 8812
rect 556 6812 956 8812
rect 1060 6812 1460 8812
rect 1564 6812 1964 8812
rect 2068 6812 2468 8812
rect -2468 4580 -2068 6580
rect -1964 4580 -1564 6580
rect -1460 4580 -1060 6580
rect -956 4580 -556 6580
rect -452 4580 -52 6580
rect 52 4580 452 6580
rect 556 4580 956 6580
rect 1060 4580 1460 6580
rect 1564 4580 1964 6580
rect 2068 4580 2468 6580
rect -2468 2348 -2068 4348
rect -1964 2348 -1564 4348
rect -1460 2348 -1060 4348
rect -956 2348 -556 4348
rect -452 2348 -52 4348
rect 52 2348 452 4348
rect 556 2348 956 4348
rect 1060 2348 1460 4348
rect 1564 2348 1964 4348
rect 2068 2348 2468 4348
rect -2468 116 -2068 2116
rect -1964 116 -1564 2116
rect -1460 116 -1060 2116
rect -956 116 -556 2116
rect -452 116 -52 2116
rect 52 116 452 2116
rect 556 116 956 2116
rect 1060 116 1460 2116
rect 1564 116 1964 2116
rect 2068 116 2468 2116
rect -2468 -2116 -2068 -116
rect -1964 -2116 -1564 -116
rect -1460 -2116 -1060 -116
rect -956 -2116 -556 -116
rect -452 -2116 -52 -116
rect 52 -2116 452 -116
rect 556 -2116 956 -116
rect 1060 -2116 1460 -116
rect 1564 -2116 1964 -116
rect 2068 -2116 2468 -116
rect -2468 -4348 -2068 -2348
rect -1964 -4348 -1564 -2348
rect -1460 -4348 -1060 -2348
rect -956 -4348 -556 -2348
rect -452 -4348 -52 -2348
rect 52 -4348 452 -2348
rect 556 -4348 956 -2348
rect 1060 -4348 1460 -2348
rect 1564 -4348 1964 -2348
rect 2068 -4348 2468 -2348
rect -2468 -6580 -2068 -4580
rect -1964 -6580 -1564 -4580
rect -1460 -6580 -1060 -4580
rect -956 -6580 -556 -4580
rect -452 -6580 -52 -4580
rect 52 -6580 452 -4580
rect 556 -6580 956 -4580
rect 1060 -6580 1460 -4580
rect 1564 -6580 1964 -4580
rect 2068 -6580 2468 -4580
rect -2468 -8812 -2068 -6812
rect -1964 -8812 -1564 -6812
rect -1460 -8812 -1060 -6812
rect -956 -8812 -556 -6812
rect -452 -8812 -52 -6812
rect 52 -8812 452 -6812
rect 556 -8812 956 -6812
rect 1060 -8812 1460 -6812
rect 1564 -8812 1964 -6812
rect 2068 -8812 2468 -6812
rect -2468 -11044 -2068 -9044
rect -1964 -11044 -1564 -9044
rect -1460 -11044 -1060 -9044
rect -956 -11044 -556 -9044
rect -452 -11044 -52 -9044
rect 52 -11044 452 -9044
rect 556 -11044 956 -9044
rect 1060 -11044 1460 -9044
rect 1564 -11044 1964 -9044
rect 2068 -11044 2468 -9044
rect -2468 -13276 -2068 -11276
rect -1964 -13276 -1564 -11276
rect -1460 -13276 -1060 -11276
rect -956 -13276 -556 -11276
rect -452 -13276 -52 -11276
rect 52 -13276 452 -11276
rect 556 -13276 956 -11276
rect 1060 -13276 1460 -11276
rect 1564 -13276 1964 -11276
rect 2068 -13276 2468 -11276
rect -2468 -15508 -2068 -13508
rect -1964 -15508 -1564 -13508
rect -1460 -15508 -1060 -13508
rect -956 -15508 -556 -13508
rect -452 -15508 -52 -13508
rect 52 -15508 452 -13508
rect 556 -15508 956 -13508
rect 1060 -15508 1460 -13508
rect 1564 -15508 1964 -13508
rect 2068 -15508 2468 -13508
rect -2468 -17740 -2068 -15740
rect -1964 -17740 -1564 -15740
rect -1460 -17740 -1060 -15740
rect -956 -17740 -556 -15740
rect -452 -17740 -52 -15740
rect 52 -17740 452 -15740
rect 556 -17740 956 -15740
rect 1060 -17740 1460 -15740
rect 1564 -17740 1964 -15740
rect 2068 -17740 2468 -15740
rect -2468 -19972 -2068 -17972
rect -1964 -19972 -1564 -17972
rect -1460 -19972 -1060 -17972
rect -956 -19972 -556 -17972
rect -452 -19972 -52 -17972
rect 52 -19972 452 -17972
rect 556 -19972 956 -17972
rect 1060 -19972 1460 -17972
rect 1564 -19972 1964 -17972
rect 2068 -19972 2468 -17972
rect -2468 -22204 -2068 -20204
rect -1964 -22204 -1564 -20204
rect -1460 -22204 -1060 -20204
rect -956 -22204 -556 -20204
rect -452 -22204 -52 -20204
rect 52 -22204 452 -20204
rect 556 -22204 956 -20204
rect 1060 -22204 1460 -20204
rect 1564 -22204 1964 -20204
rect 2068 -22204 2468 -20204
rect -2468 -24436 -2068 -22436
rect -1964 -24436 -1564 -22436
rect -1460 -24436 -1060 -22436
rect -956 -24436 -556 -22436
rect -452 -24436 -52 -22436
rect 52 -24436 452 -22436
rect 556 -24436 956 -22436
rect 1060 -24436 1460 -22436
rect 1564 -24436 1964 -22436
rect 2068 -24436 2468 -22436
rect -2468 -26668 -2068 -24668
rect -1964 -26668 -1564 -24668
rect -1460 -26668 -1060 -24668
rect -956 -26668 -556 -24668
rect -452 -26668 -52 -24668
rect 52 -26668 452 -24668
rect 556 -26668 956 -24668
rect 1060 -26668 1460 -24668
rect 1564 -26668 1964 -24668
rect 2068 -26668 2468 -24668
rect -2468 -28900 -2068 -26900
rect -1964 -28900 -1564 -26900
rect -1460 -28900 -1060 -26900
rect -956 -28900 -556 -26900
rect -452 -28900 -52 -26900
rect 52 -28900 452 -26900
rect 556 -28900 956 -26900
rect 1060 -28900 1460 -26900
rect 1564 -28900 1964 -26900
rect 2068 -28900 2468 -26900
<< ndiff >>
rect -2556 28887 -2468 28900
rect -2556 26913 -2543 28887
rect -2497 26913 -2468 28887
rect -2556 26900 -2468 26913
rect -2068 28887 -1964 28900
rect -2068 26913 -2039 28887
rect -1993 26913 -1964 28887
rect -2068 26900 -1964 26913
rect -1564 28887 -1460 28900
rect -1564 26913 -1535 28887
rect -1489 26913 -1460 28887
rect -1564 26900 -1460 26913
rect -1060 28887 -956 28900
rect -1060 26913 -1031 28887
rect -985 26913 -956 28887
rect -1060 26900 -956 26913
rect -556 28887 -452 28900
rect -556 26913 -527 28887
rect -481 26913 -452 28887
rect -556 26900 -452 26913
rect -52 28887 52 28900
rect -52 26913 -23 28887
rect 23 26913 52 28887
rect -52 26900 52 26913
rect 452 28887 556 28900
rect 452 26913 481 28887
rect 527 26913 556 28887
rect 452 26900 556 26913
rect 956 28887 1060 28900
rect 956 26913 985 28887
rect 1031 26913 1060 28887
rect 956 26900 1060 26913
rect 1460 28887 1564 28900
rect 1460 26913 1489 28887
rect 1535 26913 1564 28887
rect 1460 26900 1564 26913
rect 1964 28887 2068 28900
rect 1964 26913 1993 28887
rect 2039 26913 2068 28887
rect 1964 26900 2068 26913
rect 2468 28887 2556 28900
rect 2468 26913 2497 28887
rect 2543 26913 2556 28887
rect 2468 26900 2556 26913
rect -2556 26655 -2468 26668
rect -2556 24681 -2543 26655
rect -2497 24681 -2468 26655
rect -2556 24668 -2468 24681
rect -2068 26655 -1964 26668
rect -2068 24681 -2039 26655
rect -1993 24681 -1964 26655
rect -2068 24668 -1964 24681
rect -1564 26655 -1460 26668
rect -1564 24681 -1535 26655
rect -1489 24681 -1460 26655
rect -1564 24668 -1460 24681
rect -1060 26655 -956 26668
rect -1060 24681 -1031 26655
rect -985 24681 -956 26655
rect -1060 24668 -956 24681
rect -556 26655 -452 26668
rect -556 24681 -527 26655
rect -481 24681 -452 26655
rect -556 24668 -452 24681
rect -52 26655 52 26668
rect -52 24681 -23 26655
rect 23 24681 52 26655
rect -52 24668 52 24681
rect 452 26655 556 26668
rect 452 24681 481 26655
rect 527 24681 556 26655
rect 452 24668 556 24681
rect 956 26655 1060 26668
rect 956 24681 985 26655
rect 1031 24681 1060 26655
rect 956 24668 1060 24681
rect 1460 26655 1564 26668
rect 1460 24681 1489 26655
rect 1535 24681 1564 26655
rect 1460 24668 1564 24681
rect 1964 26655 2068 26668
rect 1964 24681 1993 26655
rect 2039 24681 2068 26655
rect 1964 24668 2068 24681
rect 2468 26655 2556 26668
rect 2468 24681 2497 26655
rect 2543 24681 2556 26655
rect 2468 24668 2556 24681
rect -2556 24423 -2468 24436
rect -2556 22449 -2543 24423
rect -2497 22449 -2468 24423
rect -2556 22436 -2468 22449
rect -2068 24423 -1964 24436
rect -2068 22449 -2039 24423
rect -1993 22449 -1964 24423
rect -2068 22436 -1964 22449
rect -1564 24423 -1460 24436
rect -1564 22449 -1535 24423
rect -1489 22449 -1460 24423
rect -1564 22436 -1460 22449
rect -1060 24423 -956 24436
rect -1060 22449 -1031 24423
rect -985 22449 -956 24423
rect -1060 22436 -956 22449
rect -556 24423 -452 24436
rect -556 22449 -527 24423
rect -481 22449 -452 24423
rect -556 22436 -452 22449
rect -52 24423 52 24436
rect -52 22449 -23 24423
rect 23 22449 52 24423
rect -52 22436 52 22449
rect 452 24423 556 24436
rect 452 22449 481 24423
rect 527 22449 556 24423
rect 452 22436 556 22449
rect 956 24423 1060 24436
rect 956 22449 985 24423
rect 1031 22449 1060 24423
rect 956 22436 1060 22449
rect 1460 24423 1564 24436
rect 1460 22449 1489 24423
rect 1535 22449 1564 24423
rect 1460 22436 1564 22449
rect 1964 24423 2068 24436
rect 1964 22449 1993 24423
rect 2039 22449 2068 24423
rect 1964 22436 2068 22449
rect 2468 24423 2556 24436
rect 2468 22449 2497 24423
rect 2543 22449 2556 24423
rect 2468 22436 2556 22449
rect -2556 22191 -2468 22204
rect -2556 20217 -2543 22191
rect -2497 20217 -2468 22191
rect -2556 20204 -2468 20217
rect -2068 22191 -1964 22204
rect -2068 20217 -2039 22191
rect -1993 20217 -1964 22191
rect -2068 20204 -1964 20217
rect -1564 22191 -1460 22204
rect -1564 20217 -1535 22191
rect -1489 20217 -1460 22191
rect -1564 20204 -1460 20217
rect -1060 22191 -956 22204
rect -1060 20217 -1031 22191
rect -985 20217 -956 22191
rect -1060 20204 -956 20217
rect -556 22191 -452 22204
rect -556 20217 -527 22191
rect -481 20217 -452 22191
rect -556 20204 -452 20217
rect -52 22191 52 22204
rect -52 20217 -23 22191
rect 23 20217 52 22191
rect -52 20204 52 20217
rect 452 22191 556 22204
rect 452 20217 481 22191
rect 527 20217 556 22191
rect 452 20204 556 20217
rect 956 22191 1060 22204
rect 956 20217 985 22191
rect 1031 20217 1060 22191
rect 956 20204 1060 20217
rect 1460 22191 1564 22204
rect 1460 20217 1489 22191
rect 1535 20217 1564 22191
rect 1460 20204 1564 20217
rect 1964 22191 2068 22204
rect 1964 20217 1993 22191
rect 2039 20217 2068 22191
rect 1964 20204 2068 20217
rect 2468 22191 2556 22204
rect 2468 20217 2497 22191
rect 2543 20217 2556 22191
rect 2468 20204 2556 20217
rect -2556 19959 -2468 19972
rect -2556 17985 -2543 19959
rect -2497 17985 -2468 19959
rect -2556 17972 -2468 17985
rect -2068 19959 -1964 19972
rect -2068 17985 -2039 19959
rect -1993 17985 -1964 19959
rect -2068 17972 -1964 17985
rect -1564 19959 -1460 19972
rect -1564 17985 -1535 19959
rect -1489 17985 -1460 19959
rect -1564 17972 -1460 17985
rect -1060 19959 -956 19972
rect -1060 17985 -1031 19959
rect -985 17985 -956 19959
rect -1060 17972 -956 17985
rect -556 19959 -452 19972
rect -556 17985 -527 19959
rect -481 17985 -452 19959
rect -556 17972 -452 17985
rect -52 19959 52 19972
rect -52 17985 -23 19959
rect 23 17985 52 19959
rect -52 17972 52 17985
rect 452 19959 556 19972
rect 452 17985 481 19959
rect 527 17985 556 19959
rect 452 17972 556 17985
rect 956 19959 1060 19972
rect 956 17985 985 19959
rect 1031 17985 1060 19959
rect 956 17972 1060 17985
rect 1460 19959 1564 19972
rect 1460 17985 1489 19959
rect 1535 17985 1564 19959
rect 1460 17972 1564 17985
rect 1964 19959 2068 19972
rect 1964 17985 1993 19959
rect 2039 17985 2068 19959
rect 1964 17972 2068 17985
rect 2468 19959 2556 19972
rect 2468 17985 2497 19959
rect 2543 17985 2556 19959
rect 2468 17972 2556 17985
rect -2556 17727 -2468 17740
rect -2556 15753 -2543 17727
rect -2497 15753 -2468 17727
rect -2556 15740 -2468 15753
rect -2068 17727 -1964 17740
rect -2068 15753 -2039 17727
rect -1993 15753 -1964 17727
rect -2068 15740 -1964 15753
rect -1564 17727 -1460 17740
rect -1564 15753 -1535 17727
rect -1489 15753 -1460 17727
rect -1564 15740 -1460 15753
rect -1060 17727 -956 17740
rect -1060 15753 -1031 17727
rect -985 15753 -956 17727
rect -1060 15740 -956 15753
rect -556 17727 -452 17740
rect -556 15753 -527 17727
rect -481 15753 -452 17727
rect -556 15740 -452 15753
rect -52 17727 52 17740
rect -52 15753 -23 17727
rect 23 15753 52 17727
rect -52 15740 52 15753
rect 452 17727 556 17740
rect 452 15753 481 17727
rect 527 15753 556 17727
rect 452 15740 556 15753
rect 956 17727 1060 17740
rect 956 15753 985 17727
rect 1031 15753 1060 17727
rect 956 15740 1060 15753
rect 1460 17727 1564 17740
rect 1460 15753 1489 17727
rect 1535 15753 1564 17727
rect 1460 15740 1564 15753
rect 1964 17727 2068 17740
rect 1964 15753 1993 17727
rect 2039 15753 2068 17727
rect 1964 15740 2068 15753
rect 2468 17727 2556 17740
rect 2468 15753 2497 17727
rect 2543 15753 2556 17727
rect 2468 15740 2556 15753
rect -2556 15495 -2468 15508
rect -2556 13521 -2543 15495
rect -2497 13521 -2468 15495
rect -2556 13508 -2468 13521
rect -2068 15495 -1964 15508
rect -2068 13521 -2039 15495
rect -1993 13521 -1964 15495
rect -2068 13508 -1964 13521
rect -1564 15495 -1460 15508
rect -1564 13521 -1535 15495
rect -1489 13521 -1460 15495
rect -1564 13508 -1460 13521
rect -1060 15495 -956 15508
rect -1060 13521 -1031 15495
rect -985 13521 -956 15495
rect -1060 13508 -956 13521
rect -556 15495 -452 15508
rect -556 13521 -527 15495
rect -481 13521 -452 15495
rect -556 13508 -452 13521
rect -52 15495 52 15508
rect -52 13521 -23 15495
rect 23 13521 52 15495
rect -52 13508 52 13521
rect 452 15495 556 15508
rect 452 13521 481 15495
rect 527 13521 556 15495
rect 452 13508 556 13521
rect 956 15495 1060 15508
rect 956 13521 985 15495
rect 1031 13521 1060 15495
rect 956 13508 1060 13521
rect 1460 15495 1564 15508
rect 1460 13521 1489 15495
rect 1535 13521 1564 15495
rect 1460 13508 1564 13521
rect 1964 15495 2068 15508
rect 1964 13521 1993 15495
rect 2039 13521 2068 15495
rect 1964 13508 2068 13521
rect 2468 15495 2556 15508
rect 2468 13521 2497 15495
rect 2543 13521 2556 15495
rect 2468 13508 2556 13521
rect -2556 13263 -2468 13276
rect -2556 11289 -2543 13263
rect -2497 11289 -2468 13263
rect -2556 11276 -2468 11289
rect -2068 13263 -1964 13276
rect -2068 11289 -2039 13263
rect -1993 11289 -1964 13263
rect -2068 11276 -1964 11289
rect -1564 13263 -1460 13276
rect -1564 11289 -1535 13263
rect -1489 11289 -1460 13263
rect -1564 11276 -1460 11289
rect -1060 13263 -956 13276
rect -1060 11289 -1031 13263
rect -985 11289 -956 13263
rect -1060 11276 -956 11289
rect -556 13263 -452 13276
rect -556 11289 -527 13263
rect -481 11289 -452 13263
rect -556 11276 -452 11289
rect -52 13263 52 13276
rect -52 11289 -23 13263
rect 23 11289 52 13263
rect -52 11276 52 11289
rect 452 13263 556 13276
rect 452 11289 481 13263
rect 527 11289 556 13263
rect 452 11276 556 11289
rect 956 13263 1060 13276
rect 956 11289 985 13263
rect 1031 11289 1060 13263
rect 956 11276 1060 11289
rect 1460 13263 1564 13276
rect 1460 11289 1489 13263
rect 1535 11289 1564 13263
rect 1460 11276 1564 11289
rect 1964 13263 2068 13276
rect 1964 11289 1993 13263
rect 2039 11289 2068 13263
rect 1964 11276 2068 11289
rect 2468 13263 2556 13276
rect 2468 11289 2497 13263
rect 2543 11289 2556 13263
rect 2468 11276 2556 11289
rect -2556 11031 -2468 11044
rect -2556 9057 -2543 11031
rect -2497 9057 -2468 11031
rect -2556 9044 -2468 9057
rect -2068 11031 -1964 11044
rect -2068 9057 -2039 11031
rect -1993 9057 -1964 11031
rect -2068 9044 -1964 9057
rect -1564 11031 -1460 11044
rect -1564 9057 -1535 11031
rect -1489 9057 -1460 11031
rect -1564 9044 -1460 9057
rect -1060 11031 -956 11044
rect -1060 9057 -1031 11031
rect -985 9057 -956 11031
rect -1060 9044 -956 9057
rect -556 11031 -452 11044
rect -556 9057 -527 11031
rect -481 9057 -452 11031
rect -556 9044 -452 9057
rect -52 11031 52 11044
rect -52 9057 -23 11031
rect 23 9057 52 11031
rect -52 9044 52 9057
rect 452 11031 556 11044
rect 452 9057 481 11031
rect 527 9057 556 11031
rect 452 9044 556 9057
rect 956 11031 1060 11044
rect 956 9057 985 11031
rect 1031 9057 1060 11031
rect 956 9044 1060 9057
rect 1460 11031 1564 11044
rect 1460 9057 1489 11031
rect 1535 9057 1564 11031
rect 1460 9044 1564 9057
rect 1964 11031 2068 11044
rect 1964 9057 1993 11031
rect 2039 9057 2068 11031
rect 1964 9044 2068 9057
rect 2468 11031 2556 11044
rect 2468 9057 2497 11031
rect 2543 9057 2556 11031
rect 2468 9044 2556 9057
rect -2556 8799 -2468 8812
rect -2556 6825 -2543 8799
rect -2497 6825 -2468 8799
rect -2556 6812 -2468 6825
rect -2068 8799 -1964 8812
rect -2068 6825 -2039 8799
rect -1993 6825 -1964 8799
rect -2068 6812 -1964 6825
rect -1564 8799 -1460 8812
rect -1564 6825 -1535 8799
rect -1489 6825 -1460 8799
rect -1564 6812 -1460 6825
rect -1060 8799 -956 8812
rect -1060 6825 -1031 8799
rect -985 6825 -956 8799
rect -1060 6812 -956 6825
rect -556 8799 -452 8812
rect -556 6825 -527 8799
rect -481 6825 -452 8799
rect -556 6812 -452 6825
rect -52 8799 52 8812
rect -52 6825 -23 8799
rect 23 6825 52 8799
rect -52 6812 52 6825
rect 452 8799 556 8812
rect 452 6825 481 8799
rect 527 6825 556 8799
rect 452 6812 556 6825
rect 956 8799 1060 8812
rect 956 6825 985 8799
rect 1031 6825 1060 8799
rect 956 6812 1060 6825
rect 1460 8799 1564 8812
rect 1460 6825 1489 8799
rect 1535 6825 1564 8799
rect 1460 6812 1564 6825
rect 1964 8799 2068 8812
rect 1964 6825 1993 8799
rect 2039 6825 2068 8799
rect 1964 6812 2068 6825
rect 2468 8799 2556 8812
rect 2468 6825 2497 8799
rect 2543 6825 2556 8799
rect 2468 6812 2556 6825
rect -2556 6567 -2468 6580
rect -2556 4593 -2543 6567
rect -2497 4593 -2468 6567
rect -2556 4580 -2468 4593
rect -2068 6567 -1964 6580
rect -2068 4593 -2039 6567
rect -1993 4593 -1964 6567
rect -2068 4580 -1964 4593
rect -1564 6567 -1460 6580
rect -1564 4593 -1535 6567
rect -1489 4593 -1460 6567
rect -1564 4580 -1460 4593
rect -1060 6567 -956 6580
rect -1060 4593 -1031 6567
rect -985 4593 -956 6567
rect -1060 4580 -956 4593
rect -556 6567 -452 6580
rect -556 4593 -527 6567
rect -481 4593 -452 6567
rect -556 4580 -452 4593
rect -52 6567 52 6580
rect -52 4593 -23 6567
rect 23 4593 52 6567
rect -52 4580 52 4593
rect 452 6567 556 6580
rect 452 4593 481 6567
rect 527 4593 556 6567
rect 452 4580 556 4593
rect 956 6567 1060 6580
rect 956 4593 985 6567
rect 1031 4593 1060 6567
rect 956 4580 1060 4593
rect 1460 6567 1564 6580
rect 1460 4593 1489 6567
rect 1535 4593 1564 6567
rect 1460 4580 1564 4593
rect 1964 6567 2068 6580
rect 1964 4593 1993 6567
rect 2039 4593 2068 6567
rect 1964 4580 2068 4593
rect 2468 6567 2556 6580
rect 2468 4593 2497 6567
rect 2543 4593 2556 6567
rect 2468 4580 2556 4593
rect -2556 4335 -2468 4348
rect -2556 2361 -2543 4335
rect -2497 2361 -2468 4335
rect -2556 2348 -2468 2361
rect -2068 4335 -1964 4348
rect -2068 2361 -2039 4335
rect -1993 2361 -1964 4335
rect -2068 2348 -1964 2361
rect -1564 4335 -1460 4348
rect -1564 2361 -1535 4335
rect -1489 2361 -1460 4335
rect -1564 2348 -1460 2361
rect -1060 4335 -956 4348
rect -1060 2361 -1031 4335
rect -985 2361 -956 4335
rect -1060 2348 -956 2361
rect -556 4335 -452 4348
rect -556 2361 -527 4335
rect -481 2361 -452 4335
rect -556 2348 -452 2361
rect -52 4335 52 4348
rect -52 2361 -23 4335
rect 23 2361 52 4335
rect -52 2348 52 2361
rect 452 4335 556 4348
rect 452 2361 481 4335
rect 527 2361 556 4335
rect 452 2348 556 2361
rect 956 4335 1060 4348
rect 956 2361 985 4335
rect 1031 2361 1060 4335
rect 956 2348 1060 2361
rect 1460 4335 1564 4348
rect 1460 2361 1489 4335
rect 1535 2361 1564 4335
rect 1460 2348 1564 2361
rect 1964 4335 2068 4348
rect 1964 2361 1993 4335
rect 2039 2361 2068 4335
rect 1964 2348 2068 2361
rect 2468 4335 2556 4348
rect 2468 2361 2497 4335
rect 2543 2361 2556 4335
rect 2468 2348 2556 2361
rect -2556 2103 -2468 2116
rect -2556 129 -2543 2103
rect -2497 129 -2468 2103
rect -2556 116 -2468 129
rect -2068 2103 -1964 2116
rect -2068 129 -2039 2103
rect -1993 129 -1964 2103
rect -2068 116 -1964 129
rect -1564 2103 -1460 2116
rect -1564 129 -1535 2103
rect -1489 129 -1460 2103
rect -1564 116 -1460 129
rect -1060 2103 -956 2116
rect -1060 129 -1031 2103
rect -985 129 -956 2103
rect -1060 116 -956 129
rect -556 2103 -452 2116
rect -556 129 -527 2103
rect -481 129 -452 2103
rect -556 116 -452 129
rect -52 2103 52 2116
rect -52 129 -23 2103
rect 23 129 52 2103
rect -52 116 52 129
rect 452 2103 556 2116
rect 452 129 481 2103
rect 527 129 556 2103
rect 452 116 556 129
rect 956 2103 1060 2116
rect 956 129 985 2103
rect 1031 129 1060 2103
rect 956 116 1060 129
rect 1460 2103 1564 2116
rect 1460 129 1489 2103
rect 1535 129 1564 2103
rect 1460 116 1564 129
rect 1964 2103 2068 2116
rect 1964 129 1993 2103
rect 2039 129 2068 2103
rect 1964 116 2068 129
rect 2468 2103 2556 2116
rect 2468 129 2497 2103
rect 2543 129 2556 2103
rect 2468 116 2556 129
rect -2556 -129 -2468 -116
rect -2556 -2103 -2543 -129
rect -2497 -2103 -2468 -129
rect -2556 -2116 -2468 -2103
rect -2068 -129 -1964 -116
rect -2068 -2103 -2039 -129
rect -1993 -2103 -1964 -129
rect -2068 -2116 -1964 -2103
rect -1564 -129 -1460 -116
rect -1564 -2103 -1535 -129
rect -1489 -2103 -1460 -129
rect -1564 -2116 -1460 -2103
rect -1060 -129 -956 -116
rect -1060 -2103 -1031 -129
rect -985 -2103 -956 -129
rect -1060 -2116 -956 -2103
rect -556 -129 -452 -116
rect -556 -2103 -527 -129
rect -481 -2103 -452 -129
rect -556 -2116 -452 -2103
rect -52 -129 52 -116
rect -52 -2103 -23 -129
rect 23 -2103 52 -129
rect -52 -2116 52 -2103
rect 452 -129 556 -116
rect 452 -2103 481 -129
rect 527 -2103 556 -129
rect 452 -2116 556 -2103
rect 956 -129 1060 -116
rect 956 -2103 985 -129
rect 1031 -2103 1060 -129
rect 956 -2116 1060 -2103
rect 1460 -129 1564 -116
rect 1460 -2103 1489 -129
rect 1535 -2103 1564 -129
rect 1460 -2116 1564 -2103
rect 1964 -129 2068 -116
rect 1964 -2103 1993 -129
rect 2039 -2103 2068 -129
rect 1964 -2116 2068 -2103
rect 2468 -129 2556 -116
rect 2468 -2103 2497 -129
rect 2543 -2103 2556 -129
rect 2468 -2116 2556 -2103
rect -2556 -2361 -2468 -2348
rect -2556 -4335 -2543 -2361
rect -2497 -4335 -2468 -2361
rect -2556 -4348 -2468 -4335
rect -2068 -2361 -1964 -2348
rect -2068 -4335 -2039 -2361
rect -1993 -4335 -1964 -2361
rect -2068 -4348 -1964 -4335
rect -1564 -2361 -1460 -2348
rect -1564 -4335 -1535 -2361
rect -1489 -4335 -1460 -2361
rect -1564 -4348 -1460 -4335
rect -1060 -2361 -956 -2348
rect -1060 -4335 -1031 -2361
rect -985 -4335 -956 -2361
rect -1060 -4348 -956 -4335
rect -556 -2361 -452 -2348
rect -556 -4335 -527 -2361
rect -481 -4335 -452 -2361
rect -556 -4348 -452 -4335
rect -52 -2361 52 -2348
rect -52 -4335 -23 -2361
rect 23 -4335 52 -2361
rect -52 -4348 52 -4335
rect 452 -2361 556 -2348
rect 452 -4335 481 -2361
rect 527 -4335 556 -2361
rect 452 -4348 556 -4335
rect 956 -2361 1060 -2348
rect 956 -4335 985 -2361
rect 1031 -4335 1060 -2361
rect 956 -4348 1060 -4335
rect 1460 -2361 1564 -2348
rect 1460 -4335 1489 -2361
rect 1535 -4335 1564 -2361
rect 1460 -4348 1564 -4335
rect 1964 -2361 2068 -2348
rect 1964 -4335 1993 -2361
rect 2039 -4335 2068 -2361
rect 1964 -4348 2068 -4335
rect 2468 -2361 2556 -2348
rect 2468 -4335 2497 -2361
rect 2543 -4335 2556 -2361
rect 2468 -4348 2556 -4335
rect -2556 -4593 -2468 -4580
rect -2556 -6567 -2543 -4593
rect -2497 -6567 -2468 -4593
rect -2556 -6580 -2468 -6567
rect -2068 -4593 -1964 -4580
rect -2068 -6567 -2039 -4593
rect -1993 -6567 -1964 -4593
rect -2068 -6580 -1964 -6567
rect -1564 -4593 -1460 -4580
rect -1564 -6567 -1535 -4593
rect -1489 -6567 -1460 -4593
rect -1564 -6580 -1460 -6567
rect -1060 -4593 -956 -4580
rect -1060 -6567 -1031 -4593
rect -985 -6567 -956 -4593
rect -1060 -6580 -956 -6567
rect -556 -4593 -452 -4580
rect -556 -6567 -527 -4593
rect -481 -6567 -452 -4593
rect -556 -6580 -452 -6567
rect -52 -4593 52 -4580
rect -52 -6567 -23 -4593
rect 23 -6567 52 -4593
rect -52 -6580 52 -6567
rect 452 -4593 556 -4580
rect 452 -6567 481 -4593
rect 527 -6567 556 -4593
rect 452 -6580 556 -6567
rect 956 -4593 1060 -4580
rect 956 -6567 985 -4593
rect 1031 -6567 1060 -4593
rect 956 -6580 1060 -6567
rect 1460 -4593 1564 -4580
rect 1460 -6567 1489 -4593
rect 1535 -6567 1564 -4593
rect 1460 -6580 1564 -6567
rect 1964 -4593 2068 -4580
rect 1964 -6567 1993 -4593
rect 2039 -6567 2068 -4593
rect 1964 -6580 2068 -6567
rect 2468 -4593 2556 -4580
rect 2468 -6567 2497 -4593
rect 2543 -6567 2556 -4593
rect 2468 -6580 2556 -6567
rect -2556 -6825 -2468 -6812
rect -2556 -8799 -2543 -6825
rect -2497 -8799 -2468 -6825
rect -2556 -8812 -2468 -8799
rect -2068 -6825 -1964 -6812
rect -2068 -8799 -2039 -6825
rect -1993 -8799 -1964 -6825
rect -2068 -8812 -1964 -8799
rect -1564 -6825 -1460 -6812
rect -1564 -8799 -1535 -6825
rect -1489 -8799 -1460 -6825
rect -1564 -8812 -1460 -8799
rect -1060 -6825 -956 -6812
rect -1060 -8799 -1031 -6825
rect -985 -8799 -956 -6825
rect -1060 -8812 -956 -8799
rect -556 -6825 -452 -6812
rect -556 -8799 -527 -6825
rect -481 -8799 -452 -6825
rect -556 -8812 -452 -8799
rect -52 -6825 52 -6812
rect -52 -8799 -23 -6825
rect 23 -8799 52 -6825
rect -52 -8812 52 -8799
rect 452 -6825 556 -6812
rect 452 -8799 481 -6825
rect 527 -8799 556 -6825
rect 452 -8812 556 -8799
rect 956 -6825 1060 -6812
rect 956 -8799 985 -6825
rect 1031 -8799 1060 -6825
rect 956 -8812 1060 -8799
rect 1460 -6825 1564 -6812
rect 1460 -8799 1489 -6825
rect 1535 -8799 1564 -6825
rect 1460 -8812 1564 -8799
rect 1964 -6825 2068 -6812
rect 1964 -8799 1993 -6825
rect 2039 -8799 2068 -6825
rect 1964 -8812 2068 -8799
rect 2468 -6825 2556 -6812
rect 2468 -8799 2497 -6825
rect 2543 -8799 2556 -6825
rect 2468 -8812 2556 -8799
rect -2556 -9057 -2468 -9044
rect -2556 -11031 -2543 -9057
rect -2497 -11031 -2468 -9057
rect -2556 -11044 -2468 -11031
rect -2068 -9057 -1964 -9044
rect -2068 -11031 -2039 -9057
rect -1993 -11031 -1964 -9057
rect -2068 -11044 -1964 -11031
rect -1564 -9057 -1460 -9044
rect -1564 -11031 -1535 -9057
rect -1489 -11031 -1460 -9057
rect -1564 -11044 -1460 -11031
rect -1060 -9057 -956 -9044
rect -1060 -11031 -1031 -9057
rect -985 -11031 -956 -9057
rect -1060 -11044 -956 -11031
rect -556 -9057 -452 -9044
rect -556 -11031 -527 -9057
rect -481 -11031 -452 -9057
rect -556 -11044 -452 -11031
rect -52 -9057 52 -9044
rect -52 -11031 -23 -9057
rect 23 -11031 52 -9057
rect -52 -11044 52 -11031
rect 452 -9057 556 -9044
rect 452 -11031 481 -9057
rect 527 -11031 556 -9057
rect 452 -11044 556 -11031
rect 956 -9057 1060 -9044
rect 956 -11031 985 -9057
rect 1031 -11031 1060 -9057
rect 956 -11044 1060 -11031
rect 1460 -9057 1564 -9044
rect 1460 -11031 1489 -9057
rect 1535 -11031 1564 -9057
rect 1460 -11044 1564 -11031
rect 1964 -9057 2068 -9044
rect 1964 -11031 1993 -9057
rect 2039 -11031 2068 -9057
rect 1964 -11044 2068 -11031
rect 2468 -9057 2556 -9044
rect 2468 -11031 2497 -9057
rect 2543 -11031 2556 -9057
rect 2468 -11044 2556 -11031
rect -2556 -11289 -2468 -11276
rect -2556 -13263 -2543 -11289
rect -2497 -13263 -2468 -11289
rect -2556 -13276 -2468 -13263
rect -2068 -11289 -1964 -11276
rect -2068 -13263 -2039 -11289
rect -1993 -13263 -1964 -11289
rect -2068 -13276 -1964 -13263
rect -1564 -11289 -1460 -11276
rect -1564 -13263 -1535 -11289
rect -1489 -13263 -1460 -11289
rect -1564 -13276 -1460 -13263
rect -1060 -11289 -956 -11276
rect -1060 -13263 -1031 -11289
rect -985 -13263 -956 -11289
rect -1060 -13276 -956 -13263
rect -556 -11289 -452 -11276
rect -556 -13263 -527 -11289
rect -481 -13263 -452 -11289
rect -556 -13276 -452 -13263
rect -52 -11289 52 -11276
rect -52 -13263 -23 -11289
rect 23 -13263 52 -11289
rect -52 -13276 52 -13263
rect 452 -11289 556 -11276
rect 452 -13263 481 -11289
rect 527 -13263 556 -11289
rect 452 -13276 556 -13263
rect 956 -11289 1060 -11276
rect 956 -13263 985 -11289
rect 1031 -13263 1060 -11289
rect 956 -13276 1060 -13263
rect 1460 -11289 1564 -11276
rect 1460 -13263 1489 -11289
rect 1535 -13263 1564 -11289
rect 1460 -13276 1564 -13263
rect 1964 -11289 2068 -11276
rect 1964 -13263 1993 -11289
rect 2039 -13263 2068 -11289
rect 1964 -13276 2068 -13263
rect 2468 -11289 2556 -11276
rect 2468 -13263 2497 -11289
rect 2543 -13263 2556 -11289
rect 2468 -13276 2556 -13263
rect -2556 -13521 -2468 -13508
rect -2556 -15495 -2543 -13521
rect -2497 -15495 -2468 -13521
rect -2556 -15508 -2468 -15495
rect -2068 -13521 -1964 -13508
rect -2068 -15495 -2039 -13521
rect -1993 -15495 -1964 -13521
rect -2068 -15508 -1964 -15495
rect -1564 -13521 -1460 -13508
rect -1564 -15495 -1535 -13521
rect -1489 -15495 -1460 -13521
rect -1564 -15508 -1460 -15495
rect -1060 -13521 -956 -13508
rect -1060 -15495 -1031 -13521
rect -985 -15495 -956 -13521
rect -1060 -15508 -956 -15495
rect -556 -13521 -452 -13508
rect -556 -15495 -527 -13521
rect -481 -15495 -452 -13521
rect -556 -15508 -452 -15495
rect -52 -13521 52 -13508
rect -52 -15495 -23 -13521
rect 23 -15495 52 -13521
rect -52 -15508 52 -15495
rect 452 -13521 556 -13508
rect 452 -15495 481 -13521
rect 527 -15495 556 -13521
rect 452 -15508 556 -15495
rect 956 -13521 1060 -13508
rect 956 -15495 985 -13521
rect 1031 -15495 1060 -13521
rect 956 -15508 1060 -15495
rect 1460 -13521 1564 -13508
rect 1460 -15495 1489 -13521
rect 1535 -15495 1564 -13521
rect 1460 -15508 1564 -15495
rect 1964 -13521 2068 -13508
rect 1964 -15495 1993 -13521
rect 2039 -15495 2068 -13521
rect 1964 -15508 2068 -15495
rect 2468 -13521 2556 -13508
rect 2468 -15495 2497 -13521
rect 2543 -15495 2556 -13521
rect 2468 -15508 2556 -15495
rect -2556 -15753 -2468 -15740
rect -2556 -17727 -2543 -15753
rect -2497 -17727 -2468 -15753
rect -2556 -17740 -2468 -17727
rect -2068 -15753 -1964 -15740
rect -2068 -17727 -2039 -15753
rect -1993 -17727 -1964 -15753
rect -2068 -17740 -1964 -17727
rect -1564 -15753 -1460 -15740
rect -1564 -17727 -1535 -15753
rect -1489 -17727 -1460 -15753
rect -1564 -17740 -1460 -17727
rect -1060 -15753 -956 -15740
rect -1060 -17727 -1031 -15753
rect -985 -17727 -956 -15753
rect -1060 -17740 -956 -17727
rect -556 -15753 -452 -15740
rect -556 -17727 -527 -15753
rect -481 -17727 -452 -15753
rect -556 -17740 -452 -17727
rect -52 -15753 52 -15740
rect -52 -17727 -23 -15753
rect 23 -17727 52 -15753
rect -52 -17740 52 -17727
rect 452 -15753 556 -15740
rect 452 -17727 481 -15753
rect 527 -17727 556 -15753
rect 452 -17740 556 -17727
rect 956 -15753 1060 -15740
rect 956 -17727 985 -15753
rect 1031 -17727 1060 -15753
rect 956 -17740 1060 -17727
rect 1460 -15753 1564 -15740
rect 1460 -17727 1489 -15753
rect 1535 -17727 1564 -15753
rect 1460 -17740 1564 -17727
rect 1964 -15753 2068 -15740
rect 1964 -17727 1993 -15753
rect 2039 -17727 2068 -15753
rect 1964 -17740 2068 -17727
rect 2468 -15753 2556 -15740
rect 2468 -17727 2497 -15753
rect 2543 -17727 2556 -15753
rect 2468 -17740 2556 -17727
rect -2556 -17985 -2468 -17972
rect -2556 -19959 -2543 -17985
rect -2497 -19959 -2468 -17985
rect -2556 -19972 -2468 -19959
rect -2068 -17985 -1964 -17972
rect -2068 -19959 -2039 -17985
rect -1993 -19959 -1964 -17985
rect -2068 -19972 -1964 -19959
rect -1564 -17985 -1460 -17972
rect -1564 -19959 -1535 -17985
rect -1489 -19959 -1460 -17985
rect -1564 -19972 -1460 -19959
rect -1060 -17985 -956 -17972
rect -1060 -19959 -1031 -17985
rect -985 -19959 -956 -17985
rect -1060 -19972 -956 -19959
rect -556 -17985 -452 -17972
rect -556 -19959 -527 -17985
rect -481 -19959 -452 -17985
rect -556 -19972 -452 -19959
rect -52 -17985 52 -17972
rect -52 -19959 -23 -17985
rect 23 -19959 52 -17985
rect -52 -19972 52 -19959
rect 452 -17985 556 -17972
rect 452 -19959 481 -17985
rect 527 -19959 556 -17985
rect 452 -19972 556 -19959
rect 956 -17985 1060 -17972
rect 956 -19959 985 -17985
rect 1031 -19959 1060 -17985
rect 956 -19972 1060 -19959
rect 1460 -17985 1564 -17972
rect 1460 -19959 1489 -17985
rect 1535 -19959 1564 -17985
rect 1460 -19972 1564 -19959
rect 1964 -17985 2068 -17972
rect 1964 -19959 1993 -17985
rect 2039 -19959 2068 -17985
rect 1964 -19972 2068 -19959
rect 2468 -17985 2556 -17972
rect 2468 -19959 2497 -17985
rect 2543 -19959 2556 -17985
rect 2468 -19972 2556 -19959
rect -2556 -20217 -2468 -20204
rect -2556 -22191 -2543 -20217
rect -2497 -22191 -2468 -20217
rect -2556 -22204 -2468 -22191
rect -2068 -20217 -1964 -20204
rect -2068 -22191 -2039 -20217
rect -1993 -22191 -1964 -20217
rect -2068 -22204 -1964 -22191
rect -1564 -20217 -1460 -20204
rect -1564 -22191 -1535 -20217
rect -1489 -22191 -1460 -20217
rect -1564 -22204 -1460 -22191
rect -1060 -20217 -956 -20204
rect -1060 -22191 -1031 -20217
rect -985 -22191 -956 -20217
rect -1060 -22204 -956 -22191
rect -556 -20217 -452 -20204
rect -556 -22191 -527 -20217
rect -481 -22191 -452 -20217
rect -556 -22204 -452 -22191
rect -52 -20217 52 -20204
rect -52 -22191 -23 -20217
rect 23 -22191 52 -20217
rect -52 -22204 52 -22191
rect 452 -20217 556 -20204
rect 452 -22191 481 -20217
rect 527 -22191 556 -20217
rect 452 -22204 556 -22191
rect 956 -20217 1060 -20204
rect 956 -22191 985 -20217
rect 1031 -22191 1060 -20217
rect 956 -22204 1060 -22191
rect 1460 -20217 1564 -20204
rect 1460 -22191 1489 -20217
rect 1535 -22191 1564 -20217
rect 1460 -22204 1564 -22191
rect 1964 -20217 2068 -20204
rect 1964 -22191 1993 -20217
rect 2039 -22191 2068 -20217
rect 1964 -22204 2068 -22191
rect 2468 -20217 2556 -20204
rect 2468 -22191 2497 -20217
rect 2543 -22191 2556 -20217
rect 2468 -22204 2556 -22191
rect -2556 -22449 -2468 -22436
rect -2556 -24423 -2543 -22449
rect -2497 -24423 -2468 -22449
rect -2556 -24436 -2468 -24423
rect -2068 -22449 -1964 -22436
rect -2068 -24423 -2039 -22449
rect -1993 -24423 -1964 -22449
rect -2068 -24436 -1964 -24423
rect -1564 -22449 -1460 -22436
rect -1564 -24423 -1535 -22449
rect -1489 -24423 -1460 -22449
rect -1564 -24436 -1460 -24423
rect -1060 -22449 -956 -22436
rect -1060 -24423 -1031 -22449
rect -985 -24423 -956 -22449
rect -1060 -24436 -956 -24423
rect -556 -22449 -452 -22436
rect -556 -24423 -527 -22449
rect -481 -24423 -452 -22449
rect -556 -24436 -452 -24423
rect -52 -22449 52 -22436
rect -52 -24423 -23 -22449
rect 23 -24423 52 -22449
rect -52 -24436 52 -24423
rect 452 -22449 556 -22436
rect 452 -24423 481 -22449
rect 527 -24423 556 -22449
rect 452 -24436 556 -24423
rect 956 -22449 1060 -22436
rect 956 -24423 985 -22449
rect 1031 -24423 1060 -22449
rect 956 -24436 1060 -24423
rect 1460 -22449 1564 -22436
rect 1460 -24423 1489 -22449
rect 1535 -24423 1564 -22449
rect 1460 -24436 1564 -24423
rect 1964 -22449 2068 -22436
rect 1964 -24423 1993 -22449
rect 2039 -24423 2068 -22449
rect 1964 -24436 2068 -24423
rect 2468 -22449 2556 -22436
rect 2468 -24423 2497 -22449
rect 2543 -24423 2556 -22449
rect 2468 -24436 2556 -24423
rect -2556 -24681 -2468 -24668
rect -2556 -26655 -2543 -24681
rect -2497 -26655 -2468 -24681
rect -2556 -26668 -2468 -26655
rect -2068 -24681 -1964 -24668
rect -2068 -26655 -2039 -24681
rect -1993 -26655 -1964 -24681
rect -2068 -26668 -1964 -26655
rect -1564 -24681 -1460 -24668
rect -1564 -26655 -1535 -24681
rect -1489 -26655 -1460 -24681
rect -1564 -26668 -1460 -26655
rect -1060 -24681 -956 -24668
rect -1060 -26655 -1031 -24681
rect -985 -26655 -956 -24681
rect -1060 -26668 -956 -26655
rect -556 -24681 -452 -24668
rect -556 -26655 -527 -24681
rect -481 -26655 -452 -24681
rect -556 -26668 -452 -26655
rect -52 -24681 52 -24668
rect -52 -26655 -23 -24681
rect 23 -26655 52 -24681
rect -52 -26668 52 -26655
rect 452 -24681 556 -24668
rect 452 -26655 481 -24681
rect 527 -26655 556 -24681
rect 452 -26668 556 -26655
rect 956 -24681 1060 -24668
rect 956 -26655 985 -24681
rect 1031 -26655 1060 -24681
rect 956 -26668 1060 -26655
rect 1460 -24681 1564 -24668
rect 1460 -26655 1489 -24681
rect 1535 -26655 1564 -24681
rect 1460 -26668 1564 -26655
rect 1964 -24681 2068 -24668
rect 1964 -26655 1993 -24681
rect 2039 -26655 2068 -24681
rect 1964 -26668 2068 -26655
rect 2468 -24681 2556 -24668
rect 2468 -26655 2497 -24681
rect 2543 -26655 2556 -24681
rect 2468 -26668 2556 -26655
rect -2556 -26913 -2468 -26900
rect -2556 -28887 -2543 -26913
rect -2497 -28887 -2468 -26913
rect -2556 -28900 -2468 -28887
rect -2068 -26913 -1964 -26900
rect -2068 -28887 -2039 -26913
rect -1993 -28887 -1964 -26913
rect -2068 -28900 -1964 -28887
rect -1564 -26913 -1460 -26900
rect -1564 -28887 -1535 -26913
rect -1489 -28887 -1460 -26913
rect -1564 -28900 -1460 -28887
rect -1060 -26913 -956 -26900
rect -1060 -28887 -1031 -26913
rect -985 -28887 -956 -26913
rect -1060 -28900 -956 -28887
rect -556 -26913 -452 -26900
rect -556 -28887 -527 -26913
rect -481 -28887 -452 -26913
rect -556 -28900 -452 -28887
rect -52 -26913 52 -26900
rect -52 -28887 -23 -26913
rect 23 -28887 52 -26913
rect -52 -28900 52 -28887
rect 452 -26913 556 -26900
rect 452 -28887 481 -26913
rect 527 -28887 556 -26913
rect 452 -28900 556 -28887
rect 956 -26913 1060 -26900
rect 956 -28887 985 -26913
rect 1031 -28887 1060 -26913
rect 956 -28900 1060 -28887
rect 1460 -26913 1564 -26900
rect 1460 -28887 1489 -26913
rect 1535 -28887 1564 -26913
rect 1460 -28900 1564 -28887
rect 1964 -26913 2068 -26900
rect 1964 -28887 1993 -26913
rect 2039 -28887 2068 -26913
rect 1964 -28900 2068 -28887
rect 2468 -26913 2556 -26900
rect 2468 -28887 2497 -26913
rect 2543 -28887 2556 -26913
rect 2468 -28900 2556 -28887
<< ndiffc >>
rect -2543 26913 -2497 28887
rect -2039 26913 -1993 28887
rect -1535 26913 -1489 28887
rect -1031 26913 -985 28887
rect -527 26913 -481 28887
rect -23 26913 23 28887
rect 481 26913 527 28887
rect 985 26913 1031 28887
rect 1489 26913 1535 28887
rect 1993 26913 2039 28887
rect 2497 26913 2543 28887
rect -2543 24681 -2497 26655
rect -2039 24681 -1993 26655
rect -1535 24681 -1489 26655
rect -1031 24681 -985 26655
rect -527 24681 -481 26655
rect -23 24681 23 26655
rect 481 24681 527 26655
rect 985 24681 1031 26655
rect 1489 24681 1535 26655
rect 1993 24681 2039 26655
rect 2497 24681 2543 26655
rect -2543 22449 -2497 24423
rect -2039 22449 -1993 24423
rect -1535 22449 -1489 24423
rect -1031 22449 -985 24423
rect -527 22449 -481 24423
rect -23 22449 23 24423
rect 481 22449 527 24423
rect 985 22449 1031 24423
rect 1489 22449 1535 24423
rect 1993 22449 2039 24423
rect 2497 22449 2543 24423
rect -2543 20217 -2497 22191
rect -2039 20217 -1993 22191
rect -1535 20217 -1489 22191
rect -1031 20217 -985 22191
rect -527 20217 -481 22191
rect -23 20217 23 22191
rect 481 20217 527 22191
rect 985 20217 1031 22191
rect 1489 20217 1535 22191
rect 1993 20217 2039 22191
rect 2497 20217 2543 22191
rect -2543 17985 -2497 19959
rect -2039 17985 -1993 19959
rect -1535 17985 -1489 19959
rect -1031 17985 -985 19959
rect -527 17985 -481 19959
rect -23 17985 23 19959
rect 481 17985 527 19959
rect 985 17985 1031 19959
rect 1489 17985 1535 19959
rect 1993 17985 2039 19959
rect 2497 17985 2543 19959
rect -2543 15753 -2497 17727
rect -2039 15753 -1993 17727
rect -1535 15753 -1489 17727
rect -1031 15753 -985 17727
rect -527 15753 -481 17727
rect -23 15753 23 17727
rect 481 15753 527 17727
rect 985 15753 1031 17727
rect 1489 15753 1535 17727
rect 1993 15753 2039 17727
rect 2497 15753 2543 17727
rect -2543 13521 -2497 15495
rect -2039 13521 -1993 15495
rect -1535 13521 -1489 15495
rect -1031 13521 -985 15495
rect -527 13521 -481 15495
rect -23 13521 23 15495
rect 481 13521 527 15495
rect 985 13521 1031 15495
rect 1489 13521 1535 15495
rect 1993 13521 2039 15495
rect 2497 13521 2543 15495
rect -2543 11289 -2497 13263
rect -2039 11289 -1993 13263
rect -1535 11289 -1489 13263
rect -1031 11289 -985 13263
rect -527 11289 -481 13263
rect -23 11289 23 13263
rect 481 11289 527 13263
rect 985 11289 1031 13263
rect 1489 11289 1535 13263
rect 1993 11289 2039 13263
rect 2497 11289 2543 13263
rect -2543 9057 -2497 11031
rect -2039 9057 -1993 11031
rect -1535 9057 -1489 11031
rect -1031 9057 -985 11031
rect -527 9057 -481 11031
rect -23 9057 23 11031
rect 481 9057 527 11031
rect 985 9057 1031 11031
rect 1489 9057 1535 11031
rect 1993 9057 2039 11031
rect 2497 9057 2543 11031
rect -2543 6825 -2497 8799
rect -2039 6825 -1993 8799
rect -1535 6825 -1489 8799
rect -1031 6825 -985 8799
rect -527 6825 -481 8799
rect -23 6825 23 8799
rect 481 6825 527 8799
rect 985 6825 1031 8799
rect 1489 6825 1535 8799
rect 1993 6825 2039 8799
rect 2497 6825 2543 8799
rect -2543 4593 -2497 6567
rect -2039 4593 -1993 6567
rect -1535 4593 -1489 6567
rect -1031 4593 -985 6567
rect -527 4593 -481 6567
rect -23 4593 23 6567
rect 481 4593 527 6567
rect 985 4593 1031 6567
rect 1489 4593 1535 6567
rect 1993 4593 2039 6567
rect 2497 4593 2543 6567
rect -2543 2361 -2497 4335
rect -2039 2361 -1993 4335
rect -1535 2361 -1489 4335
rect -1031 2361 -985 4335
rect -527 2361 -481 4335
rect -23 2361 23 4335
rect 481 2361 527 4335
rect 985 2361 1031 4335
rect 1489 2361 1535 4335
rect 1993 2361 2039 4335
rect 2497 2361 2543 4335
rect -2543 129 -2497 2103
rect -2039 129 -1993 2103
rect -1535 129 -1489 2103
rect -1031 129 -985 2103
rect -527 129 -481 2103
rect -23 129 23 2103
rect 481 129 527 2103
rect 985 129 1031 2103
rect 1489 129 1535 2103
rect 1993 129 2039 2103
rect 2497 129 2543 2103
rect -2543 -2103 -2497 -129
rect -2039 -2103 -1993 -129
rect -1535 -2103 -1489 -129
rect -1031 -2103 -985 -129
rect -527 -2103 -481 -129
rect -23 -2103 23 -129
rect 481 -2103 527 -129
rect 985 -2103 1031 -129
rect 1489 -2103 1535 -129
rect 1993 -2103 2039 -129
rect 2497 -2103 2543 -129
rect -2543 -4335 -2497 -2361
rect -2039 -4335 -1993 -2361
rect -1535 -4335 -1489 -2361
rect -1031 -4335 -985 -2361
rect -527 -4335 -481 -2361
rect -23 -4335 23 -2361
rect 481 -4335 527 -2361
rect 985 -4335 1031 -2361
rect 1489 -4335 1535 -2361
rect 1993 -4335 2039 -2361
rect 2497 -4335 2543 -2361
rect -2543 -6567 -2497 -4593
rect -2039 -6567 -1993 -4593
rect -1535 -6567 -1489 -4593
rect -1031 -6567 -985 -4593
rect -527 -6567 -481 -4593
rect -23 -6567 23 -4593
rect 481 -6567 527 -4593
rect 985 -6567 1031 -4593
rect 1489 -6567 1535 -4593
rect 1993 -6567 2039 -4593
rect 2497 -6567 2543 -4593
rect -2543 -8799 -2497 -6825
rect -2039 -8799 -1993 -6825
rect -1535 -8799 -1489 -6825
rect -1031 -8799 -985 -6825
rect -527 -8799 -481 -6825
rect -23 -8799 23 -6825
rect 481 -8799 527 -6825
rect 985 -8799 1031 -6825
rect 1489 -8799 1535 -6825
rect 1993 -8799 2039 -6825
rect 2497 -8799 2543 -6825
rect -2543 -11031 -2497 -9057
rect -2039 -11031 -1993 -9057
rect -1535 -11031 -1489 -9057
rect -1031 -11031 -985 -9057
rect -527 -11031 -481 -9057
rect -23 -11031 23 -9057
rect 481 -11031 527 -9057
rect 985 -11031 1031 -9057
rect 1489 -11031 1535 -9057
rect 1993 -11031 2039 -9057
rect 2497 -11031 2543 -9057
rect -2543 -13263 -2497 -11289
rect -2039 -13263 -1993 -11289
rect -1535 -13263 -1489 -11289
rect -1031 -13263 -985 -11289
rect -527 -13263 -481 -11289
rect -23 -13263 23 -11289
rect 481 -13263 527 -11289
rect 985 -13263 1031 -11289
rect 1489 -13263 1535 -11289
rect 1993 -13263 2039 -11289
rect 2497 -13263 2543 -11289
rect -2543 -15495 -2497 -13521
rect -2039 -15495 -1993 -13521
rect -1535 -15495 -1489 -13521
rect -1031 -15495 -985 -13521
rect -527 -15495 -481 -13521
rect -23 -15495 23 -13521
rect 481 -15495 527 -13521
rect 985 -15495 1031 -13521
rect 1489 -15495 1535 -13521
rect 1993 -15495 2039 -13521
rect 2497 -15495 2543 -13521
rect -2543 -17727 -2497 -15753
rect -2039 -17727 -1993 -15753
rect -1535 -17727 -1489 -15753
rect -1031 -17727 -985 -15753
rect -527 -17727 -481 -15753
rect -23 -17727 23 -15753
rect 481 -17727 527 -15753
rect 985 -17727 1031 -15753
rect 1489 -17727 1535 -15753
rect 1993 -17727 2039 -15753
rect 2497 -17727 2543 -15753
rect -2543 -19959 -2497 -17985
rect -2039 -19959 -1993 -17985
rect -1535 -19959 -1489 -17985
rect -1031 -19959 -985 -17985
rect -527 -19959 -481 -17985
rect -23 -19959 23 -17985
rect 481 -19959 527 -17985
rect 985 -19959 1031 -17985
rect 1489 -19959 1535 -17985
rect 1993 -19959 2039 -17985
rect 2497 -19959 2543 -17985
rect -2543 -22191 -2497 -20217
rect -2039 -22191 -1993 -20217
rect -1535 -22191 -1489 -20217
rect -1031 -22191 -985 -20217
rect -527 -22191 -481 -20217
rect -23 -22191 23 -20217
rect 481 -22191 527 -20217
rect 985 -22191 1031 -20217
rect 1489 -22191 1535 -20217
rect 1993 -22191 2039 -20217
rect 2497 -22191 2543 -20217
rect -2543 -24423 -2497 -22449
rect -2039 -24423 -1993 -22449
rect -1535 -24423 -1489 -22449
rect -1031 -24423 -985 -22449
rect -527 -24423 -481 -22449
rect -23 -24423 23 -22449
rect 481 -24423 527 -22449
rect 985 -24423 1031 -22449
rect 1489 -24423 1535 -22449
rect 1993 -24423 2039 -22449
rect 2497 -24423 2543 -22449
rect -2543 -26655 -2497 -24681
rect -2039 -26655 -1993 -24681
rect -1535 -26655 -1489 -24681
rect -1031 -26655 -985 -24681
rect -527 -26655 -481 -24681
rect -23 -26655 23 -24681
rect 481 -26655 527 -24681
rect 985 -26655 1031 -24681
rect 1489 -26655 1535 -24681
rect 1993 -26655 2039 -24681
rect 2497 -26655 2543 -24681
rect -2543 -28887 -2497 -26913
rect -2039 -28887 -1993 -26913
rect -1535 -28887 -1489 -26913
rect -1031 -28887 -985 -26913
rect -527 -28887 -481 -26913
rect -23 -28887 23 -26913
rect 481 -28887 527 -26913
rect 985 -28887 1031 -26913
rect 1489 -28887 1535 -26913
rect 1993 -28887 2039 -26913
rect 2497 -28887 2543 -26913
<< psubdiff >>
rect -2694 29014 2694 29086
rect -2694 28970 -2622 29014
rect -2694 -28970 -2681 28970
rect -2635 -28970 -2622 28970
rect 2622 28970 2694 29014
rect -2694 -29014 -2622 -28970
rect 2622 -28970 2635 28970
rect 2681 -28970 2694 28970
rect 2622 -29014 2694 -28970
rect -2694 -29086 2694 -29014
<< psubdiffcont >>
rect -2681 -28970 -2635 28970
rect 2635 -28970 2681 28970
<< polysilicon >>
rect -2468 28979 -2068 28992
rect -2468 28933 -2455 28979
rect -2081 28933 -2068 28979
rect -2468 28900 -2068 28933
rect -1964 28979 -1564 28992
rect -1964 28933 -1951 28979
rect -1577 28933 -1564 28979
rect -1964 28900 -1564 28933
rect -1460 28979 -1060 28992
rect -1460 28933 -1447 28979
rect -1073 28933 -1060 28979
rect -1460 28900 -1060 28933
rect -956 28979 -556 28992
rect -956 28933 -943 28979
rect -569 28933 -556 28979
rect -956 28900 -556 28933
rect -452 28979 -52 28992
rect -452 28933 -439 28979
rect -65 28933 -52 28979
rect -452 28900 -52 28933
rect 52 28979 452 28992
rect 52 28933 65 28979
rect 439 28933 452 28979
rect 52 28900 452 28933
rect 556 28979 956 28992
rect 556 28933 569 28979
rect 943 28933 956 28979
rect 556 28900 956 28933
rect 1060 28979 1460 28992
rect 1060 28933 1073 28979
rect 1447 28933 1460 28979
rect 1060 28900 1460 28933
rect 1564 28979 1964 28992
rect 1564 28933 1577 28979
rect 1951 28933 1964 28979
rect 1564 28900 1964 28933
rect 2068 28979 2468 28992
rect 2068 28933 2081 28979
rect 2455 28933 2468 28979
rect 2068 28900 2468 28933
rect -2468 26867 -2068 26900
rect -2468 26821 -2455 26867
rect -2081 26821 -2068 26867
rect -2468 26808 -2068 26821
rect -1964 26867 -1564 26900
rect -1964 26821 -1951 26867
rect -1577 26821 -1564 26867
rect -1964 26808 -1564 26821
rect -1460 26867 -1060 26900
rect -1460 26821 -1447 26867
rect -1073 26821 -1060 26867
rect -1460 26808 -1060 26821
rect -956 26867 -556 26900
rect -956 26821 -943 26867
rect -569 26821 -556 26867
rect -956 26808 -556 26821
rect -452 26867 -52 26900
rect -452 26821 -439 26867
rect -65 26821 -52 26867
rect -452 26808 -52 26821
rect 52 26867 452 26900
rect 52 26821 65 26867
rect 439 26821 452 26867
rect 52 26808 452 26821
rect 556 26867 956 26900
rect 556 26821 569 26867
rect 943 26821 956 26867
rect 556 26808 956 26821
rect 1060 26867 1460 26900
rect 1060 26821 1073 26867
rect 1447 26821 1460 26867
rect 1060 26808 1460 26821
rect 1564 26867 1964 26900
rect 1564 26821 1577 26867
rect 1951 26821 1964 26867
rect 1564 26808 1964 26821
rect 2068 26867 2468 26900
rect 2068 26821 2081 26867
rect 2455 26821 2468 26867
rect 2068 26808 2468 26821
rect -2468 26747 -2068 26760
rect -2468 26701 -2455 26747
rect -2081 26701 -2068 26747
rect -2468 26668 -2068 26701
rect -1964 26747 -1564 26760
rect -1964 26701 -1951 26747
rect -1577 26701 -1564 26747
rect -1964 26668 -1564 26701
rect -1460 26747 -1060 26760
rect -1460 26701 -1447 26747
rect -1073 26701 -1060 26747
rect -1460 26668 -1060 26701
rect -956 26747 -556 26760
rect -956 26701 -943 26747
rect -569 26701 -556 26747
rect -956 26668 -556 26701
rect -452 26747 -52 26760
rect -452 26701 -439 26747
rect -65 26701 -52 26747
rect -452 26668 -52 26701
rect 52 26747 452 26760
rect 52 26701 65 26747
rect 439 26701 452 26747
rect 52 26668 452 26701
rect 556 26747 956 26760
rect 556 26701 569 26747
rect 943 26701 956 26747
rect 556 26668 956 26701
rect 1060 26747 1460 26760
rect 1060 26701 1073 26747
rect 1447 26701 1460 26747
rect 1060 26668 1460 26701
rect 1564 26747 1964 26760
rect 1564 26701 1577 26747
rect 1951 26701 1964 26747
rect 1564 26668 1964 26701
rect 2068 26747 2468 26760
rect 2068 26701 2081 26747
rect 2455 26701 2468 26747
rect 2068 26668 2468 26701
rect -2468 24635 -2068 24668
rect -2468 24589 -2455 24635
rect -2081 24589 -2068 24635
rect -2468 24576 -2068 24589
rect -1964 24635 -1564 24668
rect -1964 24589 -1951 24635
rect -1577 24589 -1564 24635
rect -1964 24576 -1564 24589
rect -1460 24635 -1060 24668
rect -1460 24589 -1447 24635
rect -1073 24589 -1060 24635
rect -1460 24576 -1060 24589
rect -956 24635 -556 24668
rect -956 24589 -943 24635
rect -569 24589 -556 24635
rect -956 24576 -556 24589
rect -452 24635 -52 24668
rect -452 24589 -439 24635
rect -65 24589 -52 24635
rect -452 24576 -52 24589
rect 52 24635 452 24668
rect 52 24589 65 24635
rect 439 24589 452 24635
rect 52 24576 452 24589
rect 556 24635 956 24668
rect 556 24589 569 24635
rect 943 24589 956 24635
rect 556 24576 956 24589
rect 1060 24635 1460 24668
rect 1060 24589 1073 24635
rect 1447 24589 1460 24635
rect 1060 24576 1460 24589
rect 1564 24635 1964 24668
rect 1564 24589 1577 24635
rect 1951 24589 1964 24635
rect 1564 24576 1964 24589
rect 2068 24635 2468 24668
rect 2068 24589 2081 24635
rect 2455 24589 2468 24635
rect 2068 24576 2468 24589
rect -2468 24515 -2068 24528
rect -2468 24469 -2455 24515
rect -2081 24469 -2068 24515
rect -2468 24436 -2068 24469
rect -1964 24515 -1564 24528
rect -1964 24469 -1951 24515
rect -1577 24469 -1564 24515
rect -1964 24436 -1564 24469
rect -1460 24515 -1060 24528
rect -1460 24469 -1447 24515
rect -1073 24469 -1060 24515
rect -1460 24436 -1060 24469
rect -956 24515 -556 24528
rect -956 24469 -943 24515
rect -569 24469 -556 24515
rect -956 24436 -556 24469
rect -452 24515 -52 24528
rect -452 24469 -439 24515
rect -65 24469 -52 24515
rect -452 24436 -52 24469
rect 52 24515 452 24528
rect 52 24469 65 24515
rect 439 24469 452 24515
rect 52 24436 452 24469
rect 556 24515 956 24528
rect 556 24469 569 24515
rect 943 24469 956 24515
rect 556 24436 956 24469
rect 1060 24515 1460 24528
rect 1060 24469 1073 24515
rect 1447 24469 1460 24515
rect 1060 24436 1460 24469
rect 1564 24515 1964 24528
rect 1564 24469 1577 24515
rect 1951 24469 1964 24515
rect 1564 24436 1964 24469
rect 2068 24515 2468 24528
rect 2068 24469 2081 24515
rect 2455 24469 2468 24515
rect 2068 24436 2468 24469
rect -2468 22403 -2068 22436
rect -2468 22357 -2455 22403
rect -2081 22357 -2068 22403
rect -2468 22344 -2068 22357
rect -1964 22403 -1564 22436
rect -1964 22357 -1951 22403
rect -1577 22357 -1564 22403
rect -1964 22344 -1564 22357
rect -1460 22403 -1060 22436
rect -1460 22357 -1447 22403
rect -1073 22357 -1060 22403
rect -1460 22344 -1060 22357
rect -956 22403 -556 22436
rect -956 22357 -943 22403
rect -569 22357 -556 22403
rect -956 22344 -556 22357
rect -452 22403 -52 22436
rect -452 22357 -439 22403
rect -65 22357 -52 22403
rect -452 22344 -52 22357
rect 52 22403 452 22436
rect 52 22357 65 22403
rect 439 22357 452 22403
rect 52 22344 452 22357
rect 556 22403 956 22436
rect 556 22357 569 22403
rect 943 22357 956 22403
rect 556 22344 956 22357
rect 1060 22403 1460 22436
rect 1060 22357 1073 22403
rect 1447 22357 1460 22403
rect 1060 22344 1460 22357
rect 1564 22403 1964 22436
rect 1564 22357 1577 22403
rect 1951 22357 1964 22403
rect 1564 22344 1964 22357
rect 2068 22403 2468 22436
rect 2068 22357 2081 22403
rect 2455 22357 2468 22403
rect 2068 22344 2468 22357
rect -2468 22283 -2068 22296
rect -2468 22237 -2455 22283
rect -2081 22237 -2068 22283
rect -2468 22204 -2068 22237
rect -1964 22283 -1564 22296
rect -1964 22237 -1951 22283
rect -1577 22237 -1564 22283
rect -1964 22204 -1564 22237
rect -1460 22283 -1060 22296
rect -1460 22237 -1447 22283
rect -1073 22237 -1060 22283
rect -1460 22204 -1060 22237
rect -956 22283 -556 22296
rect -956 22237 -943 22283
rect -569 22237 -556 22283
rect -956 22204 -556 22237
rect -452 22283 -52 22296
rect -452 22237 -439 22283
rect -65 22237 -52 22283
rect -452 22204 -52 22237
rect 52 22283 452 22296
rect 52 22237 65 22283
rect 439 22237 452 22283
rect 52 22204 452 22237
rect 556 22283 956 22296
rect 556 22237 569 22283
rect 943 22237 956 22283
rect 556 22204 956 22237
rect 1060 22283 1460 22296
rect 1060 22237 1073 22283
rect 1447 22237 1460 22283
rect 1060 22204 1460 22237
rect 1564 22283 1964 22296
rect 1564 22237 1577 22283
rect 1951 22237 1964 22283
rect 1564 22204 1964 22237
rect 2068 22283 2468 22296
rect 2068 22237 2081 22283
rect 2455 22237 2468 22283
rect 2068 22204 2468 22237
rect -2468 20171 -2068 20204
rect -2468 20125 -2455 20171
rect -2081 20125 -2068 20171
rect -2468 20112 -2068 20125
rect -1964 20171 -1564 20204
rect -1964 20125 -1951 20171
rect -1577 20125 -1564 20171
rect -1964 20112 -1564 20125
rect -1460 20171 -1060 20204
rect -1460 20125 -1447 20171
rect -1073 20125 -1060 20171
rect -1460 20112 -1060 20125
rect -956 20171 -556 20204
rect -956 20125 -943 20171
rect -569 20125 -556 20171
rect -956 20112 -556 20125
rect -452 20171 -52 20204
rect -452 20125 -439 20171
rect -65 20125 -52 20171
rect -452 20112 -52 20125
rect 52 20171 452 20204
rect 52 20125 65 20171
rect 439 20125 452 20171
rect 52 20112 452 20125
rect 556 20171 956 20204
rect 556 20125 569 20171
rect 943 20125 956 20171
rect 556 20112 956 20125
rect 1060 20171 1460 20204
rect 1060 20125 1073 20171
rect 1447 20125 1460 20171
rect 1060 20112 1460 20125
rect 1564 20171 1964 20204
rect 1564 20125 1577 20171
rect 1951 20125 1964 20171
rect 1564 20112 1964 20125
rect 2068 20171 2468 20204
rect 2068 20125 2081 20171
rect 2455 20125 2468 20171
rect 2068 20112 2468 20125
rect -2468 20051 -2068 20064
rect -2468 20005 -2455 20051
rect -2081 20005 -2068 20051
rect -2468 19972 -2068 20005
rect -1964 20051 -1564 20064
rect -1964 20005 -1951 20051
rect -1577 20005 -1564 20051
rect -1964 19972 -1564 20005
rect -1460 20051 -1060 20064
rect -1460 20005 -1447 20051
rect -1073 20005 -1060 20051
rect -1460 19972 -1060 20005
rect -956 20051 -556 20064
rect -956 20005 -943 20051
rect -569 20005 -556 20051
rect -956 19972 -556 20005
rect -452 20051 -52 20064
rect -452 20005 -439 20051
rect -65 20005 -52 20051
rect -452 19972 -52 20005
rect 52 20051 452 20064
rect 52 20005 65 20051
rect 439 20005 452 20051
rect 52 19972 452 20005
rect 556 20051 956 20064
rect 556 20005 569 20051
rect 943 20005 956 20051
rect 556 19972 956 20005
rect 1060 20051 1460 20064
rect 1060 20005 1073 20051
rect 1447 20005 1460 20051
rect 1060 19972 1460 20005
rect 1564 20051 1964 20064
rect 1564 20005 1577 20051
rect 1951 20005 1964 20051
rect 1564 19972 1964 20005
rect 2068 20051 2468 20064
rect 2068 20005 2081 20051
rect 2455 20005 2468 20051
rect 2068 19972 2468 20005
rect -2468 17939 -2068 17972
rect -2468 17893 -2455 17939
rect -2081 17893 -2068 17939
rect -2468 17880 -2068 17893
rect -1964 17939 -1564 17972
rect -1964 17893 -1951 17939
rect -1577 17893 -1564 17939
rect -1964 17880 -1564 17893
rect -1460 17939 -1060 17972
rect -1460 17893 -1447 17939
rect -1073 17893 -1060 17939
rect -1460 17880 -1060 17893
rect -956 17939 -556 17972
rect -956 17893 -943 17939
rect -569 17893 -556 17939
rect -956 17880 -556 17893
rect -452 17939 -52 17972
rect -452 17893 -439 17939
rect -65 17893 -52 17939
rect -452 17880 -52 17893
rect 52 17939 452 17972
rect 52 17893 65 17939
rect 439 17893 452 17939
rect 52 17880 452 17893
rect 556 17939 956 17972
rect 556 17893 569 17939
rect 943 17893 956 17939
rect 556 17880 956 17893
rect 1060 17939 1460 17972
rect 1060 17893 1073 17939
rect 1447 17893 1460 17939
rect 1060 17880 1460 17893
rect 1564 17939 1964 17972
rect 1564 17893 1577 17939
rect 1951 17893 1964 17939
rect 1564 17880 1964 17893
rect 2068 17939 2468 17972
rect 2068 17893 2081 17939
rect 2455 17893 2468 17939
rect 2068 17880 2468 17893
rect -2468 17819 -2068 17832
rect -2468 17773 -2455 17819
rect -2081 17773 -2068 17819
rect -2468 17740 -2068 17773
rect -1964 17819 -1564 17832
rect -1964 17773 -1951 17819
rect -1577 17773 -1564 17819
rect -1964 17740 -1564 17773
rect -1460 17819 -1060 17832
rect -1460 17773 -1447 17819
rect -1073 17773 -1060 17819
rect -1460 17740 -1060 17773
rect -956 17819 -556 17832
rect -956 17773 -943 17819
rect -569 17773 -556 17819
rect -956 17740 -556 17773
rect -452 17819 -52 17832
rect -452 17773 -439 17819
rect -65 17773 -52 17819
rect -452 17740 -52 17773
rect 52 17819 452 17832
rect 52 17773 65 17819
rect 439 17773 452 17819
rect 52 17740 452 17773
rect 556 17819 956 17832
rect 556 17773 569 17819
rect 943 17773 956 17819
rect 556 17740 956 17773
rect 1060 17819 1460 17832
rect 1060 17773 1073 17819
rect 1447 17773 1460 17819
rect 1060 17740 1460 17773
rect 1564 17819 1964 17832
rect 1564 17773 1577 17819
rect 1951 17773 1964 17819
rect 1564 17740 1964 17773
rect 2068 17819 2468 17832
rect 2068 17773 2081 17819
rect 2455 17773 2468 17819
rect 2068 17740 2468 17773
rect -2468 15707 -2068 15740
rect -2468 15661 -2455 15707
rect -2081 15661 -2068 15707
rect -2468 15648 -2068 15661
rect -1964 15707 -1564 15740
rect -1964 15661 -1951 15707
rect -1577 15661 -1564 15707
rect -1964 15648 -1564 15661
rect -1460 15707 -1060 15740
rect -1460 15661 -1447 15707
rect -1073 15661 -1060 15707
rect -1460 15648 -1060 15661
rect -956 15707 -556 15740
rect -956 15661 -943 15707
rect -569 15661 -556 15707
rect -956 15648 -556 15661
rect -452 15707 -52 15740
rect -452 15661 -439 15707
rect -65 15661 -52 15707
rect -452 15648 -52 15661
rect 52 15707 452 15740
rect 52 15661 65 15707
rect 439 15661 452 15707
rect 52 15648 452 15661
rect 556 15707 956 15740
rect 556 15661 569 15707
rect 943 15661 956 15707
rect 556 15648 956 15661
rect 1060 15707 1460 15740
rect 1060 15661 1073 15707
rect 1447 15661 1460 15707
rect 1060 15648 1460 15661
rect 1564 15707 1964 15740
rect 1564 15661 1577 15707
rect 1951 15661 1964 15707
rect 1564 15648 1964 15661
rect 2068 15707 2468 15740
rect 2068 15661 2081 15707
rect 2455 15661 2468 15707
rect 2068 15648 2468 15661
rect -2468 15587 -2068 15600
rect -2468 15541 -2455 15587
rect -2081 15541 -2068 15587
rect -2468 15508 -2068 15541
rect -1964 15587 -1564 15600
rect -1964 15541 -1951 15587
rect -1577 15541 -1564 15587
rect -1964 15508 -1564 15541
rect -1460 15587 -1060 15600
rect -1460 15541 -1447 15587
rect -1073 15541 -1060 15587
rect -1460 15508 -1060 15541
rect -956 15587 -556 15600
rect -956 15541 -943 15587
rect -569 15541 -556 15587
rect -956 15508 -556 15541
rect -452 15587 -52 15600
rect -452 15541 -439 15587
rect -65 15541 -52 15587
rect -452 15508 -52 15541
rect 52 15587 452 15600
rect 52 15541 65 15587
rect 439 15541 452 15587
rect 52 15508 452 15541
rect 556 15587 956 15600
rect 556 15541 569 15587
rect 943 15541 956 15587
rect 556 15508 956 15541
rect 1060 15587 1460 15600
rect 1060 15541 1073 15587
rect 1447 15541 1460 15587
rect 1060 15508 1460 15541
rect 1564 15587 1964 15600
rect 1564 15541 1577 15587
rect 1951 15541 1964 15587
rect 1564 15508 1964 15541
rect 2068 15587 2468 15600
rect 2068 15541 2081 15587
rect 2455 15541 2468 15587
rect 2068 15508 2468 15541
rect -2468 13475 -2068 13508
rect -2468 13429 -2455 13475
rect -2081 13429 -2068 13475
rect -2468 13416 -2068 13429
rect -1964 13475 -1564 13508
rect -1964 13429 -1951 13475
rect -1577 13429 -1564 13475
rect -1964 13416 -1564 13429
rect -1460 13475 -1060 13508
rect -1460 13429 -1447 13475
rect -1073 13429 -1060 13475
rect -1460 13416 -1060 13429
rect -956 13475 -556 13508
rect -956 13429 -943 13475
rect -569 13429 -556 13475
rect -956 13416 -556 13429
rect -452 13475 -52 13508
rect -452 13429 -439 13475
rect -65 13429 -52 13475
rect -452 13416 -52 13429
rect 52 13475 452 13508
rect 52 13429 65 13475
rect 439 13429 452 13475
rect 52 13416 452 13429
rect 556 13475 956 13508
rect 556 13429 569 13475
rect 943 13429 956 13475
rect 556 13416 956 13429
rect 1060 13475 1460 13508
rect 1060 13429 1073 13475
rect 1447 13429 1460 13475
rect 1060 13416 1460 13429
rect 1564 13475 1964 13508
rect 1564 13429 1577 13475
rect 1951 13429 1964 13475
rect 1564 13416 1964 13429
rect 2068 13475 2468 13508
rect 2068 13429 2081 13475
rect 2455 13429 2468 13475
rect 2068 13416 2468 13429
rect -2468 13355 -2068 13368
rect -2468 13309 -2455 13355
rect -2081 13309 -2068 13355
rect -2468 13276 -2068 13309
rect -1964 13355 -1564 13368
rect -1964 13309 -1951 13355
rect -1577 13309 -1564 13355
rect -1964 13276 -1564 13309
rect -1460 13355 -1060 13368
rect -1460 13309 -1447 13355
rect -1073 13309 -1060 13355
rect -1460 13276 -1060 13309
rect -956 13355 -556 13368
rect -956 13309 -943 13355
rect -569 13309 -556 13355
rect -956 13276 -556 13309
rect -452 13355 -52 13368
rect -452 13309 -439 13355
rect -65 13309 -52 13355
rect -452 13276 -52 13309
rect 52 13355 452 13368
rect 52 13309 65 13355
rect 439 13309 452 13355
rect 52 13276 452 13309
rect 556 13355 956 13368
rect 556 13309 569 13355
rect 943 13309 956 13355
rect 556 13276 956 13309
rect 1060 13355 1460 13368
rect 1060 13309 1073 13355
rect 1447 13309 1460 13355
rect 1060 13276 1460 13309
rect 1564 13355 1964 13368
rect 1564 13309 1577 13355
rect 1951 13309 1964 13355
rect 1564 13276 1964 13309
rect 2068 13355 2468 13368
rect 2068 13309 2081 13355
rect 2455 13309 2468 13355
rect 2068 13276 2468 13309
rect -2468 11243 -2068 11276
rect -2468 11197 -2455 11243
rect -2081 11197 -2068 11243
rect -2468 11184 -2068 11197
rect -1964 11243 -1564 11276
rect -1964 11197 -1951 11243
rect -1577 11197 -1564 11243
rect -1964 11184 -1564 11197
rect -1460 11243 -1060 11276
rect -1460 11197 -1447 11243
rect -1073 11197 -1060 11243
rect -1460 11184 -1060 11197
rect -956 11243 -556 11276
rect -956 11197 -943 11243
rect -569 11197 -556 11243
rect -956 11184 -556 11197
rect -452 11243 -52 11276
rect -452 11197 -439 11243
rect -65 11197 -52 11243
rect -452 11184 -52 11197
rect 52 11243 452 11276
rect 52 11197 65 11243
rect 439 11197 452 11243
rect 52 11184 452 11197
rect 556 11243 956 11276
rect 556 11197 569 11243
rect 943 11197 956 11243
rect 556 11184 956 11197
rect 1060 11243 1460 11276
rect 1060 11197 1073 11243
rect 1447 11197 1460 11243
rect 1060 11184 1460 11197
rect 1564 11243 1964 11276
rect 1564 11197 1577 11243
rect 1951 11197 1964 11243
rect 1564 11184 1964 11197
rect 2068 11243 2468 11276
rect 2068 11197 2081 11243
rect 2455 11197 2468 11243
rect 2068 11184 2468 11197
rect -2468 11123 -2068 11136
rect -2468 11077 -2455 11123
rect -2081 11077 -2068 11123
rect -2468 11044 -2068 11077
rect -1964 11123 -1564 11136
rect -1964 11077 -1951 11123
rect -1577 11077 -1564 11123
rect -1964 11044 -1564 11077
rect -1460 11123 -1060 11136
rect -1460 11077 -1447 11123
rect -1073 11077 -1060 11123
rect -1460 11044 -1060 11077
rect -956 11123 -556 11136
rect -956 11077 -943 11123
rect -569 11077 -556 11123
rect -956 11044 -556 11077
rect -452 11123 -52 11136
rect -452 11077 -439 11123
rect -65 11077 -52 11123
rect -452 11044 -52 11077
rect 52 11123 452 11136
rect 52 11077 65 11123
rect 439 11077 452 11123
rect 52 11044 452 11077
rect 556 11123 956 11136
rect 556 11077 569 11123
rect 943 11077 956 11123
rect 556 11044 956 11077
rect 1060 11123 1460 11136
rect 1060 11077 1073 11123
rect 1447 11077 1460 11123
rect 1060 11044 1460 11077
rect 1564 11123 1964 11136
rect 1564 11077 1577 11123
rect 1951 11077 1964 11123
rect 1564 11044 1964 11077
rect 2068 11123 2468 11136
rect 2068 11077 2081 11123
rect 2455 11077 2468 11123
rect 2068 11044 2468 11077
rect -2468 9011 -2068 9044
rect -2468 8965 -2455 9011
rect -2081 8965 -2068 9011
rect -2468 8952 -2068 8965
rect -1964 9011 -1564 9044
rect -1964 8965 -1951 9011
rect -1577 8965 -1564 9011
rect -1964 8952 -1564 8965
rect -1460 9011 -1060 9044
rect -1460 8965 -1447 9011
rect -1073 8965 -1060 9011
rect -1460 8952 -1060 8965
rect -956 9011 -556 9044
rect -956 8965 -943 9011
rect -569 8965 -556 9011
rect -956 8952 -556 8965
rect -452 9011 -52 9044
rect -452 8965 -439 9011
rect -65 8965 -52 9011
rect -452 8952 -52 8965
rect 52 9011 452 9044
rect 52 8965 65 9011
rect 439 8965 452 9011
rect 52 8952 452 8965
rect 556 9011 956 9044
rect 556 8965 569 9011
rect 943 8965 956 9011
rect 556 8952 956 8965
rect 1060 9011 1460 9044
rect 1060 8965 1073 9011
rect 1447 8965 1460 9011
rect 1060 8952 1460 8965
rect 1564 9011 1964 9044
rect 1564 8965 1577 9011
rect 1951 8965 1964 9011
rect 1564 8952 1964 8965
rect 2068 9011 2468 9044
rect 2068 8965 2081 9011
rect 2455 8965 2468 9011
rect 2068 8952 2468 8965
rect -2468 8891 -2068 8904
rect -2468 8845 -2455 8891
rect -2081 8845 -2068 8891
rect -2468 8812 -2068 8845
rect -1964 8891 -1564 8904
rect -1964 8845 -1951 8891
rect -1577 8845 -1564 8891
rect -1964 8812 -1564 8845
rect -1460 8891 -1060 8904
rect -1460 8845 -1447 8891
rect -1073 8845 -1060 8891
rect -1460 8812 -1060 8845
rect -956 8891 -556 8904
rect -956 8845 -943 8891
rect -569 8845 -556 8891
rect -956 8812 -556 8845
rect -452 8891 -52 8904
rect -452 8845 -439 8891
rect -65 8845 -52 8891
rect -452 8812 -52 8845
rect 52 8891 452 8904
rect 52 8845 65 8891
rect 439 8845 452 8891
rect 52 8812 452 8845
rect 556 8891 956 8904
rect 556 8845 569 8891
rect 943 8845 956 8891
rect 556 8812 956 8845
rect 1060 8891 1460 8904
rect 1060 8845 1073 8891
rect 1447 8845 1460 8891
rect 1060 8812 1460 8845
rect 1564 8891 1964 8904
rect 1564 8845 1577 8891
rect 1951 8845 1964 8891
rect 1564 8812 1964 8845
rect 2068 8891 2468 8904
rect 2068 8845 2081 8891
rect 2455 8845 2468 8891
rect 2068 8812 2468 8845
rect -2468 6779 -2068 6812
rect -2468 6733 -2455 6779
rect -2081 6733 -2068 6779
rect -2468 6720 -2068 6733
rect -1964 6779 -1564 6812
rect -1964 6733 -1951 6779
rect -1577 6733 -1564 6779
rect -1964 6720 -1564 6733
rect -1460 6779 -1060 6812
rect -1460 6733 -1447 6779
rect -1073 6733 -1060 6779
rect -1460 6720 -1060 6733
rect -956 6779 -556 6812
rect -956 6733 -943 6779
rect -569 6733 -556 6779
rect -956 6720 -556 6733
rect -452 6779 -52 6812
rect -452 6733 -439 6779
rect -65 6733 -52 6779
rect -452 6720 -52 6733
rect 52 6779 452 6812
rect 52 6733 65 6779
rect 439 6733 452 6779
rect 52 6720 452 6733
rect 556 6779 956 6812
rect 556 6733 569 6779
rect 943 6733 956 6779
rect 556 6720 956 6733
rect 1060 6779 1460 6812
rect 1060 6733 1073 6779
rect 1447 6733 1460 6779
rect 1060 6720 1460 6733
rect 1564 6779 1964 6812
rect 1564 6733 1577 6779
rect 1951 6733 1964 6779
rect 1564 6720 1964 6733
rect 2068 6779 2468 6812
rect 2068 6733 2081 6779
rect 2455 6733 2468 6779
rect 2068 6720 2468 6733
rect -2468 6659 -2068 6672
rect -2468 6613 -2455 6659
rect -2081 6613 -2068 6659
rect -2468 6580 -2068 6613
rect -1964 6659 -1564 6672
rect -1964 6613 -1951 6659
rect -1577 6613 -1564 6659
rect -1964 6580 -1564 6613
rect -1460 6659 -1060 6672
rect -1460 6613 -1447 6659
rect -1073 6613 -1060 6659
rect -1460 6580 -1060 6613
rect -956 6659 -556 6672
rect -956 6613 -943 6659
rect -569 6613 -556 6659
rect -956 6580 -556 6613
rect -452 6659 -52 6672
rect -452 6613 -439 6659
rect -65 6613 -52 6659
rect -452 6580 -52 6613
rect 52 6659 452 6672
rect 52 6613 65 6659
rect 439 6613 452 6659
rect 52 6580 452 6613
rect 556 6659 956 6672
rect 556 6613 569 6659
rect 943 6613 956 6659
rect 556 6580 956 6613
rect 1060 6659 1460 6672
rect 1060 6613 1073 6659
rect 1447 6613 1460 6659
rect 1060 6580 1460 6613
rect 1564 6659 1964 6672
rect 1564 6613 1577 6659
rect 1951 6613 1964 6659
rect 1564 6580 1964 6613
rect 2068 6659 2468 6672
rect 2068 6613 2081 6659
rect 2455 6613 2468 6659
rect 2068 6580 2468 6613
rect -2468 4547 -2068 4580
rect -2468 4501 -2455 4547
rect -2081 4501 -2068 4547
rect -2468 4488 -2068 4501
rect -1964 4547 -1564 4580
rect -1964 4501 -1951 4547
rect -1577 4501 -1564 4547
rect -1964 4488 -1564 4501
rect -1460 4547 -1060 4580
rect -1460 4501 -1447 4547
rect -1073 4501 -1060 4547
rect -1460 4488 -1060 4501
rect -956 4547 -556 4580
rect -956 4501 -943 4547
rect -569 4501 -556 4547
rect -956 4488 -556 4501
rect -452 4547 -52 4580
rect -452 4501 -439 4547
rect -65 4501 -52 4547
rect -452 4488 -52 4501
rect 52 4547 452 4580
rect 52 4501 65 4547
rect 439 4501 452 4547
rect 52 4488 452 4501
rect 556 4547 956 4580
rect 556 4501 569 4547
rect 943 4501 956 4547
rect 556 4488 956 4501
rect 1060 4547 1460 4580
rect 1060 4501 1073 4547
rect 1447 4501 1460 4547
rect 1060 4488 1460 4501
rect 1564 4547 1964 4580
rect 1564 4501 1577 4547
rect 1951 4501 1964 4547
rect 1564 4488 1964 4501
rect 2068 4547 2468 4580
rect 2068 4501 2081 4547
rect 2455 4501 2468 4547
rect 2068 4488 2468 4501
rect -2468 4427 -2068 4440
rect -2468 4381 -2455 4427
rect -2081 4381 -2068 4427
rect -2468 4348 -2068 4381
rect -1964 4427 -1564 4440
rect -1964 4381 -1951 4427
rect -1577 4381 -1564 4427
rect -1964 4348 -1564 4381
rect -1460 4427 -1060 4440
rect -1460 4381 -1447 4427
rect -1073 4381 -1060 4427
rect -1460 4348 -1060 4381
rect -956 4427 -556 4440
rect -956 4381 -943 4427
rect -569 4381 -556 4427
rect -956 4348 -556 4381
rect -452 4427 -52 4440
rect -452 4381 -439 4427
rect -65 4381 -52 4427
rect -452 4348 -52 4381
rect 52 4427 452 4440
rect 52 4381 65 4427
rect 439 4381 452 4427
rect 52 4348 452 4381
rect 556 4427 956 4440
rect 556 4381 569 4427
rect 943 4381 956 4427
rect 556 4348 956 4381
rect 1060 4427 1460 4440
rect 1060 4381 1073 4427
rect 1447 4381 1460 4427
rect 1060 4348 1460 4381
rect 1564 4427 1964 4440
rect 1564 4381 1577 4427
rect 1951 4381 1964 4427
rect 1564 4348 1964 4381
rect 2068 4427 2468 4440
rect 2068 4381 2081 4427
rect 2455 4381 2468 4427
rect 2068 4348 2468 4381
rect -2468 2315 -2068 2348
rect -2468 2269 -2455 2315
rect -2081 2269 -2068 2315
rect -2468 2256 -2068 2269
rect -1964 2315 -1564 2348
rect -1964 2269 -1951 2315
rect -1577 2269 -1564 2315
rect -1964 2256 -1564 2269
rect -1460 2315 -1060 2348
rect -1460 2269 -1447 2315
rect -1073 2269 -1060 2315
rect -1460 2256 -1060 2269
rect -956 2315 -556 2348
rect -956 2269 -943 2315
rect -569 2269 -556 2315
rect -956 2256 -556 2269
rect -452 2315 -52 2348
rect -452 2269 -439 2315
rect -65 2269 -52 2315
rect -452 2256 -52 2269
rect 52 2315 452 2348
rect 52 2269 65 2315
rect 439 2269 452 2315
rect 52 2256 452 2269
rect 556 2315 956 2348
rect 556 2269 569 2315
rect 943 2269 956 2315
rect 556 2256 956 2269
rect 1060 2315 1460 2348
rect 1060 2269 1073 2315
rect 1447 2269 1460 2315
rect 1060 2256 1460 2269
rect 1564 2315 1964 2348
rect 1564 2269 1577 2315
rect 1951 2269 1964 2315
rect 1564 2256 1964 2269
rect 2068 2315 2468 2348
rect 2068 2269 2081 2315
rect 2455 2269 2468 2315
rect 2068 2256 2468 2269
rect -2468 2195 -2068 2208
rect -2468 2149 -2455 2195
rect -2081 2149 -2068 2195
rect -2468 2116 -2068 2149
rect -1964 2195 -1564 2208
rect -1964 2149 -1951 2195
rect -1577 2149 -1564 2195
rect -1964 2116 -1564 2149
rect -1460 2195 -1060 2208
rect -1460 2149 -1447 2195
rect -1073 2149 -1060 2195
rect -1460 2116 -1060 2149
rect -956 2195 -556 2208
rect -956 2149 -943 2195
rect -569 2149 -556 2195
rect -956 2116 -556 2149
rect -452 2195 -52 2208
rect -452 2149 -439 2195
rect -65 2149 -52 2195
rect -452 2116 -52 2149
rect 52 2195 452 2208
rect 52 2149 65 2195
rect 439 2149 452 2195
rect 52 2116 452 2149
rect 556 2195 956 2208
rect 556 2149 569 2195
rect 943 2149 956 2195
rect 556 2116 956 2149
rect 1060 2195 1460 2208
rect 1060 2149 1073 2195
rect 1447 2149 1460 2195
rect 1060 2116 1460 2149
rect 1564 2195 1964 2208
rect 1564 2149 1577 2195
rect 1951 2149 1964 2195
rect 1564 2116 1964 2149
rect 2068 2195 2468 2208
rect 2068 2149 2081 2195
rect 2455 2149 2468 2195
rect 2068 2116 2468 2149
rect -2468 83 -2068 116
rect -2468 37 -2455 83
rect -2081 37 -2068 83
rect -2468 24 -2068 37
rect -1964 83 -1564 116
rect -1964 37 -1951 83
rect -1577 37 -1564 83
rect -1964 24 -1564 37
rect -1460 83 -1060 116
rect -1460 37 -1447 83
rect -1073 37 -1060 83
rect -1460 24 -1060 37
rect -956 83 -556 116
rect -956 37 -943 83
rect -569 37 -556 83
rect -956 24 -556 37
rect -452 83 -52 116
rect -452 37 -439 83
rect -65 37 -52 83
rect -452 24 -52 37
rect 52 83 452 116
rect 52 37 65 83
rect 439 37 452 83
rect 52 24 452 37
rect 556 83 956 116
rect 556 37 569 83
rect 943 37 956 83
rect 556 24 956 37
rect 1060 83 1460 116
rect 1060 37 1073 83
rect 1447 37 1460 83
rect 1060 24 1460 37
rect 1564 83 1964 116
rect 1564 37 1577 83
rect 1951 37 1964 83
rect 1564 24 1964 37
rect 2068 83 2468 116
rect 2068 37 2081 83
rect 2455 37 2468 83
rect 2068 24 2468 37
rect -2468 -37 -2068 -24
rect -2468 -83 -2455 -37
rect -2081 -83 -2068 -37
rect -2468 -116 -2068 -83
rect -1964 -37 -1564 -24
rect -1964 -83 -1951 -37
rect -1577 -83 -1564 -37
rect -1964 -116 -1564 -83
rect -1460 -37 -1060 -24
rect -1460 -83 -1447 -37
rect -1073 -83 -1060 -37
rect -1460 -116 -1060 -83
rect -956 -37 -556 -24
rect -956 -83 -943 -37
rect -569 -83 -556 -37
rect -956 -116 -556 -83
rect -452 -37 -52 -24
rect -452 -83 -439 -37
rect -65 -83 -52 -37
rect -452 -116 -52 -83
rect 52 -37 452 -24
rect 52 -83 65 -37
rect 439 -83 452 -37
rect 52 -116 452 -83
rect 556 -37 956 -24
rect 556 -83 569 -37
rect 943 -83 956 -37
rect 556 -116 956 -83
rect 1060 -37 1460 -24
rect 1060 -83 1073 -37
rect 1447 -83 1460 -37
rect 1060 -116 1460 -83
rect 1564 -37 1964 -24
rect 1564 -83 1577 -37
rect 1951 -83 1964 -37
rect 1564 -116 1964 -83
rect 2068 -37 2468 -24
rect 2068 -83 2081 -37
rect 2455 -83 2468 -37
rect 2068 -116 2468 -83
rect -2468 -2149 -2068 -2116
rect -2468 -2195 -2455 -2149
rect -2081 -2195 -2068 -2149
rect -2468 -2208 -2068 -2195
rect -1964 -2149 -1564 -2116
rect -1964 -2195 -1951 -2149
rect -1577 -2195 -1564 -2149
rect -1964 -2208 -1564 -2195
rect -1460 -2149 -1060 -2116
rect -1460 -2195 -1447 -2149
rect -1073 -2195 -1060 -2149
rect -1460 -2208 -1060 -2195
rect -956 -2149 -556 -2116
rect -956 -2195 -943 -2149
rect -569 -2195 -556 -2149
rect -956 -2208 -556 -2195
rect -452 -2149 -52 -2116
rect -452 -2195 -439 -2149
rect -65 -2195 -52 -2149
rect -452 -2208 -52 -2195
rect 52 -2149 452 -2116
rect 52 -2195 65 -2149
rect 439 -2195 452 -2149
rect 52 -2208 452 -2195
rect 556 -2149 956 -2116
rect 556 -2195 569 -2149
rect 943 -2195 956 -2149
rect 556 -2208 956 -2195
rect 1060 -2149 1460 -2116
rect 1060 -2195 1073 -2149
rect 1447 -2195 1460 -2149
rect 1060 -2208 1460 -2195
rect 1564 -2149 1964 -2116
rect 1564 -2195 1577 -2149
rect 1951 -2195 1964 -2149
rect 1564 -2208 1964 -2195
rect 2068 -2149 2468 -2116
rect 2068 -2195 2081 -2149
rect 2455 -2195 2468 -2149
rect 2068 -2208 2468 -2195
rect -2468 -2269 -2068 -2256
rect -2468 -2315 -2455 -2269
rect -2081 -2315 -2068 -2269
rect -2468 -2348 -2068 -2315
rect -1964 -2269 -1564 -2256
rect -1964 -2315 -1951 -2269
rect -1577 -2315 -1564 -2269
rect -1964 -2348 -1564 -2315
rect -1460 -2269 -1060 -2256
rect -1460 -2315 -1447 -2269
rect -1073 -2315 -1060 -2269
rect -1460 -2348 -1060 -2315
rect -956 -2269 -556 -2256
rect -956 -2315 -943 -2269
rect -569 -2315 -556 -2269
rect -956 -2348 -556 -2315
rect -452 -2269 -52 -2256
rect -452 -2315 -439 -2269
rect -65 -2315 -52 -2269
rect -452 -2348 -52 -2315
rect 52 -2269 452 -2256
rect 52 -2315 65 -2269
rect 439 -2315 452 -2269
rect 52 -2348 452 -2315
rect 556 -2269 956 -2256
rect 556 -2315 569 -2269
rect 943 -2315 956 -2269
rect 556 -2348 956 -2315
rect 1060 -2269 1460 -2256
rect 1060 -2315 1073 -2269
rect 1447 -2315 1460 -2269
rect 1060 -2348 1460 -2315
rect 1564 -2269 1964 -2256
rect 1564 -2315 1577 -2269
rect 1951 -2315 1964 -2269
rect 1564 -2348 1964 -2315
rect 2068 -2269 2468 -2256
rect 2068 -2315 2081 -2269
rect 2455 -2315 2468 -2269
rect 2068 -2348 2468 -2315
rect -2468 -4381 -2068 -4348
rect -2468 -4427 -2455 -4381
rect -2081 -4427 -2068 -4381
rect -2468 -4440 -2068 -4427
rect -1964 -4381 -1564 -4348
rect -1964 -4427 -1951 -4381
rect -1577 -4427 -1564 -4381
rect -1964 -4440 -1564 -4427
rect -1460 -4381 -1060 -4348
rect -1460 -4427 -1447 -4381
rect -1073 -4427 -1060 -4381
rect -1460 -4440 -1060 -4427
rect -956 -4381 -556 -4348
rect -956 -4427 -943 -4381
rect -569 -4427 -556 -4381
rect -956 -4440 -556 -4427
rect -452 -4381 -52 -4348
rect -452 -4427 -439 -4381
rect -65 -4427 -52 -4381
rect -452 -4440 -52 -4427
rect 52 -4381 452 -4348
rect 52 -4427 65 -4381
rect 439 -4427 452 -4381
rect 52 -4440 452 -4427
rect 556 -4381 956 -4348
rect 556 -4427 569 -4381
rect 943 -4427 956 -4381
rect 556 -4440 956 -4427
rect 1060 -4381 1460 -4348
rect 1060 -4427 1073 -4381
rect 1447 -4427 1460 -4381
rect 1060 -4440 1460 -4427
rect 1564 -4381 1964 -4348
rect 1564 -4427 1577 -4381
rect 1951 -4427 1964 -4381
rect 1564 -4440 1964 -4427
rect 2068 -4381 2468 -4348
rect 2068 -4427 2081 -4381
rect 2455 -4427 2468 -4381
rect 2068 -4440 2468 -4427
rect -2468 -4501 -2068 -4488
rect -2468 -4547 -2455 -4501
rect -2081 -4547 -2068 -4501
rect -2468 -4580 -2068 -4547
rect -1964 -4501 -1564 -4488
rect -1964 -4547 -1951 -4501
rect -1577 -4547 -1564 -4501
rect -1964 -4580 -1564 -4547
rect -1460 -4501 -1060 -4488
rect -1460 -4547 -1447 -4501
rect -1073 -4547 -1060 -4501
rect -1460 -4580 -1060 -4547
rect -956 -4501 -556 -4488
rect -956 -4547 -943 -4501
rect -569 -4547 -556 -4501
rect -956 -4580 -556 -4547
rect -452 -4501 -52 -4488
rect -452 -4547 -439 -4501
rect -65 -4547 -52 -4501
rect -452 -4580 -52 -4547
rect 52 -4501 452 -4488
rect 52 -4547 65 -4501
rect 439 -4547 452 -4501
rect 52 -4580 452 -4547
rect 556 -4501 956 -4488
rect 556 -4547 569 -4501
rect 943 -4547 956 -4501
rect 556 -4580 956 -4547
rect 1060 -4501 1460 -4488
rect 1060 -4547 1073 -4501
rect 1447 -4547 1460 -4501
rect 1060 -4580 1460 -4547
rect 1564 -4501 1964 -4488
rect 1564 -4547 1577 -4501
rect 1951 -4547 1964 -4501
rect 1564 -4580 1964 -4547
rect 2068 -4501 2468 -4488
rect 2068 -4547 2081 -4501
rect 2455 -4547 2468 -4501
rect 2068 -4580 2468 -4547
rect -2468 -6613 -2068 -6580
rect -2468 -6659 -2455 -6613
rect -2081 -6659 -2068 -6613
rect -2468 -6672 -2068 -6659
rect -1964 -6613 -1564 -6580
rect -1964 -6659 -1951 -6613
rect -1577 -6659 -1564 -6613
rect -1964 -6672 -1564 -6659
rect -1460 -6613 -1060 -6580
rect -1460 -6659 -1447 -6613
rect -1073 -6659 -1060 -6613
rect -1460 -6672 -1060 -6659
rect -956 -6613 -556 -6580
rect -956 -6659 -943 -6613
rect -569 -6659 -556 -6613
rect -956 -6672 -556 -6659
rect -452 -6613 -52 -6580
rect -452 -6659 -439 -6613
rect -65 -6659 -52 -6613
rect -452 -6672 -52 -6659
rect 52 -6613 452 -6580
rect 52 -6659 65 -6613
rect 439 -6659 452 -6613
rect 52 -6672 452 -6659
rect 556 -6613 956 -6580
rect 556 -6659 569 -6613
rect 943 -6659 956 -6613
rect 556 -6672 956 -6659
rect 1060 -6613 1460 -6580
rect 1060 -6659 1073 -6613
rect 1447 -6659 1460 -6613
rect 1060 -6672 1460 -6659
rect 1564 -6613 1964 -6580
rect 1564 -6659 1577 -6613
rect 1951 -6659 1964 -6613
rect 1564 -6672 1964 -6659
rect 2068 -6613 2468 -6580
rect 2068 -6659 2081 -6613
rect 2455 -6659 2468 -6613
rect 2068 -6672 2468 -6659
rect -2468 -6733 -2068 -6720
rect -2468 -6779 -2455 -6733
rect -2081 -6779 -2068 -6733
rect -2468 -6812 -2068 -6779
rect -1964 -6733 -1564 -6720
rect -1964 -6779 -1951 -6733
rect -1577 -6779 -1564 -6733
rect -1964 -6812 -1564 -6779
rect -1460 -6733 -1060 -6720
rect -1460 -6779 -1447 -6733
rect -1073 -6779 -1060 -6733
rect -1460 -6812 -1060 -6779
rect -956 -6733 -556 -6720
rect -956 -6779 -943 -6733
rect -569 -6779 -556 -6733
rect -956 -6812 -556 -6779
rect -452 -6733 -52 -6720
rect -452 -6779 -439 -6733
rect -65 -6779 -52 -6733
rect -452 -6812 -52 -6779
rect 52 -6733 452 -6720
rect 52 -6779 65 -6733
rect 439 -6779 452 -6733
rect 52 -6812 452 -6779
rect 556 -6733 956 -6720
rect 556 -6779 569 -6733
rect 943 -6779 956 -6733
rect 556 -6812 956 -6779
rect 1060 -6733 1460 -6720
rect 1060 -6779 1073 -6733
rect 1447 -6779 1460 -6733
rect 1060 -6812 1460 -6779
rect 1564 -6733 1964 -6720
rect 1564 -6779 1577 -6733
rect 1951 -6779 1964 -6733
rect 1564 -6812 1964 -6779
rect 2068 -6733 2468 -6720
rect 2068 -6779 2081 -6733
rect 2455 -6779 2468 -6733
rect 2068 -6812 2468 -6779
rect -2468 -8845 -2068 -8812
rect -2468 -8891 -2455 -8845
rect -2081 -8891 -2068 -8845
rect -2468 -8904 -2068 -8891
rect -1964 -8845 -1564 -8812
rect -1964 -8891 -1951 -8845
rect -1577 -8891 -1564 -8845
rect -1964 -8904 -1564 -8891
rect -1460 -8845 -1060 -8812
rect -1460 -8891 -1447 -8845
rect -1073 -8891 -1060 -8845
rect -1460 -8904 -1060 -8891
rect -956 -8845 -556 -8812
rect -956 -8891 -943 -8845
rect -569 -8891 -556 -8845
rect -956 -8904 -556 -8891
rect -452 -8845 -52 -8812
rect -452 -8891 -439 -8845
rect -65 -8891 -52 -8845
rect -452 -8904 -52 -8891
rect 52 -8845 452 -8812
rect 52 -8891 65 -8845
rect 439 -8891 452 -8845
rect 52 -8904 452 -8891
rect 556 -8845 956 -8812
rect 556 -8891 569 -8845
rect 943 -8891 956 -8845
rect 556 -8904 956 -8891
rect 1060 -8845 1460 -8812
rect 1060 -8891 1073 -8845
rect 1447 -8891 1460 -8845
rect 1060 -8904 1460 -8891
rect 1564 -8845 1964 -8812
rect 1564 -8891 1577 -8845
rect 1951 -8891 1964 -8845
rect 1564 -8904 1964 -8891
rect 2068 -8845 2468 -8812
rect 2068 -8891 2081 -8845
rect 2455 -8891 2468 -8845
rect 2068 -8904 2468 -8891
rect -2468 -8965 -2068 -8952
rect -2468 -9011 -2455 -8965
rect -2081 -9011 -2068 -8965
rect -2468 -9044 -2068 -9011
rect -1964 -8965 -1564 -8952
rect -1964 -9011 -1951 -8965
rect -1577 -9011 -1564 -8965
rect -1964 -9044 -1564 -9011
rect -1460 -8965 -1060 -8952
rect -1460 -9011 -1447 -8965
rect -1073 -9011 -1060 -8965
rect -1460 -9044 -1060 -9011
rect -956 -8965 -556 -8952
rect -956 -9011 -943 -8965
rect -569 -9011 -556 -8965
rect -956 -9044 -556 -9011
rect -452 -8965 -52 -8952
rect -452 -9011 -439 -8965
rect -65 -9011 -52 -8965
rect -452 -9044 -52 -9011
rect 52 -8965 452 -8952
rect 52 -9011 65 -8965
rect 439 -9011 452 -8965
rect 52 -9044 452 -9011
rect 556 -8965 956 -8952
rect 556 -9011 569 -8965
rect 943 -9011 956 -8965
rect 556 -9044 956 -9011
rect 1060 -8965 1460 -8952
rect 1060 -9011 1073 -8965
rect 1447 -9011 1460 -8965
rect 1060 -9044 1460 -9011
rect 1564 -8965 1964 -8952
rect 1564 -9011 1577 -8965
rect 1951 -9011 1964 -8965
rect 1564 -9044 1964 -9011
rect 2068 -8965 2468 -8952
rect 2068 -9011 2081 -8965
rect 2455 -9011 2468 -8965
rect 2068 -9044 2468 -9011
rect -2468 -11077 -2068 -11044
rect -2468 -11123 -2455 -11077
rect -2081 -11123 -2068 -11077
rect -2468 -11136 -2068 -11123
rect -1964 -11077 -1564 -11044
rect -1964 -11123 -1951 -11077
rect -1577 -11123 -1564 -11077
rect -1964 -11136 -1564 -11123
rect -1460 -11077 -1060 -11044
rect -1460 -11123 -1447 -11077
rect -1073 -11123 -1060 -11077
rect -1460 -11136 -1060 -11123
rect -956 -11077 -556 -11044
rect -956 -11123 -943 -11077
rect -569 -11123 -556 -11077
rect -956 -11136 -556 -11123
rect -452 -11077 -52 -11044
rect -452 -11123 -439 -11077
rect -65 -11123 -52 -11077
rect -452 -11136 -52 -11123
rect 52 -11077 452 -11044
rect 52 -11123 65 -11077
rect 439 -11123 452 -11077
rect 52 -11136 452 -11123
rect 556 -11077 956 -11044
rect 556 -11123 569 -11077
rect 943 -11123 956 -11077
rect 556 -11136 956 -11123
rect 1060 -11077 1460 -11044
rect 1060 -11123 1073 -11077
rect 1447 -11123 1460 -11077
rect 1060 -11136 1460 -11123
rect 1564 -11077 1964 -11044
rect 1564 -11123 1577 -11077
rect 1951 -11123 1964 -11077
rect 1564 -11136 1964 -11123
rect 2068 -11077 2468 -11044
rect 2068 -11123 2081 -11077
rect 2455 -11123 2468 -11077
rect 2068 -11136 2468 -11123
rect -2468 -11197 -2068 -11184
rect -2468 -11243 -2455 -11197
rect -2081 -11243 -2068 -11197
rect -2468 -11276 -2068 -11243
rect -1964 -11197 -1564 -11184
rect -1964 -11243 -1951 -11197
rect -1577 -11243 -1564 -11197
rect -1964 -11276 -1564 -11243
rect -1460 -11197 -1060 -11184
rect -1460 -11243 -1447 -11197
rect -1073 -11243 -1060 -11197
rect -1460 -11276 -1060 -11243
rect -956 -11197 -556 -11184
rect -956 -11243 -943 -11197
rect -569 -11243 -556 -11197
rect -956 -11276 -556 -11243
rect -452 -11197 -52 -11184
rect -452 -11243 -439 -11197
rect -65 -11243 -52 -11197
rect -452 -11276 -52 -11243
rect 52 -11197 452 -11184
rect 52 -11243 65 -11197
rect 439 -11243 452 -11197
rect 52 -11276 452 -11243
rect 556 -11197 956 -11184
rect 556 -11243 569 -11197
rect 943 -11243 956 -11197
rect 556 -11276 956 -11243
rect 1060 -11197 1460 -11184
rect 1060 -11243 1073 -11197
rect 1447 -11243 1460 -11197
rect 1060 -11276 1460 -11243
rect 1564 -11197 1964 -11184
rect 1564 -11243 1577 -11197
rect 1951 -11243 1964 -11197
rect 1564 -11276 1964 -11243
rect 2068 -11197 2468 -11184
rect 2068 -11243 2081 -11197
rect 2455 -11243 2468 -11197
rect 2068 -11276 2468 -11243
rect -2468 -13309 -2068 -13276
rect -2468 -13355 -2455 -13309
rect -2081 -13355 -2068 -13309
rect -2468 -13368 -2068 -13355
rect -1964 -13309 -1564 -13276
rect -1964 -13355 -1951 -13309
rect -1577 -13355 -1564 -13309
rect -1964 -13368 -1564 -13355
rect -1460 -13309 -1060 -13276
rect -1460 -13355 -1447 -13309
rect -1073 -13355 -1060 -13309
rect -1460 -13368 -1060 -13355
rect -956 -13309 -556 -13276
rect -956 -13355 -943 -13309
rect -569 -13355 -556 -13309
rect -956 -13368 -556 -13355
rect -452 -13309 -52 -13276
rect -452 -13355 -439 -13309
rect -65 -13355 -52 -13309
rect -452 -13368 -52 -13355
rect 52 -13309 452 -13276
rect 52 -13355 65 -13309
rect 439 -13355 452 -13309
rect 52 -13368 452 -13355
rect 556 -13309 956 -13276
rect 556 -13355 569 -13309
rect 943 -13355 956 -13309
rect 556 -13368 956 -13355
rect 1060 -13309 1460 -13276
rect 1060 -13355 1073 -13309
rect 1447 -13355 1460 -13309
rect 1060 -13368 1460 -13355
rect 1564 -13309 1964 -13276
rect 1564 -13355 1577 -13309
rect 1951 -13355 1964 -13309
rect 1564 -13368 1964 -13355
rect 2068 -13309 2468 -13276
rect 2068 -13355 2081 -13309
rect 2455 -13355 2468 -13309
rect 2068 -13368 2468 -13355
rect -2468 -13429 -2068 -13416
rect -2468 -13475 -2455 -13429
rect -2081 -13475 -2068 -13429
rect -2468 -13508 -2068 -13475
rect -1964 -13429 -1564 -13416
rect -1964 -13475 -1951 -13429
rect -1577 -13475 -1564 -13429
rect -1964 -13508 -1564 -13475
rect -1460 -13429 -1060 -13416
rect -1460 -13475 -1447 -13429
rect -1073 -13475 -1060 -13429
rect -1460 -13508 -1060 -13475
rect -956 -13429 -556 -13416
rect -956 -13475 -943 -13429
rect -569 -13475 -556 -13429
rect -956 -13508 -556 -13475
rect -452 -13429 -52 -13416
rect -452 -13475 -439 -13429
rect -65 -13475 -52 -13429
rect -452 -13508 -52 -13475
rect 52 -13429 452 -13416
rect 52 -13475 65 -13429
rect 439 -13475 452 -13429
rect 52 -13508 452 -13475
rect 556 -13429 956 -13416
rect 556 -13475 569 -13429
rect 943 -13475 956 -13429
rect 556 -13508 956 -13475
rect 1060 -13429 1460 -13416
rect 1060 -13475 1073 -13429
rect 1447 -13475 1460 -13429
rect 1060 -13508 1460 -13475
rect 1564 -13429 1964 -13416
rect 1564 -13475 1577 -13429
rect 1951 -13475 1964 -13429
rect 1564 -13508 1964 -13475
rect 2068 -13429 2468 -13416
rect 2068 -13475 2081 -13429
rect 2455 -13475 2468 -13429
rect 2068 -13508 2468 -13475
rect -2468 -15541 -2068 -15508
rect -2468 -15587 -2455 -15541
rect -2081 -15587 -2068 -15541
rect -2468 -15600 -2068 -15587
rect -1964 -15541 -1564 -15508
rect -1964 -15587 -1951 -15541
rect -1577 -15587 -1564 -15541
rect -1964 -15600 -1564 -15587
rect -1460 -15541 -1060 -15508
rect -1460 -15587 -1447 -15541
rect -1073 -15587 -1060 -15541
rect -1460 -15600 -1060 -15587
rect -956 -15541 -556 -15508
rect -956 -15587 -943 -15541
rect -569 -15587 -556 -15541
rect -956 -15600 -556 -15587
rect -452 -15541 -52 -15508
rect -452 -15587 -439 -15541
rect -65 -15587 -52 -15541
rect -452 -15600 -52 -15587
rect 52 -15541 452 -15508
rect 52 -15587 65 -15541
rect 439 -15587 452 -15541
rect 52 -15600 452 -15587
rect 556 -15541 956 -15508
rect 556 -15587 569 -15541
rect 943 -15587 956 -15541
rect 556 -15600 956 -15587
rect 1060 -15541 1460 -15508
rect 1060 -15587 1073 -15541
rect 1447 -15587 1460 -15541
rect 1060 -15600 1460 -15587
rect 1564 -15541 1964 -15508
rect 1564 -15587 1577 -15541
rect 1951 -15587 1964 -15541
rect 1564 -15600 1964 -15587
rect 2068 -15541 2468 -15508
rect 2068 -15587 2081 -15541
rect 2455 -15587 2468 -15541
rect 2068 -15600 2468 -15587
rect -2468 -15661 -2068 -15648
rect -2468 -15707 -2455 -15661
rect -2081 -15707 -2068 -15661
rect -2468 -15740 -2068 -15707
rect -1964 -15661 -1564 -15648
rect -1964 -15707 -1951 -15661
rect -1577 -15707 -1564 -15661
rect -1964 -15740 -1564 -15707
rect -1460 -15661 -1060 -15648
rect -1460 -15707 -1447 -15661
rect -1073 -15707 -1060 -15661
rect -1460 -15740 -1060 -15707
rect -956 -15661 -556 -15648
rect -956 -15707 -943 -15661
rect -569 -15707 -556 -15661
rect -956 -15740 -556 -15707
rect -452 -15661 -52 -15648
rect -452 -15707 -439 -15661
rect -65 -15707 -52 -15661
rect -452 -15740 -52 -15707
rect 52 -15661 452 -15648
rect 52 -15707 65 -15661
rect 439 -15707 452 -15661
rect 52 -15740 452 -15707
rect 556 -15661 956 -15648
rect 556 -15707 569 -15661
rect 943 -15707 956 -15661
rect 556 -15740 956 -15707
rect 1060 -15661 1460 -15648
rect 1060 -15707 1073 -15661
rect 1447 -15707 1460 -15661
rect 1060 -15740 1460 -15707
rect 1564 -15661 1964 -15648
rect 1564 -15707 1577 -15661
rect 1951 -15707 1964 -15661
rect 1564 -15740 1964 -15707
rect 2068 -15661 2468 -15648
rect 2068 -15707 2081 -15661
rect 2455 -15707 2468 -15661
rect 2068 -15740 2468 -15707
rect -2468 -17773 -2068 -17740
rect -2468 -17819 -2455 -17773
rect -2081 -17819 -2068 -17773
rect -2468 -17832 -2068 -17819
rect -1964 -17773 -1564 -17740
rect -1964 -17819 -1951 -17773
rect -1577 -17819 -1564 -17773
rect -1964 -17832 -1564 -17819
rect -1460 -17773 -1060 -17740
rect -1460 -17819 -1447 -17773
rect -1073 -17819 -1060 -17773
rect -1460 -17832 -1060 -17819
rect -956 -17773 -556 -17740
rect -956 -17819 -943 -17773
rect -569 -17819 -556 -17773
rect -956 -17832 -556 -17819
rect -452 -17773 -52 -17740
rect -452 -17819 -439 -17773
rect -65 -17819 -52 -17773
rect -452 -17832 -52 -17819
rect 52 -17773 452 -17740
rect 52 -17819 65 -17773
rect 439 -17819 452 -17773
rect 52 -17832 452 -17819
rect 556 -17773 956 -17740
rect 556 -17819 569 -17773
rect 943 -17819 956 -17773
rect 556 -17832 956 -17819
rect 1060 -17773 1460 -17740
rect 1060 -17819 1073 -17773
rect 1447 -17819 1460 -17773
rect 1060 -17832 1460 -17819
rect 1564 -17773 1964 -17740
rect 1564 -17819 1577 -17773
rect 1951 -17819 1964 -17773
rect 1564 -17832 1964 -17819
rect 2068 -17773 2468 -17740
rect 2068 -17819 2081 -17773
rect 2455 -17819 2468 -17773
rect 2068 -17832 2468 -17819
rect -2468 -17893 -2068 -17880
rect -2468 -17939 -2455 -17893
rect -2081 -17939 -2068 -17893
rect -2468 -17972 -2068 -17939
rect -1964 -17893 -1564 -17880
rect -1964 -17939 -1951 -17893
rect -1577 -17939 -1564 -17893
rect -1964 -17972 -1564 -17939
rect -1460 -17893 -1060 -17880
rect -1460 -17939 -1447 -17893
rect -1073 -17939 -1060 -17893
rect -1460 -17972 -1060 -17939
rect -956 -17893 -556 -17880
rect -956 -17939 -943 -17893
rect -569 -17939 -556 -17893
rect -956 -17972 -556 -17939
rect -452 -17893 -52 -17880
rect -452 -17939 -439 -17893
rect -65 -17939 -52 -17893
rect -452 -17972 -52 -17939
rect 52 -17893 452 -17880
rect 52 -17939 65 -17893
rect 439 -17939 452 -17893
rect 52 -17972 452 -17939
rect 556 -17893 956 -17880
rect 556 -17939 569 -17893
rect 943 -17939 956 -17893
rect 556 -17972 956 -17939
rect 1060 -17893 1460 -17880
rect 1060 -17939 1073 -17893
rect 1447 -17939 1460 -17893
rect 1060 -17972 1460 -17939
rect 1564 -17893 1964 -17880
rect 1564 -17939 1577 -17893
rect 1951 -17939 1964 -17893
rect 1564 -17972 1964 -17939
rect 2068 -17893 2468 -17880
rect 2068 -17939 2081 -17893
rect 2455 -17939 2468 -17893
rect 2068 -17972 2468 -17939
rect -2468 -20005 -2068 -19972
rect -2468 -20051 -2455 -20005
rect -2081 -20051 -2068 -20005
rect -2468 -20064 -2068 -20051
rect -1964 -20005 -1564 -19972
rect -1964 -20051 -1951 -20005
rect -1577 -20051 -1564 -20005
rect -1964 -20064 -1564 -20051
rect -1460 -20005 -1060 -19972
rect -1460 -20051 -1447 -20005
rect -1073 -20051 -1060 -20005
rect -1460 -20064 -1060 -20051
rect -956 -20005 -556 -19972
rect -956 -20051 -943 -20005
rect -569 -20051 -556 -20005
rect -956 -20064 -556 -20051
rect -452 -20005 -52 -19972
rect -452 -20051 -439 -20005
rect -65 -20051 -52 -20005
rect -452 -20064 -52 -20051
rect 52 -20005 452 -19972
rect 52 -20051 65 -20005
rect 439 -20051 452 -20005
rect 52 -20064 452 -20051
rect 556 -20005 956 -19972
rect 556 -20051 569 -20005
rect 943 -20051 956 -20005
rect 556 -20064 956 -20051
rect 1060 -20005 1460 -19972
rect 1060 -20051 1073 -20005
rect 1447 -20051 1460 -20005
rect 1060 -20064 1460 -20051
rect 1564 -20005 1964 -19972
rect 1564 -20051 1577 -20005
rect 1951 -20051 1964 -20005
rect 1564 -20064 1964 -20051
rect 2068 -20005 2468 -19972
rect 2068 -20051 2081 -20005
rect 2455 -20051 2468 -20005
rect 2068 -20064 2468 -20051
rect -2468 -20125 -2068 -20112
rect -2468 -20171 -2455 -20125
rect -2081 -20171 -2068 -20125
rect -2468 -20204 -2068 -20171
rect -1964 -20125 -1564 -20112
rect -1964 -20171 -1951 -20125
rect -1577 -20171 -1564 -20125
rect -1964 -20204 -1564 -20171
rect -1460 -20125 -1060 -20112
rect -1460 -20171 -1447 -20125
rect -1073 -20171 -1060 -20125
rect -1460 -20204 -1060 -20171
rect -956 -20125 -556 -20112
rect -956 -20171 -943 -20125
rect -569 -20171 -556 -20125
rect -956 -20204 -556 -20171
rect -452 -20125 -52 -20112
rect -452 -20171 -439 -20125
rect -65 -20171 -52 -20125
rect -452 -20204 -52 -20171
rect 52 -20125 452 -20112
rect 52 -20171 65 -20125
rect 439 -20171 452 -20125
rect 52 -20204 452 -20171
rect 556 -20125 956 -20112
rect 556 -20171 569 -20125
rect 943 -20171 956 -20125
rect 556 -20204 956 -20171
rect 1060 -20125 1460 -20112
rect 1060 -20171 1073 -20125
rect 1447 -20171 1460 -20125
rect 1060 -20204 1460 -20171
rect 1564 -20125 1964 -20112
rect 1564 -20171 1577 -20125
rect 1951 -20171 1964 -20125
rect 1564 -20204 1964 -20171
rect 2068 -20125 2468 -20112
rect 2068 -20171 2081 -20125
rect 2455 -20171 2468 -20125
rect 2068 -20204 2468 -20171
rect -2468 -22237 -2068 -22204
rect -2468 -22283 -2455 -22237
rect -2081 -22283 -2068 -22237
rect -2468 -22296 -2068 -22283
rect -1964 -22237 -1564 -22204
rect -1964 -22283 -1951 -22237
rect -1577 -22283 -1564 -22237
rect -1964 -22296 -1564 -22283
rect -1460 -22237 -1060 -22204
rect -1460 -22283 -1447 -22237
rect -1073 -22283 -1060 -22237
rect -1460 -22296 -1060 -22283
rect -956 -22237 -556 -22204
rect -956 -22283 -943 -22237
rect -569 -22283 -556 -22237
rect -956 -22296 -556 -22283
rect -452 -22237 -52 -22204
rect -452 -22283 -439 -22237
rect -65 -22283 -52 -22237
rect -452 -22296 -52 -22283
rect 52 -22237 452 -22204
rect 52 -22283 65 -22237
rect 439 -22283 452 -22237
rect 52 -22296 452 -22283
rect 556 -22237 956 -22204
rect 556 -22283 569 -22237
rect 943 -22283 956 -22237
rect 556 -22296 956 -22283
rect 1060 -22237 1460 -22204
rect 1060 -22283 1073 -22237
rect 1447 -22283 1460 -22237
rect 1060 -22296 1460 -22283
rect 1564 -22237 1964 -22204
rect 1564 -22283 1577 -22237
rect 1951 -22283 1964 -22237
rect 1564 -22296 1964 -22283
rect 2068 -22237 2468 -22204
rect 2068 -22283 2081 -22237
rect 2455 -22283 2468 -22237
rect 2068 -22296 2468 -22283
rect -2468 -22357 -2068 -22344
rect -2468 -22403 -2455 -22357
rect -2081 -22403 -2068 -22357
rect -2468 -22436 -2068 -22403
rect -1964 -22357 -1564 -22344
rect -1964 -22403 -1951 -22357
rect -1577 -22403 -1564 -22357
rect -1964 -22436 -1564 -22403
rect -1460 -22357 -1060 -22344
rect -1460 -22403 -1447 -22357
rect -1073 -22403 -1060 -22357
rect -1460 -22436 -1060 -22403
rect -956 -22357 -556 -22344
rect -956 -22403 -943 -22357
rect -569 -22403 -556 -22357
rect -956 -22436 -556 -22403
rect -452 -22357 -52 -22344
rect -452 -22403 -439 -22357
rect -65 -22403 -52 -22357
rect -452 -22436 -52 -22403
rect 52 -22357 452 -22344
rect 52 -22403 65 -22357
rect 439 -22403 452 -22357
rect 52 -22436 452 -22403
rect 556 -22357 956 -22344
rect 556 -22403 569 -22357
rect 943 -22403 956 -22357
rect 556 -22436 956 -22403
rect 1060 -22357 1460 -22344
rect 1060 -22403 1073 -22357
rect 1447 -22403 1460 -22357
rect 1060 -22436 1460 -22403
rect 1564 -22357 1964 -22344
rect 1564 -22403 1577 -22357
rect 1951 -22403 1964 -22357
rect 1564 -22436 1964 -22403
rect 2068 -22357 2468 -22344
rect 2068 -22403 2081 -22357
rect 2455 -22403 2468 -22357
rect 2068 -22436 2468 -22403
rect -2468 -24469 -2068 -24436
rect -2468 -24515 -2455 -24469
rect -2081 -24515 -2068 -24469
rect -2468 -24528 -2068 -24515
rect -1964 -24469 -1564 -24436
rect -1964 -24515 -1951 -24469
rect -1577 -24515 -1564 -24469
rect -1964 -24528 -1564 -24515
rect -1460 -24469 -1060 -24436
rect -1460 -24515 -1447 -24469
rect -1073 -24515 -1060 -24469
rect -1460 -24528 -1060 -24515
rect -956 -24469 -556 -24436
rect -956 -24515 -943 -24469
rect -569 -24515 -556 -24469
rect -956 -24528 -556 -24515
rect -452 -24469 -52 -24436
rect -452 -24515 -439 -24469
rect -65 -24515 -52 -24469
rect -452 -24528 -52 -24515
rect 52 -24469 452 -24436
rect 52 -24515 65 -24469
rect 439 -24515 452 -24469
rect 52 -24528 452 -24515
rect 556 -24469 956 -24436
rect 556 -24515 569 -24469
rect 943 -24515 956 -24469
rect 556 -24528 956 -24515
rect 1060 -24469 1460 -24436
rect 1060 -24515 1073 -24469
rect 1447 -24515 1460 -24469
rect 1060 -24528 1460 -24515
rect 1564 -24469 1964 -24436
rect 1564 -24515 1577 -24469
rect 1951 -24515 1964 -24469
rect 1564 -24528 1964 -24515
rect 2068 -24469 2468 -24436
rect 2068 -24515 2081 -24469
rect 2455 -24515 2468 -24469
rect 2068 -24528 2468 -24515
rect -2468 -24589 -2068 -24576
rect -2468 -24635 -2455 -24589
rect -2081 -24635 -2068 -24589
rect -2468 -24668 -2068 -24635
rect -1964 -24589 -1564 -24576
rect -1964 -24635 -1951 -24589
rect -1577 -24635 -1564 -24589
rect -1964 -24668 -1564 -24635
rect -1460 -24589 -1060 -24576
rect -1460 -24635 -1447 -24589
rect -1073 -24635 -1060 -24589
rect -1460 -24668 -1060 -24635
rect -956 -24589 -556 -24576
rect -956 -24635 -943 -24589
rect -569 -24635 -556 -24589
rect -956 -24668 -556 -24635
rect -452 -24589 -52 -24576
rect -452 -24635 -439 -24589
rect -65 -24635 -52 -24589
rect -452 -24668 -52 -24635
rect 52 -24589 452 -24576
rect 52 -24635 65 -24589
rect 439 -24635 452 -24589
rect 52 -24668 452 -24635
rect 556 -24589 956 -24576
rect 556 -24635 569 -24589
rect 943 -24635 956 -24589
rect 556 -24668 956 -24635
rect 1060 -24589 1460 -24576
rect 1060 -24635 1073 -24589
rect 1447 -24635 1460 -24589
rect 1060 -24668 1460 -24635
rect 1564 -24589 1964 -24576
rect 1564 -24635 1577 -24589
rect 1951 -24635 1964 -24589
rect 1564 -24668 1964 -24635
rect 2068 -24589 2468 -24576
rect 2068 -24635 2081 -24589
rect 2455 -24635 2468 -24589
rect 2068 -24668 2468 -24635
rect -2468 -26701 -2068 -26668
rect -2468 -26747 -2455 -26701
rect -2081 -26747 -2068 -26701
rect -2468 -26760 -2068 -26747
rect -1964 -26701 -1564 -26668
rect -1964 -26747 -1951 -26701
rect -1577 -26747 -1564 -26701
rect -1964 -26760 -1564 -26747
rect -1460 -26701 -1060 -26668
rect -1460 -26747 -1447 -26701
rect -1073 -26747 -1060 -26701
rect -1460 -26760 -1060 -26747
rect -956 -26701 -556 -26668
rect -956 -26747 -943 -26701
rect -569 -26747 -556 -26701
rect -956 -26760 -556 -26747
rect -452 -26701 -52 -26668
rect -452 -26747 -439 -26701
rect -65 -26747 -52 -26701
rect -452 -26760 -52 -26747
rect 52 -26701 452 -26668
rect 52 -26747 65 -26701
rect 439 -26747 452 -26701
rect 52 -26760 452 -26747
rect 556 -26701 956 -26668
rect 556 -26747 569 -26701
rect 943 -26747 956 -26701
rect 556 -26760 956 -26747
rect 1060 -26701 1460 -26668
rect 1060 -26747 1073 -26701
rect 1447 -26747 1460 -26701
rect 1060 -26760 1460 -26747
rect 1564 -26701 1964 -26668
rect 1564 -26747 1577 -26701
rect 1951 -26747 1964 -26701
rect 1564 -26760 1964 -26747
rect 2068 -26701 2468 -26668
rect 2068 -26747 2081 -26701
rect 2455 -26747 2468 -26701
rect 2068 -26760 2468 -26747
rect -2468 -26821 -2068 -26808
rect -2468 -26867 -2455 -26821
rect -2081 -26867 -2068 -26821
rect -2468 -26900 -2068 -26867
rect -1964 -26821 -1564 -26808
rect -1964 -26867 -1951 -26821
rect -1577 -26867 -1564 -26821
rect -1964 -26900 -1564 -26867
rect -1460 -26821 -1060 -26808
rect -1460 -26867 -1447 -26821
rect -1073 -26867 -1060 -26821
rect -1460 -26900 -1060 -26867
rect -956 -26821 -556 -26808
rect -956 -26867 -943 -26821
rect -569 -26867 -556 -26821
rect -956 -26900 -556 -26867
rect -452 -26821 -52 -26808
rect -452 -26867 -439 -26821
rect -65 -26867 -52 -26821
rect -452 -26900 -52 -26867
rect 52 -26821 452 -26808
rect 52 -26867 65 -26821
rect 439 -26867 452 -26821
rect 52 -26900 452 -26867
rect 556 -26821 956 -26808
rect 556 -26867 569 -26821
rect 943 -26867 956 -26821
rect 556 -26900 956 -26867
rect 1060 -26821 1460 -26808
rect 1060 -26867 1073 -26821
rect 1447 -26867 1460 -26821
rect 1060 -26900 1460 -26867
rect 1564 -26821 1964 -26808
rect 1564 -26867 1577 -26821
rect 1951 -26867 1964 -26821
rect 1564 -26900 1964 -26867
rect 2068 -26821 2468 -26808
rect 2068 -26867 2081 -26821
rect 2455 -26867 2468 -26821
rect 2068 -26900 2468 -26867
rect -2468 -28933 -2068 -28900
rect -2468 -28979 -2455 -28933
rect -2081 -28979 -2068 -28933
rect -2468 -28992 -2068 -28979
rect -1964 -28933 -1564 -28900
rect -1964 -28979 -1951 -28933
rect -1577 -28979 -1564 -28933
rect -1964 -28992 -1564 -28979
rect -1460 -28933 -1060 -28900
rect -1460 -28979 -1447 -28933
rect -1073 -28979 -1060 -28933
rect -1460 -28992 -1060 -28979
rect -956 -28933 -556 -28900
rect -956 -28979 -943 -28933
rect -569 -28979 -556 -28933
rect -956 -28992 -556 -28979
rect -452 -28933 -52 -28900
rect -452 -28979 -439 -28933
rect -65 -28979 -52 -28933
rect -452 -28992 -52 -28979
rect 52 -28933 452 -28900
rect 52 -28979 65 -28933
rect 439 -28979 452 -28933
rect 52 -28992 452 -28979
rect 556 -28933 956 -28900
rect 556 -28979 569 -28933
rect 943 -28979 956 -28933
rect 556 -28992 956 -28979
rect 1060 -28933 1460 -28900
rect 1060 -28979 1073 -28933
rect 1447 -28979 1460 -28933
rect 1060 -28992 1460 -28979
rect 1564 -28933 1964 -28900
rect 1564 -28979 1577 -28933
rect 1951 -28979 1964 -28933
rect 1564 -28992 1964 -28979
rect 2068 -28933 2468 -28900
rect 2068 -28979 2081 -28933
rect 2455 -28979 2468 -28933
rect 2068 -28992 2468 -28979
<< polycontact >>
rect -2455 28933 -2081 28979
rect -1951 28933 -1577 28979
rect -1447 28933 -1073 28979
rect -943 28933 -569 28979
rect -439 28933 -65 28979
rect 65 28933 439 28979
rect 569 28933 943 28979
rect 1073 28933 1447 28979
rect 1577 28933 1951 28979
rect 2081 28933 2455 28979
rect -2455 26821 -2081 26867
rect -1951 26821 -1577 26867
rect -1447 26821 -1073 26867
rect -943 26821 -569 26867
rect -439 26821 -65 26867
rect 65 26821 439 26867
rect 569 26821 943 26867
rect 1073 26821 1447 26867
rect 1577 26821 1951 26867
rect 2081 26821 2455 26867
rect -2455 26701 -2081 26747
rect -1951 26701 -1577 26747
rect -1447 26701 -1073 26747
rect -943 26701 -569 26747
rect -439 26701 -65 26747
rect 65 26701 439 26747
rect 569 26701 943 26747
rect 1073 26701 1447 26747
rect 1577 26701 1951 26747
rect 2081 26701 2455 26747
rect -2455 24589 -2081 24635
rect -1951 24589 -1577 24635
rect -1447 24589 -1073 24635
rect -943 24589 -569 24635
rect -439 24589 -65 24635
rect 65 24589 439 24635
rect 569 24589 943 24635
rect 1073 24589 1447 24635
rect 1577 24589 1951 24635
rect 2081 24589 2455 24635
rect -2455 24469 -2081 24515
rect -1951 24469 -1577 24515
rect -1447 24469 -1073 24515
rect -943 24469 -569 24515
rect -439 24469 -65 24515
rect 65 24469 439 24515
rect 569 24469 943 24515
rect 1073 24469 1447 24515
rect 1577 24469 1951 24515
rect 2081 24469 2455 24515
rect -2455 22357 -2081 22403
rect -1951 22357 -1577 22403
rect -1447 22357 -1073 22403
rect -943 22357 -569 22403
rect -439 22357 -65 22403
rect 65 22357 439 22403
rect 569 22357 943 22403
rect 1073 22357 1447 22403
rect 1577 22357 1951 22403
rect 2081 22357 2455 22403
rect -2455 22237 -2081 22283
rect -1951 22237 -1577 22283
rect -1447 22237 -1073 22283
rect -943 22237 -569 22283
rect -439 22237 -65 22283
rect 65 22237 439 22283
rect 569 22237 943 22283
rect 1073 22237 1447 22283
rect 1577 22237 1951 22283
rect 2081 22237 2455 22283
rect -2455 20125 -2081 20171
rect -1951 20125 -1577 20171
rect -1447 20125 -1073 20171
rect -943 20125 -569 20171
rect -439 20125 -65 20171
rect 65 20125 439 20171
rect 569 20125 943 20171
rect 1073 20125 1447 20171
rect 1577 20125 1951 20171
rect 2081 20125 2455 20171
rect -2455 20005 -2081 20051
rect -1951 20005 -1577 20051
rect -1447 20005 -1073 20051
rect -943 20005 -569 20051
rect -439 20005 -65 20051
rect 65 20005 439 20051
rect 569 20005 943 20051
rect 1073 20005 1447 20051
rect 1577 20005 1951 20051
rect 2081 20005 2455 20051
rect -2455 17893 -2081 17939
rect -1951 17893 -1577 17939
rect -1447 17893 -1073 17939
rect -943 17893 -569 17939
rect -439 17893 -65 17939
rect 65 17893 439 17939
rect 569 17893 943 17939
rect 1073 17893 1447 17939
rect 1577 17893 1951 17939
rect 2081 17893 2455 17939
rect -2455 17773 -2081 17819
rect -1951 17773 -1577 17819
rect -1447 17773 -1073 17819
rect -943 17773 -569 17819
rect -439 17773 -65 17819
rect 65 17773 439 17819
rect 569 17773 943 17819
rect 1073 17773 1447 17819
rect 1577 17773 1951 17819
rect 2081 17773 2455 17819
rect -2455 15661 -2081 15707
rect -1951 15661 -1577 15707
rect -1447 15661 -1073 15707
rect -943 15661 -569 15707
rect -439 15661 -65 15707
rect 65 15661 439 15707
rect 569 15661 943 15707
rect 1073 15661 1447 15707
rect 1577 15661 1951 15707
rect 2081 15661 2455 15707
rect -2455 15541 -2081 15587
rect -1951 15541 -1577 15587
rect -1447 15541 -1073 15587
rect -943 15541 -569 15587
rect -439 15541 -65 15587
rect 65 15541 439 15587
rect 569 15541 943 15587
rect 1073 15541 1447 15587
rect 1577 15541 1951 15587
rect 2081 15541 2455 15587
rect -2455 13429 -2081 13475
rect -1951 13429 -1577 13475
rect -1447 13429 -1073 13475
rect -943 13429 -569 13475
rect -439 13429 -65 13475
rect 65 13429 439 13475
rect 569 13429 943 13475
rect 1073 13429 1447 13475
rect 1577 13429 1951 13475
rect 2081 13429 2455 13475
rect -2455 13309 -2081 13355
rect -1951 13309 -1577 13355
rect -1447 13309 -1073 13355
rect -943 13309 -569 13355
rect -439 13309 -65 13355
rect 65 13309 439 13355
rect 569 13309 943 13355
rect 1073 13309 1447 13355
rect 1577 13309 1951 13355
rect 2081 13309 2455 13355
rect -2455 11197 -2081 11243
rect -1951 11197 -1577 11243
rect -1447 11197 -1073 11243
rect -943 11197 -569 11243
rect -439 11197 -65 11243
rect 65 11197 439 11243
rect 569 11197 943 11243
rect 1073 11197 1447 11243
rect 1577 11197 1951 11243
rect 2081 11197 2455 11243
rect -2455 11077 -2081 11123
rect -1951 11077 -1577 11123
rect -1447 11077 -1073 11123
rect -943 11077 -569 11123
rect -439 11077 -65 11123
rect 65 11077 439 11123
rect 569 11077 943 11123
rect 1073 11077 1447 11123
rect 1577 11077 1951 11123
rect 2081 11077 2455 11123
rect -2455 8965 -2081 9011
rect -1951 8965 -1577 9011
rect -1447 8965 -1073 9011
rect -943 8965 -569 9011
rect -439 8965 -65 9011
rect 65 8965 439 9011
rect 569 8965 943 9011
rect 1073 8965 1447 9011
rect 1577 8965 1951 9011
rect 2081 8965 2455 9011
rect -2455 8845 -2081 8891
rect -1951 8845 -1577 8891
rect -1447 8845 -1073 8891
rect -943 8845 -569 8891
rect -439 8845 -65 8891
rect 65 8845 439 8891
rect 569 8845 943 8891
rect 1073 8845 1447 8891
rect 1577 8845 1951 8891
rect 2081 8845 2455 8891
rect -2455 6733 -2081 6779
rect -1951 6733 -1577 6779
rect -1447 6733 -1073 6779
rect -943 6733 -569 6779
rect -439 6733 -65 6779
rect 65 6733 439 6779
rect 569 6733 943 6779
rect 1073 6733 1447 6779
rect 1577 6733 1951 6779
rect 2081 6733 2455 6779
rect -2455 6613 -2081 6659
rect -1951 6613 -1577 6659
rect -1447 6613 -1073 6659
rect -943 6613 -569 6659
rect -439 6613 -65 6659
rect 65 6613 439 6659
rect 569 6613 943 6659
rect 1073 6613 1447 6659
rect 1577 6613 1951 6659
rect 2081 6613 2455 6659
rect -2455 4501 -2081 4547
rect -1951 4501 -1577 4547
rect -1447 4501 -1073 4547
rect -943 4501 -569 4547
rect -439 4501 -65 4547
rect 65 4501 439 4547
rect 569 4501 943 4547
rect 1073 4501 1447 4547
rect 1577 4501 1951 4547
rect 2081 4501 2455 4547
rect -2455 4381 -2081 4427
rect -1951 4381 -1577 4427
rect -1447 4381 -1073 4427
rect -943 4381 -569 4427
rect -439 4381 -65 4427
rect 65 4381 439 4427
rect 569 4381 943 4427
rect 1073 4381 1447 4427
rect 1577 4381 1951 4427
rect 2081 4381 2455 4427
rect -2455 2269 -2081 2315
rect -1951 2269 -1577 2315
rect -1447 2269 -1073 2315
rect -943 2269 -569 2315
rect -439 2269 -65 2315
rect 65 2269 439 2315
rect 569 2269 943 2315
rect 1073 2269 1447 2315
rect 1577 2269 1951 2315
rect 2081 2269 2455 2315
rect -2455 2149 -2081 2195
rect -1951 2149 -1577 2195
rect -1447 2149 -1073 2195
rect -943 2149 -569 2195
rect -439 2149 -65 2195
rect 65 2149 439 2195
rect 569 2149 943 2195
rect 1073 2149 1447 2195
rect 1577 2149 1951 2195
rect 2081 2149 2455 2195
rect -2455 37 -2081 83
rect -1951 37 -1577 83
rect -1447 37 -1073 83
rect -943 37 -569 83
rect -439 37 -65 83
rect 65 37 439 83
rect 569 37 943 83
rect 1073 37 1447 83
rect 1577 37 1951 83
rect 2081 37 2455 83
rect -2455 -83 -2081 -37
rect -1951 -83 -1577 -37
rect -1447 -83 -1073 -37
rect -943 -83 -569 -37
rect -439 -83 -65 -37
rect 65 -83 439 -37
rect 569 -83 943 -37
rect 1073 -83 1447 -37
rect 1577 -83 1951 -37
rect 2081 -83 2455 -37
rect -2455 -2195 -2081 -2149
rect -1951 -2195 -1577 -2149
rect -1447 -2195 -1073 -2149
rect -943 -2195 -569 -2149
rect -439 -2195 -65 -2149
rect 65 -2195 439 -2149
rect 569 -2195 943 -2149
rect 1073 -2195 1447 -2149
rect 1577 -2195 1951 -2149
rect 2081 -2195 2455 -2149
rect -2455 -2315 -2081 -2269
rect -1951 -2315 -1577 -2269
rect -1447 -2315 -1073 -2269
rect -943 -2315 -569 -2269
rect -439 -2315 -65 -2269
rect 65 -2315 439 -2269
rect 569 -2315 943 -2269
rect 1073 -2315 1447 -2269
rect 1577 -2315 1951 -2269
rect 2081 -2315 2455 -2269
rect -2455 -4427 -2081 -4381
rect -1951 -4427 -1577 -4381
rect -1447 -4427 -1073 -4381
rect -943 -4427 -569 -4381
rect -439 -4427 -65 -4381
rect 65 -4427 439 -4381
rect 569 -4427 943 -4381
rect 1073 -4427 1447 -4381
rect 1577 -4427 1951 -4381
rect 2081 -4427 2455 -4381
rect -2455 -4547 -2081 -4501
rect -1951 -4547 -1577 -4501
rect -1447 -4547 -1073 -4501
rect -943 -4547 -569 -4501
rect -439 -4547 -65 -4501
rect 65 -4547 439 -4501
rect 569 -4547 943 -4501
rect 1073 -4547 1447 -4501
rect 1577 -4547 1951 -4501
rect 2081 -4547 2455 -4501
rect -2455 -6659 -2081 -6613
rect -1951 -6659 -1577 -6613
rect -1447 -6659 -1073 -6613
rect -943 -6659 -569 -6613
rect -439 -6659 -65 -6613
rect 65 -6659 439 -6613
rect 569 -6659 943 -6613
rect 1073 -6659 1447 -6613
rect 1577 -6659 1951 -6613
rect 2081 -6659 2455 -6613
rect -2455 -6779 -2081 -6733
rect -1951 -6779 -1577 -6733
rect -1447 -6779 -1073 -6733
rect -943 -6779 -569 -6733
rect -439 -6779 -65 -6733
rect 65 -6779 439 -6733
rect 569 -6779 943 -6733
rect 1073 -6779 1447 -6733
rect 1577 -6779 1951 -6733
rect 2081 -6779 2455 -6733
rect -2455 -8891 -2081 -8845
rect -1951 -8891 -1577 -8845
rect -1447 -8891 -1073 -8845
rect -943 -8891 -569 -8845
rect -439 -8891 -65 -8845
rect 65 -8891 439 -8845
rect 569 -8891 943 -8845
rect 1073 -8891 1447 -8845
rect 1577 -8891 1951 -8845
rect 2081 -8891 2455 -8845
rect -2455 -9011 -2081 -8965
rect -1951 -9011 -1577 -8965
rect -1447 -9011 -1073 -8965
rect -943 -9011 -569 -8965
rect -439 -9011 -65 -8965
rect 65 -9011 439 -8965
rect 569 -9011 943 -8965
rect 1073 -9011 1447 -8965
rect 1577 -9011 1951 -8965
rect 2081 -9011 2455 -8965
rect -2455 -11123 -2081 -11077
rect -1951 -11123 -1577 -11077
rect -1447 -11123 -1073 -11077
rect -943 -11123 -569 -11077
rect -439 -11123 -65 -11077
rect 65 -11123 439 -11077
rect 569 -11123 943 -11077
rect 1073 -11123 1447 -11077
rect 1577 -11123 1951 -11077
rect 2081 -11123 2455 -11077
rect -2455 -11243 -2081 -11197
rect -1951 -11243 -1577 -11197
rect -1447 -11243 -1073 -11197
rect -943 -11243 -569 -11197
rect -439 -11243 -65 -11197
rect 65 -11243 439 -11197
rect 569 -11243 943 -11197
rect 1073 -11243 1447 -11197
rect 1577 -11243 1951 -11197
rect 2081 -11243 2455 -11197
rect -2455 -13355 -2081 -13309
rect -1951 -13355 -1577 -13309
rect -1447 -13355 -1073 -13309
rect -943 -13355 -569 -13309
rect -439 -13355 -65 -13309
rect 65 -13355 439 -13309
rect 569 -13355 943 -13309
rect 1073 -13355 1447 -13309
rect 1577 -13355 1951 -13309
rect 2081 -13355 2455 -13309
rect -2455 -13475 -2081 -13429
rect -1951 -13475 -1577 -13429
rect -1447 -13475 -1073 -13429
rect -943 -13475 -569 -13429
rect -439 -13475 -65 -13429
rect 65 -13475 439 -13429
rect 569 -13475 943 -13429
rect 1073 -13475 1447 -13429
rect 1577 -13475 1951 -13429
rect 2081 -13475 2455 -13429
rect -2455 -15587 -2081 -15541
rect -1951 -15587 -1577 -15541
rect -1447 -15587 -1073 -15541
rect -943 -15587 -569 -15541
rect -439 -15587 -65 -15541
rect 65 -15587 439 -15541
rect 569 -15587 943 -15541
rect 1073 -15587 1447 -15541
rect 1577 -15587 1951 -15541
rect 2081 -15587 2455 -15541
rect -2455 -15707 -2081 -15661
rect -1951 -15707 -1577 -15661
rect -1447 -15707 -1073 -15661
rect -943 -15707 -569 -15661
rect -439 -15707 -65 -15661
rect 65 -15707 439 -15661
rect 569 -15707 943 -15661
rect 1073 -15707 1447 -15661
rect 1577 -15707 1951 -15661
rect 2081 -15707 2455 -15661
rect -2455 -17819 -2081 -17773
rect -1951 -17819 -1577 -17773
rect -1447 -17819 -1073 -17773
rect -943 -17819 -569 -17773
rect -439 -17819 -65 -17773
rect 65 -17819 439 -17773
rect 569 -17819 943 -17773
rect 1073 -17819 1447 -17773
rect 1577 -17819 1951 -17773
rect 2081 -17819 2455 -17773
rect -2455 -17939 -2081 -17893
rect -1951 -17939 -1577 -17893
rect -1447 -17939 -1073 -17893
rect -943 -17939 -569 -17893
rect -439 -17939 -65 -17893
rect 65 -17939 439 -17893
rect 569 -17939 943 -17893
rect 1073 -17939 1447 -17893
rect 1577 -17939 1951 -17893
rect 2081 -17939 2455 -17893
rect -2455 -20051 -2081 -20005
rect -1951 -20051 -1577 -20005
rect -1447 -20051 -1073 -20005
rect -943 -20051 -569 -20005
rect -439 -20051 -65 -20005
rect 65 -20051 439 -20005
rect 569 -20051 943 -20005
rect 1073 -20051 1447 -20005
rect 1577 -20051 1951 -20005
rect 2081 -20051 2455 -20005
rect -2455 -20171 -2081 -20125
rect -1951 -20171 -1577 -20125
rect -1447 -20171 -1073 -20125
rect -943 -20171 -569 -20125
rect -439 -20171 -65 -20125
rect 65 -20171 439 -20125
rect 569 -20171 943 -20125
rect 1073 -20171 1447 -20125
rect 1577 -20171 1951 -20125
rect 2081 -20171 2455 -20125
rect -2455 -22283 -2081 -22237
rect -1951 -22283 -1577 -22237
rect -1447 -22283 -1073 -22237
rect -943 -22283 -569 -22237
rect -439 -22283 -65 -22237
rect 65 -22283 439 -22237
rect 569 -22283 943 -22237
rect 1073 -22283 1447 -22237
rect 1577 -22283 1951 -22237
rect 2081 -22283 2455 -22237
rect -2455 -22403 -2081 -22357
rect -1951 -22403 -1577 -22357
rect -1447 -22403 -1073 -22357
rect -943 -22403 -569 -22357
rect -439 -22403 -65 -22357
rect 65 -22403 439 -22357
rect 569 -22403 943 -22357
rect 1073 -22403 1447 -22357
rect 1577 -22403 1951 -22357
rect 2081 -22403 2455 -22357
rect -2455 -24515 -2081 -24469
rect -1951 -24515 -1577 -24469
rect -1447 -24515 -1073 -24469
rect -943 -24515 -569 -24469
rect -439 -24515 -65 -24469
rect 65 -24515 439 -24469
rect 569 -24515 943 -24469
rect 1073 -24515 1447 -24469
rect 1577 -24515 1951 -24469
rect 2081 -24515 2455 -24469
rect -2455 -24635 -2081 -24589
rect -1951 -24635 -1577 -24589
rect -1447 -24635 -1073 -24589
rect -943 -24635 -569 -24589
rect -439 -24635 -65 -24589
rect 65 -24635 439 -24589
rect 569 -24635 943 -24589
rect 1073 -24635 1447 -24589
rect 1577 -24635 1951 -24589
rect 2081 -24635 2455 -24589
rect -2455 -26747 -2081 -26701
rect -1951 -26747 -1577 -26701
rect -1447 -26747 -1073 -26701
rect -943 -26747 -569 -26701
rect -439 -26747 -65 -26701
rect 65 -26747 439 -26701
rect 569 -26747 943 -26701
rect 1073 -26747 1447 -26701
rect 1577 -26747 1951 -26701
rect 2081 -26747 2455 -26701
rect -2455 -26867 -2081 -26821
rect -1951 -26867 -1577 -26821
rect -1447 -26867 -1073 -26821
rect -943 -26867 -569 -26821
rect -439 -26867 -65 -26821
rect 65 -26867 439 -26821
rect 569 -26867 943 -26821
rect 1073 -26867 1447 -26821
rect 1577 -26867 1951 -26821
rect 2081 -26867 2455 -26821
rect -2455 -28979 -2081 -28933
rect -1951 -28979 -1577 -28933
rect -1447 -28979 -1073 -28933
rect -943 -28979 -569 -28933
rect -439 -28979 -65 -28933
rect 65 -28979 439 -28933
rect 569 -28979 943 -28933
rect 1073 -28979 1447 -28933
rect 1577 -28979 1951 -28933
rect 2081 -28979 2455 -28933
<< metal1 >>
rect -2681 29027 2681 29073
rect -2681 28970 -2635 29027
rect -2466 28933 -2455 28979
rect -2081 28933 -2070 28979
rect -1962 28933 -1951 28979
rect -1577 28933 -1566 28979
rect -1458 28933 -1447 28979
rect -1073 28933 -1062 28979
rect -954 28933 -943 28979
rect -569 28933 -558 28979
rect -450 28933 -439 28979
rect -65 28933 -54 28979
rect 54 28933 65 28979
rect 439 28933 450 28979
rect 558 28933 569 28979
rect 943 28933 954 28979
rect 1062 28933 1073 28979
rect 1447 28933 1458 28979
rect 1566 28933 1577 28979
rect 1951 28933 1962 28979
rect 2070 28933 2081 28979
rect 2455 28933 2466 28979
rect 2635 28970 2681 29027
rect -2543 28887 -2497 28898
rect -2543 26902 -2497 26913
rect -2039 28887 -1993 28898
rect -2039 26902 -1993 26913
rect -1535 28887 -1489 28898
rect -1535 26902 -1489 26913
rect -1031 28887 -985 28898
rect -1031 26902 -985 26913
rect -527 28887 -481 28898
rect -527 26902 -481 26913
rect -23 28887 23 28898
rect -23 26902 23 26913
rect 481 28887 527 28898
rect 481 26902 527 26913
rect 985 28887 1031 28898
rect 985 26902 1031 26913
rect 1489 28887 1535 28898
rect 1489 26902 1535 26913
rect 1993 28887 2039 28898
rect 1993 26902 2039 26913
rect 2497 28887 2543 28898
rect 2497 26902 2543 26913
rect -2466 26821 -2455 26867
rect -2081 26821 -2070 26867
rect -1962 26821 -1951 26867
rect -1577 26821 -1566 26867
rect -1458 26821 -1447 26867
rect -1073 26821 -1062 26867
rect -954 26821 -943 26867
rect -569 26821 -558 26867
rect -450 26821 -439 26867
rect -65 26821 -54 26867
rect 54 26821 65 26867
rect 439 26821 450 26867
rect 558 26821 569 26867
rect 943 26821 954 26867
rect 1062 26821 1073 26867
rect 1447 26821 1458 26867
rect 1566 26821 1577 26867
rect 1951 26821 1962 26867
rect 2070 26821 2081 26867
rect 2455 26821 2466 26867
rect -2466 26701 -2455 26747
rect -2081 26701 -2070 26747
rect -1962 26701 -1951 26747
rect -1577 26701 -1566 26747
rect -1458 26701 -1447 26747
rect -1073 26701 -1062 26747
rect -954 26701 -943 26747
rect -569 26701 -558 26747
rect -450 26701 -439 26747
rect -65 26701 -54 26747
rect 54 26701 65 26747
rect 439 26701 450 26747
rect 558 26701 569 26747
rect 943 26701 954 26747
rect 1062 26701 1073 26747
rect 1447 26701 1458 26747
rect 1566 26701 1577 26747
rect 1951 26701 1962 26747
rect 2070 26701 2081 26747
rect 2455 26701 2466 26747
rect -2543 26655 -2497 26666
rect -2543 24670 -2497 24681
rect -2039 26655 -1993 26666
rect -2039 24670 -1993 24681
rect -1535 26655 -1489 26666
rect -1535 24670 -1489 24681
rect -1031 26655 -985 26666
rect -1031 24670 -985 24681
rect -527 26655 -481 26666
rect -527 24670 -481 24681
rect -23 26655 23 26666
rect -23 24670 23 24681
rect 481 26655 527 26666
rect 481 24670 527 24681
rect 985 26655 1031 26666
rect 985 24670 1031 24681
rect 1489 26655 1535 26666
rect 1489 24670 1535 24681
rect 1993 26655 2039 26666
rect 1993 24670 2039 24681
rect 2497 26655 2543 26666
rect 2497 24670 2543 24681
rect -2466 24589 -2455 24635
rect -2081 24589 -2070 24635
rect -1962 24589 -1951 24635
rect -1577 24589 -1566 24635
rect -1458 24589 -1447 24635
rect -1073 24589 -1062 24635
rect -954 24589 -943 24635
rect -569 24589 -558 24635
rect -450 24589 -439 24635
rect -65 24589 -54 24635
rect 54 24589 65 24635
rect 439 24589 450 24635
rect 558 24589 569 24635
rect 943 24589 954 24635
rect 1062 24589 1073 24635
rect 1447 24589 1458 24635
rect 1566 24589 1577 24635
rect 1951 24589 1962 24635
rect 2070 24589 2081 24635
rect 2455 24589 2466 24635
rect -2466 24469 -2455 24515
rect -2081 24469 -2070 24515
rect -1962 24469 -1951 24515
rect -1577 24469 -1566 24515
rect -1458 24469 -1447 24515
rect -1073 24469 -1062 24515
rect -954 24469 -943 24515
rect -569 24469 -558 24515
rect -450 24469 -439 24515
rect -65 24469 -54 24515
rect 54 24469 65 24515
rect 439 24469 450 24515
rect 558 24469 569 24515
rect 943 24469 954 24515
rect 1062 24469 1073 24515
rect 1447 24469 1458 24515
rect 1566 24469 1577 24515
rect 1951 24469 1962 24515
rect 2070 24469 2081 24515
rect 2455 24469 2466 24515
rect -2543 24423 -2497 24434
rect -2543 22438 -2497 22449
rect -2039 24423 -1993 24434
rect -2039 22438 -1993 22449
rect -1535 24423 -1489 24434
rect -1535 22438 -1489 22449
rect -1031 24423 -985 24434
rect -1031 22438 -985 22449
rect -527 24423 -481 24434
rect -527 22438 -481 22449
rect -23 24423 23 24434
rect -23 22438 23 22449
rect 481 24423 527 24434
rect 481 22438 527 22449
rect 985 24423 1031 24434
rect 985 22438 1031 22449
rect 1489 24423 1535 24434
rect 1489 22438 1535 22449
rect 1993 24423 2039 24434
rect 1993 22438 2039 22449
rect 2497 24423 2543 24434
rect 2497 22438 2543 22449
rect -2466 22357 -2455 22403
rect -2081 22357 -2070 22403
rect -1962 22357 -1951 22403
rect -1577 22357 -1566 22403
rect -1458 22357 -1447 22403
rect -1073 22357 -1062 22403
rect -954 22357 -943 22403
rect -569 22357 -558 22403
rect -450 22357 -439 22403
rect -65 22357 -54 22403
rect 54 22357 65 22403
rect 439 22357 450 22403
rect 558 22357 569 22403
rect 943 22357 954 22403
rect 1062 22357 1073 22403
rect 1447 22357 1458 22403
rect 1566 22357 1577 22403
rect 1951 22357 1962 22403
rect 2070 22357 2081 22403
rect 2455 22357 2466 22403
rect -2466 22237 -2455 22283
rect -2081 22237 -2070 22283
rect -1962 22237 -1951 22283
rect -1577 22237 -1566 22283
rect -1458 22237 -1447 22283
rect -1073 22237 -1062 22283
rect -954 22237 -943 22283
rect -569 22237 -558 22283
rect -450 22237 -439 22283
rect -65 22237 -54 22283
rect 54 22237 65 22283
rect 439 22237 450 22283
rect 558 22237 569 22283
rect 943 22237 954 22283
rect 1062 22237 1073 22283
rect 1447 22237 1458 22283
rect 1566 22237 1577 22283
rect 1951 22237 1962 22283
rect 2070 22237 2081 22283
rect 2455 22237 2466 22283
rect -2543 22191 -2497 22202
rect -2543 20206 -2497 20217
rect -2039 22191 -1993 22202
rect -2039 20206 -1993 20217
rect -1535 22191 -1489 22202
rect -1535 20206 -1489 20217
rect -1031 22191 -985 22202
rect -1031 20206 -985 20217
rect -527 22191 -481 22202
rect -527 20206 -481 20217
rect -23 22191 23 22202
rect -23 20206 23 20217
rect 481 22191 527 22202
rect 481 20206 527 20217
rect 985 22191 1031 22202
rect 985 20206 1031 20217
rect 1489 22191 1535 22202
rect 1489 20206 1535 20217
rect 1993 22191 2039 22202
rect 1993 20206 2039 20217
rect 2497 22191 2543 22202
rect 2497 20206 2543 20217
rect -2466 20125 -2455 20171
rect -2081 20125 -2070 20171
rect -1962 20125 -1951 20171
rect -1577 20125 -1566 20171
rect -1458 20125 -1447 20171
rect -1073 20125 -1062 20171
rect -954 20125 -943 20171
rect -569 20125 -558 20171
rect -450 20125 -439 20171
rect -65 20125 -54 20171
rect 54 20125 65 20171
rect 439 20125 450 20171
rect 558 20125 569 20171
rect 943 20125 954 20171
rect 1062 20125 1073 20171
rect 1447 20125 1458 20171
rect 1566 20125 1577 20171
rect 1951 20125 1962 20171
rect 2070 20125 2081 20171
rect 2455 20125 2466 20171
rect -2466 20005 -2455 20051
rect -2081 20005 -2070 20051
rect -1962 20005 -1951 20051
rect -1577 20005 -1566 20051
rect -1458 20005 -1447 20051
rect -1073 20005 -1062 20051
rect -954 20005 -943 20051
rect -569 20005 -558 20051
rect -450 20005 -439 20051
rect -65 20005 -54 20051
rect 54 20005 65 20051
rect 439 20005 450 20051
rect 558 20005 569 20051
rect 943 20005 954 20051
rect 1062 20005 1073 20051
rect 1447 20005 1458 20051
rect 1566 20005 1577 20051
rect 1951 20005 1962 20051
rect 2070 20005 2081 20051
rect 2455 20005 2466 20051
rect -2543 19959 -2497 19970
rect -2543 17974 -2497 17985
rect -2039 19959 -1993 19970
rect -2039 17974 -1993 17985
rect -1535 19959 -1489 19970
rect -1535 17974 -1489 17985
rect -1031 19959 -985 19970
rect -1031 17974 -985 17985
rect -527 19959 -481 19970
rect -527 17974 -481 17985
rect -23 19959 23 19970
rect -23 17974 23 17985
rect 481 19959 527 19970
rect 481 17974 527 17985
rect 985 19959 1031 19970
rect 985 17974 1031 17985
rect 1489 19959 1535 19970
rect 1489 17974 1535 17985
rect 1993 19959 2039 19970
rect 1993 17974 2039 17985
rect 2497 19959 2543 19970
rect 2497 17974 2543 17985
rect -2466 17893 -2455 17939
rect -2081 17893 -2070 17939
rect -1962 17893 -1951 17939
rect -1577 17893 -1566 17939
rect -1458 17893 -1447 17939
rect -1073 17893 -1062 17939
rect -954 17893 -943 17939
rect -569 17893 -558 17939
rect -450 17893 -439 17939
rect -65 17893 -54 17939
rect 54 17893 65 17939
rect 439 17893 450 17939
rect 558 17893 569 17939
rect 943 17893 954 17939
rect 1062 17893 1073 17939
rect 1447 17893 1458 17939
rect 1566 17893 1577 17939
rect 1951 17893 1962 17939
rect 2070 17893 2081 17939
rect 2455 17893 2466 17939
rect -2466 17773 -2455 17819
rect -2081 17773 -2070 17819
rect -1962 17773 -1951 17819
rect -1577 17773 -1566 17819
rect -1458 17773 -1447 17819
rect -1073 17773 -1062 17819
rect -954 17773 -943 17819
rect -569 17773 -558 17819
rect -450 17773 -439 17819
rect -65 17773 -54 17819
rect 54 17773 65 17819
rect 439 17773 450 17819
rect 558 17773 569 17819
rect 943 17773 954 17819
rect 1062 17773 1073 17819
rect 1447 17773 1458 17819
rect 1566 17773 1577 17819
rect 1951 17773 1962 17819
rect 2070 17773 2081 17819
rect 2455 17773 2466 17819
rect -2543 17727 -2497 17738
rect -2543 15742 -2497 15753
rect -2039 17727 -1993 17738
rect -2039 15742 -1993 15753
rect -1535 17727 -1489 17738
rect -1535 15742 -1489 15753
rect -1031 17727 -985 17738
rect -1031 15742 -985 15753
rect -527 17727 -481 17738
rect -527 15742 -481 15753
rect -23 17727 23 17738
rect -23 15742 23 15753
rect 481 17727 527 17738
rect 481 15742 527 15753
rect 985 17727 1031 17738
rect 985 15742 1031 15753
rect 1489 17727 1535 17738
rect 1489 15742 1535 15753
rect 1993 17727 2039 17738
rect 1993 15742 2039 15753
rect 2497 17727 2543 17738
rect 2497 15742 2543 15753
rect -2466 15661 -2455 15707
rect -2081 15661 -2070 15707
rect -1962 15661 -1951 15707
rect -1577 15661 -1566 15707
rect -1458 15661 -1447 15707
rect -1073 15661 -1062 15707
rect -954 15661 -943 15707
rect -569 15661 -558 15707
rect -450 15661 -439 15707
rect -65 15661 -54 15707
rect 54 15661 65 15707
rect 439 15661 450 15707
rect 558 15661 569 15707
rect 943 15661 954 15707
rect 1062 15661 1073 15707
rect 1447 15661 1458 15707
rect 1566 15661 1577 15707
rect 1951 15661 1962 15707
rect 2070 15661 2081 15707
rect 2455 15661 2466 15707
rect -2466 15541 -2455 15587
rect -2081 15541 -2070 15587
rect -1962 15541 -1951 15587
rect -1577 15541 -1566 15587
rect -1458 15541 -1447 15587
rect -1073 15541 -1062 15587
rect -954 15541 -943 15587
rect -569 15541 -558 15587
rect -450 15541 -439 15587
rect -65 15541 -54 15587
rect 54 15541 65 15587
rect 439 15541 450 15587
rect 558 15541 569 15587
rect 943 15541 954 15587
rect 1062 15541 1073 15587
rect 1447 15541 1458 15587
rect 1566 15541 1577 15587
rect 1951 15541 1962 15587
rect 2070 15541 2081 15587
rect 2455 15541 2466 15587
rect -2543 15495 -2497 15506
rect -2543 13510 -2497 13521
rect -2039 15495 -1993 15506
rect -2039 13510 -1993 13521
rect -1535 15495 -1489 15506
rect -1535 13510 -1489 13521
rect -1031 15495 -985 15506
rect -1031 13510 -985 13521
rect -527 15495 -481 15506
rect -527 13510 -481 13521
rect -23 15495 23 15506
rect -23 13510 23 13521
rect 481 15495 527 15506
rect 481 13510 527 13521
rect 985 15495 1031 15506
rect 985 13510 1031 13521
rect 1489 15495 1535 15506
rect 1489 13510 1535 13521
rect 1993 15495 2039 15506
rect 1993 13510 2039 13521
rect 2497 15495 2543 15506
rect 2497 13510 2543 13521
rect -2466 13429 -2455 13475
rect -2081 13429 -2070 13475
rect -1962 13429 -1951 13475
rect -1577 13429 -1566 13475
rect -1458 13429 -1447 13475
rect -1073 13429 -1062 13475
rect -954 13429 -943 13475
rect -569 13429 -558 13475
rect -450 13429 -439 13475
rect -65 13429 -54 13475
rect 54 13429 65 13475
rect 439 13429 450 13475
rect 558 13429 569 13475
rect 943 13429 954 13475
rect 1062 13429 1073 13475
rect 1447 13429 1458 13475
rect 1566 13429 1577 13475
rect 1951 13429 1962 13475
rect 2070 13429 2081 13475
rect 2455 13429 2466 13475
rect -2466 13309 -2455 13355
rect -2081 13309 -2070 13355
rect -1962 13309 -1951 13355
rect -1577 13309 -1566 13355
rect -1458 13309 -1447 13355
rect -1073 13309 -1062 13355
rect -954 13309 -943 13355
rect -569 13309 -558 13355
rect -450 13309 -439 13355
rect -65 13309 -54 13355
rect 54 13309 65 13355
rect 439 13309 450 13355
rect 558 13309 569 13355
rect 943 13309 954 13355
rect 1062 13309 1073 13355
rect 1447 13309 1458 13355
rect 1566 13309 1577 13355
rect 1951 13309 1962 13355
rect 2070 13309 2081 13355
rect 2455 13309 2466 13355
rect -2543 13263 -2497 13274
rect -2543 11278 -2497 11289
rect -2039 13263 -1993 13274
rect -2039 11278 -1993 11289
rect -1535 13263 -1489 13274
rect -1535 11278 -1489 11289
rect -1031 13263 -985 13274
rect -1031 11278 -985 11289
rect -527 13263 -481 13274
rect -527 11278 -481 11289
rect -23 13263 23 13274
rect -23 11278 23 11289
rect 481 13263 527 13274
rect 481 11278 527 11289
rect 985 13263 1031 13274
rect 985 11278 1031 11289
rect 1489 13263 1535 13274
rect 1489 11278 1535 11289
rect 1993 13263 2039 13274
rect 1993 11278 2039 11289
rect 2497 13263 2543 13274
rect 2497 11278 2543 11289
rect -2466 11197 -2455 11243
rect -2081 11197 -2070 11243
rect -1962 11197 -1951 11243
rect -1577 11197 -1566 11243
rect -1458 11197 -1447 11243
rect -1073 11197 -1062 11243
rect -954 11197 -943 11243
rect -569 11197 -558 11243
rect -450 11197 -439 11243
rect -65 11197 -54 11243
rect 54 11197 65 11243
rect 439 11197 450 11243
rect 558 11197 569 11243
rect 943 11197 954 11243
rect 1062 11197 1073 11243
rect 1447 11197 1458 11243
rect 1566 11197 1577 11243
rect 1951 11197 1962 11243
rect 2070 11197 2081 11243
rect 2455 11197 2466 11243
rect -2466 11077 -2455 11123
rect -2081 11077 -2070 11123
rect -1962 11077 -1951 11123
rect -1577 11077 -1566 11123
rect -1458 11077 -1447 11123
rect -1073 11077 -1062 11123
rect -954 11077 -943 11123
rect -569 11077 -558 11123
rect -450 11077 -439 11123
rect -65 11077 -54 11123
rect 54 11077 65 11123
rect 439 11077 450 11123
rect 558 11077 569 11123
rect 943 11077 954 11123
rect 1062 11077 1073 11123
rect 1447 11077 1458 11123
rect 1566 11077 1577 11123
rect 1951 11077 1962 11123
rect 2070 11077 2081 11123
rect 2455 11077 2466 11123
rect -2543 11031 -2497 11042
rect -2543 9046 -2497 9057
rect -2039 11031 -1993 11042
rect -2039 9046 -1993 9057
rect -1535 11031 -1489 11042
rect -1535 9046 -1489 9057
rect -1031 11031 -985 11042
rect -1031 9046 -985 9057
rect -527 11031 -481 11042
rect -527 9046 -481 9057
rect -23 11031 23 11042
rect -23 9046 23 9057
rect 481 11031 527 11042
rect 481 9046 527 9057
rect 985 11031 1031 11042
rect 985 9046 1031 9057
rect 1489 11031 1535 11042
rect 1489 9046 1535 9057
rect 1993 11031 2039 11042
rect 1993 9046 2039 9057
rect 2497 11031 2543 11042
rect 2497 9046 2543 9057
rect -2466 8965 -2455 9011
rect -2081 8965 -2070 9011
rect -1962 8965 -1951 9011
rect -1577 8965 -1566 9011
rect -1458 8965 -1447 9011
rect -1073 8965 -1062 9011
rect -954 8965 -943 9011
rect -569 8965 -558 9011
rect -450 8965 -439 9011
rect -65 8965 -54 9011
rect 54 8965 65 9011
rect 439 8965 450 9011
rect 558 8965 569 9011
rect 943 8965 954 9011
rect 1062 8965 1073 9011
rect 1447 8965 1458 9011
rect 1566 8965 1577 9011
rect 1951 8965 1962 9011
rect 2070 8965 2081 9011
rect 2455 8965 2466 9011
rect -2466 8845 -2455 8891
rect -2081 8845 -2070 8891
rect -1962 8845 -1951 8891
rect -1577 8845 -1566 8891
rect -1458 8845 -1447 8891
rect -1073 8845 -1062 8891
rect -954 8845 -943 8891
rect -569 8845 -558 8891
rect -450 8845 -439 8891
rect -65 8845 -54 8891
rect 54 8845 65 8891
rect 439 8845 450 8891
rect 558 8845 569 8891
rect 943 8845 954 8891
rect 1062 8845 1073 8891
rect 1447 8845 1458 8891
rect 1566 8845 1577 8891
rect 1951 8845 1962 8891
rect 2070 8845 2081 8891
rect 2455 8845 2466 8891
rect -2543 8799 -2497 8810
rect -2543 6814 -2497 6825
rect -2039 8799 -1993 8810
rect -2039 6814 -1993 6825
rect -1535 8799 -1489 8810
rect -1535 6814 -1489 6825
rect -1031 8799 -985 8810
rect -1031 6814 -985 6825
rect -527 8799 -481 8810
rect -527 6814 -481 6825
rect -23 8799 23 8810
rect -23 6814 23 6825
rect 481 8799 527 8810
rect 481 6814 527 6825
rect 985 8799 1031 8810
rect 985 6814 1031 6825
rect 1489 8799 1535 8810
rect 1489 6814 1535 6825
rect 1993 8799 2039 8810
rect 1993 6814 2039 6825
rect 2497 8799 2543 8810
rect 2497 6814 2543 6825
rect -2466 6733 -2455 6779
rect -2081 6733 -2070 6779
rect -1962 6733 -1951 6779
rect -1577 6733 -1566 6779
rect -1458 6733 -1447 6779
rect -1073 6733 -1062 6779
rect -954 6733 -943 6779
rect -569 6733 -558 6779
rect -450 6733 -439 6779
rect -65 6733 -54 6779
rect 54 6733 65 6779
rect 439 6733 450 6779
rect 558 6733 569 6779
rect 943 6733 954 6779
rect 1062 6733 1073 6779
rect 1447 6733 1458 6779
rect 1566 6733 1577 6779
rect 1951 6733 1962 6779
rect 2070 6733 2081 6779
rect 2455 6733 2466 6779
rect -2466 6613 -2455 6659
rect -2081 6613 -2070 6659
rect -1962 6613 -1951 6659
rect -1577 6613 -1566 6659
rect -1458 6613 -1447 6659
rect -1073 6613 -1062 6659
rect -954 6613 -943 6659
rect -569 6613 -558 6659
rect -450 6613 -439 6659
rect -65 6613 -54 6659
rect 54 6613 65 6659
rect 439 6613 450 6659
rect 558 6613 569 6659
rect 943 6613 954 6659
rect 1062 6613 1073 6659
rect 1447 6613 1458 6659
rect 1566 6613 1577 6659
rect 1951 6613 1962 6659
rect 2070 6613 2081 6659
rect 2455 6613 2466 6659
rect -2543 6567 -2497 6578
rect -2543 4582 -2497 4593
rect -2039 6567 -1993 6578
rect -2039 4582 -1993 4593
rect -1535 6567 -1489 6578
rect -1535 4582 -1489 4593
rect -1031 6567 -985 6578
rect -1031 4582 -985 4593
rect -527 6567 -481 6578
rect -527 4582 -481 4593
rect -23 6567 23 6578
rect -23 4582 23 4593
rect 481 6567 527 6578
rect 481 4582 527 4593
rect 985 6567 1031 6578
rect 985 4582 1031 4593
rect 1489 6567 1535 6578
rect 1489 4582 1535 4593
rect 1993 6567 2039 6578
rect 1993 4582 2039 4593
rect 2497 6567 2543 6578
rect 2497 4582 2543 4593
rect -2466 4501 -2455 4547
rect -2081 4501 -2070 4547
rect -1962 4501 -1951 4547
rect -1577 4501 -1566 4547
rect -1458 4501 -1447 4547
rect -1073 4501 -1062 4547
rect -954 4501 -943 4547
rect -569 4501 -558 4547
rect -450 4501 -439 4547
rect -65 4501 -54 4547
rect 54 4501 65 4547
rect 439 4501 450 4547
rect 558 4501 569 4547
rect 943 4501 954 4547
rect 1062 4501 1073 4547
rect 1447 4501 1458 4547
rect 1566 4501 1577 4547
rect 1951 4501 1962 4547
rect 2070 4501 2081 4547
rect 2455 4501 2466 4547
rect -2466 4381 -2455 4427
rect -2081 4381 -2070 4427
rect -1962 4381 -1951 4427
rect -1577 4381 -1566 4427
rect -1458 4381 -1447 4427
rect -1073 4381 -1062 4427
rect -954 4381 -943 4427
rect -569 4381 -558 4427
rect -450 4381 -439 4427
rect -65 4381 -54 4427
rect 54 4381 65 4427
rect 439 4381 450 4427
rect 558 4381 569 4427
rect 943 4381 954 4427
rect 1062 4381 1073 4427
rect 1447 4381 1458 4427
rect 1566 4381 1577 4427
rect 1951 4381 1962 4427
rect 2070 4381 2081 4427
rect 2455 4381 2466 4427
rect -2543 4335 -2497 4346
rect -2543 2350 -2497 2361
rect -2039 4335 -1993 4346
rect -2039 2350 -1993 2361
rect -1535 4335 -1489 4346
rect -1535 2350 -1489 2361
rect -1031 4335 -985 4346
rect -1031 2350 -985 2361
rect -527 4335 -481 4346
rect -527 2350 -481 2361
rect -23 4335 23 4346
rect -23 2350 23 2361
rect 481 4335 527 4346
rect 481 2350 527 2361
rect 985 4335 1031 4346
rect 985 2350 1031 2361
rect 1489 4335 1535 4346
rect 1489 2350 1535 2361
rect 1993 4335 2039 4346
rect 1993 2350 2039 2361
rect 2497 4335 2543 4346
rect 2497 2350 2543 2361
rect -2466 2269 -2455 2315
rect -2081 2269 -2070 2315
rect -1962 2269 -1951 2315
rect -1577 2269 -1566 2315
rect -1458 2269 -1447 2315
rect -1073 2269 -1062 2315
rect -954 2269 -943 2315
rect -569 2269 -558 2315
rect -450 2269 -439 2315
rect -65 2269 -54 2315
rect 54 2269 65 2315
rect 439 2269 450 2315
rect 558 2269 569 2315
rect 943 2269 954 2315
rect 1062 2269 1073 2315
rect 1447 2269 1458 2315
rect 1566 2269 1577 2315
rect 1951 2269 1962 2315
rect 2070 2269 2081 2315
rect 2455 2269 2466 2315
rect -2466 2149 -2455 2195
rect -2081 2149 -2070 2195
rect -1962 2149 -1951 2195
rect -1577 2149 -1566 2195
rect -1458 2149 -1447 2195
rect -1073 2149 -1062 2195
rect -954 2149 -943 2195
rect -569 2149 -558 2195
rect -450 2149 -439 2195
rect -65 2149 -54 2195
rect 54 2149 65 2195
rect 439 2149 450 2195
rect 558 2149 569 2195
rect 943 2149 954 2195
rect 1062 2149 1073 2195
rect 1447 2149 1458 2195
rect 1566 2149 1577 2195
rect 1951 2149 1962 2195
rect 2070 2149 2081 2195
rect 2455 2149 2466 2195
rect -2543 2103 -2497 2114
rect -2543 118 -2497 129
rect -2039 2103 -1993 2114
rect -2039 118 -1993 129
rect -1535 2103 -1489 2114
rect -1535 118 -1489 129
rect -1031 2103 -985 2114
rect -1031 118 -985 129
rect -527 2103 -481 2114
rect -527 118 -481 129
rect -23 2103 23 2114
rect -23 118 23 129
rect 481 2103 527 2114
rect 481 118 527 129
rect 985 2103 1031 2114
rect 985 118 1031 129
rect 1489 2103 1535 2114
rect 1489 118 1535 129
rect 1993 2103 2039 2114
rect 1993 118 2039 129
rect 2497 2103 2543 2114
rect 2497 118 2543 129
rect -2466 37 -2455 83
rect -2081 37 -2070 83
rect -1962 37 -1951 83
rect -1577 37 -1566 83
rect -1458 37 -1447 83
rect -1073 37 -1062 83
rect -954 37 -943 83
rect -569 37 -558 83
rect -450 37 -439 83
rect -65 37 -54 83
rect 54 37 65 83
rect 439 37 450 83
rect 558 37 569 83
rect 943 37 954 83
rect 1062 37 1073 83
rect 1447 37 1458 83
rect 1566 37 1577 83
rect 1951 37 1962 83
rect 2070 37 2081 83
rect 2455 37 2466 83
rect -2466 -83 -2455 -37
rect -2081 -83 -2070 -37
rect -1962 -83 -1951 -37
rect -1577 -83 -1566 -37
rect -1458 -83 -1447 -37
rect -1073 -83 -1062 -37
rect -954 -83 -943 -37
rect -569 -83 -558 -37
rect -450 -83 -439 -37
rect -65 -83 -54 -37
rect 54 -83 65 -37
rect 439 -83 450 -37
rect 558 -83 569 -37
rect 943 -83 954 -37
rect 1062 -83 1073 -37
rect 1447 -83 1458 -37
rect 1566 -83 1577 -37
rect 1951 -83 1962 -37
rect 2070 -83 2081 -37
rect 2455 -83 2466 -37
rect -2543 -129 -2497 -118
rect -2543 -2114 -2497 -2103
rect -2039 -129 -1993 -118
rect -2039 -2114 -1993 -2103
rect -1535 -129 -1489 -118
rect -1535 -2114 -1489 -2103
rect -1031 -129 -985 -118
rect -1031 -2114 -985 -2103
rect -527 -129 -481 -118
rect -527 -2114 -481 -2103
rect -23 -129 23 -118
rect -23 -2114 23 -2103
rect 481 -129 527 -118
rect 481 -2114 527 -2103
rect 985 -129 1031 -118
rect 985 -2114 1031 -2103
rect 1489 -129 1535 -118
rect 1489 -2114 1535 -2103
rect 1993 -129 2039 -118
rect 1993 -2114 2039 -2103
rect 2497 -129 2543 -118
rect 2497 -2114 2543 -2103
rect -2466 -2195 -2455 -2149
rect -2081 -2195 -2070 -2149
rect -1962 -2195 -1951 -2149
rect -1577 -2195 -1566 -2149
rect -1458 -2195 -1447 -2149
rect -1073 -2195 -1062 -2149
rect -954 -2195 -943 -2149
rect -569 -2195 -558 -2149
rect -450 -2195 -439 -2149
rect -65 -2195 -54 -2149
rect 54 -2195 65 -2149
rect 439 -2195 450 -2149
rect 558 -2195 569 -2149
rect 943 -2195 954 -2149
rect 1062 -2195 1073 -2149
rect 1447 -2195 1458 -2149
rect 1566 -2195 1577 -2149
rect 1951 -2195 1962 -2149
rect 2070 -2195 2081 -2149
rect 2455 -2195 2466 -2149
rect -2466 -2315 -2455 -2269
rect -2081 -2315 -2070 -2269
rect -1962 -2315 -1951 -2269
rect -1577 -2315 -1566 -2269
rect -1458 -2315 -1447 -2269
rect -1073 -2315 -1062 -2269
rect -954 -2315 -943 -2269
rect -569 -2315 -558 -2269
rect -450 -2315 -439 -2269
rect -65 -2315 -54 -2269
rect 54 -2315 65 -2269
rect 439 -2315 450 -2269
rect 558 -2315 569 -2269
rect 943 -2315 954 -2269
rect 1062 -2315 1073 -2269
rect 1447 -2315 1458 -2269
rect 1566 -2315 1577 -2269
rect 1951 -2315 1962 -2269
rect 2070 -2315 2081 -2269
rect 2455 -2315 2466 -2269
rect -2543 -2361 -2497 -2350
rect -2543 -4346 -2497 -4335
rect -2039 -2361 -1993 -2350
rect -2039 -4346 -1993 -4335
rect -1535 -2361 -1489 -2350
rect -1535 -4346 -1489 -4335
rect -1031 -2361 -985 -2350
rect -1031 -4346 -985 -4335
rect -527 -2361 -481 -2350
rect -527 -4346 -481 -4335
rect -23 -2361 23 -2350
rect -23 -4346 23 -4335
rect 481 -2361 527 -2350
rect 481 -4346 527 -4335
rect 985 -2361 1031 -2350
rect 985 -4346 1031 -4335
rect 1489 -2361 1535 -2350
rect 1489 -4346 1535 -4335
rect 1993 -2361 2039 -2350
rect 1993 -4346 2039 -4335
rect 2497 -2361 2543 -2350
rect 2497 -4346 2543 -4335
rect -2466 -4427 -2455 -4381
rect -2081 -4427 -2070 -4381
rect -1962 -4427 -1951 -4381
rect -1577 -4427 -1566 -4381
rect -1458 -4427 -1447 -4381
rect -1073 -4427 -1062 -4381
rect -954 -4427 -943 -4381
rect -569 -4427 -558 -4381
rect -450 -4427 -439 -4381
rect -65 -4427 -54 -4381
rect 54 -4427 65 -4381
rect 439 -4427 450 -4381
rect 558 -4427 569 -4381
rect 943 -4427 954 -4381
rect 1062 -4427 1073 -4381
rect 1447 -4427 1458 -4381
rect 1566 -4427 1577 -4381
rect 1951 -4427 1962 -4381
rect 2070 -4427 2081 -4381
rect 2455 -4427 2466 -4381
rect -2466 -4547 -2455 -4501
rect -2081 -4547 -2070 -4501
rect -1962 -4547 -1951 -4501
rect -1577 -4547 -1566 -4501
rect -1458 -4547 -1447 -4501
rect -1073 -4547 -1062 -4501
rect -954 -4547 -943 -4501
rect -569 -4547 -558 -4501
rect -450 -4547 -439 -4501
rect -65 -4547 -54 -4501
rect 54 -4547 65 -4501
rect 439 -4547 450 -4501
rect 558 -4547 569 -4501
rect 943 -4547 954 -4501
rect 1062 -4547 1073 -4501
rect 1447 -4547 1458 -4501
rect 1566 -4547 1577 -4501
rect 1951 -4547 1962 -4501
rect 2070 -4547 2081 -4501
rect 2455 -4547 2466 -4501
rect -2543 -4593 -2497 -4582
rect -2543 -6578 -2497 -6567
rect -2039 -4593 -1993 -4582
rect -2039 -6578 -1993 -6567
rect -1535 -4593 -1489 -4582
rect -1535 -6578 -1489 -6567
rect -1031 -4593 -985 -4582
rect -1031 -6578 -985 -6567
rect -527 -4593 -481 -4582
rect -527 -6578 -481 -6567
rect -23 -4593 23 -4582
rect -23 -6578 23 -6567
rect 481 -4593 527 -4582
rect 481 -6578 527 -6567
rect 985 -4593 1031 -4582
rect 985 -6578 1031 -6567
rect 1489 -4593 1535 -4582
rect 1489 -6578 1535 -6567
rect 1993 -4593 2039 -4582
rect 1993 -6578 2039 -6567
rect 2497 -4593 2543 -4582
rect 2497 -6578 2543 -6567
rect -2466 -6659 -2455 -6613
rect -2081 -6659 -2070 -6613
rect -1962 -6659 -1951 -6613
rect -1577 -6659 -1566 -6613
rect -1458 -6659 -1447 -6613
rect -1073 -6659 -1062 -6613
rect -954 -6659 -943 -6613
rect -569 -6659 -558 -6613
rect -450 -6659 -439 -6613
rect -65 -6659 -54 -6613
rect 54 -6659 65 -6613
rect 439 -6659 450 -6613
rect 558 -6659 569 -6613
rect 943 -6659 954 -6613
rect 1062 -6659 1073 -6613
rect 1447 -6659 1458 -6613
rect 1566 -6659 1577 -6613
rect 1951 -6659 1962 -6613
rect 2070 -6659 2081 -6613
rect 2455 -6659 2466 -6613
rect -2466 -6779 -2455 -6733
rect -2081 -6779 -2070 -6733
rect -1962 -6779 -1951 -6733
rect -1577 -6779 -1566 -6733
rect -1458 -6779 -1447 -6733
rect -1073 -6779 -1062 -6733
rect -954 -6779 -943 -6733
rect -569 -6779 -558 -6733
rect -450 -6779 -439 -6733
rect -65 -6779 -54 -6733
rect 54 -6779 65 -6733
rect 439 -6779 450 -6733
rect 558 -6779 569 -6733
rect 943 -6779 954 -6733
rect 1062 -6779 1073 -6733
rect 1447 -6779 1458 -6733
rect 1566 -6779 1577 -6733
rect 1951 -6779 1962 -6733
rect 2070 -6779 2081 -6733
rect 2455 -6779 2466 -6733
rect -2543 -6825 -2497 -6814
rect -2543 -8810 -2497 -8799
rect -2039 -6825 -1993 -6814
rect -2039 -8810 -1993 -8799
rect -1535 -6825 -1489 -6814
rect -1535 -8810 -1489 -8799
rect -1031 -6825 -985 -6814
rect -1031 -8810 -985 -8799
rect -527 -6825 -481 -6814
rect -527 -8810 -481 -8799
rect -23 -6825 23 -6814
rect -23 -8810 23 -8799
rect 481 -6825 527 -6814
rect 481 -8810 527 -8799
rect 985 -6825 1031 -6814
rect 985 -8810 1031 -8799
rect 1489 -6825 1535 -6814
rect 1489 -8810 1535 -8799
rect 1993 -6825 2039 -6814
rect 1993 -8810 2039 -8799
rect 2497 -6825 2543 -6814
rect 2497 -8810 2543 -8799
rect -2466 -8891 -2455 -8845
rect -2081 -8891 -2070 -8845
rect -1962 -8891 -1951 -8845
rect -1577 -8891 -1566 -8845
rect -1458 -8891 -1447 -8845
rect -1073 -8891 -1062 -8845
rect -954 -8891 -943 -8845
rect -569 -8891 -558 -8845
rect -450 -8891 -439 -8845
rect -65 -8891 -54 -8845
rect 54 -8891 65 -8845
rect 439 -8891 450 -8845
rect 558 -8891 569 -8845
rect 943 -8891 954 -8845
rect 1062 -8891 1073 -8845
rect 1447 -8891 1458 -8845
rect 1566 -8891 1577 -8845
rect 1951 -8891 1962 -8845
rect 2070 -8891 2081 -8845
rect 2455 -8891 2466 -8845
rect -2466 -9011 -2455 -8965
rect -2081 -9011 -2070 -8965
rect -1962 -9011 -1951 -8965
rect -1577 -9011 -1566 -8965
rect -1458 -9011 -1447 -8965
rect -1073 -9011 -1062 -8965
rect -954 -9011 -943 -8965
rect -569 -9011 -558 -8965
rect -450 -9011 -439 -8965
rect -65 -9011 -54 -8965
rect 54 -9011 65 -8965
rect 439 -9011 450 -8965
rect 558 -9011 569 -8965
rect 943 -9011 954 -8965
rect 1062 -9011 1073 -8965
rect 1447 -9011 1458 -8965
rect 1566 -9011 1577 -8965
rect 1951 -9011 1962 -8965
rect 2070 -9011 2081 -8965
rect 2455 -9011 2466 -8965
rect -2543 -9057 -2497 -9046
rect -2543 -11042 -2497 -11031
rect -2039 -9057 -1993 -9046
rect -2039 -11042 -1993 -11031
rect -1535 -9057 -1489 -9046
rect -1535 -11042 -1489 -11031
rect -1031 -9057 -985 -9046
rect -1031 -11042 -985 -11031
rect -527 -9057 -481 -9046
rect -527 -11042 -481 -11031
rect -23 -9057 23 -9046
rect -23 -11042 23 -11031
rect 481 -9057 527 -9046
rect 481 -11042 527 -11031
rect 985 -9057 1031 -9046
rect 985 -11042 1031 -11031
rect 1489 -9057 1535 -9046
rect 1489 -11042 1535 -11031
rect 1993 -9057 2039 -9046
rect 1993 -11042 2039 -11031
rect 2497 -9057 2543 -9046
rect 2497 -11042 2543 -11031
rect -2466 -11123 -2455 -11077
rect -2081 -11123 -2070 -11077
rect -1962 -11123 -1951 -11077
rect -1577 -11123 -1566 -11077
rect -1458 -11123 -1447 -11077
rect -1073 -11123 -1062 -11077
rect -954 -11123 -943 -11077
rect -569 -11123 -558 -11077
rect -450 -11123 -439 -11077
rect -65 -11123 -54 -11077
rect 54 -11123 65 -11077
rect 439 -11123 450 -11077
rect 558 -11123 569 -11077
rect 943 -11123 954 -11077
rect 1062 -11123 1073 -11077
rect 1447 -11123 1458 -11077
rect 1566 -11123 1577 -11077
rect 1951 -11123 1962 -11077
rect 2070 -11123 2081 -11077
rect 2455 -11123 2466 -11077
rect -2466 -11243 -2455 -11197
rect -2081 -11243 -2070 -11197
rect -1962 -11243 -1951 -11197
rect -1577 -11243 -1566 -11197
rect -1458 -11243 -1447 -11197
rect -1073 -11243 -1062 -11197
rect -954 -11243 -943 -11197
rect -569 -11243 -558 -11197
rect -450 -11243 -439 -11197
rect -65 -11243 -54 -11197
rect 54 -11243 65 -11197
rect 439 -11243 450 -11197
rect 558 -11243 569 -11197
rect 943 -11243 954 -11197
rect 1062 -11243 1073 -11197
rect 1447 -11243 1458 -11197
rect 1566 -11243 1577 -11197
rect 1951 -11243 1962 -11197
rect 2070 -11243 2081 -11197
rect 2455 -11243 2466 -11197
rect -2543 -11289 -2497 -11278
rect -2543 -13274 -2497 -13263
rect -2039 -11289 -1993 -11278
rect -2039 -13274 -1993 -13263
rect -1535 -11289 -1489 -11278
rect -1535 -13274 -1489 -13263
rect -1031 -11289 -985 -11278
rect -1031 -13274 -985 -13263
rect -527 -11289 -481 -11278
rect -527 -13274 -481 -13263
rect -23 -11289 23 -11278
rect -23 -13274 23 -13263
rect 481 -11289 527 -11278
rect 481 -13274 527 -13263
rect 985 -11289 1031 -11278
rect 985 -13274 1031 -13263
rect 1489 -11289 1535 -11278
rect 1489 -13274 1535 -13263
rect 1993 -11289 2039 -11278
rect 1993 -13274 2039 -13263
rect 2497 -11289 2543 -11278
rect 2497 -13274 2543 -13263
rect -2466 -13355 -2455 -13309
rect -2081 -13355 -2070 -13309
rect -1962 -13355 -1951 -13309
rect -1577 -13355 -1566 -13309
rect -1458 -13355 -1447 -13309
rect -1073 -13355 -1062 -13309
rect -954 -13355 -943 -13309
rect -569 -13355 -558 -13309
rect -450 -13355 -439 -13309
rect -65 -13355 -54 -13309
rect 54 -13355 65 -13309
rect 439 -13355 450 -13309
rect 558 -13355 569 -13309
rect 943 -13355 954 -13309
rect 1062 -13355 1073 -13309
rect 1447 -13355 1458 -13309
rect 1566 -13355 1577 -13309
rect 1951 -13355 1962 -13309
rect 2070 -13355 2081 -13309
rect 2455 -13355 2466 -13309
rect -2466 -13475 -2455 -13429
rect -2081 -13475 -2070 -13429
rect -1962 -13475 -1951 -13429
rect -1577 -13475 -1566 -13429
rect -1458 -13475 -1447 -13429
rect -1073 -13475 -1062 -13429
rect -954 -13475 -943 -13429
rect -569 -13475 -558 -13429
rect -450 -13475 -439 -13429
rect -65 -13475 -54 -13429
rect 54 -13475 65 -13429
rect 439 -13475 450 -13429
rect 558 -13475 569 -13429
rect 943 -13475 954 -13429
rect 1062 -13475 1073 -13429
rect 1447 -13475 1458 -13429
rect 1566 -13475 1577 -13429
rect 1951 -13475 1962 -13429
rect 2070 -13475 2081 -13429
rect 2455 -13475 2466 -13429
rect -2543 -13521 -2497 -13510
rect -2543 -15506 -2497 -15495
rect -2039 -13521 -1993 -13510
rect -2039 -15506 -1993 -15495
rect -1535 -13521 -1489 -13510
rect -1535 -15506 -1489 -15495
rect -1031 -13521 -985 -13510
rect -1031 -15506 -985 -15495
rect -527 -13521 -481 -13510
rect -527 -15506 -481 -15495
rect -23 -13521 23 -13510
rect -23 -15506 23 -15495
rect 481 -13521 527 -13510
rect 481 -15506 527 -15495
rect 985 -13521 1031 -13510
rect 985 -15506 1031 -15495
rect 1489 -13521 1535 -13510
rect 1489 -15506 1535 -15495
rect 1993 -13521 2039 -13510
rect 1993 -15506 2039 -15495
rect 2497 -13521 2543 -13510
rect 2497 -15506 2543 -15495
rect -2466 -15587 -2455 -15541
rect -2081 -15587 -2070 -15541
rect -1962 -15587 -1951 -15541
rect -1577 -15587 -1566 -15541
rect -1458 -15587 -1447 -15541
rect -1073 -15587 -1062 -15541
rect -954 -15587 -943 -15541
rect -569 -15587 -558 -15541
rect -450 -15587 -439 -15541
rect -65 -15587 -54 -15541
rect 54 -15587 65 -15541
rect 439 -15587 450 -15541
rect 558 -15587 569 -15541
rect 943 -15587 954 -15541
rect 1062 -15587 1073 -15541
rect 1447 -15587 1458 -15541
rect 1566 -15587 1577 -15541
rect 1951 -15587 1962 -15541
rect 2070 -15587 2081 -15541
rect 2455 -15587 2466 -15541
rect -2466 -15707 -2455 -15661
rect -2081 -15707 -2070 -15661
rect -1962 -15707 -1951 -15661
rect -1577 -15707 -1566 -15661
rect -1458 -15707 -1447 -15661
rect -1073 -15707 -1062 -15661
rect -954 -15707 -943 -15661
rect -569 -15707 -558 -15661
rect -450 -15707 -439 -15661
rect -65 -15707 -54 -15661
rect 54 -15707 65 -15661
rect 439 -15707 450 -15661
rect 558 -15707 569 -15661
rect 943 -15707 954 -15661
rect 1062 -15707 1073 -15661
rect 1447 -15707 1458 -15661
rect 1566 -15707 1577 -15661
rect 1951 -15707 1962 -15661
rect 2070 -15707 2081 -15661
rect 2455 -15707 2466 -15661
rect -2543 -15753 -2497 -15742
rect -2543 -17738 -2497 -17727
rect -2039 -15753 -1993 -15742
rect -2039 -17738 -1993 -17727
rect -1535 -15753 -1489 -15742
rect -1535 -17738 -1489 -17727
rect -1031 -15753 -985 -15742
rect -1031 -17738 -985 -17727
rect -527 -15753 -481 -15742
rect -527 -17738 -481 -17727
rect -23 -15753 23 -15742
rect -23 -17738 23 -17727
rect 481 -15753 527 -15742
rect 481 -17738 527 -17727
rect 985 -15753 1031 -15742
rect 985 -17738 1031 -17727
rect 1489 -15753 1535 -15742
rect 1489 -17738 1535 -17727
rect 1993 -15753 2039 -15742
rect 1993 -17738 2039 -17727
rect 2497 -15753 2543 -15742
rect 2497 -17738 2543 -17727
rect -2466 -17819 -2455 -17773
rect -2081 -17819 -2070 -17773
rect -1962 -17819 -1951 -17773
rect -1577 -17819 -1566 -17773
rect -1458 -17819 -1447 -17773
rect -1073 -17819 -1062 -17773
rect -954 -17819 -943 -17773
rect -569 -17819 -558 -17773
rect -450 -17819 -439 -17773
rect -65 -17819 -54 -17773
rect 54 -17819 65 -17773
rect 439 -17819 450 -17773
rect 558 -17819 569 -17773
rect 943 -17819 954 -17773
rect 1062 -17819 1073 -17773
rect 1447 -17819 1458 -17773
rect 1566 -17819 1577 -17773
rect 1951 -17819 1962 -17773
rect 2070 -17819 2081 -17773
rect 2455 -17819 2466 -17773
rect -2466 -17939 -2455 -17893
rect -2081 -17939 -2070 -17893
rect -1962 -17939 -1951 -17893
rect -1577 -17939 -1566 -17893
rect -1458 -17939 -1447 -17893
rect -1073 -17939 -1062 -17893
rect -954 -17939 -943 -17893
rect -569 -17939 -558 -17893
rect -450 -17939 -439 -17893
rect -65 -17939 -54 -17893
rect 54 -17939 65 -17893
rect 439 -17939 450 -17893
rect 558 -17939 569 -17893
rect 943 -17939 954 -17893
rect 1062 -17939 1073 -17893
rect 1447 -17939 1458 -17893
rect 1566 -17939 1577 -17893
rect 1951 -17939 1962 -17893
rect 2070 -17939 2081 -17893
rect 2455 -17939 2466 -17893
rect -2543 -17985 -2497 -17974
rect -2543 -19970 -2497 -19959
rect -2039 -17985 -1993 -17974
rect -2039 -19970 -1993 -19959
rect -1535 -17985 -1489 -17974
rect -1535 -19970 -1489 -19959
rect -1031 -17985 -985 -17974
rect -1031 -19970 -985 -19959
rect -527 -17985 -481 -17974
rect -527 -19970 -481 -19959
rect -23 -17985 23 -17974
rect -23 -19970 23 -19959
rect 481 -17985 527 -17974
rect 481 -19970 527 -19959
rect 985 -17985 1031 -17974
rect 985 -19970 1031 -19959
rect 1489 -17985 1535 -17974
rect 1489 -19970 1535 -19959
rect 1993 -17985 2039 -17974
rect 1993 -19970 2039 -19959
rect 2497 -17985 2543 -17974
rect 2497 -19970 2543 -19959
rect -2466 -20051 -2455 -20005
rect -2081 -20051 -2070 -20005
rect -1962 -20051 -1951 -20005
rect -1577 -20051 -1566 -20005
rect -1458 -20051 -1447 -20005
rect -1073 -20051 -1062 -20005
rect -954 -20051 -943 -20005
rect -569 -20051 -558 -20005
rect -450 -20051 -439 -20005
rect -65 -20051 -54 -20005
rect 54 -20051 65 -20005
rect 439 -20051 450 -20005
rect 558 -20051 569 -20005
rect 943 -20051 954 -20005
rect 1062 -20051 1073 -20005
rect 1447 -20051 1458 -20005
rect 1566 -20051 1577 -20005
rect 1951 -20051 1962 -20005
rect 2070 -20051 2081 -20005
rect 2455 -20051 2466 -20005
rect -2466 -20171 -2455 -20125
rect -2081 -20171 -2070 -20125
rect -1962 -20171 -1951 -20125
rect -1577 -20171 -1566 -20125
rect -1458 -20171 -1447 -20125
rect -1073 -20171 -1062 -20125
rect -954 -20171 -943 -20125
rect -569 -20171 -558 -20125
rect -450 -20171 -439 -20125
rect -65 -20171 -54 -20125
rect 54 -20171 65 -20125
rect 439 -20171 450 -20125
rect 558 -20171 569 -20125
rect 943 -20171 954 -20125
rect 1062 -20171 1073 -20125
rect 1447 -20171 1458 -20125
rect 1566 -20171 1577 -20125
rect 1951 -20171 1962 -20125
rect 2070 -20171 2081 -20125
rect 2455 -20171 2466 -20125
rect -2543 -20217 -2497 -20206
rect -2543 -22202 -2497 -22191
rect -2039 -20217 -1993 -20206
rect -2039 -22202 -1993 -22191
rect -1535 -20217 -1489 -20206
rect -1535 -22202 -1489 -22191
rect -1031 -20217 -985 -20206
rect -1031 -22202 -985 -22191
rect -527 -20217 -481 -20206
rect -527 -22202 -481 -22191
rect -23 -20217 23 -20206
rect -23 -22202 23 -22191
rect 481 -20217 527 -20206
rect 481 -22202 527 -22191
rect 985 -20217 1031 -20206
rect 985 -22202 1031 -22191
rect 1489 -20217 1535 -20206
rect 1489 -22202 1535 -22191
rect 1993 -20217 2039 -20206
rect 1993 -22202 2039 -22191
rect 2497 -20217 2543 -20206
rect 2497 -22202 2543 -22191
rect -2466 -22283 -2455 -22237
rect -2081 -22283 -2070 -22237
rect -1962 -22283 -1951 -22237
rect -1577 -22283 -1566 -22237
rect -1458 -22283 -1447 -22237
rect -1073 -22283 -1062 -22237
rect -954 -22283 -943 -22237
rect -569 -22283 -558 -22237
rect -450 -22283 -439 -22237
rect -65 -22283 -54 -22237
rect 54 -22283 65 -22237
rect 439 -22283 450 -22237
rect 558 -22283 569 -22237
rect 943 -22283 954 -22237
rect 1062 -22283 1073 -22237
rect 1447 -22283 1458 -22237
rect 1566 -22283 1577 -22237
rect 1951 -22283 1962 -22237
rect 2070 -22283 2081 -22237
rect 2455 -22283 2466 -22237
rect -2466 -22403 -2455 -22357
rect -2081 -22403 -2070 -22357
rect -1962 -22403 -1951 -22357
rect -1577 -22403 -1566 -22357
rect -1458 -22403 -1447 -22357
rect -1073 -22403 -1062 -22357
rect -954 -22403 -943 -22357
rect -569 -22403 -558 -22357
rect -450 -22403 -439 -22357
rect -65 -22403 -54 -22357
rect 54 -22403 65 -22357
rect 439 -22403 450 -22357
rect 558 -22403 569 -22357
rect 943 -22403 954 -22357
rect 1062 -22403 1073 -22357
rect 1447 -22403 1458 -22357
rect 1566 -22403 1577 -22357
rect 1951 -22403 1962 -22357
rect 2070 -22403 2081 -22357
rect 2455 -22403 2466 -22357
rect -2543 -22449 -2497 -22438
rect -2543 -24434 -2497 -24423
rect -2039 -22449 -1993 -22438
rect -2039 -24434 -1993 -24423
rect -1535 -22449 -1489 -22438
rect -1535 -24434 -1489 -24423
rect -1031 -22449 -985 -22438
rect -1031 -24434 -985 -24423
rect -527 -22449 -481 -22438
rect -527 -24434 -481 -24423
rect -23 -22449 23 -22438
rect -23 -24434 23 -24423
rect 481 -22449 527 -22438
rect 481 -24434 527 -24423
rect 985 -22449 1031 -22438
rect 985 -24434 1031 -24423
rect 1489 -22449 1535 -22438
rect 1489 -24434 1535 -24423
rect 1993 -22449 2039 -22438
rect 1993 -24434 2039 -24423
rect 2497 -22449 2543 -22438
rect 2497 -24434 2543 -24423
rect -2466 -24515 -2455 -24469
rect -2081 -24515 -2070 -24469
rect -1962 -24515 -1951 -24469
rect -1577 -24515 -1566 -24469
rect -1458 -24515 -1447 -24469
rect -1073 -24515 -1062 -24469
rect -954 -24515 -943 -24469
rect -569 -24515 -558 -24469
rect -450 -24515 -439 -24469
rect -65 -24515 -54 -24469
rect 54 -24515 65 -24469
rect 439 -24515 450 -24469
rect 558 -24515 569 -24469
rect 943 -24515 954 -24469
rect 1062 -24515 1073 -24469
rect 1447 -24515 1458 -24469
rect 1566 -24515 1577 -24469
rect 1951 -24515 1962 -24469
rect 2070 -24515 2081 -24469
rect 2455 -24515 2466 -24469
rect -2466 -24635 -2455 -24589
rect -2081 -24635 -2070 -24589
rect -1962 -24635 -1951 -24589
rect -1577 -24635 -1566 -24589
rect -1458 -24635 -1447 -24589
rect -1073 -24635 -1062 -24589
rect -954 -24635 -943 -24589
rect -569 -24635 -558 -24589
rect -450 -24635 -439 -24589
rect -65 -24635 -54 -24589
rect 54 -24635 65 -24589
rect 439 -24635 450 -24589
rect 558 -24635 569 -24589
rect 943 -24635 954 -24589
rect 1062 -24635 1073 -24589
rect 1447 -24635 1458 -24589
rect 1566 -24635 1577 -24589
rect 1951 -24635 1962 -24589
rect 2070 -24635 2081 -24589
rect 2455 -24635 2466 -24589
rect -2543 -24681 -2497 -24670
rect -2543 -26666 -2497 -26655
rect -2039 -24681 -1993 -24670
rect -2039 -26666 -1993 -26655
rect -1535 -24681 -1489 -24670
rect -1535 -26666 -1489 -26655
rect -1031 -24681 -985 -24670
rect -1031 -26666 -985 -26655
rect -527 -24681 -481 -24670
rect -527 -26666 -481 -26655
rect -23 -24681 23 -24670
rect -23 -26666 23 -26655
rect 481 -24681 527 -24670
rect 481 -26666 527 -26655
rect 985 -24681 1031 -24670
rect 985 -26666 1031 -26655
rect 1489 -24681 1535 -24670
rect 1489 -26666 1535 -26655
rect 1993 -24681 2039 -24670
rect 1993 -26666 2039 -26655
rect 2497 -24681 2543 -24670
rect 2497 -26666 2543 -26655
rect -2466 -26747 -2455 -26701
rect -2081 -26747 -2070 -26701
rect -1962 -26747 -1951 -26701
rect -1577 -26747 -1566 -26701
rect -1458 -26747 -1447 -26701
rect -1073 -26747 -1062 -26701
rect -954 -26747 -943 -26701
rect -569 -26747 -558 -26701
rect -450 -26747 -439 -26701
rect -65 -26747 -54 -26701
rect 54 -26747 65 -26701
rect 439 -26747 450 -26701
rect 558 -26747 569 -26701
rect 943 -26747 954 -26701
rect 1062 -26747 1073 -26701
rect 1447 -26747 1458 -26701
rect 1566 -26747 1577 -26701
rect 1951 -26747 1962 -26701
rect 2070 -26747 2081 -26701
rect 2455 -26747 2466 -26701
rect -2466 -26867 -2455 -26821
rect -2081 -26867 -2070 -26821
rect -1962 -26867 -1951 -26821
rect -1577 -26867 -1566 -26821
rect -1458 -26867 -1447 -26821
rect -1073 -26867 -1062 -26821
rect -954 -26867 -943 -26821
rect -569 -26867 -558 -26821
rect -450 -26867 -439 -26821
rect -65 -26867 -54 -26821
rect 54 -26867 65 -26821
rect 439 -26867 450 -26821
rect 558 -26867 569 -26821
rect 943 -26867 954 -26821
rect 1062 -26867 1073 -26821
rect 1447 -26867 1458 -26821
rect 1566 -26867 1577 -26821
rect 1951 -26867 1962 -26821
rect 2070 -26867 2081 -26821
rect 2455 -26867 2466 -26821
rect -2543 -26913 -2497 -26902
rect -2543 -28898 -2497 -28887
rect -2039 -26913 -1993 -26902
rect -2039 -28898 -1993 -28887
rect -1535 -26913 -1489 -26902
rect -1535 -28898 -1489 -28887
rect -1031 -26913 -985 -26902
rect -1031 -28898 -985 -28887
rect -527 -26913 -481 -26902
rect -527 -28898 -481 -28887
rect -23 -26913 23 -26902
rect -23 -28898 23 -28887
rect 481 -26913 527 -26902
rect 481 -28898 527 -28887
rect 985 -26913 1031 -26902
rect 985 -28898 1031 -28887
rect 1489 -26913 1535 -26902
rect 1489 -28898 1535 -28887
rect 1993 -26913 2039 -26902
rect 1993 -28898 2039 -28887
rect 2497 -26913 2543 -26902
rect 2497 -28898 2543 -28887
rect -2681 -29027 -2635 -28970
rect -2466 -28979 -2455 -28933
rect -2081 -28979 -2070 -28933
rect -1962 -28979 -1951 -28933
rect -1577 -28979 -1566 -28933
rect -1458 -28979 -1447 -28933
rect -1073 -28979 -1062 -28933
rect -954 -28979 -943 -28933
rect -569 -28979 -558 -28933
rect -450 -28979 -439 -28933
rect -65 -28979 -54 -28933
rect 54 -28979 65 -28933
rect 439 -28979 450 -28933
rect 558 -28979 569 -28933
rect 943 -28979 954 -28933
rect 1062 -28979 1073 -28933
rect 1447 -28979 1458 -28933
rect 1566 -28979 1577 -28933
rect 1951 -28979 1962 -28933
rect 2070 -28979 2081 -28933
rect 2455 -28979 2466 -28933
rect 2635 -29027 2681 -28970
rect -2681 -29073 2681 -29027
<< properties >>
string FIXED_BBOX -2658 -29050 2658 29050
string gencell nfet_03v3
string library gf180mcu
string parameters w 10.0 l 2.0 m 26 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
