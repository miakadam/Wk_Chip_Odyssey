magic
tech gf180mcuD
magscale 1 10
timestamp 1757668360
<< error_p >>
rect -130 118 -119 164
rect 54 118 65 164
rect -130 -164 -119 -118
rect 54 -164 65 -118
<< pwell >>
rect -382 -295 382 295
<< nmos >>
rect -132 -85 -52 85
rect 52 -85 132 85
<< ndiff >>
rect -220 72 -132 85
rect -220 -72 -207 72
rect -161 -72 -132 72
rect -220 -85 -132 -72
rect -52 72 52 85
rect -52 -72 -23 72
rect 23 -72 52 72
rect -52 -85 52 -72
rect 132 72 220 85
rect 132 -72 161 72
rect 207 -72 220 72
rect 132 -85 220 -72
<< ndiffc >>
rect -207 -72 -161 72
rect -23 -72 23 72
rect 161 -72 207 72
<< psubdiff >>
rect -358 199 358 271
rect -358 155 -286 199
rect -358 -155 -345 155
rect -299 -155 -286 155
rect 286 155 358 199
rect -358 -199 -286 -155
rect 286 -155 299 155
rect 345 -155 358 155
rect 286 -199 358 -155
rect -358 -271 358 -199
<< psubdiffcont >>
rect -345 -155 -299 155
rect 299 -155 345 155
<< polysilicon >>
rect -132 164 -52 177
rect -132 118 -119 164
rect -65 118 -52 164
rect -132 85 -52 118
rect 52 164 132 177
rect 52 118 65 164
rect 119 118 132 164
rect 52 85 132 118
rect -132 -118 -52 -85
rect -132 -164 -119 -118
rect -65 -164 -52 -118
rect -132 -177 -52 -164
rect 52 -118 132 -85
rect 52 -164 65 -118
rect 119 -164 132 -118
rect 52 -177 132 -164
<< polycontact >>
rect -119 118 -65 164
rect 65 118 119 164
rect -119 -164 -65 -118
rect 65 -164 119 -118
<< metal1 >>
rect -345 212 345 258
rect -345 155 -299 212
rect -130 118 -119 164
rect -65 118 -54 164
rect 54 118 65 164
rect 119 118 130 164
rect 299 155 345 212
rect -207 72 -161 83
rect -207 -83 -161 -72
rect -23 72 23 83
rect -23 -83 23 -72
rect 161 72 207 83
rect 161 -83 207 -72
rect -345 -212 -299 -155
rect -130 -164 -119 -118
rect -65 -164 -54 -118
rect 54 -164 65 -118
rect 119 -164 130 -118
rect 299 -212 345 -155
rect -345 -258 345 -212
<< properties >>
string FIXED_BBOX -322 -235 322 235
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.85 l 0.4 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
