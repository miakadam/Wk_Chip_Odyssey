magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< nwell >>
rect -954 -40494 954 40494
<< pmos >>
rect -704 37284 -304 40284
rect -200 37284 200 40284
rect 304 37284 704 40284
rect -704 34052 -304 37052
rect -200 34052 200 37052
rect 304 34052 704 37052
rect -704 30820 -304 33820
rect -200 30820 200 33820
rect 304 30820 704 33820
rect -704 27588 -304 30588
rect -200 27588 200 30588
rect 304 27588 704 30588
rect -704 24356 -304 27356
rect -200 24356 200 27356
rect 304 24356 704 27356
rect -704 21124 -304 24124
rect -200 21124 200 24124
rect 304 21124 704 24124
rect -704 17892 -304 20892
rect -200 17892 200 20892
rect 304 17892 704 20892
rect -704 14660 -304 17660
rect -200 14660 200 17660
rect 304 14660 704 17660
rect -704 11428 -304 14428
rect -200 11428 200 14428
rect 304 11428 704 14428
rect -704 8196 -304 11196
rect -200 8196 200 11196
rect 304 8196 704 11196
rect -704 4964 -304 7964
rect -200 4964 200 7964
rect 304 4964 704 7964
rect -704 1732 -304 4732
rect -200 1732 200 4732
rect 304 1732 704 4732
rect -704 -1500 -304 1500
rect -200 -1500 200 1500
rect 304 -1500 704 1500
rect -704 -4732 -304 -1732
rect -200 -4732 200 -1732
rect 304 -4732 704 -1732
rect -704 -7964 -304 -4964
rect -200 -7964 200 -4964
rect 304 -7964 704 -4964
rect -704 -11196 -304 -8196
rect -200 -11196 200 -8196
rect 304 -11196 704 -8196
rect -704 -14428 -304 -11428
rect -200 -14428 200 -11428
rect 304 -14428 704 -11428
rect -704 -17660 -304 -14660
rect -200 -17660 200 -14660
rect 304 -17660 704 -14660
rect -704 -20892 -304 -17892
rect -200 -20892 200 -17892
rect 304 -20892 704 -17892
rect -704 -24124 -304 -21124
rect -200 -24124 200 -21124
rect 304 -24124 704 -21124
rect -704 -27356 -304 -24356
rect -200 -27356 200 -24356
rect 304 -27356 704 -24356
rect -704 -30588 -304 -27588
rect -200 -30588 200 -27588
rect 304 -30588 704 -27588
rect -704 -33820 -304 -30820
rect -200 -33820 200 -30820
rect 304 -33820 704 -30820
rect -704 -37052 -304 -34052
rect -200 -37052 200 -34052
rect 304 -37052 704 -34052
rect -704 -40284 -304 -37284
rect -200 -40284 200 -37284
rect 304 -40284 704 -37284
<< pdiff >>
rect -792 40271 -704 40284
rect -792 37297 -779 40271
rect -733 37297 -704 40271
rect -792 37284 -704 37297
rect -304 40271 -200 40284
rect -304 37297 -275 40271
rect -229 37297 -200 40271
rect -304 37284 -200 37297
rect 200 40271 304 40284
rect 200 37297 229 40271
rect 275 37297 304 40271
rect 200 37284 304 37297
rect 704 40271 792 40284
rect 704 37297 733 40271
rect 779 37297 792 40271
rect 704 37284 792 37297
rect -792 37039 -704 37052
rect -792 34065 -779 37039
rect -733 34065 -704 37039
rect -792 34052 -704 34065
rect -304 37039 -200 37052
rect -304 34065 -275 37039
rect -229 34065 -200 37039
rect -304 34052 -200 34065
rect 200 37039 304 37052
rect 200 34065 229 37039
rect 275 34065 304 37039
rect 200 34052 304 34065
rect 704 37039 792 37052
rect 704 34065 733 37039
rect 779 34065 792 37039
rect 704 34052 792 34065
rect -792 33807 -704 33820
rect -792 30833 -779 33807
rect -733 30833 -704 33807
rect -792 30820 -704 30833
rect -304 33807 -200 33820
rect -304 30833 -275 33807
rect -229 30833 -200 33807
rect -304 30820 -200 30833
rect 200 33807 304 33820
rect 200 30833 229 33807
rect 275 30833 304 33807
rect 200 30820 304 30833
rect 704 33807 792 33820
rect 704 30833 733 33807
rect 779 30833 792 33807
rect 704 30820 792 30833
rect -792 30575 -704 30588
rect -792 27601 -779 30575
rect -733 27601 -704 30575
rect -792 27588 -704 27601
rect -304 30575 -200 30588
rect -304 27601 -275 30575
rect -229 27601 -200 30575
rect -304 27588 -200 27601
rect 200 30575 304 30588
rect 200 27601 229 30575
rect 275 27601 304 30575
rect 200 27588 304 27601
rect 704 30575 792 30588
rect 704 27601 733 30575
rect 779 27601 792 30575
rect 704 27588 792 27601
rect -792 27343 -704 27356
rect -792 24369 -779 27343
rect -733 24369 -704 27343
rect -792 24356 -704 24369
rect -304 27343 -200 27356
rect -304 24369 -275 27343
rect -229 24369 -200 27343
rect -304 24356 -200 24369
rect 200 27343 304 27356
rect 200 24369 229 27343
rect 275 24369 304 27343
rect 200 24356 304 24369
rect 704 27343 792 27356
rect 704 24369 733 27343
rect 779 24369 792 27343
rect 704 24356 792 24369
rect -792 24111 -704 24124
rect -792 21137 -779 24111
rect -733 21137 -704 24111
rect -792 21124 -704 21137
rect -304 24111 -200 24124
rect -304 21137 -275 24111
rect -229 21137 -200 24111
rect -304 21124 -200 21137
rect 200 24111 304 24124
rect 200 21137 229 24111
rect 275 21137 304 24111
rect 200 21124 304 21137
rect 704 24111 792 24124
rect 704 21137 733 24111
rect 779 21137 792 24111
rect 704 21124 792 21137
rect -792 20879 -704 20892
rect -792 17905 -779 20879
rect -733 17905 -704 20879
rect -792 17892 -704 17905
rect -304 20879 -200 20892
rect -304 17905 -275 20879
rect -229 17905 -200 20879
rect -304 17892 -200 17905
rect 200 20879 304 20892
rect 200 17905 229 20879
rect 275 17905 304 20879
rect 200 17892 304 17905
rect 704 20879 792 20892
rect 704 17905 733 20879
rect 779 17905 792 20879
rect 704 17892 792 17905
rect -792 17647 -704 17660
rect -792 14673 -779 17647
rect -733 14673 -704 17647
rect -792 14660 -704 14673
rect -304 17647 -200 17660
rect -304 14673 -275 17647
rect -229 14673 -200 17647
rect -304 14660 -200 14673
rect 200 17647 304 17660
rect 200 14673 229 17647
rect 275 14673 304 17647
rect 200 14660 304 14673
rect 704 17647 792 17660
rect 704 14673 733 17647
rect 779 14673 792 17647
rect 704 14660 792 14673
rect -792 14415 -704 14428
rect -792 11441 -779 14415
rect -733 11441 -704 14415
rect -792 11428 -704 11441
rect -304 14415 -200 14428
rect -304 11441 -275 14415
rect -229 11441 -200 14415
rect -304 11428 -200 11441
rect 200 14415 304 14428
rect 200 11441 229 14415
rect 275 11441 304 14415
rect 200 11428 304 11441
rect 704 14415 792 14428
rect 704 11441 733 14415
rect 779 11441 792 14415
rect 704 11428 792 11441
rect -792 11183 -704 11196
rect -792 8209 -779 11183
rect -733 8209 -704 11183
rect -792 8196 -704 8209
rect -304 11183 -200 11196
rect -304 8209 -275 11183
rect -229 8209 -200 11183
rect -304 8196 -200 8209
rect 200 11183 304 11196
rect 200 8209 229 11183
rect 275 8209 304 11183
rect 200 8196 304 8209
rect 704 11183 792 11196
rect 704 8209 733 11183
rect 779 8209 792 11183
rect 704 8196 792 8209
rect -792 7951 -704 7964
rect -792 4977 -779 7951
rect -733 4977 -704 7951
rect -792 4964 -704 4977
rect -304 7951 -200 7964
rect -304 4977 -275 7951
rect -229 4977 -200 7951
rect -304 4964 -200 4977
rect 200 7951 304 7964
rect 200 4977 229 7951
rect 275 4977 304 7951
rect 200 4964 304 4977
rect 704 7951 792 7964
rect 704 4977 733 7951
rect 779 4977 792 7951
rect 704 4964 792 4977
rect -792 4719 -704 4732
rect -792 1745 -779 4719
rect -733 1745 -704 4719
rect -792 1732 -704 1745
rect -304 4719 -200 4732
rect -304 1745 -275 4719
rect -229 1745 -200 4719
rect -304 1732 -200 1745
rect 200 4719 304 4732
rect 200 1745 229 4719
rect 275 1745 304 4719
rect 200 1732 304 1745
rect 704 4719 792 4732
rect 704 1745 733 4719
rect 779 1745 792 4719
rect 704 1732 792 1745
rect -792 1487 -704 1500
rect -792 -1487 -779 1487
rect -733 -1487 -704 1487
rect -792 -1500 -704 -1487
rect -304 1487 -200 1500
rect -304 -1487 -275 1487
rect -229 -1487 -200 1487
rect -304 -1500 -200 -1487
rect 200 1487 304 1500
rect 200 -1487 229 1487
rect 275 -1487 304 1487
rect 200 -1500 304 -1487
rect 704 1487 792 1500
rect 704 -1487 733 1487
rect 779 -1487 792 1487
rect 704 -1500 792 -1487
rect -792 -1745 -704 -1732
rect -792 -4719 -779 -1745
rect -733 -4719 -704 -1745
rect -792 -4732 -704 -4719
rect -304 -1745 -200 -1732
rect -304 -4719 -275 -1745
rect -229 -4719 -200 -1745
rect -304 -4732 -200 -4719
rect 200 -1745 304 -1732
rect 200 -4719 229 -1745
rect 275 -4719 304 -1745
rect 200 -4732 304 -4719
rect 704 -1745 792 -1732
rect 704 -4719 733 -1745
rect 779 -4719 792 -1745
rect 704 -4732 792 -4719
rect -792 -4977 -704 -4964
rect -792 -7951 -779 -4977
rect -733 -7951 -704 -4977
rect -792 -7964 -704 -7951
rect -304 -4977 -200 -4964
rect -304 -7951 -275 -4977
rect -229 -7951 -200 -4977
rect -304 -7964 -200 -7951
rect 200 -4977 304 -4964
rect 200 -7951 229 -4977
rect 275 -7951 304 -4977
rect 200 -7964 304 -7951
rect 704 -4977 792 -4964
rect 704 -7951 733 -4977
rect 779 -7951 792 -4977
rect 704 -7964 792 -7951
rect -792 -8209 -704 -8196
rect -792 -11183 -779 -8209
rect -733 -11183 -704 -8209
rect -792 -11196 -704 -11183
rect -304 -8209 -200 -8196
rect -304 -11183 -275 -8209
rect -229 -11183 -200 -8209
rect -304 -11196 -200 -11183
rect 200 -8209 304 -8196
rect 200 -11183 229 -8209
rect 275 -11183 304 -8209
rect 200 -11196 304 -11183
rect 704 -8209 792 -8196
rect 704 -11183 733 -8209
rect 779 -11183 792 -8209
rect 704 -11196 792 -11183
rect -792 -11441 -704 -11428
rect -792 -14415 -779 -11441
rect -733 -14415 -704 -11441
rect -792 -14428 -704 -14415
rect -304 -11441 -200 -11428
rect -304 -14415 -275 -11441
rect -229 -14415 -200 -11441
rect -304 -14428 -200 -14415
rect 200 -11441 304 -11428
rect 200 -14415 229 -11441
rect 275 -14415 304 -11441
rect 200 -14428 304 -14415
rect 704 -11441 792 -11428
rect 704 -14415 733 -11441
rect 779 -14415 792 -11441
rect 704 -14428 792 -14415
rect -792 -14673 -704 -14660
rect -792 -17647 -779 -14673
rect -733 -17647 -704 -14673
rect -792 -17660 -704 -17647
rect -304 -14673 -200 -14660
rect -304 -17647 -275 -14673
rect -229 -17647 -200 -14673
rect -304 -17660 -200 -17647
rect 200 -14673 304 -14660
rect 200 -17647 229 -14673
rect 275 -17647 304 -14673
rect 200 -17660 304 -17647
rect 704 -14673 792 -14660
rect 704 -17647 733 -14673
rect 779 -17647 792 -14673
rect 704 -17660 792 -17647
rect -792 -17905 -704 -17892
rect -792 -20879 -779 -17905
rect -733 -20879 -704 -17905
rect -792 -20892 -704 -20879
rect -304 -17905 -200 -17892
rect -304 -20879 -275 -17905
rect -229 -20879 -200 -17905
rect -304 -20892 -200 -20879
rect 200 -17905 304 -17892
rect 200 -20879 229 -17905
rect 275 -20879 304 -17905
rect 200 -20892 304 -20879
rect 704 -17905 792 -17892
rect 704 -20879 733 -17905
rect 779 -20879 792 -17905
rect 704 -20892 792 -20879
rect -792 -21137 -704 -21124
rect -792 -24111 -779 -21137
rect -733 -24111 -704 -21137
rect -792 -24124 -704 -24111
rect -304 -21137 -200 -21124
rect -304 -24111 -275 -21137
rect -229 -24111 -200 -21137
rect -304 -24124 -200 -24111
rect 200 -21137 304 -21124
rect 200 -24111 229 -21137
rect 275 -24111 304 -21137
rect 200 -24124 304 -24111
rect 704 -21137 792 -21124
rect 704 -24111 733 -21137
rect 779 -24111 792 -21137
rect 704 -24124 792 -24111
rect -792 -24369 -704 -24356
rect -792 -27343 -779 -24369
rect -733 -27343 -704 -24369
rect -792 -27356 -704 -27343
rect -304 -24369 -200 -24356
rect -304 -27343 -275 -24369
rect -229 -27343 -200 -24369
rect -304 -27356 -200 -27343
rect 200 -24369 304 -24356
rect 200 -27343 229 -24369
rect 275 -27343 304 -24369
rect 200 -27356 304 -27343
rect 704 -24369 792 -24356
rect 704 -27343 733 -24369
rect 779 -27343 792 -24369
rect 704 -27356 792 -27343
rect -792 -27601 -704 -27588
rect -792 -30575 -779 -27601
rect -733 -30575 -704 -27601
rect -792 -30588 -704 -30575
rect -304 -27601 -200 -27588
rect -304 -30575 -275 -27601
rect -229 -30575 -200 -27601
rect -304 -30588 -200 -30575
rect 200 -27601 304 -27588
rect 200 -30575 229 -27601
rect 275 -30575 304 -27601
rect 200 -30588 304 -30575
rect 704 -27601 792 -27588
rect 704 -30575 733 -27601
rect 779 -30575 792 -27601
rect 704 -30588 792 -30575
rect -792 -30833 -704 -30820
rect -792 -33807 -779 -30833
rect -733 -33807 -704 -30833
rect -792 -33820 -704 -33807
rect -304 -30833 -200 -30820
rect -304 -33807 -275 -30833
rect -229 -33807 -200 -30833
rect -304 -33820 -200 -33807
rect 200 -30833 304 -30820
rect 200 -33807 229 -30833
rect 275 -33807 304 -30833
rect 200 -33820 304 -33807
rect 704 -30833 792 -30820
rect 704 -33807 733 -30833
rect 779 -33807 792 -30833
rect 704 -33820 792 -33807
rect -792 -34065 -704 -34052
rect -792 -37039 -779 -34065
rect -733 -37039 -704 -34065
rect -792 -37052 -704 -37039
rect -304 -34065 -200 -34052
rect -304 -37039 -275 -34065
rect -229 -37039 -200 -34065
rect -304 -37052 -200 -37039
rect 200 -34065 304 -34052
rect 200 -37039 229 -34065
rect 275 -37039 304 -34065
rect 200 -37052 304 -37039
rect 704 -34065 792 -34052
rect 704 -37039 733 -34065
rect 779 -37039 792 -34065
rect 704 -37052 792 -37039
rect -792 -37297 -704 -37284
rect -792 -40271 -779 -37297
rect -733 -40271 -704 -37297
rect -792 -40284 -704 -40271
rect -304 -37297 -200 -37284
rect -304 -40271 -275 -37297
rect -229 -40271 -200 -37297
rect -304 -40284 -200 -40271
rect 200 -37297 304 -37284
rect 200 -40271 229 -37297
rect 275 -40271 304 -37297
rect 200 -40284 304 -40271
rect 704 -37297 792 -37284
rect 704 -40271 733 -37297
rect 779 -40271 792 -37297
rect 704 -40284 792 -40271
<< pdiffc >>
rect -779 37297 -733 40271
rect -275 37297 -229 40271
rect 229 37297 275 40271
rect 733 37297 779 40271
rect -779 34065 -733 37039
rect -275 34065 -229 37039
rect 229 34065 275 37039
rect 733 34065 779 37039
rect -779 30833 -733 33807
rect -275 30833 -229 33807
rect 229 30833 275 33807
rect 733 30833 779 33807
rect -779 27601 -733 30575
rect -275 27601 -229 30575
rect 229 27601 275 30575
rect 733 27601 779 30575
rect -779 24369 -733 27343
rect -275 24369 -229 27343
rect 229 24369 275 27343
rect 733 24369 779 27343
rect -779 21137 -733 24111
rect -275 21137 -229 24111
rect 229 21137 275 24111
rect 733 21137 779 24111
rect -779 17905 -733 20879
rect -275 17905 -229 20879
rect 229 17905 275 20879
rect 733 17905 779 20879
rect -779 14673 -733 17647
rect -275 14673 -229 17647
rect 229 14673 275 17647
rect 733 14673 779 17647
rect -779 11441 -733 14415
rect -275 11441 -229 14415
rect 229 11441 275 14415
rect 733 11441 779 14415
rect -779 8209 -733 11183
rect -275 8209 -229 11183
rect 229 8209 275 11183
rect 733 8209 779 11183
rect -779 4977 -733 7951
rect -275 4977 -229 7951
rect 229 4977 275 7951
rect 733 4977 779 7951
rect -779 1745 -733 4719
rect -275 1745 -229 4719
rect 229 1745 275 4719
rect 733 1745 779 4719
rect -779 -1487 -733 1487
rect -275 -1487 -229 1487
rect 229 -1487 275 1487
rect 733 -1487 779 1487
rect -779 -4719 -733 -1745
rect -275 -4719 -229 -1745
rect 229 -4719 275 -1745
rect 733 -4719 779 -1745
rect -779 -7951 -733 -4977
rect -275 -7951 -229 -4977
rect 229 -7951 275 -4977
rect 733 -7951 779 -4977
rect -779 -11183 -733 -8209
rect -275 -11183 -229 -8209
rect 229 -11183 275 -8209
rect 733 -11183 779 -8209
rect -779 -14415 -733 -11441
rect -275 -14415 -229 -11441
rect 229 -14415 275 -11441
rect 733 -14415 779 -11441
rect -779 -17647 -733 -14673
rect -275 -17647 -229 -14673
rect 229 -17647 275 -14673
rect 733 -17647 779 -14673
rect -779 -20879 -733 -17905
rect -275 -20879 -229 -17905
rect 229 -20879 275 -17905
rect 733 -20879 779 -17905
rect -779 -24111 -733 -21137
rect -275 -24111 -229 -21137
rect 229 -24111 275 -21137
rect 733 -24111 779 -21137
rect -779 -27343 -733 -24369
rect -275 -27343 -229 -24369
rect 229 -27343 275 -24369
rect 733 -27343 779 -24369
rect -779 -30575 -733 -27601
rect -275 -30575 -229 -27601
rect 229 -30575 275 -27601
rect 733 -30575 779 -27601
rect -779 -33807 -733 -30833
rect -275 -33807 -229 -30833
rect 229 -33807 275 -30833
rect 733 -33807 779 -30833
rect -779 -37039 -733 -34065
rect -275 -37039 -229 -34065
rect 229 -37039 275 -34065
rect 733 -37039 779 -34065
rect -779 -40271 -733 -37297
rect -275 -40271 -229 -37297
rect 229 -40271 275 -37297
rect 733 -40271 779 -37297
<< nsubdiff >>
rect -930 40398 930 40470
rect -930 40354 -858 40398
rect -930 -40354 -917 40354
rect -871 -40354 -858 40354
rect 858 40354 930 40398
rect -930 -40398 -858 -40354
rect 858 -40354 871 40354
rect 917 -40354 930 40354
rect 858 -40398 930 -40354
rect -930 -40470 930 -40398
<< nsubdiffcont >>
rect -917 -40354 -871 40354
rect 871 -40354 917 40354
<< polysilicon >>
rect -704 40363 -304 40376
rect -704 40317 -691 40363
rect -317 40317 -304 40363
rect -704 40284 -304 40317
rect -200 40363 200 40376
rect -200 40317 -187 40363
rect 187 40317 200 40363
rect -200 40284 200 40317
rect 304 40363 704 40376
rect 304 40317 317 40363
rect 691 40317 704 40363
rect 304 40284 704 40317
rect -704 37251 -304 37284
rect -704 37205 -691 37251
rect -317 37205 -304 37251
rect -704 37192 -304 37205
rect -200 37251 200 37284
rect -200 37205 -187 37251
rect 187 37205 200 37251
rect -200 37192 200 37205
rect 304 37251 704 37284
rect 304 37205 317 37251
rect 691 37205 704 37251
rect 304 37192 704 37205
rect -704 37131 -304 37144
rect -704 37085 -691 37131
rect -317 37085 -304 37131
rect -704 37052 -304 37085
rect -200 37131 200 37144
rect -200 37085 -187 37131
rect 187 37085 200 37131
rect -200 37052 200 37085
rect 304 37131 704 37144
rect 304 37085 317 37131
rect 691 37085 704 37131
rect 304 37052 704 37085
rect -704 34019 -304 34052
rect -704 33973 -691 34019
rect -317 33973 -304 34019
rect -704 33960 -304 33973
rect -200 34019 200 34052
rect -200 33973 -187 34019
rect 187 33973 200 34019
rect -200 33960 200 33973
rect 304 34019 704 34052
rect 304 33973 317 34019
rect 691 33973 704 34019
rect 304 33960 704 33973
rect -704 33899 -304 33912
rect -704 33853 -691 33899
rect -317 33853 -304 33899
rect -704 33820 -304 33853
rect -200 33899 200 33912
rect -200 33853 -187 33899
rect 187 33853 200 33899
rect -200 33820 200 33853
rect 304 33899 704 33912
rect 304 33853 317 33899
rect 691 33853 704 33899
rect 304 33820 704 33853
rect -704 30787 -304 30820
rect -704 30741 -691 30787
rect -317 30741 -304 30787
rect -704 30728 -304 30741
rect -200 30787 200 30820
rect -200 30741 -187 30787
rect 187 30741 200 30787
rect -200 30728 200 30741
rect 304 30787 704 30820
rect 304 30741 317 30787
rect 691 30741 704 30787
rect 304 30728 704 30741
rect -704 30667 -304 30680
rect -704 30621 -691 30667
rect -317 30621 -304 30667
rect -704 30588 -304 30621
rect -200 30667 200 30680
rect -200 30621 -187 30667
rect 187 30621 200 30667
rect -200 30588 200 30621
rect 304 30667 704 30680
rect 304 30621 317 30667
rect 691 30621 704 30667
rect 304 30588 704 30621
rect -704 27555 -304 27588
rect -704 27509 -691 27555
rect -317 27509 -304 27555
rect -704 27496 -304 27509
rect -200 27555 200 27588
rect -200 27509 -187 27555
rect 187 27509 200 27555
rect -200 27496 200 27509
rect 304 27555 704 27588
rect 304 27509 317 27555
rect 691 27509 704 27555
rect 304 27496 704 27509
rect -704 27435 -304 27448
rect -704 27389 -691 27435
rect -317 27389 -304 27435
rect -704 27356 -304 27389
rect -200 27435 200 27448
rect -200 27389 -187 27435
rect 187 27389 200 27435
rect -200 27356 200 27389
rect 304 27435 704 27448
rect 304 27389 317 27435
rect 691 27389 704 27435
rect 304 27356 704 27389
rect -704 24323 -304 24356
rect -704 24277 -691 24323
rect -317 24277 -304 24323
rect -704 24264 -304 24277
rect -200 24323 200 24356
rect -200 24277 -187 24323
rect 187 24277 200 24323
rect -200 24264 200 24277
rect 304 24323 704 24356
rect 304 24277 317 24323
rect 691 24277 704 24323
rect 304 24264 704 24277
rect -704 24203 -304 24216
rect -704 24157 -691 24203
rect -317 24157 -304 24203
rect -704 24124 -304 24157
rect -200 24203 200 24216
rect -200 24157 -187 24203
rect 187 24157 200 24203
rect -200 24124 200 24157
rect 304 24203 704 24216
rect 304 24157 317 24203
rect 691 24157 704 24203
rect 304 24124 704 24157
rect -704 21091 -304 21124
rect -704 21045 -691 21091
rect -317 21045 -304 21091
rect -704 21032 -304 21045
rect -200 21091 200 21124
rect -200 21045 -187 21091
rect 187 21045 200 21091
rect -200 21032 200 21045
rect 304 21091 704 21124
rect 304 21045 317 21091
rect 691 21045 704 21091
rect 304 21032 704 21045
rect -704 20971 -304 20984
rect -704 20925 -691 20971
rect -317 20925 -304 20971
rect -704 20892 -304 20925
rect -200 20971 200 20984
rect -200 20925 -187 20971
rect 187 20925 200 20971
rect -200 20892 200 20925
rect 304 20971 704 20984
rect 304 20925 317 20971
rect 691 20925 704 20971
rect 304 20892 704 20925
rect -704 17859 -304 17892
rect -704 17813 -691 17859
rect -317 17813 -304 17859
rect -704 17800 -304 17813
rect -200 17859 200 17892
rect -200 17813 -187 17859
rect 187 17813 200 17859
rect -200 17800 200 17813
rect 304 17859 704 17892
rect 304 17813 317 17859
rect 691 17813 704 17859
rect 304 17800 704 17813
rect -704 17739 -304 17752
rect -704 17693 -691 17739
rect -317 17693 -304 17739
rect -704 17660 -304 17693
rect -200 17739 200 17752
rect -200 17693 -187 17739
rect 187 17693 200 17739
rect -200 17660 200 17693
rect 304 17739 704 17752
rect 304 17693 317 17739
rect 691 17693 704 17739
rect 304 17660 704 17693
rect -704 14627 -304 14660
rect -704 14581 -691 14627
rect -317 14581 -304 14627
rect -704 14568 -304 14581
rect -200 14627 200 14660
rect -200 14581 -187 14627
rect 187 14581 200 14627
rect -200 14568 200 14581
rect 304 14627 704 14660
rect 304 14581 317 14627
rect 691 14581 704 14627
rect 304 14568 704 14581
rect -704 14507 -304 14520
rect -704 14461 -691 14507
rect -317 14461 -304 14507
rect -704 14428 -304 14461
rect -200 14507 200 14520
rect -200 14461 -187 14507
rect 187 14461 200 14507
rect -200 14428 200 14461
rect 304 14507 704 14520
rect 304 14461 317 14507
rect 691 14461 704 14507
rect 304 14428 704 14461
rect -704 11395 -304 11428
rect -704 11349 -691 11395
rect -317 11349 -304 11395
rect -704 11336 -304 11349
rect -200 11395 200 11428
rect -200 11349 -187 11395
rect 187 11349 200 11395
rect -200 11336 200 11349
rect 304 11395 704 11428
rect 304 11349 317 11395
rect 691 11349 704 11395
rect 304 11336 704 11349
rect -704 11275 -304 11288
rect -704 11229 -691 11275
rect -317 11229 -304 11275
rect -704 11196 -304 11229
rect -200 11275 200 11288
rect -200 11229 -187 11275
rect 187 11229 200 11275
rect -200 11196 200 11229
rect 304 11275 704 11288
rect 304 11229 317 11275
rect 691 11229 704 11275
rect 304 11196 704 11229
rect -704 8163 -304 8196
rect -704 8117 -691 8163
rect -317 8117 -304 8163
rect -704 8104 -304 8117
rect -200 8163 200 8196
rect -200 8117 -187 8163
rect 187 8117 200 8163
rect -200 8104 200 8117
rect 304 8163 704 8196
rect 304 8117 317 8163
rect 691 8117 704 8163
rect 304 8104 704 8117
rect -704 8043 -304 8056
rect -704 7997 -691 8043
rect -317 7997 -304 8043
rect -704 7964 -304 7997
rect -200 8043 200 8056
rect -200 7997 -187 8043
rect 187 7997 200 8043
rect -200 7964 200 7997
rect 304 8043 704 8056
rect 304 7997 317 8043
rect 691 7997 704 8043
rect 304 7964 704 7997
rect -704 4931 -304 4964
rect -704 4885 -691 4931
rect -317 4885 -304 4931
rect -704 4872 -304 4885
rect -200 4931 200 4964
rect -200 4885 -187 4931
rect 187 4885 200 4931
rect -200 4872 200 4885
rect 304 4931 704 4964
rect 304 4885 317 4931
rect 691 4885 704 4931
rect 304 4872 704 4885
rect -704 4811 -304 4824
rect -704 4765 -691 4811
rect -317 4765 -304 4811
rect -704 4732 -304 4765
rect -200 4811 200 4824
rect -200 4765 -187 4811
rect 187 4765 200 4811
rect -200 4732 200 4765
rect 304 4811 704 4824
rect 304 4765 317 4811
rect 691 4765 704 4811
rect 304 4732 704 4765
rect -704 1699 -304 1732
rect -704 1653 -691 1699
rect -317 1653 -304 1699
rect -704 1640 -304 1653
rect -200 1699 200 1732
rect -200 1653 -187 1699
rect 187 1653 200 1699
rect -200 1640 200 1653
rect 304 1699 704 1732
rect 304 1653 317 1699
rect 691 1653 704 1699
rect 304 1640 704 1653
rect -704 1579 -304 1592
rect -704 1533 -691 1579
rect -317 1533 -304 1579
rect -704 1500 -304 1533
rect -200 1579 200 1592
rect -200 1533 -187 1579
rect 187 1533 200 1579
rect -200 1500 200 1533
rect 304 1579 704 1592
rect 304 1533 317 1579
rect 691 1533 704 1579
rect 304 1500 704 1533
rect -704 -1533 -304 -1500
rect -704 -1579 -691 -1533
rect -317 -1579 -304 -1533
rect -704 -1592 -304 -1579
rect -200 -1533 200 -1500
rect -200 -1579 -187 -1533
rect 187 -1579 200 -1533
rect -200 -1592 200 -1579
rect 304 -1533 704 -1500
rect 304 -1579 317 -1533
rect 691 -1579 704 -1533
rect 304 -1592 704 -1579
rect -704 -1653 -304 -1640
rect -704 -1699 -691 -1653
rect -317 -1699 -304 -1653
rect -704 -1732 -304 -1699
rect -200 -1653 200 -1640
rect -200 -1699 -187 -1653
rect 187 -1699 200 -1653
rect -200 -1732 200 -1699
rect 304 -1653 704 -1640
rect 304 -1699 317 -1653
rect 691 -1699 704 -1653
rect 304 -1732 704 -1699
rect -704 -4765 -304 -4732
rect -704 -4811 -691 -4765
rect -317 -4811 -304 -4765
rect -704 -4824 -304 -4811
rect -200 -4765 200 -4732
rect -200 -4811 -187 -4765
rect 187 -4811 200 -4765
rect -200 -4824 200 -4811
rect 304 -4765 704 -4732
rect 304 -4811 317 -4765
rect 691 -4811 704 -4765
rect 304 -4824 704 -4811
rect -704 -4885 -304 -4872
rect -704 -4931 -691 -4885
rect -317 -4931 -304 -4885
rect -704 -4964 -304 -4931
rect -200 -4885 200 -4872
rect -200 -4931 -187 -4885
rect 187 -4931 200 -4885
rect -200 -4964 200 -4931
rect 304 -4885 704 -4872
rect 304 -4931 317 -4885
rect 691 -4931 704 -4885
rect 304 -4964 704 -4931
rect -704 -7997 -304 -7964
rect -704 -8043 -691 -7997
rect -317 -8043 -304 -7997
rect -704 -8056 -304 -8043
rect -200 -7997 200 -7964
rect -200 -8043 -187 -7997
rect 187 -8043 200 -7997
rect -200 -8056 200 -8043
rect 304 -7997 704 -7964
rect 304 -8043 317 -7997
rect 691 -8043 704 -7997
rect 304 -8056 704 -8043
rect -704 -8117 -304 -8104
rect -704 -8163 -691 -8117
rect -317 -8163 -304 -8117
rect -704 -8196 -304 -8163
rect -200 -8117 200 -8104
rect -200 -8163 -187 -8117
rect 187 -8163 200 -8117
rect -200 -8196 200 -8163
rect 304 -8117 704 -8104
rect 304 -8163 317 -8117
rect 691 -8163 704 -8117
rect 304 -8196 704 -8163
rect -704 -11229 -304 -11196
rect -704 -11275 -691 -11229
rect -317 -11275 -304 -11229
rect -704 -11288 -304 -11275
rect -200 -11229 200 -11196
rect -200 -11275 -187 -11229
rect 187 -11275 200 -11229
rect -200 -11288 200 -11275
rect 304 -11229 704 -11196
rect 304 -11275 317 -11229
rect 691 -11275 704 -11229
rect 304 -11288 704 -11275
rect -704 -11349 -304 -11336
rect -704 -11395 -691 -11349
rect -317 -11395 -304 -11349
rect -704 -11428 -304 -11395
rect -200 -11349 200 -11336
rect -200 -11395 -187 -11349
rect 187 -11395 200 -11349
rect -200 -11428 200 -11395
rect 304 -11349 704 -11336
rect 304 -11395 317 -11349
rect 691 -11395 704 -11349
rect 304 -11428 704 -11395
rect -704 -14461 -304 -14428
rect -704 -14507 -691 -14461
rect -317 -14507 -304 -14461
rect -704 -14520 -304 -14507
rect -200 -14461 200 -14428
rect -200 -14507 -187 -14461
rect 187 -14507 200 -14461
rect -200 -14520 200 -14507
rect 304 -14461 704 -14428
rect 304 -14507 317 -14461
rect 691 -14507 704 -14461
rect 304 -14520 704 -14507
rect -704 -14581 -304 -14568
rect -704 -14627 -691 -14581
rect -317 -14627 -304 -14581
rect -704 -14660 -304 -14627
rect -200 -14581 200 -14568
rect -200 -14627 -187 -14581
rect 187 -14627 200 -14581
rect -200 -14660 200 -14627
rect 304 -14581 704 -14568
rect 304 -14627 317 -14581
rect 691 -14627 704 -14581
rect 304 -14660 704 -14627
rect -704 -17693 -304 -17660
rect -704 -17739 -691 -17693
rect -317 -17739 -304 -17693
rect -704 -17752 -304 -17739
rect -200 -17693 200 -17660
rect -200 -17739 -187 -17693
rect 187 -17739 200 -17693
rect -200 -17752 200 -17739
rect 304 -17693 704 -17660
rect 304 -17739 317 -17693
rect 691 -17739 704 -17693
rect 304 -17752 704 -17739
rect -704 -17813 -304 -17800
rect -704 -17859 -691 -17813
rect -317 -17859 -304 -17813
rect -704 -17892 -304 -17859
rect -200 -17813 200 -17800
rect -200 -17859 -187 -17813
rect 187 -17859 200 -17813
rect -200 -17892 200 -17859
rect 304 -17813 704 -17800
rect 304 -17859 317 -17813
rect 691 -17859 704 -17813
rect 304 -17892 704 -17859
rect -704 -20925 -304 -20892
rect -704 -20971 -691 -20925
rect -317 -20971 -304 -20925
rect -704 -20984 -304 -20971
rect -200 -20925 200 -20892
rect -200 -20971 -187 -20925
rect 187 -20971 200 -20925
rect -200 -20984 200 -20971
rect 304 -20925 704 -20892
rect 304 -20971 317 -20925
rect 691 -20971 704 -20925
rect 304 -20984 704 -20971
rect -704 -21045 -304 -21032
rect -704 -21091 -691 -21045
rect -317 -21091 -304 -21045
rect -704 -21124 -304 -21091
rect -200 -21045 200 -21032
rect -200 -21091 -187 -21045
rect 187 -21091 200 -21045
rect -200 -21124 200 -21091
rect 304 -21045 704 -21032
rect 304 -21091 317 -21045
rect 691 -21091 704 -21045
rect 304 -21124 704 -21091
rect -704 -24157 -304 -24124
rect -704 -24203 -691 -24157
rect -317 -24203 -304 -24157
rect -704 -24216 -304 -24203
rect -200 -24157 200 -24124
rect -200 -24203 -187 -24157
rect 187 -24203 200 -24157
rect -200 -24216 200 -24203
rect 304 -24157 704 -24124
rect 304 -24203 317 -24157
rect 691 -24203 704 -24157
rect 304 -24216 704 -24203
rect -704 -24277 -304 -24264
rect -704 -24323 -691 -24277
rect -317 -24323 -304 -24277
rect -704 -24356 -304 -24323
rect -200 -24277 200 -24264
rect -200 -24323 -187 -24277
rect 187 -24323 200 -24277
rect -200 -24356 200 -24323
rect 304 -24277 704 -24264
rect 304 -24323 317 -24277
rect 691 -24323 704 -24277
rect 304 -24356 704 -24323
rect -704 -27389 -304 -27356
rect -704 -27435 -691 -27389
rect -317 -27435 -304 -27389
rect -704 -27448 -304 -27435
rect -200 -27389 200 -27356
rect -200 -27435 -187 -27389
rect 187 -27435 200 -27389
rect -200 -27448 200 -27435
rect 304 -27389 704 -27356
rect 304 -27435 317 -27389
rect 691 -27435 704 -27389
rect 304 -27448 704 -27435
rect -704 -27509 -304 -27496
rect -704 -27555 -691 -27509
rect -317 -27555 -304 -27509
rect -704 -27588 -304 -27555
rect -200 -27509 200 -27496
rect -200 -27555 -187 -27509
rect 187 -27555 200 -27509
rect -200 -27588 200 -27555
rect 304 -27509 704 -27496
rect 304 -27555 317 -27509
rect 691 -27555 704 -27509
rect 304 -27588 704 -27555
rect -704 -30621 -304 -30588
rect -704 -30667 -691 -30621
rect -317 -30667 -304 -30621
rect -704 -30680 -304 -30667
rect -200 -30621 200 -30588
rect -200 -30667 -187 -30621
rect 187 -30667 200 -30621
rect -200 -30680 200 -30667
rect 304 -30621 704 -30588
rect 304 -30667 317 -30621
rect 691 -30667 704 -30621
rect 304 -30680 704 -30667
rect -704 -30741 -304 -30728
rect -704 -30787 -691 -30741
rect -317 -30787 -304 -30741
rect -704 -30820 -304 -30787
rect -200 -30741 200 -30728
rect -200 -30787 -187 -30741
rect 187 -30787 200 -30741
rect -200 -30820 200 -30787
rect 304 -30741 704 -30728
rect 304 -30787 317 -30741
rect 691 -30787 704 -30741
rect 304 -30820 704 -30787
rect -704 -33853 -304 -33820
rect -704 -33899 -691 -33853
rect -317 -33899 -304 -33853
rect -704 -33912 -304 -33899
rect -200 -33853 200 -33820
rect -200 -33899 -187 -33853
rect 187 -33899 200 -33853
rect -200 -33912 200 -33899
rect 304 -33853 704 -33820
rect 304 -33899 317 -33853
rect 691 -33899 704 -33853
rect 304 -33912 704 -33899
rect -704 -33973 -304 -33960
rect -704 -34019 -691 -33973
rect -317 -34019 -304 -33973
rect -704 -34052 -304 -34019
rect -200 -33973 200 -33960
rect -200 -34019 -187 -33973
rect 187 -34019 200 -33973
rect -200 -34052 200 -34019
rect 304 -33973 704 -33960
rect 304 -34019 317 -33973
rect 691 -34019 704 -33973
rect 304 -34052 704 -34019
rect -704 -37085 -304 -37052
rect -704 -37131 -691 -37085
rect -317 -37131 -304 -37085
rect -704 -37144 -304 -37131
rect -200 -37085 200 -37052
rect -200 -37131 -187 -37085
rect 187 -37131 200 -37085
rect -200 -37144 200 -37131
rect 304 -37085 704 -37052
rect 304 -37131 317 -37085
rect 691 -37131 704 -37085
rect 304 -37144 704 -37131
rect -704 -37205 -304 -37192
rect -704 -37251 -691 -37205
rect -317 -37251 -304 -37205
rect -704 -37284 -304 -37251
rect -200 -37205 200 -37192
rect -200 -37251 -187 -37205
rect 187 -37251 200 -37205
rect -200 -37284 200 -37251
rect 304 -37205 704 -37192
rect 304 -37251 317 -37205
rect 691 -37251 704 -37205
rect 304 -37284 704 -37251
rect -704 -40317 -304 -40284
rect -704 -40363 -691 -40317
rect -317 -40363 -304 -40317
rect -704 -40376 -304 -40363
rect -200 -40317 200 -40284
rect -200 -40363 -187 -40317
rect 187 -40363 200 -40317
rect -200 -40376 200 -40363
rect 304 -40317 704 -40284
rect 304 -40363 317 -40317
rect 691 -40363 704 -40317
rect 304 -40376 704 -40363
<< polycontact >>
rect -691 40317 -317 40363
rect -187 40317 187 40363
rect 317 40317 691 40363
rect -691 37205 -317 37251
rect -187 37205 187 37251
rect 317 37205 691 37251
rect -691 37085 -317 37131
rect -187 37085 187 37131
rect 317 37085 691 37131
rect -691 33973 -317 34019
rect -187 33973 187 34019
rect 317 33973 691 34019
rect -691 33853 -317 33899
rect -187 33853 187 33899
rect 317 33853 691 33899
rect -691 30741 -317 30787
rect -187 30741 187 30787
rect 317 30741 691 30787
rect -691 30621 -317 30667
rect -187 30621 187 30667
rect 317 30621 691 30667
rect -691 27509 -317 27555
rect -187 27509 187 27555
rect 317 27509 691 27555
rect -691 27389 -317 27435
rect -187 27389 187 27435
rect 317 27389 691 27435
rect -691 24277 -317 24323
rect -187 24277 187 24323
rect 317 24277 691 24323
rect -691 24157 -317 24203
rect -187 24157 187 24203
rect 317 24157 691 24203
rect -691 21045 -317 21091
rect -187 21045 187 21091
rect 317 21045 691 21091
rect -691 20925 -317 20971
rect -187 20925 187 20971
rect 317 20925 691 20971
rect -691 17813 -317 17859
rect -187 17813 187 17859
rect 317 17813 691 17859
rect -691 17693 -317 17739
rect -187 17693 187 17739
rect 317 17693 691 17739
rect -691 14581 -317 14627
rect -187 14581 187 14627
rect 317 14581 691 14627
rect -691 14461 -317 14507
rect -187 14461 187 14507
rect 317 14461 691 14507
rect -691 11349 -317 11395
rect -187 11349 187 11395
rect 317 11349 691 11395
rect -691 11229 -317 11275
rect -187 11229 187 11275
rect 317 11229 691 11275
rect -691 8117 -317 8163
rect -187 8117 187 8163
rect 317 8117 691 8163
rect -691 7997 -317 8043
rect -187 7997 187 8043
rect 317 7997 691 8043
rect -691 4885 -317 4931
rect -187 4885 187 4931
rect 317 4885 691 4931
rect -691 4765 -317 4811
rect -187 4765 187 4811
rect 317 4765 691 4811
rect -691 1653 -317 1699
rect -187 1653 187 1699
rect 317 1653 691 1699
rect -691 1533 -317 1579
rect -187 1533 187 1579
rect 317 1533 691 1579
rect -691 -1579 -317 -1533
rect -187 -1579 187 -1533
rect 317 -1579 691 -1533
rect -691 -1699 -317 -1653
rect -187 -1699 187 -1653
rect 317 -1699 691 -1653
rect -691 -4811 -317 -4765
rect -187 -4811 187 -4765
rect 317 -4811 691 -4765
rect -691 -4931 -317 -4885
rect -187 -4931 187 -4885
rect 317 -4931 691 -4885
rect -691 -8043 -317 -7997
rect -187 -8043 187 -7997
rect 317 -8043 691 -7997
rect -691 -8163 -317 -8117
rect -187 -8163 187 -8117
rect 317 -8163 691 -8117
rect -691 -11275 -317 -11229
rect -187 -11275 187 -11229
rect 317 -11275 691 -11229
rect -691 -11395 -317 -11349
rect -187 -11395 187 -11349
rect 317 -11395 691 -11349
rect -691 -14507 -317 -14461
rect -187 -14507 187 -14461
rect 317 -14507 691 -14461
rect -691 -14627 -317 -14581
rect -187 -14627 187 -14581
rect 317 -14627 691 -14581
rect -691 -17739 -317 -17693
rect -187 -17739 187 -17693
rect 317 -17739 691 -17693
rect -691 -17859 -317 -17813
rect -187 -17859 187 -17813
rect 317 -17859 691 -17813
rect -691 -20971 -317 -20925
rect -187 -20971 187 -20925
rect 317 -20971 691 -20925
rect -691 -21091 -317 -21045
rect -187 -21091 187 -21045
rect 317 -21091 691 -21045
rect -691 -24203 -317 -24157
rect -187 -24203 187 -24157
rect 317 -24203 691 -24157
rect -691 -24323 -317 -24277
rect -187 -24323 187 -24277
rect 317 -24323 691 -24277
rect -691 -27435 -317 -27389
rect -187 -27435 187 -27389
rect 317 -27435 691 -27389
rect -691 -27555 -317 -27509
rect -187 -27555 187 -27509
rect 317 -27555 691 -27509
rect -691 -30667 -317 -30621
rect -187 -30667 187 -30621
rect 317 -30667 691 -30621
rect -691 -30787 -317 -30741
rect -187 -30787 187 -30741
rect 317 -30787 691 -30741
rect -691 -33899 -317 -33853
rect -187 -33899 187 -33853
rect 317 -33899 691 -33853
rect -691 -34019 -317 -33973
rect -187 -34019 187 -33973
rect 317 -34019 691 -33973
rect -691 -37131 -317 -37085
rect -187 -37131 187 -37085
rect 317 -37131 691 -37085
rect -691 -37251 -317 -37205
rect -187 -37251 187 -37205
rect 317 -37251 691 -37205
rect -691 -40363 -317 -40317
rect -187 -40363 187 -40317
rect 317 -40363 691 -40317
<< metal1 >>
rect -917 40411 917 40457
rect -917 40354 -871 40411
rect -702 40317 -691 40363
rect -317 40317 -306 40363
rect -198 40317 -187 40363
rect 187 40317 198 40363
rect 306 40317 317 40363
rect 691 40317 702 40363
rect 871 40354 917 40411
rect -779 40271 -733 40282
rect -779 37286 -733 37297
rect -275 40271 -229 40282
rect -275 37286 -229 37297
rect 229 40271 275 40282
rect 229 37286 275 37297
rect 733 40271 779 40282
rect 733 37286 779 37297
rect -702 37205 -691 37251
rect -317 37205 -306 37251
rect -198 37205 -187 37251
rect 187 37205 198 37251
rect 306 37205 317 37251
rect 691 37205 702 37251
rect -702 37085 -691 37131
rect -317 37085 -306 37131
rect -198 37085 -187 37131
rect 187 37085 198 37131
rect 306 37085 317 37131
rect 691 37085 702 37131
rect -779 37039 -733 37050
rect -779 34054 -733 34065
rect -275 37039 -229 37050
rect -275 34054 -229 34065
rect 229 37039 275 37050
rect 229 34054 275 34065
rect 733 37039 779 37050
rect 733 34054 779 34065
rect -702 33973 -691 34019
rect -317 33973 -306 34019
rect -198 33973 -187 34019
rect 187 33973 198 34019
rect 306 33973 317 34019
rect 691 33973 702 34019
rect -702 33853 -691 33899
rect -317 33853 -306 33899
rect -198 33853 -187 33899
rect 187 33853 198 33899
rect 306 33853 317 33899
rect 691 33853 702 33899
rect -779 33807 -733 33818
rect -779 30822 -733 30833
rect -275 33807 -229 33818
rect -275 30822 -229 30833
rect 229 33807 275 33818
rect 229 30822 275 30833
rect 733 33807 779 33818
rect 733 30822 779 30833
rect -702 30741 -691 30787
rect -317 30741 -306 30787
rect -198 30741 -187 30787
rect 187 30741 198 30787
rect 306 30741 317 30787
rect 691 30741 702 30787
rect -702 30621 -691 30667
rect -317 30621 -306 30667
rect -198 30621 -187 30667
rect 187 30621 198 30667
rect 306 30621 317 30667
rect 691 30621 702 30667
rect -779 30575 -733 30586
rect -779 27590 -733 27601
rect -275 30575 -229 30586
rect -275 27590 -229 27601
rect 229 30575 275 30586
rect 229 27590 275 27601
rect 733 30575 779 30586
rect 733 27590 779 27601
rect -702 27509 -691 27555
rect -317 27509 -306 27555
rect -198 27509 -187 27555
rect 187 27509 198 27555
rect 306 27509 317 27555
rect 691 27509 702 27555
rect -702 27389 -691 27435
rect -317 27389 -306 27435
rect -198 27389 -187 27435
rect 187 27389 198 27435
rect 306 27389 317 27435
rect 691 27389 702 27435
rect -779 27343 -733 27354
rect -779 24358 -733 24369
rect -275 27343 -229 27354
rect -275 24358 -229 24369
rect 229 27343 275 27354
rect 229 24358 275 24369
rect 733 27343 779 27354
rect 733 24358 779 24369
rect -702 24277 -691 24323
rect -317 24277 -306 24323
rect -198 24277 -187 24323
rect 187 24277 198 24323
rect 306 24277 317 24323
rect 691 24277 702 24323
rect -702 24157 -691 24203
rect -317 24157 -306 24203
rect -198 24157 -187 24203
rect 187 24157 198 24203
rect 306 24157 317 24203
rect 691 24157 702 24203
rect -779 24111 -733 24122
rect -779 21126 -733 21137
rect -275 24111 -229 24122
rect -275 21126 -229 21137
rect 229 24111 275 24122
rect 229 21126 275 21137
rect 733 24111 779 24122
rect 733 21126 779 21137
rect -702 21045 -691 21091
rect -317 21045 -306 21091
rect -198 21045 -187 21091
rect 187 21045 198 21091
rect 306 21045 317 21091
rect 691 21045 702 21091
rect -702 20925 -691 20971
rect -317 20925 -306 20971
rect -198 20925 -187 20971
rect 187 20925 198 20971
rect 306 20925 317 20971
rect 691 20925 702 20971
rect -779 20879 -733 20890
rect -779 17894 -733 17905
rect -275 20879 -229 20890
rect -275 17894 -229 17905
rect 229 20879 275 20890
rect 229 17894 275 17905
rect 733 20879 779 20890
rect 733 17894 779 17905
rect -702 17813 -691 17859
rect -317 17813 -306 17859
rect -198 17813 -187 17859
rect 187 17813 198 17859
rect 306 17813 317 17859
rect 691 17813 702 17859
rect -702 17693 -691 17739
rect -317 17693 -306 17739
rect -198 17693 -187 17739
rect 187 17693 198 17739
rect 306 17693 317 17739
rect 691 17693 702 17739
rect -779 17647 -733 17658
rect -779 14662 -733 14673
rect -275 17647 -229 17658
rect -275 14662 -229 14673
rect 229 17647 275 17658
rect 229 14662 275 14673
rect 733 17647 779 17658
rect 733 14662 779 14673
rect -702 14581 -691 14627
rect -317 14581 -306 14627
rect -198 14581 -187 14627
rect 187 14581 198 14627
rect 306 14581 317 14627
rect 691 14581 702 14627
rect -702 14461 -691 14507
rect -317 14461 -306 14507
rect -198 14461 -187 14507
rect 187 14461 198 14507
rect 306 14461 317 14507
rect 691 14461 702 14507
rect -779 14415 -733 14426
rect -779 11430 -733 11441
rect -275 14415 -229 14426
rect -275 11430 -229 11441
rect 229 14415 275 14426
rect 229 11430 275 11441
rect 733 14415 779 14426
rect 733 11430 779 11441
rect -702 11349 -691 11395
rect -317 11349 -306 11395
rect -198 11349 -187 11395
rect 187 11349 198 11395
rect 306 11349 317 11395
rect 691 11349 702 11395
rect -702 11229 -691 11275
rect -317 11229 -306 11275
rect -198 11229 -187 11275
rect 187 11229 198 11275
rect 306 11229 317 11275
rect 691 11229 702 11275
rect -779 11183 -733 11194
rect -779 8198 -733 8209
rect -275 11183 -229 11194
rect -275 8198 -229 8209
rect 229 11183 275 11194
rect 229 8198 275 8209
rect 733 11183 779 11194
rect 733 8198 779 8209
rect -702 8117 -691 8163
rect -317 8117 -306 8163
rect -198 8117 -187 8163
rect 187 8117 198 8163
rect 306 8117 317 8163
rect 691 8117 702 8163
rect -702 7997 -691 8043
rect -317 7997 -306 8043
rect -198 7997 -187 8043
rect 187 7997 198 8043
rect 306 7997 317 8043
rect 691 7997 702 8043
rect -779 7951 -733 7962
rect -779 4966 -733 4977
rect -275 7951 -229 7962
rect -275 4966 -229 4977
rect 229 7951 275 7962
rect 229 4966 275 4977
rect 733 7951 779 7962
rect 733 4966 779 4977
rect -702 4885 -691 4931
rect -317 4885 -306 4931
rect -198 4885 -187 4931
rect 187 4885 198 4931
rect 306 4885 317 4931
rect 691 4885 702 4931
rect -702 4765 -691 4811
rect -317 4765 -306 4811
rect -198 4765 -187 4811
rect 187 4765 198 4811
rect 306 4765 317 4811
rect 691 4765 702 4811
rect -779 4719 -733 4730
rect -779 1734 -733 1745
rect -275 4719 -229 4730
rect -275 1734 -229 1745
rect 229 4719 275 4730
rect 229 1734 275 1745
rect 733 4719 779 4730
rect 733 1734 779 1745
rect -702 1653 -691 1699
rect -317 1653 -306 1699
rect -198 1653 -187 1699
rect 187 1653 198 1699
rect 306 1653 317 1699
rect 691 1653 702 1699
rect -702 1533 -691 1579
rect -317 1533 -306 1579
rect -198 1533 -187 1579
rect 187 1533 198 1579
rect 306 1533 317 1579
rect 691 1533 702 1579
rect -779 1487 -733 1498
rect -779 -1498 -733 -1487
rect -275 1487 -229 1498
rect -275 -1498 -229 -1487
rect 229 1487 275 1498
rect 229 -1498 275 -1487
rect 733 1487 779 1498
rect 733 -1498 779 -1487
rect -702 -1579 -691 -1533
rect -317 -1579 -306 -1533
rect -198 -1579 -187 -1533
rect 187 -1579 198 -1533
rect 306 -1579 317 -1533
rect 691 -1579 702 -1533
rect -702 -1699 -691 -1653
rect -317 -1699 -306 -1653
rect -198 -1699 -187 -1653
rect 187 -1699 198 -1653
rect 306 -1699 317 -1653
rect 691 -1699 702 -1653
rect -779 -1745 -733 -1734
rect -779 -4730 -733 -4719
rect -275 -1745 -229 -1734
rect -275 -4730 -229 -4719
rect 229 -1745 275 -1734
rect 229 -4730 275 -4719
rect 733 -1745 779 -1734
rect 733 -4730 779 -4719
rect -702 -4811 -691 -4765
rect -317 -4811 -306 -4765
rect -198 -4811 -187 -4765
rect 187 -4811 198 -4765
rect 306 -4811 317 -4765
rect 691 -4811 702 -4765
rect -702 -4931 -691 -4885
rect -317 -4931 -306 -4885
rect -198 -4931 -187 -4885
rect 187 -4931 198 -4885
rect 306 -4931 317 -4885
rect 691 -4931 702 -4885
rect -779 -4977 -733 -4966
rect -779 -7962 -733 -7951
rect -275 -4977 -229 -4966
rect -275 -7962 -229 -7951
rect 229 -4977 275 -4966
rect 229 -7962 275 -7951
rect 733 -4977 779 -4966
rect 733 -7962 779 -7951
rect -702 -8043 -691 -7997
rect -317 -8043 -306 -7997
rect -198 -8043 -187 -7997
rect 187 -8043 198 -7997
rect 306 -8043 317 -7997
rect 691 -8043 702 -7997
rect -702 -8163 -691 -8117
rect -317 -8163 -306 -8117
rect -198 -8163 -187 -8117
rect 187 -8163 198 -8117
rect 306 -8163 317 -8117
rect 691 -8163 702 -8117
rect -779 -8209 -733 -8198
rect -779 -11194 -733 -11183
rect -275 -8209 -229 -8198
rect -275 -11194 -229 -11183
rect 229 -8209 275 -8198
rect 229 -11194 275 -11183
rect 733 -8209 779 -8198
rect 733 -11194 779 -11183
rect -702 -11275 -691 -11229
rect -317 -11275 -306 -11229
rect -198 -11275 -187 -11229
rect 187 -11275 198 -11229
rect 306 -11275 317 -11229
rect 691 -11275 702 -11229
rect -702 -11395 -691 -11349
rect -317 -11395 -306 -11349
rect -198 -11395 -187 -11349
rect 187 -11395 198 -11349
rect 306 -11395 317 -11349
rect 691 -11395 702 -11349
rect -779 -11441 -733 -11430
rect -779 -14426 -733 -14415
rect -275 -11441 -229 -11430
rect -275 -14426 -229 -14415
rect 229 -11441 275 -11430
rect 229 -14426 275 -14415
rect 733 -11441 779 -11430
rect 733 -14426 779 -14415
rect -702 -14507 -691 -14461
rect -317 -14507 -306 -14461
rect -198 -14507 -187 -14461
rect 187 -14507 198 -14461
rect 306 -14507 317 -14461
rect 691 -14507 702 -14461
rect -702 -14627 -691 -14581
rect -317 -14627 -306 -14581
rect -198 -14627 -187 -14581
rect 187 -14627 198 -14581
rect 306 -14627 317 -14581
rect 691 -14627 702 -14581
rect -779 -14673 -733 -14662
rect -779 -17658 -733 -17647
rect -275 -14673 -229 -14662
rect -275 -17658 -229 -17647
rect 229 -14673 275 -14662
rect 229 -17658 275 -17647
rect 733 -14673 779 -14662
rect 733 -17658 779 -17647
rect -702 -17739 -691 -17693
rect -317 -17739 -306 -17693
rect -198 -17739 -187 -17693
rect 187 -17739 198 -17693
rect 306 -17739 317 -17693
rect 691 -17739 702 -17693
rect -702 -17859 -691 -17813
rect -317 -17859 -306 -17813
rect -198 -17859 -187 -17813
rect 187 -17859 198 -17813
rect 306 -17859 317 -17813
rect 691 -17859 702 -17813
rect -779 -17905 -733 -17894
rect -779 -20890 -733 -20879
rect -275 -17905 -229 -17894
rect -275 -20890 -229 -20879
rect 229 -17905 275 -17894
rect 229 -20890 275 -20879
rect 733 -17905 779 -17894
rect 733 -20890 779 -20879
rect -702 -20971 -691 -20925
rect -317 -20971 -306 -20925
rect -198 -20971 -187 -20925
rect 187 -20971 198 -20925
rect 306 -20971 317 -20925
rect 691 -20971 702 -20925
rect -702 -21091 -691 -21045
rect -317 -21091 -306 -21045
rect -198 -21091 -187 -21045
rect 187 -21091 198 -21045
rect 306 -21091 317 -21045
rect 691 -21091 702 -21045
rect -779 -21137 -733 -21126
rect -779 -24122 -733 -24111
rect -275 -21137 -229 -21126
rect -275 -24122 -229 -24111
rect 229 -21137 275 -21126
rect 229 -24122 275 -24111
rect 733 -21137 779 -21126
rect 733 -24122 779 -24111
rect -702 -24203 -691 -24157
rect -317 -24203 -306 -24157
rect -198 -24203 -187 -24157
rect 187 -24203 198 -24157
rect 306 -24203 317 -24157
rect 691 -24203 702 -24157
rect -702 -24323 -691 -24277
rect -317 -24323 -306 -24277
rect -198 -24323 -187 -24277
rect 187 -24323 198 -24277
rect 306 -24323 317 -24277
rect 691 -24323 702 -24277
rect -779 -24369 -733 -24358
rect -779 -27354 -733 -27343
rect -275 -24369 -229 -24358
rect -275 -27354 -229 -27343
rect 229 -24369 275 -24358
rect 229 -27354 275 -27343
rect 733 -24369 779 -24358
rect 733 -27354 779 -27343
rect -702 -27435 -691 -27389
rect -317 -27435 -306 -27389
rect -198 -27435 -187 -27389
rect 187 -27435 198 -27389
rect 306 -27435 317 -27389
rect 691 -27435 702 -27389
rect -702 -27555 -691 -27509
rect -317 -27555 -306 -27509
rect -198 -27555 -187 -27509
rect 187 -27555 198 -27509
rect 306 -27555 317 -27509
rect 691 -27555 702 -27509
rect -779 -27601 -733 -27590
rect -779 -30586 -733 -30575
rect -275 -27601 -229 -27590
rect -275 -30586 -229 -30575
rect 229 -27601 275 -27590
rect 229 -30586 275 -30575
rect 733 -27601 779 -27590
rect 733 -30586 779 -30575
rect -702 -30667 -691 -30621
rect -317 -30667 -306 -30621
rect -198 -30667 -187 -30621
rect 187 -30667 198 -30621
rect 306 -30667 317 -30621
rect 691 -30667 702 -30621
rect -702 -30787 -691 -30741
rect -317 -30787 -306 -30741
rect -198 -30787 -187 -30741
rect 187 -30787 198 -30741
rect 306 -30787 317 -30741
rect 691 -30787 702 -30741
rect -779 -30833 -733 -30822
rect -779 -33818 -733 -33807
rect -275 -30833 -229 -30822
rect -275 -33818 -229 -33807
rect 229 -30833 275 -30822
rect 229 -33818 275 -33807
rect 733 -30833 779 -30822
rect 733 -33818 779 -33807
rect -702 -33899 -691 -33853
rect -317 -33899 -306 -33853
rect -198 -33899 -187 -33853
rect 187 -33899 198 -33853
rect 306 -33899 317 -33853
rect 691 -33899 702 -33853
rect -702 -34019 -691 -33973
rect -317 -34019 -306 -33973
rect -198 -34019 -187 -33973
rect 187 -34019 198 -33973
rect 306 -34019 317 -33973
rect 691 -34019 702 -33973
rect -779 -34065 -733 -34054
rect -779 -37050 -733 -37039
rect -275 -34065 -229 -34054
rect -275 -37050 -229 -37039
rect 229 -34065 275 -34054
rect 229 -37050 275 -37039
rect 733 -34065 779 -34054
rect 733 -37050 779 -37039
rect -702 -37131 -691 -37085
rect -317 -37131 -306 -37085
rect -198 -37131 -187 -37085
rect 187 -37131 198 -37085
rect 306 -37131 317 -37085
rect 691 -37131 702 -37085
rect -702 -37251 -691 -37205
rect -317 -37251 -306 -37205
rect -198 -37251 -187 -37205
rect 187 -37251 198 -37205
rect 306 -37251 317 -37205
rect 691 -37251 702 -37205
rect -779 -37297 -733 -37286
rect -779 -40282 -733 -40271
rect -275 -37297 -229 -37286
rect -275 -40282 -229 -40271
rect 229 -37297 275 -37286
rect 229 -40282 275 -40271
rect 733 -37297 779 -37286
rect 733 -40282 779 -40271
rect -917 -40411 -871 -40354
rect -702 -40363 -691 -40317
rect -317 -40363 -306 -40317
rect -198 -40363 -187 -40317
rect 187 -40363 198 -40317
rect 306 -40363 317 -40317
rect 691 -40363 702 -40317
rect 871 -40411 917 -40354
rect -917 -40457 917 -40411
<< properties >>
string FIXED_BBOX -894 -40434 894 40434
string gencell pfet_03v3
string library gf180mcu
string parameters w 15.0 l 2.0 m 25 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
