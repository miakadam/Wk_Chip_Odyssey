magic
tech gf180mcuD
magscale 1 10
timestamp 1757845275
<< error_p >>
rect -38 433 -27 479
rect -38 -479 -27 -433
<< nwell >>
rect -290 -610 290 610
<< pmos >>
rect -40 -400 40 400
<< pdiff >>
rect -128 387 -40 400
rect -128 -387 -115 387
rect -69 -387 -40 387
rect -128 -400 -40 -387
rect 40 387 128 400
rect 40 -387 69 387
rect 115 -387 128 387
rect 40 -400 128 -387
<< pdiffc >>
rect -115 -387 -69 387
rect 69 -387 115 387
<< nsubdiff >>
rect -266 514 266 586
rect -266 470 -194 514
rect -266 -470 -253 470
rect -207 -470 -194 470
rect 194 470 266 514
rect -266 -514 -194 -470
rect 194 -470 207 470
rect 253 -470 266 470
rect 194 -514 266 -470
rect -266 -586 266 -514
<< nsubdiffcont >>
rect -253 -470 -207 470
rect 207 -470 253 470
<< polysilicon >>
rect -40 479 40 492
rect -40 433 -27 479
rect 27 433 40 479
rect -40 400 40 433
rect -40 -433 40 -400
rect -40 -479 -27 -433
rect 27 -479 40 -433
rect -40 -492 40 -479
<< polycontact >>
rect -27 433 27 479
rect -27 -479 27 -433
<< metal1 >>
rect -253 527 253 573
rect -253 470 -207 527
rect -38 433 -27 479
rect 27 433 38 479
rect 207 470 253 527
rect -115 387 -69 398
rect -115 -398 -69 -387
rect 69 387 115 398
rect 69 -398 115 -387
rect -253 -527 -207 -470
rect -38 -479 -27 -433
rect 27 -479 38 -433
rect 207 -527 253 -470
rect -253 -573 253 -527
<< properties >>
string FIXED_BBOX -230 -550 230 550
string gencell pfet_03v3
string library gf180mcu
string parameters w 4.0 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
