magic
tech gf180mcuD
magscale 1 10
timestamp 1758272505
<< nwell >>
rect 39851 38453 40991 39093
rect -4881 36574 -3933 37494
rect 4591 36574 5539 37494
rect 14063 36575 15011 37495
rect 23535 36575 24483 37495
rect 33007 36575 33955 37495
rect 42479 36575 43427 37495
rect -4881 34369 -3933 35289
rect -3395 34369 -2447 35289
rect 4591 34369 5539 35289
rect 6077 34369 7025 35289
rect 14063 34370 15011 35290
rect 15549 34370 16497 35290
rect 23535 34370 24483 35290
rect 25021 34370 25969 35290
rect 33007 34370 33955 35290
rect 34493 34370 35441 35290
rect 42479 34370 43427 35290
rect 43965 34370 44913 35290
rect -4881 32164 -3933 33084
rect -3395 32165 -2447 33085
rect -10023 30949 -9423 31969
rect -9135 30949 -8055 31969
rect 4591 32164 5539 33084
rect 6077 32165 7025 33085
rect 14063 32165 15011 33085
rect 15549 32166 16497 33086
rect -551 30949 49 31969
rect 337 30949 1417 31969
rect 8921 30950 9521 31970
rect 9809 30950 10889 31970
rect 23535 32165 24483 33085
rect 25021 32166 25969 33086
rect 18393 30950 18993 31970
rect 19281 30950 20361 31970
rect 33007 32165 33955 33085
rect 34493 32166 35441 33086
rect 27865 30950 28465 31970
rect 28753 30950 29833 31970
rect 42479 32165 43427 33085
rect 43965 32166 44913 33086
rect 37337 30950 37937 31970
rect 38225 30950 39305 31970
rect -10917 29529 -10317 30549
rect -7795 29773 -5827 30793
rect -4881 29959 -3933 30879
rect -12630 27599 -12030 28619
rect -10023 28609 -9423 29629
rect -9135 28609 -8055 29629
rect -1445 29529 -845 30549
rect 1677 29773 3645 30793
rect 4591 29959 5539 30879
rect -551 28609 49 29629
rect 337 28609 1417 29629
rect 8027 29530 8627 30550
rect 11149 29774 13117 30794
rect 14063 29960 15011 30880
rect 8921 28610 9521 29630
rect 9809 28610 10889 29630
rect 17499 29530 18099 30550
rect 20621 29774 22589 30794
rect 23535 29960 24483 30880
rect 18393 28610 18993 29630
rect 19281 28610 20361 29630
rect 26971 29530 27571 30550
rect 30093 29774 32061 30794
rect 33007 29960 33955 30880
rect 27865 28610 28465 29630
rect 28753 28610 29833 29630
rect 36443 29530 37043 30550
rect 39565 29774 41533 30794
rect 42479 29960 43427 30880
rect 37337 28610 37937 29630
rect 38225 28610 39305 29630
rect -8139 24272 -7191 25192
rect -4097 24269 -3149 25189
rect -55 24269 893 25189
rect 3987 24269 4935 25189
rect 8029 24269 8977 25189
rect 12071 24269 13019 25189
rect 16113 24269 17061 25189
rect -8139 22067 -7191 22987
rect -6653 22067 -5705 22987
rect -4097 22064 -3149 22984
rect -2611 22064 -1663 22984
rect -55 22064 893 22984
rect 1431 22064 2379 22984
rect 3987 22064 4935 22984
rect 5473 22064 6421 22984
rect 8029 22064 8977 22984
rect 9515 22064 10463 22984
rect 12071 22064 13019 22984
rect 13557 22064 14505 22984
rect 16113 22064 17061 22984
rect 17599 22064 18547 22984
rect -8139 19862 -7191 20782
rect -6653 19863 -5705 20783
rect -4097 19859 -3149 20779
rect -2611 19860 -1663 20780
rect -55 19859 893 20779
rect 1431 19860 2379 20780
rect 3987 19859 4935 20779
rect 5473 19860 6421 20780
rect 8029 19859 8977 20779
rect 9515 19860 10463 20780
rect 12071 19859 13019 20779
rect 13557 19860 14505 20780
rect 16113 19859 17061 20779
rect 17599 19860 18547 20780
rect -8139 17657 -7191 18577
rect -4097 17654 -3149 18574
rect -55 17654 893 18574
rect 3987 17654 4935 18574
rect 8029 17654 8977 18574
rect 12071 17654 13019 18574
rect 16113 17654 17061 18574
rect -12151 14693 -11203 15613
rect -8139 14693 -7191 15613
rect -4097 14693 -3149 15613
rect -55 14693 893 15613
rect 3987 14693 4935 15613
rect 8029 14693 8977 15613
rect 12071 14693 13019 15613
rect -12151 12488 -11203 13408
rect -10665 12488 -9717 13408
rect -8139 12488 -7191 13408
rect -6653 12488 -5705 13408
rect -4097 12488 -3149 13408
rect -2611 12488 -1663 13408
rect -55 12488 893 13408
rect 1431 12488 2379 13408
rect 3987 12488 4935 13408
rect 5473 12488 6421 13408
rect 8029 12488 8977 13408
rect 9515 12488 10463 13408
rect 12071 12488 13019 13408
rect 13557 12488 14505 13408
rect -12151 10283 -11203 11203
rect -10665 10284 -9717 11204
rect -8139 10283 -7191 11203
rect -6653 10284 -5705 11204
rect -4097 10283 -3149 11203
rect -2611 10284 -1663 11204
rect -55 10283 893 11203
rect 1431 10284 2379 11204
rect 3987 10283 4935 11203
rect 5473 10284 6421 11204
rect 8029 10283 8977 11203
rect 9515 10284 10463 11204
rect 12071 10283 13019 11203
rect 13557 10284 14505 11204
rect -12151 8078 -11203 8998
rect -8139 8078 -7191 8998
rect -4097 8078 -3149 8998
rect -55 8078 893 8998
rect 3987 8078 4935 8998
rect 8029 8078 8977 8998
rect 12071 8078 13019 8998
rect -11031 4790 -9891 5430
rect -9651 3352 -9071 4524
rect -8681 4457 -7641 5077
rect -7251 3352 -6671 4524
rect -9879 1887 -6443 1907
rect -11199 1307 -10619 1887
rect -10339 1307 -5983 1887
rect -5703 1307 -5123 1887
rect -9879 1287 -6443 1307
<< pwell >>
rect -4118 36334 -4050 36574
rect 5354 36334 5422 36574
rect 14826 36335 14894 36575
rect 24298 36335 24366 36575
rect 33770 36335 33838 36575
rect 43242 36335 43310 36575
rect -4881 35714 -3933 36334
rect 4591 35714 5539 36334
rect 14063 35715 15011 36335
rect 23535 35715 24483 36335
rect 33007 35715 33955 36335
rect 42479 35715 43427 36335
rect -4118 34129 -4050 34369
rect -2632 34129 -2564 34369
rect 5354 34129 5422 34369
rect 6840 34129 6908 34369
rect 14826 34130 14894 34370
rect 16312 34130 16380 34370
rect 24298 34130 24366 34370
rect 25784 34130 25852 34370
rect 33770 34130 33838 34370
rect 35256 34130 35324 34370
rect 43242 34130 43310 34370
rect 44728 34130 44796 34370
rect -4881 33509 -3933 34129
rect -3395 33509 -2447 34129
rect 4591 33509 5539 34129
rect 6077 33509 7025 34129
rect 14063 33510 15011 34130
rect 15549 33510 16497 34130
rect 23535 33510 24483 34130
rect 25021 33510 25969 34130
rect 33007 33510 33955 34130
rect 34493 33510 35441 34130
rect 42479 33510 43427 34130
rect 43965 33510 44913 34130
rect -4118 31924 -4050 32164
rect -2632 31925 -2564 32165
rect -4881 31304 -3933 31924
rect -3395 31305 -2447 31925
rect 5354 31924 5422 32164
rect 6840 31925 6908 32165
rect 4591 31304 5539 31924
rect 6077 31305 7025 31925
rect 14826 31925 14894 32165
rect 16312 31926 16380 32166
rect 14063 31305 15011 31925
rect 15549 31306 16497 31926
rect 24298 31925 24366 32165
rect 25784 31926 25852 32166
rect 23535 31305 24483 31925
rect 25021 31306 25969 31926
rect 33770 31925 33838 32165
rect 35256 31926 35324 32166
rect 33007 31305 33955 31925
rect 34493 31306 35441 31926
rect 43242 31925 43310 32165
rect 44728 31926 44796 32166
rect 42479 31305 43427 31925
rect 43965 31306 44913 31926
rect -8403 30860 -8317 30940
rect -10023 30229 -8055 30849
rect 1069 30860 1155 30940
rect -6175 29684 -6089 29764
rect -4118 29719 -4050 29959
rect -10665 29440 -10579 29520
rect -10917 28809 -10317 29429
rect -7795 29053 -7195 29673
rect -7111 29583 -6511 29673
rect -7111 29325 -6465 29583
rect -7111 29053 -6511 29325
rect -6427 29053 -5827 29673
rect -4881 29099 -3933 29719
rect -551 30229 1417 30849
rect 10541 30861 10627 30941
rect 3297 29684 3383 29764
rect 5354 29719 5422 29959
rect -1193 29440 -1107 29520
rect -1445 28809 -845 29429
rect 1677 29053 2277 29673
rect 2361 29583 2961 29673
rect 2361 29325 3007 29583
rect 2361 29053 2961 29325
rect 3045 29053 3645 29673
rect 4591 29099 5539 29719
rect 8921 30230 10889 30850
rect 20013 30861 20099 30941
rect 12769 29685 12855 29765
rect 14826 29720 14894 29960
rect 8279 29441 8365 29521
rect 8027 28810 8627 29430
rect 11149 29054 11749 29674
rect 11833 29584 12433 29674
rect 11833 29326 12479 29584
rect 11833 29054 12433 29326
rect 12517 29054 13117 29674
rect 14063 29100 15011 29720
rect 18393 30230 20361 30850
rect 29485 30861 29571 30941
rect 22241 29685 22327 29765
rect 24298 29720 24366 29960
rect 17751 29441 17837 29521
rect 17499 28810 18099 29430
rect 20621 29054 21221 29674
rect 21305 29584 21905 29674
rect 21305 29326 21951 29584
rect 21305 29054 21905 29326
rect 21989 29054 22589 29674
rect 23535 29100 24483 29720
rect 27865 30230 29833 30850
rect 38957 30861 39043 30941
rect 31713 29685 31799 29765
rect 33770 29720 33838 29960
rect 27223 29441 27309 29521
rect 26971 28810 27571 29430
rect 30093 29054 30693 29674
rect 30777 29584 31377 29674
rect 30777 29326 31423 29584
rect 30777 29054 31377 29326
rect 31461 29054 32061 29674
rect 33007 29100 33955 29720
rect 37337 30230 39305 30850
rect 41185 29685 41271 29765
rect 43242 29720 43310 29960
rect 36695 29441 36781 29521
rect 36443 28810 37043 29430
rect 39565 29054 40165 29674
rect 40249 29584 40849 29674
rect 40249 29326 40895 29584
rect 40249 29054 40849 29326
rect 40933 29054 41533 29674
rect 42479 29100 43427 29720
rect -8403 28520 -8317 28600
rect 1069 28520 1155 28600
rect 10541 28521 10627 28601
rect 20013 28521 20099 28601
rect 29485 28521 29571 28601
rect 38957 28521 39043 28601
rect -10023 27889 -8055 28509
rect -551 27889 1417 28509
rect 8921 27890 10889 28510
rect 18393 27890 20361 28510
rect 27865 27890 29833 28510
rect 37337 27890 39305 28510
rect -12378 27510 -12292 27590
rect -12630 26879 -12030 27499
rect -7376 24032 -7308 24272
rect -8139 23412 -7191 24032
rect -3334 24029 -3266 24269
rect 708 24029 776 24269
rect 4750 24029 4818 24269
rect 8792 24029 8860 24269
rect 12834 24029 12902 24269
rect 16876 24029 16944 24269
rect -4097 23409 -3149 24029
rect -55 23409 893 24029
rect 3987 23409 4935 24029
rect 8029 23409 8977 24029
rect 12071 23409 13019 24029
rect 16113 23409 17061 24029
rect -7376 21827 -7308 22067
rect -5890 21827 -5822 22067
rect -8139 21207 -7191 21827
rect -6653 21207 -5705 21827
rect -3334 21824 -3266 22064
rect -1848 21824 -1780 22064
rect 708 21824 776 22064
rect 2194 21824 2262 22064
rect 4750 21824 4818 22064
rect 6236 21824 6304 22064
rect 8792 21824 8860 22064
rect 10278 21824 10346 22064
rect 12834 21824 12902 22064
rect 14320 21824 14388 22064
rect 16876 21824 16944 22064
rect 18362 21824 18430 22064
rect -4097 21204 -3149 21824
rect -2611 21204 -1663 21824
rect -55 21204 893 21824
rect 1431 21204 2379 21824
rect 3987 21204 4935 21824
rect 5473 21204 6421 21824
rect 8029 21204 8977 21824
rect 9515 21204 10463 21824
rect 12071 21204 13019 21824
rect 13557 21204 14505 21824
rect 16113 21204 17061 21824
rect 17599 21204 18547 21824
rect -7376 19622 -7308 19862
rect -5890 19623 -5822 19863
rect -8139 19002 -7191 19622
rect -6653 19003 -5705 19623
rect -3334 19619 -3266 19859
rect -1848 19620 -1780 19860
rect -4097 18999 -3149 19619
rect -2611 19000 -1663 19620
rect 708 19619 776 19859
rect 2194 19620 2262 19860
rect -55 18999 893 19619
rect 1431 19000 2379 19620
rect 4750 19619 4818 19859
rect 6236 19620 6304 19860
rect 3987 18999 4935 19619
rect 5473 19000 6421 19620
rect 8792 19619 8860 19859
rect 10278 19620 10346 19860
rect 8029 18999 8977 19619
rect 9515 19000 10463 19620
rect 12834 19619 12902 19859
rect 14320 19620 14388 19860
rect 12071 18999 13019 19619
rect 13557 19000 14505 19620
rect 16876 19619 16944 19859
rect 18362 19620 18430 19860
rect 16113 18999 17061 19619
rect 17599 19000 18547 19620
rect -7376 17417 -7308 17657
rect -8139 16797 -7191 17417
rect -3334 17414 -3266 17654
rect 708 17414 776 17654
rect 4750 17414 4818 17654
rect 8792 17414 8860 17654
rect 12834 17414 12902 17654
rect 16876 17414 16944 17654
rect -4097 16794 -3149 17414
rect -55 16794 893 17414
rect 3987 16794 4935 17414
rect 8029 16794 8977 17414
rect 12071 16794 13019 17414
rect 16113 16794 17061 17414
rect -11388 14453 -11320 14693
rect -7376 14453 -7308 14693
rect -3334 14453 -3266 14693
rect 708 14453 776 14693
rect 4750 14453 4818 14693
rect 8792 14453 8860 14693
rect 12834 14453 12902 14693
rect -12151 13833 -11203 14453
rect -8139 13833 -7191 14453
rect -4097 13833 -3149 14453
rect -55 13833 893 14453
rect 3987 13833 4935 14453
rect 8029 13833 8977 14453
rect 12071 13833 13019 14453
rect -11388 12248 -11320 12488
rect -9902 12248 -9834 12488
rect -7376 12248 -7308 12488
rect -5890 12248 -5822 12488
rect -3334 12248 -3266 12488
rect -1848 12248 -1780 12488
rect 708 12248 776 12488
rect 2194 12248 2262 12488
rect 4750 12248 4818 12488
rect 6236 12248 6304 12488
rect 8792 12248 8860 12488
rect 10278 12248 10346 12488
rect 12834 12248 12902 12488
rect 14320 12248 14388 12488
rect -12151 11628 -11203 12248
rect -10665 11628 -9717 12248
rect -8139 11628 -7191 12248
rect -6653 11628 -5705 12248
rect -4097 11628 -3149 12248
rect -2611 11628 -1663 12248
rect -55 11628 893 12248
rect 1431 11628 2379 12248
rect 3987 11628 4935 12248
rect 5473 11628 6421 12248
rect 8029 11628 8977 12248
rect 9515 11628 10463 12248
rect 12071 11628 13019 12248
rect 13557 11628 14505 12248
rect -11388 10043 -11320 10283
rect -9902 10044 -9834 10284
rect -12151 9423 -11203 10043
rect -10665 9424 -9717 10044
rect -7376 10043 -7308 10283
rect -5890 10044 -5822 10284
rect -8139 9423 -7191 10043
rect -6653 9424 -5705 10044
rect -3334 10043 -3266 10283
rect -1848 10044 -1780 10284
rect -4097 9423 -3149 10043
rect -2611 9424 -1663 10044
rect 708 10043 776 10283
rect 2194 10044 2262 10284
rect -55 9423 893 10043
rect 1431 9424 2379 10044
rect 4750 10043 4818 10283
rect 6236 10044 6304 10284
rect 3987 9423 4935 10043
rect 5473 9424 6421 10044
rect 8792 10043 8860 10283
rect 10278 10044 10346 10284
rect 8029 9423 8977 10043
rect 9515 9424 10463 10044
rect 12834 10043 12902 10283
rect 14320 10044 14388 10284
rect 12071 9423 13019 10043
rect 13557 9424 14505 10044
rect -11388 7838 -11320 8078
rect -7376 7838 -7308 8078
rect -3334 7838 -3266 8078
rect 708 7838 776 8078
rect 4750 7838 4818 8078
rect 8792 7838 8860 8078
rect 12834 7838 12902 8078
rect -12151 7218 -11203 7838
rect -8139 7218 -7191 7838
rect -4097 7218 -3149 7838
rect -55 7218 893 7838
rect 3987 7218 4935 7838
rect 8029 7218 8977 7838
rect 12071 7218 13019 7838
rect -8681 3637 -7641 4257
rect -9651 2552 -9071 3324
rect -7251 2552 -6671 3324
rect -10017 131 -6305 951
rect -6681 -207 -6601 -85
rect -10379 -3003 -5943 -207
<< nmos >>
rect 40051 38033 40111 38203
rect 40221 38033 40281 38203
rect 40391 38033 40451 38203
rect 40561 38033 40621 38203
rect 40731 38033 40791 38203
rect -4631 35924 -4551 36124
rect -4447 35924 -4367 36124
rect -4263 35924 -4183 36124
rect 4841 35924 4921 36124
rect 5025 35924 5105 36124
rect 5209 35924 5289 36124
rect 14313 35925 14393 36125
rect 14497 35925 14577 36125
rect 14681 35925 14761 36125
rect 23785 35925 23865 36125
rect 23969 35925 24049 36125
rect 24153 35925 24233 36125
rect 33257 35925 33337 36125
rect 33441 35925 33521 36125
rect 33625 35925 33705 36125
rect 42729 35925 42809 36125
rect 42913 35925 42993 36125
rect 43097 35925 43177 36125
rect -4631 33719 -4551 33919
rect -4447 33719 -4367 33919
rect -4263 33719 -4183 33919
rect -3145 33719 -3065 33919
rect -2961 33719 -2881 33919
rect -2777 33719 -2697 33919
rect 4841 33719 4921 33919
rect 5025 33719 5105 33919
rect 5209 33719 5289 33919
rect 6327 33719 6407 33919
rect 6511 33719 6591 33919
rect 6695 33719 6775 33919
rect 14313 33720 14393 33920
rect 14497 33720 14577 33920
rect 14681 33720 14761 33920
rect 15799 33720 15879 33920
rect 15983 33720 16063 33920
rect 16167 33720 16247 33920
rect 23785 33720 23865 33920
rect 23969 33720 24049 33920
rect 24153 33720 24233 33920
rect 25271 33720 25351 33920
rect 25455 33720 25535 33920
rect 25639 33720 25719 33920
rect 33257 33720 33337 33920
rect 33441 33720 33521 33920
rect 33625 33720 33705 33920
rect 34743 33720 34823 33920
rect 34927 33720 35007 33920
rect 35111 33720 35191 33920
rect 42729 33720 42809 33920
rect 42913 33720 42993 33920
rect 43097 33720 43177 33920
rect 44215 33720 44295 33920
rect 44399 33720 44479 33920
rect 44583 33720 44663 33920
rect -4631 31514 -4551 31714
rect -4447 31514 -4367 31714
rect -4263 31514 -4183 31714
rect -3145 31515 -3065 31715
rect -2961 31515 -2881 31715
rect -2777 31515 -2697 31715
rect 4841 31514 4921 31714
rect 5025 31514 5105 31714
rect 5209 31514 5289 31714
rect 6327 31515 6407 31715
rect 6511 31515 6591 31715
rect 6695 31515 6775 31715
rect 14313 31515 14393 31715
rect 14497 31515 14577 31715
rect 14681 31515 14761 31715
rect 15799 31516 15879 31716
rect 15983 31516 16063 31716
rect 16167 31516 16247 31716
rect 23785 31515 23865 31715
rect 23969 31515 24049 31715
rect 24153 31515 24233 31715
rect 25271 31516 25351 31716
rect 25455 31516 25535 31716
rect 25639 31516 25719 31716
rect 33257 31515 33337 31715
rect 33441 31515 33521 31715
rect 33625 31515 33705 31715
rect 34743 31516 34823 31716
rect 34927 31516 35007 31716
rect 35111 31516 35191 31716
rect 42729 31515 42809 31715
rect 42913 31515 42993 31715
rect 43097 31515 43177 31715
rect 44215 31516 44295 31716
rect 44399 31516 44479 31716
rect 44583 31516 44663 31716
rect -9773 30439 -9673 30639
rect -9569 30439 -9469 30639
rect -9089 30439 -8989 30639
rect -8885 30439 -8785 30639
rect -8405 30439 -8305 30639
rect -10667 29019 -10567 29219
rect -7545 29263 -7445 29463
rect -6861 29263 -6761 29463
rect -6177 29263 -6077 29463
rect -4631 29309 -4551 29509
rect -4447 29309 -4367 29509
rect -4263 29309 -4183 29509
rect -301 30439 -201 30639
rect -97 30439 3 30639
rect 383 30439 483 30639
rect 587 30439 687 30639
rect 1067 30439 1167 30639
rect -1195 29019 -1095 29219
rect 1927 29263 2027 29463
rect 2611 29263 2711 29463
rect 3295 29263 3395 29463
rect 4841 29309 4921 29509
rect 5025 29309 5105 29509
rect 5209 29309 5289 29509
rect 9171 30440 9271 30640
rect 9375 30440 9475 30640
rect 9855 30440 9955 30640
rect 10059 30440 10159 30640
rect 10539 30440 10639 30640
rect 8277 29020 8377 29220
rect 11399 29264 11499 29464
rect 12083 29264 12183 29464
rect 12767 29264 12867 29464
rect 14313 29310 14393 29510
rect 14497 29310 14577 29510
rect 14681 29310 14761 29510
rect 18643 30440 18743 30640
rect 18847 30440 18947 30640
rect 19327 30440 19427 30640
rect 19531 30440 19631 30640
rect 20011 30440 20111 30640
rect 17749 29020 17849 29220
rect 20871 29264 20971 29464
rect 21555 29264 21655 29464
rect 22239 29264 22339 29464
rect 23785 29310 23865 29510
rect 23969 29310 24049 29510
rect 24153 29310 24233 29510
rect 28115 30440 28215 30640
rect 28319 30440 28419 30640
rect 28799 30440 28899 30640
rect 29003 30440 29103 30640
rect 29483 30440 29583 30640
rect 27221 29020 27321 29220
rect 30343 29264 30443 29464
rect 31027 29264 31127 29464
rect 31711 29264 31811 29464
rect 33257 29310 33337 29510
rect 33441 29310 33521 29510
rect 33625 29310 33705 29510
rect 37587 30440 37687 30640
rect 37791 30440 37891 30640
rect 38271 30440 38371 30640
rect 38475 30440 38575 30640
rect 38955 30440 39055 30640
rect 36693 29020 36793 29220
rect 39815 29264 39915 29464
rect 40499 29264 40599 29464
rect 41183 29264 41283 29464
rect 42729 29310 42809 29510
rect 42913 29310 42993 29510
rect 43097 29310 43177 29510
rect -9773 28099 -9673 28299
rect -9569 28099 -9469 28299
rect -9089 28099 -8989 28299
rect -8885 28099 -8785 28299
rect -8405 28099 -8305 28299
rect -301 28099 -201 28299
rect -97 28099 3 28299
rect 383 28099 483 28299
rect 587 28099 687 28299
rect 1067 28099 1167 28299
rect 9171 28100 9271 28300
rect 9375 28100 9475 28300
rect 9855 28100 9955 28300
rect 10059 28100 10159 28300
rect 10539 28100 10639 28300
rect 18643 28100 18743 28300
rect 18847 28100 18947 28300
rect 19327 28100 19427 28300
rect 19531 28100 19631 28300
rect 20011 28100 20111 28300
rect 28115 28100 28215 28300
rect 28319 28100 28419 28300
rect 28799 28100 28899 28300
rect 29003 28100 29103 28300
rect 29483 28100 29583 28300
rect 37587 28100 37687 28300
rect 37791 28100 37891 28300
rect 38271 28100 38371 28300
rect 38475 28100 38575 28300
rect 38955 28100 39055 28300
rect -12380 27089 -12280 27289
rect -7889 23622 -7809 23822
rect -7705 23622 -7625 23822
rect -7521 23622 -7441 23822
rect -3847 23619 -3767 23819
rect -3663 23619 -3583 23819
rect -3479 23619 -3399 23819
rect 195 23619 275 23819
rect 379 23619 459 23819
rect 563 23619 643 23819
rect 4237 23619 4317 23819
rect 4421 23619 4501 23819
rect 4605 23619 4685 23819
rect 8279 23619 8359 23819
rect 8463 23619 8543 23819
rect 8647 23619 8727 23819
rect 12321 23619 12401 23819
rect 12505 23619 12585 23819
rect 12689 23619 12769 23819
rect 16363 23619 16443 23819
rect 16547 23619 16627 23819
rect 16731 23619 16811 23819
rect -7889 21417 -7809 21617
rect -7705 21417 -7625 21617
rect -7521 21417 -7441 21617
rect -6403 21417 -6323 21617
rect -6219 21417 -6139 21617
rect -6035 21417 -5955 21617
rect -3847 21414 -3767 21614
rect -3663 21414 -3583 21614
rect -3479 21414 -3399 21614
rect -2361 21414 -2281 21614
rect -2177 21414 -2097 21614
rect -1993 21414 -1913 21614
rect 195 21414 275 21614
rect 379 21414 459 21614
rect 563 21414 643 21614
rect 1681 21414 1761 21614
rect 1865 21414 1945 21614
rect 2049 21414 2129 21614
rect 4237 21414 4317 21614
rect 4421 21414 4501 21614
rect 4605 21414 4685 21614
rect 5723 21414 5803 21614
rect 5907 21414 5987 21614
rect 6091 21414 6171 21614
rect 8279 21414 8359 21614
rect 8463 21414 8543 21614
rect 8647 21414 8727 21614
rect 9765 21414 9845 21614
rect 9949 21414 10029 21614
rect 10133 21414 10213 21614
rect 12321 21414 12401 21614
rect 12505 21414 12585 21614
rect 12689 21414 12769 21614
rect 13807 21414 13887 21614
rect 13991 21414 14071 21614
rect 14175 21414 14255 21614
rect 16363 21414 16443 21614
rect 16547 21414 16627 21614
rect 16731 21414 16811 21614
rect 17849 21414 17929 21614
rect 18033 21414 18113 21614
rect 18217 21414 18297 21614
rect -7889 19212 -7809 19412
rect -7705 19212 -7625 19412
rect -7521 19212 -7441 19412
rect -6403 19213 -6323 19413
rect -6219 19213 -6139 19413
rect -6035 19213 -5955 19413
rect -3847 19209 -3767 19409
rect -3663 19209 -3583 19409
rect -3479 19209 -3399 19409
rect -2361 19210 -2281 19410
rect -2177 19210 -2097 19410
rect -1993 19210 -1913 19410
rect 195 19209 275 19409
rect 379 19209 459 19409
rect 563 19209 643 19409
rect 1681 19210 1761 19410
rect 1865 19210 1945 19410
rect 2049 19210 2129 19410
rect 4237 19209 4317 19409
rect 4421 19209 4501 19409
rect 4605 19209 4685 19409
rect 5723 19210 5803 19410
rect 5907 19210 5987 19410
rect 6091 19210 6171 19410
rect 8279 19209 8359 19409
rect 8463 19209 8543 19409
rect 8647 19209 8727 19409
rect 9765 19210 9845 19410
rect 9949 19210 10029 19410
rect 10133 19210 10213 19410
rect 12321 19209 12401 19409
rect 12505 19209 12585 19409
rect 12689 19209 12769 19409
rect 13807 19210 13887 19410
rect 13991 19210 14071 19410
rect 14175 19210 14255 19410
rect 16363 19209 16443 19409
rect 16547 19209 16627 19409
rect 16731 19209 16811 19409
rect 17849 19210 17929 19410
rect 18033 19210 18113 19410
rect 18217 19210 18297 19410
rect -7889 17007 -7809 17207
rect -7705 17007 -7625 17207
rect -7521 17007 -7441 17207
rect -3847 17004 -3767 17204
rect -3663 17004 -3583 17204
rect -3479 17004 -3399 17204
rect 195 17004 275 17204
rect 379 17004 459 17204
rect 563 17004 643 17204
rect 4237 17004 4317 17204
rect 4421 17004 4501 17204
rect 4605 17004 4685 17204
rect 8279 17004 8359 17204
rect 8463 17004 8543 17204
rect 8647 17004 8727 17204
rect 12321 17004 12401 17204
rect 12505 17004 12585 17204
rect 12689 17004 12769 17204
rect 16363 17004 16443 17204
rect 16547 17004 16627 17204
rect 16731 17004 16811 17204
rect -11901 14043 -11821 14243
rect -11717 14043 -11637 14243
rect -11533 14043 -11453 14243
rect -7889 14043 -7809 14243
rect -7705 14043 -7625 14243
rect -7521 14043 -7441 14243
rect -3847 14043 -3767 14243
rect -3663 14043 -3583 14243
rect -3479 14043 -3399 14243
rect 195 14043 275 14243
rect 379 14043 459 14243
rect 563 14043 643 14243
rect 4237 14043 4317 14243
rect 4421 14043 4501 14243
rect 4605 14043 4685 14243
rect 8279 14043 8359 14243
rect 8463 14043 8543 14243
rect 8647 14043 8727 14243
rect 12321 14043 12401 14243
rect 12505 14043 12585 14243
rect 12689 14043 12769 14243
rect -11901 11838 -11821 12038
rect -11717 11838 -11637 12038
rect -11533 11838 -11453 12038
rect -10415 11838 -10335 12038
rect -10231 11838 -10151 12038
rect -10047 11838 -9967 12038
rect -7889 11838 -7809 12038
rect -7705 11838 -7625 12038
rect -7521 11838 -7441 12038
rect -6403 11838 -6323 12038
rect -6219 11838 -6139 12038
rect -6035 11838 -5955 12038
rect -3847 11838 -3767 12038
rect -3663 11838 -3583 12038
rect -3479 11838 -3399 12038
rect -2361 11838 -2281 12038
rect -2177 11838 -2097 12038
rect -1993 11838 -1913 12038
rect 195 11838 275 12038
rect 379 11838 459 12038
rect 563 11838 643 12038
rect 1681 11838 1761 12038
rect 1865 11838 1945 12038
rect 2049 11838 2129 12038
rect 4237 11838 4317 12038
rect 4421 11838 4501 12038
rect 4605 11838 4685 12038
rect 5723 11838 5803 12038
rect 5907 11838 5987 12038
rect 6091 11838 6171 12038
rect 8279 11838 8359 12038
rect 8463 11838 8543 12038
rect 8647 11838 8727 12038
rect 9765 11838 9845 12038
rect 9949 11838 10029 12038
rect 10133 11838 10213 12038
rect 12321 11838 12401 12038
rect 12505 11838 12585 12038
rect 12689 11838 12769 12038
rect 13807 11838 13887 12038
rect 13991 11838 14071 12038
rect 14175 11838 14255 12038
rect -11901 9633 -11821 9833
rect -11717 9633 -11637 9833
rect -11533 9633 -11453 9833
rect -10415 9634 -10335 9834
rect -10231 9634 -10151 9834
rect -10047 9634 -9967 9834
rect -7889 9633 -7809 9833
rect -7705 9633 -7625 9833
rect -7521 9633 -7441 9833
rect -6403 9634 -6323 9834
rect -6219 9634 -6139 9834
rect -6035 9634 -5955 9834
rect -3847 9633 -3767 9833
rect -3663 9633 -3583 9833
rect -3479 9633 -3399 9833
rect -2361 9634 -2281 9834
rect -2177 9634 -2097 9834
rect -1993 9634 -1913 9834
rect 195 9633 275 9833
rect 379 9633 459 9833
rect 563 9633 643 9833
rect 1681 9634 1761 9834
rect 1865 9634 1945 9834
rect 2049 9634 2129 9834
rect 4237 9633 4317 9833
rect 4421 9633 4501 9833
rect 4605 9633 4685 9833
rect 5723 9634 5803 9834
rect 5907 9634 5987 9834
rect 6091 9634 6171 9834
rect 8279 9633 8359 9833
rect 8463 9633 8543 9833
rect 8647 9633 8727 9833
rect 9765 9634 9845 9834
rect 9949 9634 10029 9834
rect 10133 9634 10213 9834
rect 12321 9633 12401 9833
rect 12505 9633 12585 9833
rect 12689 9633 12769 9833
rect 13807 9634 13887 9834
rect 13991 9634 14071 9834
rect 14175 9634 14255 9834
rect -11901 7428 -11821 7628
rect -11717 7428 -11637 7628
rect -11533 7428 -11453 7628
rect -7889 7428 -7809 7628
rect -7705 7428 -7625 7628
rect -7521 7428 -7441 7628
rect -3847 7428 -3767 7628
rect -3663 7428 -3583 7628
rect -3479 7428 -3399 7628
rect 195 7428 275 7628
rect 379 7428 459 7628
rect 563 7428 643 7628
rect 4237 7428 4317 7628
rect 4421 7428 4501 7628
rect 4605 7428 4685 7628
rect 8279 7428 8359 7628
rect 8463 7428 8543 7628
rect 8647 7428 8727 7628
rect 12321 7428 12401 7628
rect 12505 7428 12585 7628
rect 12689 7428 12769 7628
rect -10831 4370 -10771 4540
rect -10661 4370 -10601 4540
rect -10491 4370 -10431 4540
rect -10321 4370 -10261 4540
rect -10151 4370 -10091 4540
rect -8431 3847 -8351 4047
rect -7971 3847 -7891 4047
rect -9401 2714 -9321 3114
rect -7001 2714 -6921 3114
rect -9767 341 -9567 741
rect -9463 341 -9263 741
rect -9159 341 -8959 741
rect -8855 341 -8655 741
rect -8551 341 -8351 741
rect -7971 341 -7771 741
rect -7667 341 -7467 741
rect -7363 341 -7163 741
rect -7059 341 -6859 741
rect -6755 341 -6555 741
rect -9933 -1044 -9733 -744
rect -9629 -1044 -9429 -744
rect -9325 -1044 -9125 -744
rect -9021 -1044 -8821 -744
rect -8717 -1044 -8517 -744
rect -8413 -1044 -8213 -744
rect -8109 -1044 -7909 -744
rect -7805 -1044 -7605 -744
rect -7501 -1044 -7301 -744
rect -7197 -1044 -6997 -744
rect -6893 -1044 -6693 -744
rect -6589 -1044 -6389 -744
rect -9933 -2007 -9733 -1707
rect -9629 -2007 -9429 -1707
rect -9325 -2007 -9125 -1707
rect -9021 -2007 -8821 -1707
rect -8717 -2007 -8517 -1707
rect -8413 -2007 -8213 -1707
rect -8109 -2007 -7909 -1707
rect -7805 -2007 -7605 -1707
rect -7501 -2007 -7301 -1707
rect -7197 -2007 -6997 -1707
rect -6893 -2007 -6693 -1707
rect -6589 -2007 -6389 -1707
rect -8385 -2793 -8305 -2633
rect -8201 -2793 -8121 -2633
rect -8017 -2793 -7937 -2633
<< pmos >>
rect 40051 38543 40111 38883
rect 40221 38543 40281 38883
rect 40391 38543 40451 38883
rect 40561 38543 40621 38883
rect 40731 38543 40791 38883
rect -4631 36784 -4551 37284
rect -4447 36784 -4367 37284
rect -4263 36784 -4183 37284
rect 4841 36784 4921 37284
rect 5025 36784 5105 37284
rect 5209 36784 5289 37284
rect 14313 36785 14393 37285
rect 14497 36785 14577 37285
rect 14681 36785 14761 37285
rect 23785 36785 23865 37285
rect 23969 36785 24049 37285
rect 24153 36785 24233 37285
rect 33257 36785 33337 37285
rect 33441 36785 33521 37285
rect 33625 36785 33705 37285
rect 42729 36785 42809 37285
rect 42913 36785 42993 37285
rect 43097 36785 43177 37285
rect -4631 34579 -4551 35079
rect -4447 34579 -4367 35079
rect -4263 34579 -4183 35079
rect -3145 34579 -3065 35079
rect -2961 34579 -2881 35079
rect -2777 34579 -2697 35079
rect 4841 34579 4921 35079
rect 5025 34579 5105 35079
rect 5209 34579 5289 35079
rect 6327 34579 6407 35079
rect 6511 34579 6591 35079
rect 6695 34579 6775 35079
rect 14313 34580 14393 35080
rect 14497 34580 14577 35080
rect 14681 34580 14761 35080
rect 15799 34580 15879 35080
rect 15983 34580 16063 35080
rect 16167 34580 16247 35080
rect 23785 34580 23865 35080
rect 23969 34580 24049 35080
rect 24153 34580 24233 35080
rect 25271 34580 25351 35080
rect 25455 34580 25535 35080
rect 25639 34580 25719 35080
rect 33257 34580 33337 35080
rect 33441 34580 33521 35080
rect 33625 34580 33705 35080
rect 34743 34580 34823 35080
rect 34927 34580 35007 35080
rect 35111 34580 35191 35080
rect 42729 34580 42809 35080
rect 42913 34580 42993 35080
rect 43097 34580 43177 35080
rect 44215 34580 44295 35080
rect 44399 34580 44479 35080
rect 44583 34580 44663 35080
rect -4631 32374 -4551 32874
rect -4447 32374 -4367 32874
rect -4263 32374 -4183 32874
rect -3145 32375 -3065 32875
rect -2961 32375 -2881 32875
rect -2777 32375 -2697 32875
rect 4841 32374 4921 32874
rect 5025 32374 5105 32874
rect 5209 32374 5289 32874
rect 6327 32375 6407 32875
rect 6511 32375 6591 32875
rect 6695 32375 6775 32875
rect 14313 32375 14393 32875
rect 14497 32375 14577 32875
rect 14681 32375 14761 32875
rect 15799 32376 15879 32876
rect 15983 32376 16063 32876
rect 16167 32376 16247 32876
rect 23785 32375 23865 32875
rect 23969 32375 24049 32875
rect 24153 32375 24233 32875
rect 25271 32376 25351 32876
rect 25455 32376 25535 32876
rect 25639 32376 25719 32876
rect 33257 32375 33337 32875
rect 33441 32375 33521 32875
rect 33625 32375 33705 32875
rect 34743 32376 34823 32876
rect 34927 32376 35007 32876
rect 35111 32376 35191 32876
rect 42729 32375 42809 32875
rect 42913 32375 42993 32875
rect 43097 32375 43177 32875
rect 44215 32376 44295 32876
rect 44399 32376 44479 32876
rect 44583 32376 44663 32876
rect -9773 31159 -9673 31759
rect -8885 31159 -8785 31759
rect -8405 31159 -8305 31759
rect -301 31159 -201 31759
rect 587 31159 687 31759
rect 1067 31159 1167 31759
rect 9171 31160 9271 31760
rect 10059 31160 10159 31760
rect 10539 31160 10639 31760
rect 18643 31160 18743 31760
rect 19531 31160 19631 31760
rect 20011 31160 20111 31760
rect 28115 31160 28215 31760
rect 29003 31160 29103 31760
rect 29483 31160 29583 31760
rect 37587 31160 37687 31760
rect 38475 31160 38575 31760
rect 38955 31160 39055 31760
rect -10667 29739 -10567 30339
rect -7545 29983 -7445 30583
rect -7341 29983 -7241 30583
rect -6861 29983 -6761 30583
rect -6657 29983 -6557 30583
rect -6177 29983 -6077 30583
rect -4631 30169 -4551 30669
rect -4447 30169 -4367 30669
rect -4263 30169 -4183 30669
rect -9773 28819 -9673 29419
rect -8885 28819 -8785 29419
rect -8405 28819 -8305 29419
rect -1195 29739 -1095 30339
rect 1927 29983 2027 30583
rect 2131 29983 2231 30583
rect 2611 29983 2711 30583
rect 2815 29983 2915 30583
rect 3295 29983 3395 30583
rect 4841 30169 4921 30669
rect 5025 30169 5105 30669
rect 5209 30169 5289 30669
rect -301 28819 -201 29419
rect 587 28819 687 29419
rect 1067 28819 1167 29419
rect 8277 29740 8377 30340
rect 11399 29984 11499 30584
rect 11603 29984 11703 30584
rect 12083 29984 12183 30584
rect 12287 29984 12387 30584
rect 12767 29984 12867 30584
rect 14313 30170 14393 30670
rect 14497 30170 14577 30670
rect 14681 30170 14761 30670
rect 9171 28820 9271 29420
rect 10059 28820 10159 29420
rect 10539 28820 10639 29420
rect 17749 29740 17849 30340
rect 20871 29984 20971 30584
rect 21075 29984 21175 30584
rect 21555 29984 21655 30584
rect 21759 29984 21859 30584
rect 22239 29984 22339 30584
rect 23785 30170 23865 30670
rect 23969 30170 24049 30670
rect 24153 30170 24233 30670
rect 18643 28820 18743 29420
rect 19531 28820 19631 29420
rect 20011 28820 20111 29420
rect 27221 29740 27321 30340
rect 30343 29984 30443 30584
rect 30547 29984 30647 30584
rect 31027 29984 31127 30584
rect 31231 29984 31331 30584
rect 31711 29984 31811 30584
rect 33257 30170 33337 30670
rect 33441 30170 33521 30670
rect 33625 30170 33705 30670
rect 28115 28820 28215 29420
rect 29003 28820 29103 29420
rect 29483 28820 29583 29420
rect 36693 29740 36793 30340
rect 39815 29984 39915 30584
rect 40019 29984 40119 30584
rect 40499 29984 40599 30584
rect 40703 29984 40803 30584
rect 41183 29984 41283 30584
rect 42729 30170 42809 30670
rect 42913 30170 42993 30670
rect 43097 30170 43177 30670
rect 37587 28820 37687 29420
rect 38475 28820 38575 29420
rect 38955 28820 39055 29420
rect -12380 27809 -12280 28409
rect -7889 24482 -7809 24982
rect -7705 24482 -7625 24982
rect -7521 24482 -7441 24982
rect -3847 24479 -3767 24979
rect -3663 24479 -3583 24979
rect -3479 24479 -3399 24979
rect 195 24479 275 24979
rect 379 24479 459 24979
rect 563 24479 643 24979
rect 4237 24479 4317 24979
rect 4421 24479 4501 24979
rect 4605 24479 4685 24979
rect 8279 24479 8359 24979
rect 8463 24479 8543 24979
rect 8647 24479 8727 24979
rect 12321 24479 12401 24979
rect 12505 24479 12585 24979
rect 12689 24479 12769 24979
rect 16363 24479 16443 24979
rect 16547 24479 16627 24979
rect 16731 24479 16811 24979
rect -7889 22277 -7809 22777
rect -7705 22277 -7625 22777
rect -7521 22277 -7441 22777
rect -6403 22277 -6323 22777
rect -6219 22277 -6139 22777
rect -6035 22277 -5955 22777
rect -3847 22274 -3767 22774
rect -3663 22274 -3583 22774
rect -3479 22274 -3399 22774
rect -2361 22274 -2281 22774
rect -2177 22274 -2097 22774
rect -1993 22274 -1913 22774
rect 195 22274 275 22774
rect 379 22274 459 22774
rect 563 22274 643 22774
rect 1681 22274 1761 22774
rect 1865 22274 1945 22774
rect 2049 22274 2129 22774
rect 4237 22274 4317 22774
rect 4421 22274 4501 22774
rect 4605 22274 4685 22774
rect 5723 22274 5803 22774
rect 5907 22274 5987 22774
rect 6091 22274 6171 22774
rect 8279 22274 8359 22774
rect 8463 22274 8543 22774
rect 8647 22274 8727 22774
rect 9765 22274 9845 22774
rect 9949 22274 10029 22774
rect 10133 22274 10213 22774
rect 12321 22274 12401 22774
rect 12505 22274 12585 22774
rect 12689 22274 12769 22774
rect 13807 22274 13887 22774
rect 13991 22274 14071 22774
rect 14175 22274 14255 22774
rect 16363 22274 16443 22774
rect 16547 22274 16627 22774
rect 16731 22274 16811 22774
rect 17849 22274 17929 22774
rect 18033 22274 18113 22774
rect 18217 22274 18297 22774
rect -7889 20072 -7809 20572
rect -7705 20072 -7625 20572
rect -7521 20072 -7441 20572
rect -6403 20073 -6323 20573
rect -6219 20073 -6139 20573
rect -6035 20073 -5955 20573
rect -3847 20069 -3767 20569
rect -3663 20069 -3583 20569
rect -3479 20069 -3399 20569
rect -2361 20070 -2281 20570
rect -2177 20070 -2097 20570
rect -1993 20070 -1913 20570
rect 195 20069 275 20569
rect 379 20069 459 20569
rect 563 20069 643 20569
rect 1681 20070 1761 20570
rect 1865 20070 1945 20570
rect 2049 20070 2129 20570
rect 4237 20069 4317 20569
rect 4421 20069 4501 20569
rect 4605 20069 4685 20569
rect 5723 20070 5803 20570
rect 5907 20070 5987 20570
rect 6091 20070 6171 20570
rect 8279 20069 8359 20569
rect 8463 20069 8543 20569
rect 8647 20069 8727 20569
rect 9765 20070 9845 20570
rect 9949 20070 10029 20570
rect 10133 20070 10213 20570
rect 12321 20069 12401 20569
rect 12505 20069 12585 20569
rect 12689 20069 12769 20569
rect 13807 20070 13887 20570
rect 13991 20070 14071 20570
rect 14175 20070 14255 20570
rect 16363 20069 16443 20569
rect 16547 20069 16627 20569
rect 16731 20069 16811 20569
rect 17849 20070 17929 20570
rect 18033 20070 18113 20570
rect 18217 20070 18297 20570
rect -7889 17867 -7809 18367
rect -7705 17867 -7625 18367
rect -7521 17867 -7441 18367
rect -3847 17864 -3767 18364
rect -3663 17864 -3583 18364
rect -3479 17864 -3399 18364
rect 195 17864 275 18364
rect 379 17864 459 18364
rect 563 17864 643 18364
rect 4237 17864 4317 18364
rect 4421 17864 4501 18364
rect 4605 17864 4685 18364
rect 8279 17864 8359 18364
rect 8463 17864 8543 18364
rect 8647 17864 8727 18364
rect 12321 17864 12401 18364
rect 12505 17864 12585 18364
rect 12689 17864 12769 18364
rect 16363 17864 16443 18364
rect 16547 17864 16627 18364
rect 16731 17864 16811 18364
rect -11901 14903 -11821 15403
rect -11717 14903 -11637 15403
rect -11533 14903 -11453 15403
rect -7889 14903 -7809 15403
rect -7705 14903 -7625 15403
rect -7521 14903 -7441 15403
rect -3847 14903 -3767 15403
rect -3663 14903 -3583 15403
rect -3479 14903 -3399 15403
rect 195 14903 275 15403
rect 379 14903 459 15403
rect 563 14903 643 15403
rect 4237 14903 4317 15403
rect 4421 14903 4501 15403
rect 4605 14903 4685 15403
rect 8279 14903 8359 15403
rect 8463 14903 8543 15403
rect 8647 14903 8727 15403
rect 12321 14903 12401 15403
rect 12505 14903 12585 15403
rect 12689 14903 12769 15403
rect -11901 12698 -11821 13198
rect -11717 12698 -11637 13198
rect -11533 12698 -11453 13198
rect -10415 12698 -10335 13198
rect -10231 12698 -10151 13198
rect -10047 12698 -9967 13198
rect -7889 12698 -7809 13198
rect -7705 12698 -7625 13198
rect -7521 12698 -7441 13198
rect -6403 12698 -6323 13198
rect -6219 12698 -6139 13198
rect -6035 12698 -5955 13198
rect -3847 12698 -3767 13198
rect -3663 12698 -3583 13198
rect -3479 12698 -3399 13198
rect -2361 12698 -2281 13198
rect -2177 12698 -2097 13198
rect -1993 12698 -1913 13198
rect 195 12698 275 13198
rect 379 12698 459 13198
rect 563 12698 643 13198
rect 1681 12698 1761 13198
rect 1865 12698 1945 13198
rect 2049 12698 2129 13198
rect 4237 12698 4317 13198
rect 4421 12698 4501 13198
rect 4605 12698 4685 13198
rect 5723 12698 5803 13198
rect 5907 12698 5987 13198
rect 6091 12698 6171 13198
rect 8279 12698 8359 13198
rect 8463 12698 8543 13198
rect 8647 12698 8727 13198
rect 9765 12698 9845 13198
rect 9949 12698 10029 13198
rect 10133 12698 10213 13198
rect 12321 12698 12401 13198
rect 12505 12698 12585 13198
rect 12689 12698 12769 13198
rect 13807 12698 13887 13198
rect 13991 12698 14071 13198
rect 14175 12698 14255 13198
rect -11901 10493 -11821 10993
rect -11717 10493 -11637 10993
rect -11533 10493 -11453 10993
rect -10415 10494 -10335 10994
rect -10231 10494 -10151 10994
rect -10047 10494 -9967 10994
rect -7889 10493 -7809 10993
rect -7705 10493 -7625 10993
rect -7521 10493 -7441 10993
rect -6403 10494 -6323 10994
rect -6219 10494 -6139 10994
rect -6035 10494 -5955 10994
rect -3847 10493 -3767 10993
rect -3663 10493 -3583 10993
rect -3479 10493 -3399 10993
rect -2361 10494 -2281 10994
rect -2177 10494 -2097 10994
rect -1993 10494 -1913 10994
rect 195 10493 275 10993
rect 379 10493 459 10993
rect 563 10493 643 10993
rect 1681 10494 1761 10994
rect 1865 10494 1945 10994
rect 2049 10494 2129 10994
rect 4237 10493 4317 10993
rect 4421 10493 4501 10993
rect 4605 10493 4685 10993
rect 5723 10494 5803 10994
rect 5907 10494 5987 10994
rect 6091 10494 6171 10994
rect 8279 10493 8359 10993
rect 8463 10493 8543 10993
rect 8647 10493 8727 10993
rect 9765 10494 9845 10994
rect 9949 10494 10029 10994
rect 10133 10494 10213 10994
rect 12321 10493 12401 10993
rect 12505 10493 12585 10993
rect 12689 10493 12769 10993
rect 13807 10494 13887 10994
rect 13991 10494 14071 10994
rect 14175 10494 14255 10994
rect -11901 8288 -11821 8788
rect -11717 8288 -11637 8788
rect -11533 8288 -11453 8788
rect -7889 8288 -7809 8788
rect -7705 8288 -7625 8788
rect -7521 8288 -7441 8788
rect -3847 8288 -3767 8788
rect -3663 8288 -3583 8788
rect -3479 8288 -3399 8788
rect 195 8288 275 8788
rect 379 8288 459 8788
rect 563 8288 643 8788
rect 4237 8288 4317 8788
rect 4421 8288 4501 8788
rect 4605 8288 4685 8788
rect 8279 8288 8359 8788
rect 8463 8288 8543 8788
rect 8647 8288 8727 8788
rect 12321 8288 12401 8788
rect 12505 8288 12585 8788
rect 12689 8288 12769 8788
rect -10831 4880 -10771 5220
rect -10661 4880 -10601 5220
rect -10491 4880 -10431 5220
rect -10321 4880 -10261 5220
rect -10151 4880 -10091 5220
rect -8431 4667 -8351 4867
rect -7971 4667 -7891 4867
rect -9401 3562 -9321 4362
rect -7001 3562 -6921 4362
rect -10949 1517 -10869 1677
rect -10089 1517 -10009 1677
rect -9629 1497 -9429 1697
rect -9325 1497 -9125 1697
rect -9021 1497 -8821 1697
rect -8717 1497 -8517 1697
rect -8413 1497 -8213 1697
rect -8109 1497 -7909 1697
rect -7805 1497 -7605 1697
rect -7501 1497 -7301 1697
rect -7197 1497 -6997 1697
rect -6893 1497 -6693 1697
rect -6313 1517 -6233 1677
rect -5453 1517 -5373 1677
<< ndiff >>
rect 39951 38141 40051 38203
rect 39951 38095 39973 38141
rect 40019 38095 40051 38141
rect 39951 38033 40051 38095
rect 40111 38141 40221 38203
rect 40111 38095 40143 38141
rect 40189 38095 40221 38141
rect 40111 38033 40221 38095
rect 40281 38141 40391 38203
rect 40281 38095 40313 38141
rect 40359 38095 40391 38141
rect 40281 38033 40391 38095
rect 40451 38141 40561 38203
rect 40451 38095 40483 38141
rect 40529 38095 40561 38141
rect 40451 38033 40561 38095
rect 40621 38141 40731 38203
rect 40621 38095 40653 38141
rect 40699 38095 40731 38141
rect 40621 38033 40731 38095
rect 40791 38141 40891 38203
rect 40791 38095 40823 38141
rect 40869 38095 40891 38141
rect 40791 38033 40891 38095
rect -4719 36111 -4631 36124
rect -4719 35937 -4706 36111
rect -4660 35937 -4631 36111
rect -4719 35924 -4631 35937
rect -4551 36111 -4447 36124
rect -4551 35937 -4522 36111
rect -4476 35937 -4447 36111
rect -4551 35924 -4447 35937
rect -4367 36111 -4263 36124
rect -4367 35937 -4338 36111
rect -4292 35937 -4263 36111
rect -4367 35924 -4263 35937
rect -4183 36111 -4095 36124
rect -4183 35937 -4154 36111
rect -4108 35937 -4095 36111
rect -4183 35924 -4095 35937
rect 4753 36111 4841 36124
rect 4753 35937 4766 36111
rect 4812 35937 4841 36111
rect 4753 35924 4841 35937
rect 4921 36111 5025 36124
rect 4921 35937 4950 36111
rect 4996 35937 5025 36111
rect 4921 35924 5025 35937
rect 5105 36111 5209 36124
rect 5105 35937 5134 36111
rect 5180 35937 5209 36111
rect 5105 35924 5209 35937
rect 5289 36111 5377 36124
rect 5289 35937 5318 36111
rect 5364 35937 5377 36111
rect 5289 35924 5377 35937
rect 14225 36112 14313 36125
rect 14225 35938 14238 36112
rect 14284 35938 14313 36112
rect 14225 35925 14313 35938
rect 14393 36112 14497 36125
rect 14393 35938 14422 36112
rect 14468 35938 14497 36112
rect 14393 35925 14497 35938
rect 14577 36112 14681 36125
rect 14577 35938 14606 36112
rect 14652 35938 14681 36112
rect 14577 35925 14681 35938
rect 14761 36112 14849 36125
rect 14761 35938 14790 36112
rect 14836 35938 14849 36112
rect 14761 35925 14849 35938
rect 23697 36112 23785 36125
rect 23697 35938 23710 36112
rect 23756 35938 23785 36112
rect 23697 35925 23785 35938
rect 23865 36112 23969 36125
rect 23865 35938 23894 36112
rect 23940 35938 23969 36112
rect 23865 35925 23969 35938
rect 24049 36112 24153 36125
rect 24049 35938 24078 36112
rect 24124 35938 24153 36112
rect 24049 35925 24153 35938
rect 24233 36112 24321 36125
rect 24233 35938 24262 36112
rect 24308 35938 24321 36112
rect 24233 35925 24321 35938
rect 33169 36112 33257 36125
rect 33169 35938 33182 36112
rect 33228 35938 33257 36112
rect 33169 35925 33257 35938
rect 33337 36112 33441 36125
rect 33337 35938 33366 36112
rect 33412 35938 33441 36112
rect 33337 35925 33441 35938
rect 33521 36112 33625 36125
rect 33521 35938 33550 36112
rect 33596 35938 33625 36112
rect 33521 35925 33625 35938
rect 33705 36112 33793 36125
rect 33705 35938 33734 36112
rect 33780 35938 33793 36112
rect 33705 35925 33793 35938
rect 42641 36112 42729 36125
rect 42641 35938 42654 36112
rect 42700 35938 42729 36112
rect 42641 35925 42729 35938
rect 42809 36112 42913 36125
rect 42809 35938 42838 36112
rect 42884 35938 42913 36112
rect 42809 35925 42913 35938
rect 42993 36112 43097 36125
rect 42993 35938 43022 36112
rect 43068 35938 43097 36112
rect 42993 35925 43097 35938
rect 43177 36112 43265 36125
rect 43177 35938 43206 36112
rect 43252 35938 43265 36112
rect 43177 35925 43265 35938
rect -4719 33906 -4631 33919
rect -4719 33732 -4706 33906
rect -4660 33732 -4631 33906
rect -4719 33719 -4631 33732
rect -4551 33906 -4447 33919
rect -4551 33732 -4522 33906
rect -4476 33732 -4447 33906
rect -4551 33719 -4447 33732
rect -4367 33906 -4263 33919
rect -4367 33732 -4338 33906
rect -4292 33732 -4263 33906
rect -4367 33719 -4263 33732
rect -4183 33906 -4095 33919
rect -4183 33732 -4154 33906
rect -4108 33732 -4095 33906
rect -4183 33719 -4095 33732
rect -3233 33906 -3145 33919
rect -3233 33732 -3220 33906
rect -3174 33732 -3145 33906
rect -3233 33719 -3145 33732
rect -3065 33906 -2961 33919
rect -3065 33732 -3036 33906
rect -2990 33732 -2961 33906
rect -3065 33719 -2961 33732
rect -2881 33906 -2777 33919
rect -2881 33732 -2852 33906
rect -2806 33732 -2777 33906
rect -2881 33719 -2777 33732
rect -2697 33906 -2609 33919
rect -2697 33732 -2668 33906
rect -2622 33732 -2609 33906
rect -2697 33719 -2609 33732
rect 4753 33906 4841 33919
rect 4753 33732 4766 33906
rect 4812 33732 4841 33906
rect 4753 33719 4841 33732
rect 4921 33906 5025 33919
rect 4921 33732 4950 33906
rect 4996 33732 5025 33906
rect 4921 33719 5025 33732
rect 5105 33906 5209 33919
rect 5105 33732 5134 33906
rect 5180 33732 5209 33906
rect 5105 33719 5209 33732
rect 5289 33906 5377 33919
rect 5289 33732 5318 33906
rect 5364 33732 5377 33906
rect 5289 33719 5377 33732
rect 6239 33906 6327 33919
rect 6239 33732 6252 33906
rect 6298 33732 6327 33906
rect 6239 33719 6327 33732
rect 6407 33906 6511 33919
rect 6407 33732 6436 33906
rect 6482 33732 6511 33906
rect 6407 33719 6511 33732
rect 6591 33906 6695 33919
rect 6591 33732 6620 33906
rect 6666 33732 6695 33906
rect 6591 33719 6695 33732
rect 6775 33906 6863 33919
rect 6775 33732 6804 33906
rect 6850 33732 6863 33906
rect 6775 33719 6863 33732
rect 14225 33907 14313 33920
rect 14225 33733 14238 33907
rect 14284 33733 14313 33907
rect 14225 33720 14313 33733
rect 14393 33907 14497 33920
rect 14393 33733 14422 33907
rect 14468 33733 14497 33907
rect 14393 33720 14497 33733
rect 14577 33907 14681 33920
rect 14577 33733 14606 33907
rect 14652 33733 14681 33907
rect 14577 33720 14681 33733
rect 14761 33907 14849 33920
rect 14761 33733 14790 33907
rect 14836 33733 14849 33907
rect 14761 33720 14849 33733
rect 15711 33907 15799 33920
rect 15711 33733 15724 33907
rect 15770 33733 15799 33907
rect 15711 33720 15799 33733
rect 15879 33907 15983 33920
rect 15879 33733 15908 33907
rect 15954 33733 15983 33907
rect 15879 33720 15983 33733
rect 16063 33907 16167 33920
rect 16063 33733 16092 33907
rect 16138 33733 16167 33907
rect 16063 33720 16167 33733
rect 16247 33907 16335 33920
rect 16247 33733 16276 33907
rect 16322 33733 16335 33907
rect 16247 33720 16335 33733
rect 23697 33907 23785 33920
rect 23697 33733 23710 33907
rect 23756 33733 23785 33907
rect 23697 33720 23785 33733
rect 23865 33907 23969 33920
rect 23865 33733 23894 33907
rect 23940 33733 23969 33907
rect 23865 33720 23969 33733
rect 24049 33907 24153 33920
rect 24049 33733 24078 33907
rect 24124 33733 24153 33907
rect 24049 33720 24153 33733
rect 24233 33907 24321 33920
rect 24233 33733 24262 33907
rect 24308 33733 24321 33907
rect 24233 33720 24321 33733
rect 25183 33907 25271 33920
rect 25183 33733 25196 33907
rect 25242 33733 25271 33907
rect 25183 33720 25271 33733
rect 25351 33907 25455 33920
rect 25351 33733 25380 33907
rect 25426 33733 25455 33907
rect 25351 33720 25455 33733
rect 25535 33907 25639 33920
rect 25535 33733 25564 33907
rect 25610 33733 25639 33907
rect 25535 33720 25639 33733
rect 25719 33907 25807 33920
rect 25719 33733 25748 33907
rect 25794 33733 25807 33907
rect 25719 33720 25807 33733
rect 33169 33907 33257 33920
rect 33169 33733 33182 33907
rect 33228 33733 33257 33907
rect 33169 33720 33257 33733
rect 33337 33907 33441 33920
rect 33337 33733 33366 33907
rect 33412 33733 33441 33907
rect 33337 33720 33441 33733
rect 33521 33907 33625 33920
rect 33521 33733 33550 33907
rect 33596 33733 33625 33907
rect 33521 33720 33625 33733
rect 33705 33907 33793 33920
rect 33705 33733 33734 33907
rect 33780 33733 33793 33907
rect 33705 33720 33793 33733
rect 34655 33907 34743 33920
rect 34655 33733 34668 33907
rect 34714 33733 34743 33907
rect 34655 33720 34743 33733
rect 34823 33907 34927 33920
rect 34823 33733 34852 33907
rect 34898 33733 34927 33907
rect 34823 33720 34927 33733
rect 35007 33907 35111 33920
rect 35007 33733 35036 33907
rect 35082 33733 35111 33907
rect 35007 33720 35111 33733
rect 35191 33907 35279 33920
rect 35191 33733 35220 33907
rect 35266 33733 35279 33907
rect 35191 33720 35279 33733
rect 42641 33907 42729 33920
rect 42641 33733 42654 33907
rect 42700 33733 42729 33907
rect 42641 33720 42729 33733
rect 42809 33907 42913 33920
rect 42809 33733 42838 33907
rect 42884 33733 42913 33907
rect 42809 33720 42913 33733
rect 42993 33907 43097 33920
rect 42993 33733 43022 33907
rect 43068 33733 43097 33907
rect 42993 33720 43097 33733
rect 43177 33907 43265 33920
rect 43177 33733 43206 33907
rect 43252 33733 43265 33907
rect 43177 33720 43265 33733
rect 44127 33907 44215 33920
rect 44127 33733 44140 33907
rect 44186 33733 44215 33907
rect 44127 33720 44215 33733
rect 44295 33907 44399 33920
rect 44295 33733 44324 33907
rect 44370 33733 44399 33907
rect 44295 33720 44399 33733
rect 44479 33907 44583 33920
rect 44479 33733 44508 33907
rect 44554 33733 44583 33907
rect 44479 33720 44583 33733
rect 44663 33907 44751 33920
rect 44663 33733 44692 33907
rect 44738 33733 44751 33907
rect 44663 33720 44751 33733
rect -4719 31701 -4631 31714
rect -4719 31527 -4706 31701
rect -4660 31527 -4631 31701
rect -4719 31514 -4631 31527
rect -4551 31701 -4447 31714
rect -4551 31527 -4522 31701
rect -4476 31527 -4447 31701
rect -4551 31514 -4447 31527
rect -4367 31701 -4263 31714
rect -4367 31527 -4338 31701
rect -4292 31527 -4263 31701
rect -4367 31514 -4263 31527
rect -4183 31701 -4095 31714
rect -4183 31527 -4154 31701
rect -4108 31527 -4095 31701
rect -4183 31514 -4095 31527
rect -3233 31702 -3145 31715
rect -3233 31528 -3220 31702
rect -3174 31528 -3145 31702
rect -3233 31515 -3145 31528
rect -3065 31702 -2961 31715
rect -3065 31528 -3036 31702
rect -2990 31528 -2961 31702
rect -3065 31515 -2961 31528
rect -2881 31702 -2777 31715
rect -2881 31528 -2852 31702
rect -2806 31528 -2777 31702
rect -2881 31515 -2777 31528
rect -2697 31702 -2609 31715
rect -2697 31528 -2668 31702
rect -2622 31528 -2609 31702
rect -2697 31515 -2609 31528
rect 4753 31701 4841 31714
rect 4753 31527 4766 31701
rect 4812 31527 4841 31701
rect 4753 31514 4841 31527
rect 4921 31701 5025 31714
rect 4921 31527 4950 31701
rect 4996 31527 5025 31701
rect 4921 31514 5025 31527
rect 5105 31701 5209 31714
rect 5105 31527 5134 31701
rect 5180 31527 5209 31701
rect 5105 31514 5209 31527
rect 5289 31701 5377 31714
rect 5289 31527 5318 31701
rect 5364 31527 5377 31701
rect 5289 31514 5377 31527
rect 6239 31702 6327 31715
rect 6239 31528 6252 31702
rect 6298 31528 6327 31702
rect 6239 31515 6327 31528
rect 6407 31702 6511 31715
rect 6407 31528 6436 31702
rect 6482 31528 6511 31702
rect 6407 31515 6511 31528
rect 6591 31702 6695 31715
rect 6591 31528 6620 31702
rect 6666 31528 6695 31702
rect 6591 31515 6695 31528
rect 6775 31702 6863 31715
rect 6775 31528 6804 31702
rect 6850 31528 6863 31702
rect 6775 31515 6863 31528
rect 14225 31702 14313 31715
rect 14225 31528 14238 31702
rect 14284 31528 14313 31702
rect 14225 31515 14313 31528
rect 14393 31702 14497 31715
rect 14393 31528 14422 31702
rect 14468 31528 14497 31702
rect 14393 31515 14497 31528
rect 14577 31702 14681 31715
rect 14577 31528 14606 31702
rect 14652 31528 14681 31702
rect 14577 31515 14681 31528
rect 14761 31702 14849 31715
rect 14761 31528 14790 31702
rect 14836 31528 14849 31702
rect 14761 31515 14849 31528
rect 15711 31703 15799 31716
rect 15711 31529 15724 31703
rect 15770 31529 15799 31703
rect 15711 31516 15799 31529
rect 15879 31703 15983 31716
rect 15879 31529 15908 31703
rect 15954 31529 15983 31703
rect 15879 31516 15983 31529
rect 16063 31703 16167 31716
rect 16063 31529 16092 31703
rect 16138 31529 16167 31703
rect 16063 31516 16167 31529
rect 16247 31703 16335 31716
rect 16247 31529 16276 31703
rect 16322 31529 16335 31703
rect 16247 31516 16335 31529
rect 23697 31702 23785 31715
rect 23697 31528 23710 31702
rect 23756 31528 23785 31702
rect 23697 31515 23785 31528
rect 23865 31702 23969 31715
rect 23865 31528 23894 31702
rect 23940 31528 23969 31702
rect 23865 31515 23969 31528
rect 24049 31702 24153 31715
rect 24049 31528 24078 31702
rect 24124 31528 24153 31702
rect 24049 31515 24153 31528
rect 24233 31702 24321 31715
rect 24233 31528 24262 31702
rect 24308 31528 24321 31702
rect 24233 31515 24321 31528
rect 25183 31703 25271 31716
rect 25183 31529 25196 31703
rect 25242 31529 25271 31703
rect 25183 31516 25271 31529
rect 25351 31703 25455 31716
rect 25351 31529 25380 31703
rect 25426 31529 25455 31703
rect 25351 31516 25455 31529
rect 25535 31703 25639 31716
rect 25535 31529 25564 31703
rect 25610 31529 25639 31703
rect 25535 31516 25639 31529
rect 25719 31703 25807 31716
rect 25719 31529 25748 31703
rect 25794 31529 25807 31703
rect 25719 31516 25807 31529
rect 33169 31702 33257 31715
rect 33169 31528 33182 31702
rect 33228 31528 33257 31702
rect 33169 31515 33257 31528
rect 33337 31702 33441 31715
rect 33337 31528 33366 31702
rect 33412 31528 33441 31702
rect 33337 31515 33441 31528
rect 33521 31702 33625 31715
rect 33521 31528 33550 31702
rect 33596 31528 33625 31702
rect 33521 31515 33625 31528
rect 33705 31702 33793 31715
rect 33705 31528 33734 31702
rect 33780 31528 33793 31702
rect 33705 31515 33793 31528
rect 34655 31703 34743 31716
rect 34655 31529 34668 31703
rect 34714 31529 34743 31703
rect 34655 31516 34743 31529
rect 34823 31703 34927 31716
rect 34823 31529 34852 31703
rect 34898 31529 34927 31703
rect 34823 31516 34927 31529
rect 35007 31703 35111 31716
rect 35007 31529 35036 31703
rect 35082 31529 35111 31703
rect 35007 31516 35111 31529
rect 35191 31703 35279 31716
rect 35191 31529 35220 31703
rect 35266 31529 35279 31703
rect 35191 31516 35279 31529
rect 42641 31702 42729 31715
rect 42641 31528 42654 31702
rect 42700 31528 42729 31702
rect 42641 31515 42729 31528
rect 42809 31702 42913 31715
rect 42809 31528 42838 31702
rect 42884 31528 42913 31702
rect 42809 31515 42913 31528
rect 42993 31702 43097 31715
rect 42993 31528 43022 31702
rect 43068 31528 43097 31702
rect 42993 31515 43097 31528
rect 43177 31702 43265 31715
rect 43177 31528 43206 31702
rect 43252 31528 43265 31702
rect 43177 31515 43265 31528
rect 44127 31703 44215 31716
rect 44127 31529 44140 31703
rect 44186 31529 44215 31703
rect 44127 31516 44215 31529
rect 44295 31703 44399 31716
rect 44295 31529 44324 31703
rect 44370 31529 44399 31703
rect 44295 31516 44399 31529
rect 44479 31703 44583 31716
rect 44479 31529 44508 31703
rect 44554 31529 44583 31703
rect 44479 31516 44583 31529
rect 44663 31703 44751 31716
rect 44663 31529 44692 31703
rect 44738 31529 44751 31703
rect 44663 31516 44751 31529
rect -9861 30626 -9773 30639
rect -9861 30452 -9848 30626
rect -9802 30452 -9773 30626
rect -9861 30439 -9773 30452
rect -9673 30626 -9569 30639
rect -9673 30452 -9644 30626
rect -9598 30452 -9569 30626
rect -9673 30439 -9569 30452
rect -9469 30626 -9381 30639
rect -9469 30452 -9440 30626
rect -9394 30452 -9381 30626
rect -9469 30439 -9381 30452
rect -9177 30626 -9089 30639
rect -9177 30452 -9164 30626
rect -9118 30452 -9089 30626
rect -9177 30439 -9089 30452
rect -8989 30626 -8885 30639
rect -8989 30452 -8960 30626
rect -8914 30452 -8885 30626
rect -8989 30439 -8885 30452
rect -8785 30626 -8697 30639
rect -8785 30452 -8756 30626
rect -8710 30452 -8697 30626
rect -8785 30439 -8697 30452
rect -8493 30626 -8405 30639
rect -8493 30452 -8480 30626
rect -8434 30452 -8405 30626
rect -8493 30439 -8405 30452
rect -8305 30626 -8217 30639
rect -8305 30452 -8276 30626
rect -8230 30452 -8217 30626
rect -8305 30439 -8217 30452
rect -10755 29206 -10667 29219
rect -10755 29032 -10742 29206
rect -10696 29032 -10667 29206
rect -10755 29019 -10667 29032
rect -10567 29206 -10479 29219
rect -10567 29032 -10538 29206
rect -10492 29032 -10479 29206
rect -10567 29019 -10479 29032
rect -7633 29450 -7545 29463
rect -7633 29276 -7620 29450
rect -7574 29276 -7545 29450
rect -7633 29263 -7545 29276
rect -7445 29450 -7357 29463
rect -7445 29276 -7416 29450
rect -7370 29276 -7357 29450
rect -7445 29263 -7357 29276
rect -6949 29450 -6861 29463
rect -6949 29276 -6936 29450
rect -6890 29276 -6861 29450
rect -6949 29263 -6861 29276
rect -6761 29450 -6673 29463
rect -6761 29276 -6732 29450
rect -6686 29276 -6673 29450
rect -6761 29263 -6673 29276
rect -6265 29450 -6177 29463
rect -6265 29276 -6252 29450
rect -6206 29276 -6177 29450
rect -6265 29263 -6177 29276
rect -6077 29450 -5989 29463
rect -6077 29276 -6048 29450
rect -6002 29276 -5989 29450
rect -6077 29263 -5989 29276
rect -4719 29496 -4631 29509
rect -4719 29322 -4706 29496
rect -4660 29322 -4631 29496
rect -4719 29309 -4631 29322
rect -4551 29496 -4447 29509
rect -4551 29322 -4522 29496
rect -4476 29322 -4447 29496
rect -4551 29309 -4447 29322
rect -4367 29496 -4263 29509
rect -4367 29322 -4338 29496
rect -4292 29322 -4263 29496
rect -4367 29309 -4263 29322
rect -4183 29496 -4095 29509
rect -4183 29322 -4154 29496
rect -4108 29322 -4095 29496
rect -4183 29309 -4095 29322
rect -389 30626 -301 30639
rect -389 30452 -376 30626
rect -330 30452 -301 30626
rect -389 30439 -301 30452
rect -201 30626 -97 30639
rect -201 30452 -172 30626
rect -126 30452 -97 30626
rect -201 30439 -97 30452
rect 3 30626 91 30639
rect 3 30452 32 30626
rect 78 30452 91 30626
rect 3 30439 91 30452
rect 295 30626 383 30639
rect 295 30452 308 30626
rect 354 30452 383 30626
rect 295 30439 383 30452
rect 483 30626 587 30639
rect 483 30452 512 30626
rect 558 30452 587 30626
rect 483 30439 587 30452
rect 687 30626 775 30639
rect 687 30452 716 30626
rect 762 30452 775 30626
rect 687 30439 775 30452
rect 979 30626 1067 30639
rect 979 30452 992 30626
rect 1038 30452 1067 30626
rect 979 30439 1067 30452
rect 1167 30626 1255 30639
rect 1167 30452 1196 30626
rect 1242 30452 1255 30626
rect 1167 30439 1255 30452
rect -1283 29206 -1195 29219
rect -1283 29032 -1270 29206
rect -1224 29032 -1195 29206
rect -1283 29019 -1195 29032
rect -1095 29206 -1007 29219
rect -1095 29032 -1066 29206
rect -1020 29032 -1007 29206
rect -1095 29019 -1007 29032
rect 1839 29450 1927 29463
rect 1839 29276 1852 29450
rect 1898 29276 1927 29450
rect 1839 29263 1927 29276
rect 2027 29450 2115 29463
rect 2027 29276 2056 29450
rect 2102 29276 2115 29450
rect 2027 29263 2115 29276
rect 2523 29450 2611 29463
rect 2523 29276 2536 29450
rect 2582 29276 2611 29450
rect 2523 29263 2611 29276
rect 2711 29450 2799 29463
rect 2711 29276 2740 29450
rect 2786 29276 2799 29450
rect 2711 29263 2799 29276
rect 3207 29450 3295 29463
rect 3207 29276 3220 29450
rect 3266 29276 3295 29450
rect 3207 29263 3295 29276
rect 3395 29450 3483 29463
rect 3395 29276 3424 29450
rect 3470 29276 3483 29450
rect 3395 29263 3483 29276
rect 4753 29496 4841 29509
rect 4753 29322 4766 29496
rect 4812 29322 4841 29496
rect 4753 29309 4841 29322
rect 4921 29496 5025 29509
rect 4921 29322 4950 29496
rect 4996 29322 5025 29496
rect 4921 29309 5025 29322
rect 5105 29496 5209 29509
rect 5105 29322 5134 29496
rect 5180 29322 5209 29496
rect 5105 29309 5209 29322
rect 5289 29496 5377 29509
rect 5289 29322 5318 29496
rect 5364 29322 5377 29496
rect 5289 29309 5377 29322
rect 9083 30627 9171 30640
rect 9083 30453 9096 30627
rect 9142 30453 9171 30627
rect 9083 30440 9171 30453
rect 9271 30627 9375 30640
rect 9271 30453 9300 30627
rect 9346 30453 9375 30627
rect 9271 30440 9375 30453
rect 9475 30627 9563 30640
rect 9475 30453 9504 30627
rect 9550 30453 9563 30627
rect 9475 30440 9563 30453
rect 9767 30627 9855 30640
rect 9767 30453 9780 30627
rect 9826 30453 9855 30627
rect 9767 30440 9855 30453
rect 9955 30627 10059 30640
rect 9955 30453 9984 30627
rect 10030 30453 10059 30627
rect 9955 30440 10059 30453
rect 10159 30627 10247 30640
rect 10159 30453 10188 30627
rect 10234 30453 10247 30627
rect 10159 30440 10247 30453
rect 10451 30627 10539 30640
rect 10451 30453 10464 30627
rect 10510 30453 10539 30627
rect 10451 30440 10539 30453
rect 10639 30627 10727 30640
rect 10639 30453 10668 30627
rect 10714 30453 10727 30627
rect 10639 30440 10727 30453
rect 8189 29207 8277 29220
rect 8189 29033 8202 29207
rect 8248 29033 8277 29207
rect 8189 29020 8277 29033
rect 8377 29207 8465 29220
rect 8377 29033 8406 29207
rect 8452 29033 8465 29207
rect 8377 29020 8465 29033
rect 11311 29451 11399 29464
rect 11311 29277 11324 29451
rect 11370 29277 11399 29451
rect 11311 29264 11399 29277
rect 11499 29451 11587 29464
rect 11499 29277 11528 29451
rect 11574 29277 11587 29451
rect 11499 29264 11587 29277
rect 11995 29451 12083 29464
rect 11995 29277 12008 29451
rect 12054 29277 12083 29451
rect 11995 29264 12083 29277
rect 12183 29451 12271 29464
rect 12183 29277 12212 29451
rect 12258 29277 12271 29451
rect 12183 29264 12271 29277
rect 12679 29451 12767 29464
rect 12679 29277 12692 29451
rect 12738 29277 12767 29451
rect 12679 29264 12767 29277
rect 12867 29451 12955 29464
rect 12867 29277 12896 29451
rect 12942 29277 12955 29451
rect 12867 29264 12955 29277
rect 14225 29497 14313 29510
rect 14225 29323 14238 29497
rect 14284 29323 14313 29497
rect 14225 29310 14313 29323
rect 14393 29497 14497 29510
rect 14393 29323 14422 29497
rect 14468 29323 14497 29497
rect 14393 29310 14497 29323
rect 14577 29497 14681 29510
rect 14577 29323 14606 29497
rect 14652 29323 14681 29497
rect 14577 29310 14681 29323
rect 14761 29497 14849 29510
rect 14761 29323 14790 29497
rect 14836 29323 14849 29497
rect 14761 29310 14849 29323
rect 18555 30627 18643 30640
rect 18555 30453 18568 30627
rect 18614 30453 18643 30627
rect 18555 30440 18643 30453
rect 18743 30627 18847 30640
rect 18743 30453 18772 30627
rect 18818 30453 18847 30627
rect 18743 30440 18847 30453
rect 18947 30627 19035 30640
rect 18947 30453 18976 30627
rect 19022 30453 19035 30627
rect 18947 30440 19035 30453
rect 19239 30627 19327 30640
rect 19239 30453 19252 30627
rect 19298 30453 19327 30627
rect 19239 30440 19327 30453
rect 19427 30627 19531 30640
rect 19427 30453 19456 30627
rect 19502 30453 19531 30627
rect 19427 30440 19531 30453
rect 19631 30627 19719 30640
rect 19631 30453 19660 30627
rect 19706 30453 19719 30627
rect 19631 30440 19719 30453
rect 19923 30627 20011 30640
rect 19923 30453 19936 30627
rect 19982 30453 20011 30627
rect 19923 30440 20011 30453
rect 20111 30627 20199 30640
rect 20111 30453 20140 30627
rect 20186 30453 20199 30627
rect 20111 30440 20199 30453
rect 17661 29207 17749 29220
rect 17661 29033 17674 29207
rect 17720 29033 17749 29207
rect 17661 29020 17749 29033
rect 17849 29207 17937 29220
rect 17849 29033 17878 29207
rect 17924 29033 17937 29207
rect 17849 29020 17937 29033
rect 20783 29451 20871 29464
rect 20783 29277 20796 29451
rect 20842 29277 20871 29451
rect 20783 29264 20871 29277
rect 20971 29451 21059 29464
rect 20971 29277 21000 29451
rect 21046 29277 21059 29451
rect 20971 29264 21059 29277
rect 21467 29451 21555 29464
rect 21467 29277 21480 29451
rect 21526 29277 21555 29451
rect 21467 29264 21555 29277
rect 21655 29451 21743 29464
rect 21655 29277 21684 29451
rect 21730 29277 21743 29451
rect 21655 29264 21743 29277
rect 22151 29451 22239 29464
rect 22151 29277 22164 29451
rect 22210 29277 22239 29451
rect 22151 29264 22239 29277
rect 22339 29451 22427 29464
rect 22339 29277 22368 29451
rect 22414 29277 22427 29451
rect 22339 29264 22427 29277
rect 23697 29497 23785 29510
rect 23697 29323 23710 29497
rect 23756 29323 23785 29497
rect 23697 29310 23785 29323
rect 23865 29497 23969 29510
rect 23865 29323 23894 29497
rect 23940 29323 23969 29497
rect 23865 29310 23969 29323
rect 24049 29497 24153 29510
rect 24049 29323 24078 29497
rect 24124 29323 24153 29497
rect 24049 29310 24153 29323
rect 24233 29497 24321 29510
rect 24233 29323 24262 29497
rect 24308 29323 24321 29497
rect 24233 29310 24321 29323
rect 28027 30627 28115 30640
rect 28027 30453 28040 30627
rect 28086 30453 28115 30627
rect 28027 30440 28115 30453
rect 28215 30627 28319 30640
rect 28215 30453 28244 30627
rect 28290 30453 28319 30627
rect 28215 30440 28319 30453
rect 28419 30627 28507 30640
rect 28419 30453 28448 30627
rect 28494 30453 28507 30627
rect 28419 30440 28507 30453
rect 28711 30627 28799 30640
rect 28711 30453 28724 30627
rect 28770 30453 28799 30627
rect 28711 30440 28799 30453
rect 28899 30627 29003 30640
rect 28899 30453 28928 30627
rect 28974 30453 29003 30627
rect 28899 30440 29003 30453
rect 29103 30627 29191 30640
rect 29103 30453 29132 30627
rect 29178 30453 29191 30627
rect 29103 30440 29191 30453
rect 29395 30627 29483 30640
rect 29395 30453 29408 30627
rect 29454 30453 29483 30627
rect 29395 30440 29483 30453
rect 29583 30627 29671 30640
rect 29583 30453 29612 30627
rect 29658 30453 29671 30627
rect 29583 30440 29671 30453
rect 27133 29207 27221 29220
rect 27133 29033 27146 29207
rect 27192 29033 27221 29207
rect 27133 29020 27221 29033
rect 27321 29207 27409 29220
rect 27321 29033 27350 29207
rect 27396 29033 27409 29207
rect 27321 29020 27409 29033
rect 30255 29451 30343 29464
rect 30255 29277 30268 29451
rect 30314 29277 30343 29451
rect 30255 29264 30343 29277
rect 30443 29451 30531 29464
rect 30443 29277 30472 29451
rect 30518 29277 30531 29451
rect 30443 29264 30531 29277
rect 30939 29451 31027 29464
rect 30939 29277 30952 29451
rect 30998 29277 31027 29451
rect 30939 29264 31027 29277
rect 31127 29451 31215 29464
rect 31127 29277 31156 29451
rect 31202 29277 31215 29451
rect 31127 29264 31215 29277
rect 31623 29451 31711 29464
rect 31623 29277 31636 29451
rect 31682 29277 31711 29451
rect 31623 29264 31711 29277
rect 31811 29451 31899 29464
rect 31811 29277 31840 29451
rect 31886 29277 31899 29451
rect 31811 29264 31899 29277
rect 33169 29497 33257 29510
rect 33169 29323 33182 29497
rect 33228 29323 33257 29497
rect 33169 29310 33257 29323
rect 33337 29497 33441 29510
rect 33337 29323 33366 29497
rect 33412 29323 33441 29497
rect 33337 29310 33441 29323
rect 33521 29497 33625 29510
rect 33521 29323 33550 29497
rect 33596 29323 33625 29497
rect 33521 29310 33625 29323
rect 33705 29497 33793 29510
rect 33705 29323 33734 29497
rect 33780 29323 33793 29497
rect 33705 29310 33793 29323
rect 37499 30627 37587 30640
rect 37499 30453 37512 30627
rect 37558 30453 37587 30627
rect 37499 30440 37587 30453
rect 37687 30627 37791 30640
rect 37687 30453 37716 30627
rect 37762 30453 37791 30627
rect 37687 30440 37791 30453
rect 37891 30627 37979 30640
rect 37891 30453 37920 30627
rect 37966 30453 37979 30627
rect 37891 30440 37979 30453
rect 38183 30627 38271 30640
rect 38183 30453 38196 30627
rect 38242 30453 38271 30627
rect 38183 30440 38271 30453
rect 38371 30627 38475 30640
rect 38371 30453 38400 30627
rect 38446 30453 38475 30627
rect 38371 30440 38475 30453
rect 38575 30627 38663 30640
rect 38575 30453 38604 30627
rect 38650 30453 38663 30627
rect 38575 30440 38663 30453
rect 38867 30627 38955 30640
rect 38867 30453 38880 30627
rect 38926 30453 38955 30627
rect 38867 30440 38955 30453
rect 39055 30627 39143 30640
rect 39055 30453 39084 30627
rect 39130 30453 39143 30627
rect 39055 30440 39143 30453
rect 36605 29207 36693 29220
rect 36605 29033 36618 29207
rect 36664 29033 36693 29207
rect 36605 29020 36693 29033
rect 36793 29207 36881 29220
rect 36793 29033 36822 29207
rect 36868 29033 36881 29207
rect 36793 29020 36881 29033
rect 39727 29451 39815 29464
rect 39727 29277 39740 29451
rect 39786 29277 39815 29451
rect 39727 29264 39815 29277
rect 39915 29451 40003 29464
rect 39915 29277 39944 29451
rect 39990 29277 40003 29451
rect 39915 29264 40003 29277
rect 40411 29451 40499 29464
rect 40411 29277 40424 29451
rect 40470 29277 40499 29451
rect 40411 29264 40499 29277
rect 40599 29451 40687 29464
rect 40599 29277 40628 29451
rect 40674 29277 40687 29451
rect 40599 29264 40687 29277
rect 41095 29451 41183 29464
rect 41095 29277 41108 29451
rect 41154 29277 41183 29451
rect 41095 29264 41183 29277
rect 41283 29451 41371 29464
rect 41283 29277 41312 29451
rect 41358 29277 41371 29451
rect 41283 29264 41371 29277
rect 42641 29497 42729 29510
rect 42641 29323 42654 29497
rect 42700 29323 42729 29497
rect 42641 29310 42729 29323
rect 42809 29497 42913 29510
rect 42809 29323 42838 29497
rect 42884 29323 42913 29497
rect 42809 29310 42913 29323
rect 42993 29497 43097 29510
rect 42993 29323 43022 29497
rect 43068 29323 43097 29497
rect 42993 29310 43097 29323
rect 43177 29497 43265 29510
rect 43177 29323 43206 29497
rect 43252 29323 43265 29497
rect 43177 29310 43265 29323
rect -9861 28286 -9773 28299
rect -9861 28112 -9848 28286
rect -9802 28112 -9773 28286
rect -9861 28099 -9773 28112
rect -9673 28286 -9569 28299
rect -9673 28112 -9644 28286
rect -9598 28112 -9569 28286
rect -9673 28099 -9569 28112
rect -9469 28286 -9381 28299
rect -9469 28112 -9440 28286
rect -9394 28112 -9381 28286
rect -9469 28099 -9381 28112
rect -9177 28286 -9089 28299
rect -9177 28112 -9164 28286
rect -9118 28112 -9089 28286
rect -9177 28099 -9089 28112
rect -8989 28286 -8885 28299
rect -8989 28112 -8960 28286
rect -8914 28112 -8885 28286
rect -8989 28099 -8885 28112
rect -8785 28286 -8697 28299
rect -8785 28112 -8756 28286
rect -8710 28112 -8697 28286
rect -8785 28099 -8697 28112
rect -8493 28286 -8405 28299
rect -8493 28112 -8480 28286
rect -8434 28112 -8405 28286
rect -8493 28099 -8405 28112
rect -8305 28286 -8217 28299
rect -8305 28112 -8276 28286
rect -8230 28112 -8217 28286
rect -8305 28099 -8217 28112
rect -389 28286 -301 28299
rect -389 28112 -376 28286
rect -330 28112 -301 28286
rect -389 28099 -301 28112
rect -201 28286 -97 28299
rect -201 28112 -172 28286
rect -126 28112 -97 28286
rect -201 28099 -97 28112
rect 3 28286 91 28299
rect 3 28112 32 28286
rect 78 28112 91 28286
rect 3 28099 91 28112
rect 295 28286 383 28299
rect 295 28112 308 28286
rect 354 28112 383 28286
rect 295 28099 383 28112
rect 483 28286 587 28299
rect 483 28112 512 28286
rect 558 28112 587 28286
rect 483 28099 587 28112
rect 687 28286 775 28299
rect 687 28112 716 28286
rect 762 28112 775 28286
rect 687 28099 775 28112
rect 979 28286 1067 28299
rect 979 28112 992 28286
rect 1038 28112 1067 28286
rect 979 28099 1067 28112
rect 1167 28286 1255 28299
rect 1167 28112 1196 28286
rect 1242 28112 1255 28286
rect 1167 28099 1255 28112
rect 9083 28287 9171 28300
rect 9083 28113 9096 28287
rect 9142 28113 9171 28287
rect 9083 28100 9171 28113
rect 9271 28287 9375 28300
rect 9271 28113 9300 28287
rect 9346 28113 9375 28287
rect 9271 28100 9375 28113
rect 9475 28287 9563 28300
rect 9475 28113 9504 28287
rect 9550 28113 9563 28287
rect 9475 28100 9563 28113
rect 9767 28287 9855 28300
rect 9767 28113 9780 28287
rect 9826 28113 9855 28287
rect 9767 28100 9855 28113
rect 9955 28287 10059 28300
rect 9955 28113 9984 28287
rect 10030 28113 10059 28287
rect 9955 28100 10059 28113
rect 10159 28287 10247 28300
rect 10159 28113 10188 28287
rect 10234 28113 10247 28287
rect 10159 28100 10247 28113
rect 10451 28287 10539 28300
rect 10451 28113 10464 28287
rect 10510 28113 10539 28287
rect 10451 28100 10539 28113
rect 10639 28287 10727 28300
rect 10639 28113 10668 28287
rect 10714 28113 10727 28287
rect 10639 28100 10727 28113
rect 18555 28287 18643 28300
rect 18555 28113 18568 28287
rect 18614 28113 18643 28287
rect 18555 28100 18643 28113
rect 18743 28287 18847 28300
rect 18743 28113 18772 28287
rect 18818 28113 18847 28287
rect 18743 28100 18847 28113
rect 18947 28287 19035 28300
rect 18947 28113 18976 28287
rect 19022 28113 19035 28287
rect 18947 28100 19035 28113
rect 19239 28287 19327 28300
rect 19239 28113 19252 28287
rect 19298 28113 19327 28287
rect 19239 28100 19327 28113
rect 19427 28287 19531 28300
rect 19427 28113 19456 28287
rect 19502 28113 19531 28287
rect 19427 28100 19531 28113
rect 19631 28287 19719 28300
rect 19631 28113 19660 28287
rect 19706 28113 19719 28287
rect 19631 28100 19719 28113
rect 19923 28287 20011 28300
rect 19923 28113 19936 28287
rect 19982 28113 20011 28287
rect 19923 28100 20011 28113
rect 20111 28287 20199 28300
rect 20111 28113 20140 28287
rect 20186 28113 20199 28287
rect 20111 28100 20199 28113
rect 28027 28287 28115 28300
rect 28027 28113 28040 28287
rect 28086 28113 28115 28287
rect 28027 28100 28115 28113
rect 28215 28287 28319 28300
rect 28215 28113 28244 28287
rect 28290 28113 28319 28287
rect 28215 28100 28319 28113
rect 28419 28287 28507 28300
rect 28419 28113 28448 28287
rect 28494 28113 28507 28287
rect 28419 28100 28507 28113
rect 28711 28287 28799 28300
rect 28711 28113 28724 28287
rect 28770 28113 28799 28287
rect 28711 28100 28799 28113
rect 28899 28287 29003 28300
rect 28899 28113 28928 28287
rect 28974 28113 29003 28287
rect 28899 28100 29003 28113
rect 29103 28287 29191 28300
rect 29103 28113 29132 28287
rect 29178 28113 29191 28287
rect 29103 28100 29191 28113
rect 29395 28287 29483 28300
rect 29395 28113 29408 28287
rect 29454 28113 29483 28287
rect 29395 28100 29483 28113
rect 29583 28287 29671 28300
rect 29583 28113 29612 28287
rect 29658 28113 29671 28287
rect 29583 28100 29671 28113
rect 37499 28287 37587 28300
rect 37499 28113 37512 28287
rect 37558 28113 37587 28287
rect 37499 28100 37587 28113
rect 37687 28287 37791 28300
rect 37687 28113 37716 28287
rect 37762 28113 37791 28287
rect 37687 28100 37791 28113
rect 37891 28287 37979 28300
rect 37891 28113 37920 28287
rect 37966 28113 37979 28287
rect 37891 28100 37979 28113
rect 38183 28287 38271 28300
rect 38183 28113 38196 28287
rect 38242 28113 38271 28287
rect 38183 28100 38271 28113
rect 38371 28287 38475 28300
rect 38371 28113 38400 28287
rect 38446 28113 38475 28287
rect 38371 28100 38475 28113
rect 38575 28287 38663 28300
rect 38575 28113 38604 28287
rect 38650 28113 38663 28287
rect 38575 28100 38663 28113
rect 38867 28287 38955 28300
rect 38867 28113 38880 28287
rect 38926 28113 38955 28287
rect 38867 28100 38955 28113
rect 39055 28287 39143 28300
rect 39055 28113 39084 28287
rect 39130 28113 39143 28287
rect 39055 28100 39143 28113
rect -12468 27276 -12380 27289
rect -12468 27102 -12455 27276
rect -12409 27102 -12380 27276
rect -12468 27089 -12380 27102
rect -12280 27276 -12192 27289
rect -12280 27102 -12251 27276
rect -12205 27102 -12192 27276
rect -12280 27089 -12192 27102
rect -7977 23809 -7889 23822
rect -7977 23635 -7964 23809
rect -7918 23635 -7889 23809
rect -7977 23622 -7889 23635
rect -7809 23809 -7705 23822
rect -7809 23635 -7780 23809
rect -7734 23635 -7705 23809
rect -7809 23622 -7705 23635
rect -7625 23809 -7521 23822
rect -7625 23635 -7596 23809
rect -7550 23635 -7521 23809
rect -7625 23622 -7521 23635
rect -7441 23809 -7353 23822
rect -7441 23635 -7412 23809
rect -7366 23635 -7353 23809
rect -7441 23622 -7353 23635
rect -3935 23806 -3847 23819
rect -3935 23632 -3922 23806
rect -3876 23632 -3847 23806
rect -3935 23619 -3847 23632
rect -3767 23806 -3663 23819
rect -3767 23632 -3738 23806
rect -3692 23632 -3663 23806
rect -3767 23619 -3663 23632
rect -3583 23806 -3479 23819
rect -3583 23632 -3554 23806
rect -3508 23632 -3479 23806
rect -3583 23619 -3479 23632
rect -3399 23806 -3311 23819
rect -3399 23632 -3370 23806
rect -3324 23632 -3311 23806
rect -3399 23619 -3311 23632
rect 107 23806 195 23819
rect 107 23632 120 23806
rect 166 23632 195 23806
rect 107 23619 195 23632
rect 275 23806 379 23819
rect 275 23632 304 23806
rect 350 23632 379 23806
rect 275 23619 379 23632
rect 459 23806 563 23819
rect 459 23632 488 23806
rect 534 23632 563 23806
rect 459 23619 563 23632
rect 643 23806 731 23819
rect 643 23632 672 23806
rect 718 23632 731 23806
rect 643 23619 731 23632
rect 4149 23806 4237 23819
rect 4149 23632 4162 23806
rect 4208 23632 4237 23806
rect 4149 23619 4237 23632
rect 4317 23806 4421 23819
rect 4317 23632 4346 23806
rect 4392 23632 4421 23806
rect 4317 23619 4421 23632
rect 4501 23806 4605 23819
rect 4501 23632 4530 23806
rect 4576 23632 4605 23806
rect 4501 23619 4605 23632
rect 4685 23806 4773 23819
rect 4685 23632 4714 23806
rect 4760 23632 4773 23806
rect 4685 23619 4773 23632
rect 8191 23806 8279 23819
rect 8191 23632 8204 23806
rect 8250 23632 8279 23806
rect 8191 23619 8279 23632
rect 8359 23806 8463 23819
rect 8359 23632 8388 23806
rect 8434 23632 8463 23806
rect 8359 23619 8463 23632
rect 8543 23806 8647 23819
rect 8543 23632 8572 23806
rect 8618 23632 8647 23806
rect 8543 23619 8647 23632
rect 8727 23806 8815 23819
rect 8727 23632 8756 23806
rect 8802 23632 8815 23806
rect 8727 23619 8815 23632
rect 12233 23806 12321 23819
rect 12233 23632 12246 23806
rect 12292 23632 12321 23806
rect 12233 23619 12321 23632
rect 12401 23806 12505 23819
rect 12401 23632 12430 23806
rect 12476 23632 12505 23806
rect 12401 23619 12505 23632
rect 12585 23806 12689 23819
rect 12585 23632 12614 23806
rect 12660 23632 12689 23806
rect 12585 23619 12689 23632
rect 12769 23806 12857 23819
rect 12769 23632 12798 23806
rect 12844 23632 12857 23806
rect 12769 23619 12857 23632
rect 16275 23806 16363 23819
rect 16275 23632 16288 23806
rect 16334 23632 16363 23806
rect 16275 23619 16363 23632
rect 16443 23806 16547 23819
rect 16443 23632 16472 23806
rect 16518 23632 16547 23806
rect 16443 23619 16547 23632
rect 16627 23806 16731 23819
rect 16627 23632 16656 23806
rect 16702 23632 16731 23806
rect 16627 23619 16731 23632
rect 16811 23806 16899 23819
rect 16811 23632 16840 23806
rect 16886 23632 16899 23806
rect 16811 23619 16899 23632
rect -7977 21604 -7889 21617
rect -7977 21430 -7964 21604
rect -7918 21430 -7889 21604
rect -7977 21417 -7889 21430
rect -7809 21604 -7705 21617
rect -7809 21430 -7780 21604
rect -7734 21430 -7705 21604
rect -7809 21417 -7705 21430
rect -7625 21604 -7521 21617
rect -7625 21430 -7596 21604
rect -7550 21430 -7521 21604
rect -7625 21417 -7521 21430
rect -7441 21604 -7353 21617
rect -7441 21430 -7412 21604
rect -7366 21430 -7353 21604
rect -7441 21417 -7353 21430
rect -6491 21604 -6403 21617
rect -6491 21430 -6478 21604
rect -6432 21430 -6403 21604
rect -6491 21417 -6403 21430
rect -6323 21604 -6219 21617
rect -6323 21430 -6294 21604
rect -6248 21430 -6219 21604
rect -6323 21417 -6219 21430
rect -6139 21604 -6035 21617
rect -6139 21430 -6110 21604
rect -6064 21430 -6035 21604
rect -6139 21417 -6035 21430
rect -5955 21604 -5867 21617
rect -5955 21430 -5926 21604
rect -5880 21430 -5867 21604
rect -5955 21417 -5867 21430
rect -3935 21601 -3847 21614
rect -3935 21427 -3922 21601
rect -3876 21427 -3847 21601
rect -3935 21414 -3847 21427
rect -3767 21601 -3663 21614
rect -3767 21427 -3738 21601
rect -3692 21427 -3663 21601
rect -3767 21414 -3663 21427
rect -3583 21601 -3479 21614
rect -3583 21427 -3554 21601
rect -3508 21427 -3479 21601
rect -3583 21414 -3479 21427
rect -3399 21601 -3311 21614
rect -3399 21427 -3370 21601
rect -3324 21427 -3311 21601
rect -3399 21414 -3311 21427
rect -2449 21601 -2361 21614
rect -2449 21427 -2436 21601
rect -2390 21427 -2361 21601
rect -2449 21414 -2361 21427
rect -2281 21601 -2177 21614
rect -2281 21427 -2252 21601
rect -2206 21427 -2177 21601
rect -2281 21414 -2177 21427
rect -2097 21601 -1993 21614
rect -2097 21427 -2068 21601
rect -2022 21427 -1993 21601
rect -2097 21414 -1993 21427
rect -1913 21601 -1825 21614
rect -1913 21427 -1884 21601
rect -1838 21427 -1825 21601
rect -1913 21414 -1825 21427
rect 107 21601 195 21614
rect 107 21427 120 21601
rect 166 21427 195 21601
rect 107 21414 195 21427
rect 275 21601 379 21614
rect 275 21427 304 21601
rect 350 21427 379 21601
rect 275 21414 379 21427
rect 459 21601 563 21614
rect 459 21427 488 21601
rect 534 21427 563 21601
rect 459 21414 563 21427
rect 643 21601 731 21614
rect 643 21427 672 21601
rect 718 21427 731 21601
rect 643 21414 731 21427
rect 1593 21601 1681 21614
rect 1593 21427 1606 21601
rect 1652 21427 1681 21601
rect 1593 21414 1681 21427
rect 1761 21601 1865 21614
rect 1761 21427 1790 21601
rect 1836 21427 1865 21601
rect 1761 21414 1865 21427
rect 1945 21601 2049 21614
rect 1945 21427 1974 21601
rect 2020 21427 2049 21601
rect 1945 21414 2049 21427
rect 2129 21601 2217 21614
rect 2129 21427 2158 21601
rect 2204 21427 2217 21601
rect 2129 21414 2217 21427
rect 4149 21601 4237 21614
rect 4149 21427 4162 21601
rect 4208 21427 4237 21601
rect 4149 21414 4237 21427
rect 4317 21601 4421 21614
rect 4317 21427 4346 21601
rect 4392 21427 4421 21601
rect 4317 21414 4421 21427
rect 4501 21601 4605 21614
rect 4501 21427 4530 21601
rect 4576 21427 4605 21601
rect 4501 21414 4605 21427
rect 4685 21601 4773 21614
rect 4685 21427 4714 21601
rect 4760 21427 4773 21601
rect 4685 21414 4773 21427
rect 5635 21601 5723 21614
rect 5635 21427 5648 21601
rect 5694 21427 5723 21601
rect 5635 21414 5723 21427
rect 5803 21601 5907 21614
rect 5803 21427 5832 21601
rect 5878 21427 5907 21601
rect 5803 21414 5907 21427
rect 5987 21601 6091 21614
rect 5987 21427 6016 21601
rect 6062 21427 6091 21601
rect 5987 21414 6091 21427
rect 6171 21601 6259 21614
rect 6171 21427 6200 21601
rect 6246 21427 6259 21601
rect 6171 21414 6259 21427
rect 8191 21601 8279 21614
rect 8191 21427 8204 21601
rect 8250 21427 8279 21601
rect 8191 21414 8279 21427
rect 8359 21601 8463 21614
rect 8359 21427 8388 21601
rect 8434 21427 8463 21601
rect 8359 21414 8463 21427
rect 8543 21601 8647 21614
rect 8543 21427 8572 21601
rect 8618 21427 8647 21601
rect 8543 21414 8647 21427
rect 8727 21601 8815 21614
rect 8727 21427 8756 21601
rect 8802 21427 8815 21601
rect 8727 21414 8815 21427
rect 9677 21601 9765 21614
rect 9677 21427 9690 21601
rect 9736 21427 9765 21601
rect 9677 21414 9765 21427
rect 9845 21601 9949 21614
rect 9845 21427 9874 21601
rect 9920 21427 9949 21601
rect 9845 21414 9949 21427
rect 10029 21601 10133 21614
rect 10029 21427 10058 21601
rect 10104 21427 10133 21601
rect 10029 21414 10133 21427
rect 10213 21601 10301 21614
rect 10213 21427 10242 21601
rect 10288 21427 10301 21601
rect 10213 21414 10301 21427
rect 12233 21601 12321 21614
rect 12233 21427 12246 21601
rect 12292 21427 12321 21601
rect 12233 21414 12321 21427
rect 12401 21601 12505 21614
rect 12401 21427 12430 21601
rect 12476 21427 12505 21601
rect 12401 21414 12505 21427
rect 12585 21601 12689 21614
rect 12585 21427 12614 21601
rect 12660 21427 12689 21601
rect 12585 21414 12689 21427
rect 12769 21601 12857 21614
rect 12769 21427 12798 21601
rect 12844 21427 12857 21601
rect 12769 21414 12857 21427
rect 13719 21601 13807 21614
rect 13719 21427 13732 21601
rect 13778 21427 13807 21601
rect 13719 21414 13807 21427
rect 13887 21601 13991 21614
rect 13887 21427 13916 21601
rect 13962 21427 13991 21601
rect 13887 21414 13991 21427
rect 14071 21601 14175 21614
rect 14071 21427 14100 21601
rect 14146 21427 14175 21601
rect 14071 21414 14175 21427
rect 14255 21601 14343 21614
rect 14255 21427 14284 21601
rect 14330 21427 14343 21601
rect 14255 21414 14343 21427
rect 16275 21601 16363 21614
rect 16275 21427 16288 21601
rect 16334 21427 16363 21601
rect 16275 21414 16363 21427
rect 16443 21601 16547 21614
rect 16443 21427 16472 21601
rect 16518 21427 16547 21601
rect 16443 21414 16547 21427
rect 16627 21601 16731 21614
rect 16627 21427 16656 21601
rect 16702 21427 16731 21601
rect 16627 21414 16731 21427
rect 16811 21601 16899 21614
rect 16811 21427 16840 21601
rect 16886 21427 16899 21601
rect 16811 21414 16899 21427
rect 17761 21601 17849 21614
rect 17761 21427 17774 21601
rect 17820 21427 17849 21601
rect 17761 21414 17849 21427
rect 17929 21601 18033 21614
rect 17929 21427 17958 21601
rect 18004 21427 18033 21601
rect 17929 21414 18033 21427
rect 18113 21601 18217 21614
rect 18113 21427 18142 21601
rect 18188 21427 18217 21601
rect 18113 21414 18217 21427
rect 18297 21601 18385 21614
rect 18297 21427 18326 21601
rect 18372 21427 18385 21601
rect 18297 21414 18385 21427
rect -7977 19399 -7889 19412
rect -7977 19225 -7964 19399
rect -7918 19225 -7889 19399
rect -7977 19212 -7889 19225
rect -7809 19399 -7705 19412
rect -7809 19225 -7780 19399
rect -7734 19225 -7705 19399
rect -7809 19212 -7705 19225
rect -7625 19399 -7521 19412
rect -7625 19225 -7596 19399
rect -7550 19225 -7521 19399
rect -7625 19212 -7521 19225
rect -7441 19399 -7353 19412
rect -7441 19225 -7412 19399
rect -7366 19225 -7353 19399
rect -7441 19212 -7353 19225
rect -6491 19400 -6403 19413
rect -6491 19226 -6478 19400
rect -6432 19226 -6403 19400
rect -6491 19213 -6403 19226
rect -6323 19400 -6219 19413
rect -6323 19226 -6294 19400
rect -6248 19226 -6219 19400
rect -6323 19213 -6219 19226
rect -6139 19400 -6035 19413
rect -6139 19226 -6110 19400
rect -6064 19226 -6035 19400
rect -6139 19213 -6035 19226
rect -5955 19400 -5867 19413
rect -5955 19226 -5926 19400
rect -5880 19226 -5867 19400
rect -5955 19213 -5867 19226
rect -3935 19396 -3847 19409
rect -3935 19222 -3922 19396
rect -3876 19222 -3847 19396
rect -3935 19209 -3847 19222
rect -3767 19396 -3663 19409
rect -3767 19222 -3738 19396
rect -3692 19222 -3663 19396
rect -3767 19209 -3663 19222
rect -3583 19396 -3479 19409
rect -3583 19222 -3554 19396
rect -3508 19222 -3479 19396
rect -3583 19209 -3479 19222
rect -3399 19396 -3311 19409
rect -3399 19222 -3370 19396
rect -3324 19222 -3311 19396
rect -3399 19209 -3311 19222
rect -2449 19397 -2361 19410
rect -2449 19223 -2436 19397
rect -2390 19223 -2361 19397
rect -2449 19210 -2361 19223
rect -2281 19397 -2177 19410
rect -2281 19223 -2252 19397
rect -2206 19223 -2177 19397
rect -2281 19210 -2177 19223
rect -2097 19397 -1993 19410
rect -2097 19223 -2068 19397
rect -2022 19223 -1993 19397
rect -2097 19210 -1993 19223
rect -1913 19397 -1825 19410
rect -1913 19223 -1884 19397
rect -1838 19223 -1825 19397
rect -1913 19210 -1825 19223
rect 107 19396 195 19409
rect 107 19222 120 19396
rect 166 19222 195 19396
rect 107 19209 195 19222
rect 275 19396 379 19409
rect 275 19222 304 19396
rect 350 19222 379 19396
rect 275 19209 379 19222
rect 459 19396 563 19409
rect 459 19222 488 19396
rect 534 19222 563 19396
rect 459 19209 563 19222
rect 643 19396 731 19409
rect 643 19222 672 19396
rect 718 19222 731 19396
rect 643 19209 731 19222
rect 1593 19397 1681 19410
rect 1593 19223 1606 19397
rect 1652 19223 1681 19397
rect 1593 19210 1681 19223
rect 1761 19397 1865 19410
rect 1761 19223 1790 19397
rect 1836 19223 1865 19397
rect 1761 19210 1865 19223
rect 1945 19397 2049 19410
rect 1945 19223 1974 19397
rect 2020 19223 2049 19397
rect 1945 19210 2049 19223
rect 2129 19397 2217 19410
rect 2129 19223 2158 19397
rect 2204 19223 2217 19397
rect 2129 19210 2217 19223
rect 4149 19396 4237 19409
rect 4149 19222 4162 19396
rect 4208 19222 4237 19396
rect 4149 19209 4237 19222
rect 4317 19396 4421 19409
rect 4317 19222 4346 19396
rect 4392 19222 4421 19396
rect 4317 19209 4421 19222
rect 4501 19396 4605 19409
rect 4501 19222 4530 19396
rect 4576 19222 4605 19396
rect 4501 19209 4605 19222
rect 4685 19396 4773 19409
rect 4685 19222 4714 19396
rect 4760 19222 4773 19396
rect 4685 19209 4773 19222
rect 5635 19397 5723 19410
rect 5635 19223 5648 19397
rect 5694 19223 5723 19397
rect 5635 19210 5723 19223
rect 5803 19397 5907 19410
rect 5803 19223 5832 19397
rect 5878 19223 5907 19397
rect 5803 19210 5907 19223
rect 5987 19397 6091 19410
rect 5987 19223 6016 19397
rect 6062 19223 6091 19397
rect 5987 19210 6091 19223
rect 6171 19397 6259 19410
rect 6171 19223 6200 19397
rect 6246 19223 6259 19397
rect 6171 19210 6259 19223
rect 8191 19396 8279 19409
rect 8191 19222 8204 19396
rect 8250 19222 8279 19396
rect 8191 19209 8279 19222
rect 8359 19396 8463 19409
rect 8359 19222 8388 19396
rect 8434 19222 8463 19396
rect 8359 19209 8463 19222
rect 8543 19396 8647 19409
rect 8543 19222 8572 19396
rect 8618 19222 8647 19396
rect 8543 19209 8647 19222
rect 8727 19396 8815 19409
rect 8727 19222 8756 19396
rect 8802 19222 8815 19396
rect 8727 19209 8815 19222
rect 9677 19397 9765 19410
rect 9677 19223 9690 19397
rect 9736 19223 9765 19397
rect 9677 19210 9765 19223
rect 9845 19397 9949 19410
rect 9845 19223 9874 19397
rect 9920 19223 9949 19397
rect 9845 19210 9949 19223
rect 10029 19397 10133 19410
rect 10029 19223 10058 19397
rect 10104 19223 10133 19397
rect 10029 19210 10133 19223
rect 10213 19397 10301 19410
rect 10213 19223 10242 19397
rect 10288 19223 10301 19397
rect 10213 19210 10301 19223
rect 12233 19396 12321 19409
rect 12233 19222 12246 19396
rect 12292 19222 12321 19396
rect 12233 19209 12321 19222
rect 12401 19396 12505 19409
rect 12401 19222 12430 19396
rect 12476 19222 12505 19396
rect 12401 19209 12505 19222
rect 12585 19396 12689 19409
rect 12585 19222 12614 19396
rect 12660 19222 12689 19396
rect 12585 19209 12689 19222
rect 12769 19396 12857 19409
rect 12769 19222 12798 19396
rect 12844 19222 12857 19396
rect 12769 19209 12857 19222
rect 13719 19397 13807 19410
rect 13719 19223 13732 19397
rect 13778 19223 13807 19397
rect 13719 19210 13807 19223
rect 13887 19397 13991 19410
rect 13887 19223 13916 19397
rect 13962 19223 13991 19397
rect 13887 19210 13991 19223
rect 14071 19397 14175 19410
rect 14071 19223 14100 19397
rect 14146 19223 14175 19397
rect 14071 19210 14175 19223
rect 14255 19397 14343 19410
rect 14255 19223 14284 19397
rect 14330 19223 14343 19397
rect 14255 19210 14343 19223
rect 16275 19396 16363 19409
rect 16275 19222 16288 19396
rect 16334 19222 16363 19396
rect 16275 19209 16363 19222
rect 16443 19396 16547 19409
rect 16443 19222 16472 19396
rect 16518 19222 16547 19396
rect 16443 19209 16547 19222
rect 16627 19396 16731 19409
rect 16627 19222 16656 19396
rect 16702 19222 16731 19396
rect 16627 19209 16731 19222
rect 16811 19396 16899 19409
rect 16811 19222 16840 19396
rect 16886 19222 16899 19396
rect 16811 19209 16899 19222
rect 17761 19397 17849 19410
rect 17761 19223 17774 19397
rect 17820 19223 17849 19397
rect 17761 19210 17849 19223
rect 17929 19397 18033 19410
rect 17929 19223 17958 19397
rect 18004 19223 18033 19397
rect 17929 19210 18033 19223
rect 18113 19397 18217 19410
rect 18113 19223 18142 19397
rect 18188 19223 18217 19397
rect 18113 19210 18217 19223
rect 18297 19397 18385 19410
rect 18297 19223 18326 19397
rect 18372 19223 18385 19397
rect 18297 19210 18385 19223
rect -7977 17194 -7889 17207
rect -7977 17020 -7964 17194
rect -7918 17020 -7889 17194
rect -7977 17007 -7889 17020
rect -7809 17194 -7705 17207
rect -7809 17020 -7780 17194
rect -7734 17020 -7705 17194
rect -7809 17007 -7705 17020
rect -7625 17194 -7521 17207
rect -7625 17020 -7596 17194
rect -7550 17020 -7521 17194
rect -7625 17007 -7521 17020
rect -7441 17194 -7353 17207
rect -7441 17020 -7412 17194
rect -7366 17020 -7353 17194
rect -7441 17007 -7353 17020
rect -3935 17191 -3847 17204
rect -3935 17017 -3922 17191
rect -3876 17017 -3847 17191
rect -3935 17004 -3847 17017
rect -3767 17191 -3663 17204
rect -3767 17017 -3738 17191
rect -3692 17017 -3663 17191
rect -3767 17004 -3663 17017
rect -3583 17191 -3479 17204
rect -3583 17017 -3554 17191
rect -3508 17017 -3479 17191
rect -3583 17004 -3479 17017
rect -3399 17191 -3311 17204
rect -3399 17017 -3370 17191
rect -3324 17017 -3311 17191
rect -3399 17004 -3311 17017
rect 107 17191 195 17204
rect 107 17017 120 17191
rect 166 17017 195 17191
rect 107 17004 195 17017
rect 275 17191 379 17204
rect 275 17017 304 17191
rect 350 17017 379 17191
rect 275 17004 379 17017
rect 459 17191 563 17204
rect 459 17017 488 17191
rect 534 17017 563 17191
rect 459 17004 563 17017
rect 643 17191 731 17204
rect 643 17017 672 17191
rect 718 17017 731 17191
rect 643 17004 731 17017
rect 4149 17191 4237 17204
rect 4149 17017 4162 17191
rect 4208 17017 4237 17191
rect 4149 17004 4237 17017
rect 4317 17191 4421 17204
rect 4317 17017 4346 17191
rect 4392 17017 4421 17191
rect 4317 17004 4421 17017
rect 4501 17191 4605 17204
rect 4501 17017 4530 17191
rect 4576 17017 4605 17191
rect 4501 17004 4605 17017
rect 4685 17191 4773 17204
rect 4685 17017 4714 17191
rect 4760 17017 4773 17191
rect 4685 17004 4773 17017
rect 8191 17191 8279 17204
rect 8191 17017 8204 17191
rect 8250 17017 8279 17191
rect 8191 17004 8279 17017
rect 8359 17191 8463 17204
rect 8359 17017 8388 17191
rect 8434 17017 8463 17191
rect 8359 17004 8463 17017
rect 8543 17191 8647 17204
rect 8543 17017 8572 17191
rect 8618 17017 8647 17191
rect 8543 17004 8647 17017
rect 8727 17191 8815 17204
rect 8727 17017 8756 17191
rect 8802 17017 8815 17191
rect 8727 17004 8815 17017
rect 12233 17191 12321 17204
rect 12233 17017 12246 17191
rect 12292 17017 12321 17191
rect 12233 17004 12321 17017
rect 12401 17191 12505 17204
rect 12401 17017 12430 17191
rect 12476 17017 12505 17191
rect 12401 17004 12505 17017
rect 12585 17191 12689 17204
rect 12585 17017 12614 17191
rect 12660 17017 12689 17191
rect 12585 17004 12689 17017
rect 12769 17191 12857 17204
rect 12769 17017 12798 17191
rect 12844 17017 12857 17191
rect 12769 17004 12857 17017
rect 16275 17191 16363 17204
rect 16275 17017 16288 17191
rect 16334 17017 16363 17191
rect 16275 17004 16363 17017
rect 16443 17191 16547 17204
rect 16443 17017 16472 17191
rect 16518 17017 16547 17191
rect 16443 17004 16547 17017
rect 16627 17191 16731 17204
rect 16627 17017 16656 17191
rect 16702 17017 16731 17191
rect 16627 17004 16731 17017
rect 16811 17191 16899 17204
rect 16811 17017 16840 17191
rect 16886 17017 16899 17191
rect 16811 17004 16899 17017
rect -11989 14230 -11901 14243
rect -11989 14056 -11976 14230
rect -11930 14056 -11901 14230
rect -11989 14043 -11901 14056
rect -11821 14230 -11717 14243
rect -11821 14056 -11792 14230
rect -11746 14056 -11717 14230
rect -11821 14043 -11717 14056
rect -11637 14230 -11533 14243
rect -11637 14056 -11608 14230
rect -11562 14056 -11533 14230
rect -11637 14043 -11533 14056
rect -11453 14230 -11365 14243
rect -11453 14056 -11424 14230
rect -11378 14056 -11365 14230
rect -11453 14043 -11365 14056
rect -7977 14230 -7889 14243
rect -7977 14056 -7964 14230
rect -7918 14056 -7889 14230
rect -7977 14043 -7889 14056
rect -7809 14230 -7705 14243
rect -7809 14056 -7780 14230
rect -7734 14056 -7705 14230
rect -7809 14043 -7705 14056
rect -7625 14230 -7521 14243
rect -7625 14056 -7596 14230
rect -7550 14056 -7521 14230
rect -7625 14043 -7521 14056
rect -7441 14230 -7353 14243
rect -7441 14056 -7412 14230
rect -7366 14056 -7353 14230
rect -7441 14043 -7353 14056
rect -3935 14230 -3847 14243
rect -3935 14056 -3922 14230
rect -3876 14056 -3847 14230
rect -3935 14043 -3847 14056
rect -3767 14230 -3663 14243
rect -3767 14056 -3738 14230
rect -3692 14056 -3663 14230
rect -3767 14043 -3663 14056
rect -3583 14230 -3479 14243
rect -3583 14056 -3554 14230
rect -3508 14056 -3479 14230
rect -3583 14043 -3479 14056
rect -3399 14230 -3311 14243
rect -3399 14056 -3370 14230
rect -3324 14056 -3311 14230
rect -3399 14043 -3311 14056
rect 107 14230 195 14243
rect 107 14056 120 14230
rect 166 14056 195 14230
rect 107 14043 195 14056
rect 275 14230 379 14243
rect 275 14056 304 14230
rect 350 14056 379 14230
rect 275 14043 379 14056
rect 459 14230 563 14243
rect 459 14056 488 14230
rect 534 14056 563 14230
rect 459 14043 563 14056
rect 643 14230 731 14243
rect 643 14056 672 14230
rect 718 14056 731 14230
rect 643 14043 731 14056
rect 4149 14230 4237 14243
rect 4149 14056 4162 14230
rect 4208 14056 4237 14230
rect 4149 14043 4237 14056
rect 4317 14230 4421 14243
rect 4317 14056 4346 14230
rect 4392 14056 4421 14230
rect 4317 14043 4421 14056
rect 4501 14230 4605 14243
rect 4501 14056 4530 14230
rect 4576 14056 4605 14230
rect 4501 14043 4605 14056
rect 4685 14230 4773 14243
rect 4685 14056 4714 14230
rect 4760 14056 4773 14230
rect 4685 14043 4773 14056
rect 8191 14230 8279 14243
rect 8191 14056 8204 14230
rect 8250 14056 8279 14230
rect 8191 14043 8279 14056
rect 8359 14230 8463 14243
rect 8359 14056 8388 14230
rect 8434 14056 8463 14230
rect 8359 14043 8463 14056
rect 8543 14230 8647 14243
rect 8543 14056 8572 14230
rect 8618 14056 8647 14230
rect 8543 14043 8647 14056
rect 8727 14230 8815 14243
rect 8727 14056 8756 14230
rect 8802 14056 8815 14230
rect 8727 14043 8815 14056
rect 12233 14230 12321 14243
rect 12233 14056 12246 14230
rect 12292 14056 12321 14230
rect 12233 14043 12321 14056
rect 12401 14230 12505 14243
rect 12401 14056 12430 14230
rect 12476 14056 12505 14230
rect 12401 14043 12505 14056
rect 12585 14230 12689 14243
rect 12585 14056 12614 14230
rect 12660 14056 12689 14230
rect 12585 14043 12689 14056
rect 12769 14230 12857 14243
rect 12769 14056 12798 14230
rect 12844 14056 12857 14230
rect 12769 14043 12857 14056
rect -11989 12025 -11901 12038
rect -11989 11851 -11976 12025
rect -11930 11851 -11901 12025
rect -11989 11838 -11901 11851
rect -11821 12025 -11717 12038
rect -11821 11851 -11792 12025
rect -11746 11851 -11717 12025
rect -11821 11838 -11717 11851
rect -11637 12025 -11533 12038
rect -11637 11851 -11608 12025
rect -11562 11851 -11533 12025
rect -11637 11838 -11533 11851
rect -11453 12025 -11365 12038
rect -11453 11851 -11424 12025
rect -11378 11851 -11365 12025
rect -11453 11838 -11365 11851
rect -10503 12025 -10415 12038
rect -10503 11851 -10490 12025
rect -10444 11851 -10415 12025
rect -10503 11838 -10415 11851
rect -10335 12025 -10231 12038
rect -10335 11851 -10306 12025
rect -10260 11851 -10231 12025
rect -10335 11838 -10231 11851
rect -10151 12025 -10047 12038
rect -10151 11851 -10122 12025
rect -10076 11851 -10047 12025
rect -10151 11838 -10047 11851
rect -9967 12025 -9879 12038
rect -9967 11851 -9938 12025
rect -9892 11851 -9879 12025
rect -9967 11838 -9879 11851
rect -7977 12025 -7889 12038
rect -7977 11851 -7964 12025
rect -7918 11851 -7889 12025
rect -7977 11838 -7889 11851
rect -7809 12025 -7705 12038
rect -7809 11851 -7780 12025
rect -7734 11851 -7705 12025
rect -7809 11838 -7705 11851
rect -7625 12025 -7521 12038
rect -7625 11851 -7596 12025
rect -7550 11851 -7521 12025
rect -7625 11838 -7521 11851
rect -7441 12025 -7353 12038
rect -7441 11851 -7412 12025
rect -7366 11851 -7353 12025
rect -7441 11838 -7353 11851
rect -6491 12025 -6403 12038
rect -6491 11851 -6478 12025
rect -6432 11851 -6403 12025
rect -6491 11838 -6403 11851
rect -6323 12025 -6219 12038
rect -6323 11851 -6294 12025
rect -6248 11851 -6219 12025
rect -6323 11838 -6219 11851
rect -6139 12025 -6035 12038
rect -6139 11851 -6110 12025
rect -6064 11851 -6035 12025
rect -6139 11838 -6035 11851
rect -5955 12025 -5867 12038
rect -5955 11851 -5926 12025
rect -5880 11851 -5867 12025
rect -5955 11838 -5867 11851
rect -3935 12025 -3847 12038
rect -3935 11851 -3922 12025
rect -3876 11851 -3847 12025
rect -3935 11838 -3847 11851
rect -3767 12025 -3663 12038
rect -3767 11851 -3738 12025
rect -3692 11851 -3663 12025
rect -3767 11838 -3663 11851
rect -3583 12025 -3479 12038
rect -3583 11851 -3554 12025
rect -3508 11851 -3479 12025
rect -3583 11838 -3479 11851
rect -3399 12025 -3311 12038
rect -3399 11851 -3370 12025
rect -3324 11851 -3311 12025
rect -3399 11838 -3311 11851
rect -2449 12025 -2361 12038
rect -2449 11851 -2436 12025
rect -2390 11851 -2361 12025
rect -2449 11838 -2361 11851
rect -2281 12025 -2177 12038
rect -2281 11851 -2252 12025
rect -2206 11851 -2177 12025
rect -2281 11838 -2177 11851
rect -2097 12025 -1993 12038
rect -2097 11851 -2068 12025
rect -2022 11851 -1993 12025
rect -2097 11838 -1993 11851
rect -1913 12025 -1825 12038
rect -1913 11851 -1884 12025
rect -1838 11851 -1825 12025
rect -1913 11838 -1825 11851
rect 107 12025 195 12038
rect 107 11851 120 12025
rect 166 11851 195 12025
rect 107 11838 195 11851
rect 275 12025 379 12038
rect 275 11851 304 12025
rect 350 11851 379 12025
rect 275 11838 379 11851
rect 459 12025 563 12038
rect 459 11851 488 12025
rect 534 11851 563 12025
rect 459 11838 563 11851
rect 643 12025 731 12038
rect 643 11851 672 12025
rect 718 11851 731 12025
rect 643 11838 731 11851
rect 1593 12025 1681 12038
rect 1593 11851 1606 12025
rect 1652 11851 1681 12025
rect 1593 11838 1681 11851
rect 1761 12025 1865 12038
rect 1761 11851 1790 12025
rect 1836 11851 1865 12025
rect 1761 11838 1865 11851
rect 1945 12025 2049 12038
rect 1945 11851 1974 12025
rect 2020 11851 2049 12025
rect 1945 11838 2049 11851
rect 2129 12025 2217 12038
rect 2129 11851 2158 12025
rect 2204 11851 2217 12025
rect 2129 11838 2217 11851
rect 4149 12025 4237 12038
rect 4149 11851 4162 12025
rect 4208 11851 4237 12025
rect 4149 11838 4237 11851
rect 4317 12025 4421 12038
rect 4317 11851 4346 12025
rect 4392 11851 4421 12025
rect 4317 11838 4421 11851
rect 4501 12025 4605 12038
rect 4501 11851 4530 12025
rect 4576 11851 4605 12025
rect 4501 11838 4605 11851
rect 4685 12025 4773 12038
rect 4685 11851 4714 12025
rect 4760 11851 4773 12025
rect 4685 11838 4773 11851
rect 5635 12025 5723 12038
rect 5635 11851 5648 12025
rect 5694 11851 5723 12025
rect 5635 11838 5723 11851
rect 5803 12025 5907 12038
rect 5803 11851 5832 12025
rect 5878 11851 5907 12025
rect 5803 11838 5907 11851
rect 5987 12025 6091 12038
rect 5987 11851 6016 12025
rect 6062 11851 6091 12025
rect 5987 11838 6091 11851
rect 6171 12025 6259 12038
rect 6171 11851 6200 12025
rect 6246 11851 6259 12025
rect 6171 11838 6259 11851
rect 8191 12025 8279 12038
rect 8191 11851 8204 12025
rect 8250 11851 8279 12025
rect 8191 11838 8279 11851
rect 8359 12025 8463 12038
rect 8359 11851 8388 12025
rect 8434 11851 8463 12025
rect 8359 11838 8463 11851
rect 8543 12025 8647 12038
rect 8543 11851 8572 12025
rect 8618 11851 8647 12025
rect 8543 11838 8647 11851
rect 8727 12025 8815 12038
rect 8727 11851 8756 12025
rect 8802 11851 8815 12025
rect 8727 11838 8815 11851
rect 9677 12025 9765 12038
rect 9677 11851 9690 12025
rect 9736 11851 9765 12025
rect 9677 11838 9765 11851
rect 9845 12025 9949 12038
rect 9845 11851 9874 12025
rect 9920 11851 9949 12025
rect 9845 11838 9949 11851
rect 10029 12025 10133 12038
rect 10029 11851 10058 12025
rect 10104 11851 10133 12025
rect 10029 11838 10133 11851
rect 10213 12025 10301 12038
rect 10213 11851 10242 12025
rect 10288 11851 10301 12025
rect 10213 11838 10301 11851
rect 12233 12025 12321 12038
rect 12233 11851 12246 12025
rect 12292 11851 12321 12025
rect 12233 11838 12321 11851
rect 12401 12025 12505 12038
rect 12401 11851 12430 12025
rect 12476 11851 12505 12025
rect 12401 11838 12505 11851
rect 12585 12025 12689 12038
rect 12585 11851 12614 12025
rect 12660 11851 12689 12025
rect 12585 11838 12689 11851
rect 12769 12025 12857 12038
rect 12769 11851 12798 12025
rect 12844 11851 12857 12025
rect 12769 11838 12857 11851
rect 13719 12025 13807 12038
rect 13719 11851 13732 12025
rect 13778 11851 13807 12025
rect 13719 11838 13807 11851
rect 13887 12025 13991 12038
rect 13887 11851 13916 12025
rect 13962 11851 13991 12025
rect 13887 11838 13991 11851
rect 14071 12025 14175 12038
rect 14071 11851 14100 12025
rect 14146 11851 14175 12025
rect 14071 11838 14175 11851
rect 14255 12025 14343 12038
rect 14255 11851 14284 12025
rect 14330 11851 14343 12025
rect 14255 11838 14343 11851
rect -11989 9820 -11901 9833
rect -11989 9646 -11976 9820
rect -11930 9646 -11901 9820
rect -11989 9633 -11901 9646
rect -11821 9820 -11717 9833
rect -11821 9646 -11792 9820
rect -11746 9646 -11717 9820
rect -11821 9633 -11717 9646
rect -11637 9820 -11533 9833
rect -11637 9646 -11608 9820
rect -11562 9646 -11533 9820
rect -11637 9633 -11533 9646
rect -11453 9820 -11365 9833
rect -11453 9646 -11424 9820
rect -11378 9646 -11365 9820
rect -11453 9633 -11365 9646
rect -10503 9821 -10415 9834
rect -10503 9647 -10490 9821
rect -10444 9647 -10415 9821
rect -10503 9634 -10415 9647
rect -10335 9821 -10231 9834
rect -10335 9647 -10306 9821
rect -10260 9647 -10231 9821
rect -10335 9634 -10231 9647
rect -10151 9821 -10047 9834
rect -10151 9647 -10122 9821
rect -10076 9647 -10047 9821
rect -10151 9634 -10047 9647
rect -9967 9821 -9879 9834
rect -9967 9647 -9938 9821
rect -9892 9647 -9879 9821
rect -9967 9634 -9879 9647
rect -7977 9820 -7889 9833
rect -7977 9646 -7964 9820
rect -7918 9646 -7889 9820
rect -7977 9633 -7889 9646
rect -7809 9820 -7705 9833
rect -7809 9646 -7780 9820
rect -7734 9646 -7705 9820
rect -7809 9633 -7705 9646
rect -7625 9820 -7521 9833
rect -7625 9646 -7596 9820
rect -7550 9646 -7521 9820
rect -7625 9633 -7521 9646
rect -7441 9820 -7353 9833
rect -7441 9646 -7412 9820
rect -7366 9646 -7353 9820
rect -7441 9633 -7353 9646
rect -6491 9821 -6403 9834
rect -6491 9647 -6478 9821
rect -6432 9647 -6403 9821
rect -6491 9634 -6403 9647
rect -6323 9821 -6219 9834
rect -6323 9647 -6294 9821
rect -6248 9647 -6219 9821
rect -6323 9634 -6219 9647
rect -6139 9821 -6035 9834
rect -6139 9647 -6110 9821
rect -6064 9647 -6035 9821
rect -6139 9634 -6035 9647
rect -5955 9821 -5867 9834
rect -5955 9647 -5926 9821
rect -5880 9647 -5867 9821
rect -5955 9634 -5867 9647
rect -3935 9820 -3847 9833
rect -3935 9646 -3922 9820
rect -3876 9646 -3847 9820
rect -3935 9633 -3847 9646
rect -3767 9820 -3663 9833
rect -3767 9646 -3738 9820
rect -3692 9646 -3663 9820
rect -3767 9633 -3663 9646
rect -3583 9820 -3479 9833
rect -3583 9646 -3554 9820
rect -3508 9646 -3479 9820
rect -3583 9633 -3479 9646
rect -3399 9820 -3311 9833
rect -3399 9646 -3370 9820
rect -3324 9646 -3311 9820
rect -3399 9633 -3311 9646
rect -2449 9821 -2361 9834
rect -2449 9647 -2436 9821
rect -2390 9647 -2361 9821
rect -2449 9634 -2361 9647
rect -2281 9821 -2177 9834
rect -2281 9647 -2252 9821
rect -2206 9647 -2177 9821
rect -2281 9634 -2177 9647
rect -2097 9821 -1993 9834
rect -2097 9647 -2068 9821
rect -2022 9647 -1993 9821
rect -2097 9634 -1993 9647
rect -1913 9821 -1825 9834
rect -1913 9647 -1884 9821
rect -1838 9647 -1825 9821
rect -1913 9634 -1825 9647
rect 107 9820 195 9833
rect 107 9646 120 9820
rect 166 9646 195 9820
rect 107 9633 195 9646
rect 275 9820 379 9833
rect 275 9646 304 9820
rect 350 9646 379 9820
rect 275 9633 379 9646
rect 459 9820 563 9833
rect 459 9646 488 9820
rect 534 9646 563 9820
rect 459 9633 563 9646
rect 643 9820 731 9833
rect 643 9646 672 9820
rect 718 9646 731 9820
rect 643 9633 731 9646
rect 1593 9821 1681 9834
rect 1593 9647 1606 9821
rect 1652 9647 1681 9821
rect 1593 9634 1681 9647
rect 1761 9821 1865 9834
rect 1761 9647 1790 9821
rect 1836 9647 1865 9821
rect 1761 9634 1865 9647
rect 1945 9821 2049 9834
rect 1945 9647 1974 9821
rect 2020 9647 2049 9821
rect 1945 9634 2049 9647
rect 2129 9821 2217 9834
rect 2129 9647 2158 9821
rect 2204 9647 2217 9821
rect 2129 9634 2217 9647
rect 4149 9820 4237 9833
rect 4149 9646 4162 9820
rect 4208 9646 4237 9820
rect 4149 9633 4237 9646
rect 4317 9820 4421 9833
rect 4317 9646 4346 9820
rect 4392 9646 4421 9820
rect 4317 9633 4421 9646
rect 4501 9820 4605 9833
rect 4501 9646 4530 9820
rect 4576 9646 4605 9820
rect 4501 9633 4605 9646
rect 4685 9820 4773 9833
rect 4685 9646 4714 9820
rect 4760 9646 4773 9820
rect 4685 9633 4773 9646
rect 5635 9821 5723 9834
rect 5635 9647 5648 9821
rect 5694 9647 5723 9821
rect 5635 9634 5723 9647
rect 5803 9821 5907 9834
rect 5803 9647 5832 9821
rect 5878 9647 5907 9821
rect 5803 9634 5907 9647
rect 5987 9821 6091 9834
rect 5987 9647 6016 9821
rect 6062 9647 6091 9821
rect 5987 9634 6091 9647
rect 6171 9821 6259 9834
rect 6171 9647 6200 9821
rect 6246 9647 6259 9821
rect 6171 9634 6259 9647
rect 8191 9820 8279 9833
rect 8191 9646 8204 9820
rect 8250 9646 8279 9820
rect 8191 9633 8279 9646
rect 8359 9820 8463 9833
rect 8359 9646 8388 9820
rect 8434 9646 8463 9820
rect 8359 9633 8463 9646
rect 8543 9820 8647 9833
rect 8543 9646 8572 9820
rect 8618 9646 8647 9820
rect 8543 9633 8647 9646
rect 8727 9820 8815 9833
rect 8727 9646 8756 9820
rect 8802 9646 8815 9820
rect 8727 9633 8815 9646
rect 9677 9821 9765 9834
rect 9677 9647 9690 9821
rect 9736 9647 9765 9821
rect 9677 9634 9765 9647
rect 9845 9821 9949 9834
rect 9845 9647 9874 9821
rect 9920 9647 9949 9821
rect 9845 9634 9949 9647
rect 10029 9821 10133 9834
rect 10029 9647 10058 9821
rect 10104 9647 10133 9821
rect 10029 9634 10133 9647
rect 10213 9821 10301 9834
rect 10213 9647 10242 9821
rect 10288 9647 10301 9821
rect 10213 9634 10301 9647
rect 12233 9820 12321 9833
rect 12233 9646 12246 9820
rect 12292 9646 12321 9820
rect 12233 9633 12321 9646
rect 12401 9820 12505 9833
rect 12401 9646 12430 9820
rect 12476 9646 12505 9820
rect 12401 9633 12505 9646
rect 12585 9820 12689 9833
rect 12585 9646 12614 9820
rect 12660 9646 12689 9820
rect 12585 9633 12689 9646
rect 12769 9820 12857 9833
rect 12769 9646 12798 9820
rect 12844 9646 12857 9820
rect 12769 9633 12857 9646
rect 13719 9821 13807 9834
rect 13719 9647 13732 9821
rect 13778 9647 13807 9821
rect 13719 9634 13807 9647
rect 13887 9821 13991 9834
rect 13887 9647 13916 9821
rect 13962 9647 13991 9821
rect 13887 9634 13991 9647
rect 14071 9821 14175 9834
rect 14071 9647 14100 9821
rect 14146 9647 14175 9821
rect 14071 9634 14175 9647
rect 14255 9821 14343 9834
rect 14255 9647 14284 9821
rect 14330 9647 14343 9821
rect 14255 9634 14343 9647
rect -11989 7615 -11901 7628
rect -11989 7441 -11976 7615
rect -11930 7441 -11901 7615
rect -11989 7428 -11901 7441
rect -11821 7615 -11717 7628
rect -11821 7441 -11792 7615
rect -11746 7441 -11717 7615
rect -11821 7428 -11717 7441
rect -11637 7615 -11533 7628
rect -11637 7441 -11608 7615
rect -11562 7441 -11533 7615
rect -11637 7428 -11533 7441
rect -11453 7615 -11365 7628
rect -11453 7441 -11424 7615
rect -11378 7441 -11365 7615
rect -11453 7428 -11365 7441
rect -7977 7615 -7889 7628
rect -7977 7441 -7964 7615
rect -7918 7441 -7889 7615
rect -7977 7428 -7889 7441
rect -7809 7615 -7705 7628
rect -7809 7441 -7780 7615
rect -7734 7441 -7705 7615
rect -7809 7428 -7705 7441
rect -7625 7615 -7521 7628
rect -7625 7441 -7596 7615
rect -7550 7441 -7521 7615
rect -7625 7428 -7521 7441
rect -7441 7615 -7353 7628
rect -7441 7441 -7412 7615
rect -7366 7441 -7353 7615
rect -7441 7428 -7353 7441
rect -3935 7615 -3847 7628
rect -3935 7441 -3922 7615
rect -3876 7441 -3847 7615
rect -3935 7428 -3847 7441
rect -3767 7615 -3663 7628
rect -3767 7441 -3738 7615
rect -3692 7441 -3663 7615
rect -3767 7428 -3663 7441
rect -3583 7615 -3479 7628
rect -3583 7441 -3554 7615
rect -3508 7441 -3479 7615
rect -3583 7428 -3479 7441
rect -3399 7615 -3311 7628
rect -3399 7441 -3370 7615
rect -3324 7441 -3311 7615
rect -3399 7428 -3311 7441
rect 107 7615 195 7628
rect 107 7441 120 7615
rect 166 7441 195 7615
rect 107 7428 195 7441
rect 275 7615 379 7628
rect 275 7441 304 7615
rect 350 7441 379 7615
rect 275 7428 379 7441
rect 459 7615 563 7628
rect 459 7441 488 7615
rect 534 7441 563 7615
rect 459 7428 563 7441
rect 643 7615 731 7628
rect 643 7441 672 7615
rect 718 7441 731 7615
rect 643 7428 731 7441
rect 4149 7615 4237 7628
rect 4149 7441 4162 7615
rect 4208 7441 4237 7615
rect 4149 7428 4237 7441
rect 4317 7615 4421 7628
rect 4317 7441 4346 7615
rect 4392 7441 4421 7615
rect 4317 7428 4421 7441
rect 4501 7615 4605 7628
rect 4501 7441 4530 7615
rect 4576 7441 4605 7615
rect 4501 7428 4605 7441
rect 4685 7615 4773 7628
rect 4685 7441 4714 7615
rect 4760 7441 4773 7615
rect 4685 7428 4773 7441
rect 8191 7615 8279 7628
rect 8191 7441 8204 7615
rect 8250 7441 8279 7615
rect 8191 7428 8279 7441
rect 8359 7615 8463 7628
rect 8359 7441 8388 7615
rect 8434 7441 8463 7615
rect 8359 7428 8463 7441
rect 8543 7615 8647 7628
rect 8543 7441 8572 7615
rect 8618 7441 8647 7615
rect 8543 7428 8647 7441
rect 8727 7615 8815 7628
rect 8727 7441 8756 7615
rect 8802 7441 8815 7615
rect 8727 7428 8815 7441
rect 12233 7615 12321 7628
rect 12233 7441 12246 7615
rect 12292 7441 12321 7615
rect 12233 7428 12321 7441
rect 12401 7615 12505 7628
rect 12401 7441 12430 7615
rect 12476 7441 12505 7615
rect 12401 7428 12505 7441
rect 12585 7615 12689 7628
rect 12585 7441 12614 7615
rect 12660 7441 12689 7615
rect 12585 7428 12689 7441
rect 12769 7615 12857 7628
rect 12769 7441 12798 7615
rect 12844 7441 12857 7615
rect 12769 7428 12857 7441
rect -10931 4478 -10831 4540
rect -10931 4432 -10909 4478
rect -10863 4432 -10831 4478
rect -10931 4370 -10831 4432
rect -10771 4478 -10661 4540
rect -10771 4432 -10739 4478
rect -10693 4432 -10661 4478
rect -10771 4370 -10661 4432
rect -10601 4478 -10491 4540
rect -10601 4432 -10569 4478
rect -10523 4432 -10491 4478
rect -10601 4370 -10491 4432
rect -10431 4478 -10321 4540
rect -10431 4432 -10399 4478
rect -10353 4432 -10321 4478
rect -10431 4370 -10321 4432
rect -10261 4478 -10151 4540
rect -10261 4432 -10229 4478
rect -10183 4432 -10151 4478
rect -10261 4370 -10151 4432
rect -10091 4478 -9991 4540
rect -10091 4432 -10059 4478
rect -10013 4432 -9991 4478
rect -10091 4370 -9991 4432
rect -8519 4034 -8431 4047
rect -8519 3860 -8506 4034
rect -8460 3860 -8431 4034
rect -8519 3847 -8431 3860
rect -8351 4034 -8263 4047
rect -8351 3860 -8322 4034
rect -8276 3860 -8263 4034
rect -8351 3847 -8263 3860
rect -8059 4034 -7971 4047
rect -8059 3860 -8046 4034
rect -8000 3860 -7971 4034
rect -8059 3847 -7971 3860
rect -7891 4034 -7803 4047
rect -7891 3860 -7862 4034
rect -7816 3860 -7803 4034
rect -7891 3847 -7803 3860
rect -9489 3101 -9401 3114
rect -9489 2727 -9476 3101
rect -9430 2727 -9401 3101
rect -9489 2714 -9401 2727
rect -9321 3101 -9233 3114
rect -9321 2727 -9292 3101
rect -9246 2727 -9233 3101
rect -9321 2714 -9233 2727
rect -7089 3101 -7001 3114
rect -7089 2727 -7076 3101
rect -7030 2727 -7001 3101
rect -7089 2714 -7001 2727
rect -6921 3101 -6833 3114
rect -6921 2727 -6892 3101
rect -6846 2727 -6833 3101
rect -6921 2714 -6833 2727
rect -9855 728 -9767 741
rect -9855 354 -9842 728
rect -9796 354 -9767 728
rect -9855 341 -9767 354
rect -9567 728 -9463 741
rect -9567 354 -9538 728
rect -9492 354 -9463 728
rect -9567 341 -9463 354
rect -9263 728 -9159 741
rect -9263 354 -9234 728
rect -9188 354 -9159 728
rect -9263 341 -9159 354
rect -8959 728 -8855 741
rect -8959 354 -8930 728
rect -8884 354 -8855 728
rect -8959 341 -8855 354
rect -8655 728 -8551 741
rect -8655 354 -8626 728
rect -8580 354 -8551 728
rect -8655 341 -8551 354
rect -8351 728 -8263 741
rect -8351 354 -8322 728
rect -8276 354 -8263 728
rect -8351 341 -8263 354
rect -8059 728 -7971 741
rect -8059 354 -8046 728
rect -8000 354 -7971 728
rect -8059 341 -7971 354
rect -7771 728 -7667 741
rect -7771 354 -7742 728
rect -7696 354 -7667 728
rect -7771 341 -7667 354
rect -7467 728 -7363 741
rect -7467 354 -7438 728
rect -7392 354 -7363 728
rect -7467 341 -7363 354
rect -7163 728 -7059 741
rect -7163 354 -7134 728
rect -7088 354 -7059 728
rect -7163 341 -7059 354
rect -6859 728 -6755 741
rect -6859 354 -6830 728
rect -6784 354 -6755 728
rect -6859 341 -6755 354
rect -6555 728 -6467 741
rect -6555 354 -6526 728
rect -6480 354 -6467 728
rect -6555 341 -6467 354
rect -10021 -757 -9933 -744
rect -10021 -1031 -10008 -757
rect -9962 -1031 -9933 -757
rect -10021 -1044 -9933 -1031
rect -9733 -757 -9629 -744
rect -9733 -1031 -9704 -757
rect -9658 -1031 -9629 -757
rect -9733 -1044 -9629 -1031
rect -9429 -757 -9325 -744
rect -9429 -1031 -9400 -757
rect -9354 -1031 -9325 -757
rect -9429 -1044 -9325 -1031
rect -9125 -757 -9021 -744
rect -9125 -1031 -9096 -757
rect -9050 -1031 -9021 -757
rect -9125 -1044 -9021 -1031
rect -8821 -757 -8717 -744
rect -8821 -1031 -8792 -757
rect -8746 -1031 -8717 -757
rect -8821 -1044 -8717 -1031
rect -8517 -757 -8413 -744
rect -8517 -1031 -8488 -757
rect -8442 -1031 -8413 -757
rect -8517 -1044 -8413 -1031
rect -8213 -757 -8109 -744
rect -8213 -1031 -8184 -757
rect -8138 -1031 -8109 -757
rect -8213 -1044 -8109 -1031
rect -7909 -757 -7805 -744
rect -7909 -1031 -7880 -757
rect -7834 -1031 -7805 -757
rect -7909 -1044 -7805 -1031
rect -7605 -757 -7501 -744
rect -7605 -1031 -7576 -757
rect -7530 -1031 -7501 -757
rect -7605 -1044 -7501 -1031
rect -7301 -757 -7197 -744
rect -7301 -1031 -7272 -757
rect -7226 -1031 -7197 -757
rect -7301 -1044 -7197 -1031
rect -6997 -757 -6893 -744
rect -6997 -1031 -6968 -757
rect -6922 -1031 -6893 -757
rect -6997 -1044 -6893 -1031
rect -6693 -757 -6589 -744
rect -6693 -1031 -6664 -757
rect -6618 -1031 -6589 -757
rect -6693 -1044 -6589 -1031
rect -6389 -757 -6301 -744
rect -6389 -1031 -6360 -757
rect -6314 -1031 -6301 -757
rect -6389 -1044 -6301 -1031
rect -10021 -1720 -9933 -1707
rect -10021 -1994 -10008 -1720
rect -9962 -1994 -9933 -1720
rect -10021 -2007 -9933 -1994
rect -9733 -1720 -9629 -1707
rect -9733 -1994 -9704 -1720
rect -9658 -1994 -9629 -1720
rect -9733 -2007 -9629 -1994
rect -9429 -1720 -9325 -1707
rect -9429 -1994 -9400 -1720
rect -9354 -1994 -9325 -1720
rect -9429 -2007 -9325 -1994
rect -9125 -1720 -9021 -1707
rect -9125 -1994 -9096 -1720
rect -9050 -1994 -9021 -1720
rect -9125 -2007 -9021 -1994
rect -8821 -1720 -8717 -1707
rect -8821 -1994 -8792 -1720
rect -8746 -1994 -8717 -1720
rect -8821 -2007 -8717 -1994
rect -8517 -1720 -8413 -1707
rect -8517 -1994 -8488 -1720
rect -8442 -1994 -8413 -1720
rect -8517 -2007 -8413 -1994
rect -8213 -1720 -8109 -1707
rect -8213 -1994 -8184 -1720
rect -8138 -1994 -8109 -1720
rect -8213 -2007 -8109 -1994
rect -7909 -1720 -7805 -1707
rect -7909 -1994 -7880 -1720
rect -7834 -1994 -7805 -1720
rect -7909 -2007 -7805 -1994
rect -7605 -1720 -7501 -1707
rect -7605 -1994 -7576 -1720
rect -7530 -1994 -7501 -1720
rect -7605 -2007 -7501 -1994
rect -7301 -1720 -7197 -1707
rect -7301 -1994 -7272 -1720
rect -7226 -1994 -7197 -1720
rect -7301 -2007 -7197 -1994
rect -6997 -1720 -6893 -1707
rect -6997 -1994 -6968 -1720
rect -6922 -1994 -6893 -1720
rect -6997 -2007 -6893 -1994
rect -6693 -1720 -6589 -1707
rect -6693 -1994 -6664 -1720
rect -6618 -1994 -6589 -1720
rect -6693 -2007 -6589 -1994
rect -6389 -1720 -6301 -1707
rect -6389 -1994 -6360 -1720
rect -6314 -1994 -6301 -1720
rect -6389 -2007 -6301 -1994
rect -8473 -2646 -8385 -2633
rect -8473 -2780 -8460 -2646
rect -8414 -2780 -8385 -2646
rect -8473 -2793 -8385 -2780
rect -8305 -2646 -8201 -2633
rect -8305 -2780 -8276 -2646
rect -8230 -2780 -8201 -2646
rect -8305 -2793 -8201 -2780
rect -8121 -2646 -8017 -2633
rect -8121 -2780 -8092 -2646
rect -8046 -2780 -8017 -2646
rect -8121 -2793 -8017 -2780
rect -7937 -2646 -7849 -2633
rect -7937 -2780 -7908 -2646
rect -7862 -2780 -7849 -2646
rect -7937 -2793 -7849 -2780
<< pdiff >>
rect 39951 38830 40051 38883
rect 39951 38596 39973 38830
rect 40019 38596 40051 38830
rect 39951 38543 40051 38596
rect 40111 38855 40221 38883
rect 40111 38621 40143 38855
rect 40189 38621 40221 38855
rect 40111 38543 40221 38621
rect 40281 38830 40391 38883
rect 40281 38596 40313 38830
rect 40359 38596 40391 38830
rect 40281 38543 40391 38596
rect 40451 38855 40561 38883
rect 40451 38621 40483 38855
rect 40529 38621 40561 38855
rect 40451 38543 40561 38621
rect 40621 38830 40731 38883
rect 40621 38596 40653 38830
rect 40699 38596 40731 38830
rect 40621 38543 40731 38596
rect 40791 38830 40891 38883
rect 40791 38596 40823 38830
rect 40869 38596 40891 38830
rect 40791 38543 40891 38596
rect -4719 37271 -4631 37284
rect -4719 36797 -4706 37271
rect -4660 36797 -4631 37271
rect -4719 36784 -4631 36797
rect -4551 37271 -4447 37284
rect -4551 36797 -4522 37271
rect -4476 36797 -4447 37271
rect -4551 36784 -4447 36797
rect -4367 37271 -4263 37284
rect -4367 36797 -4338 37271
rect -4292 36797 -4263 37271
rect -4367 36784 -4263 36797
rect -4183 37271 -4095 37284
rect -4183 36797 -4154 37271
rect -4108 36797 -4095 37271
rect -4183 36784 -4095 36797
rect 4753 37271 4841 37284
rect 4753 36797 4766 37271
rect 4812 36797 4841 37271
rect 4753 36784 4841 36797
rect 4921 37271 5025 37284
rect 4921 36797 4950 37271
rect 4996 36797 5025 37271
rect 4921 36784 5025 36797
rect 5105 37271 5209 37284
rect 5105 36797 5134 37271
rect 5180 36797 5209 37271
rect 5105 36784 5209 36797
rect 5289 37271 5377 37284
rect 5289 36797 5318 37271
rect 5364 36797 5377 37271
rect 5289 36784 5377 36797
rect 14225 37272 14313 37285
rect 14225 36798 14238 37272
rect 14284 36798 14313 37272
rect 14225 36785 14313 36798
rect 14393 37272 14497 37285
rect 14393 36798 14422 37272
rect 14468 36798 14497 37272
rect 14393 36785 14497 36798
rect 14577 37272 14681 37285
rect 14577 36798 14606 37272
rect 14652 36798 14681 37272
rect 14577 36785 14681 36798
rect 14761 37272 14849 37285
rect 14761 36798 14790 37272
rect 14836 36798 14849 37272
rect 14761 36785 14849 36798
rect 23697 37272 23785 37285
rect 23697 36798 23710 37272
rect 23756 36798 23785 37272
rect 23697 36785 23785 36798
rect 23865 37272 23969 37285
rect 23865 36798 23894 37272
rect 23940 36798 23969 37272
rect 23865 36785 23969 36798
rect 24049 37272 24153 37285
rect 24049 36798 24078 37272
rect 24124 36798 24153 37272
rect 24049 36785 24153 36798
rect 24233 37272 24321 37285
rect 24233 36798 24262 37272
rect 24308 36798 24321 37272
rect 24233 36785 24321 36798
rect 33169 37272 33257 37285
rect 33169 36798 33182 37272
rect 33228 36798 33257 37272
rect 33169 36785 33257 36798
rect 33337 37272 33441 37285
rect 33337 36798 33366 37272
rect 33412 36798 33441 37272
rect 33337 36785 33441 36798
rect 33521 37272 33625 37285
rect 33521 36798 33550 37272
rect 33596 36798 33625 37272
rect 33521 36785 33625 36798
rect 33705 37272 33793 37285
rect 33705 36798 33734 37272
rect 33780 36798 33793 37272
rect 33705 36785 33793 36798
rect 42641 37272 42729 37285
rect 42641 36798 42654 37272
rect 42700 36798 42729 37272
rect 42641 36785 42729 36798
rect 42809 37272 42913 37285
rect 42809 36798 42838 37272
rect 42884 36798 42913 37272
rect 42809 36785 42913 36798
rect 42993 37272 43097 37285
rect 42993 36798 43022 37272
rect 43068 36798 43097 37272
rect 42993 36785 43097 36798
rect 43177 37272 43265 37285
rect 43177 36798 43206 37272
rect 43252 36798 43265 37272
rect 43177 36785 43265 36798
rect -4719 35066 -4631 35079
rect -4719 34592 -4706 35066
rect -4660 34592 -4631 35066
rect -4719 34579 -4631 34592
rect -4551 35066 -4447 35079
rect -4551 34592 -4522 35066
rect -4476 34592 -4447 35066
rect -4551 34579 -4447 34592
rect -4367 35066 -4263 35079
rect -4367 34592 -4338 35066
rect -4292 34592 -4263 35066
rect -4367 34579 -4263 34592
rect -4183 35066 -4095 35079
rect -4183 34592 -4154 35066
rect -4108 34592 -4095 35066
rect -4183 34579 -4095 34592
rect -3233 35066 -3145 35079
rect -3233 34592 -3220 35066
rect -3174 34592 -3145 35066
rect -3233 34579 -3145 34592
rect -3065 35066 -2961 35079
rect -3065 34592 -3036 35066
rect -2990 34592 -2961 35066
rect -3065 34579 -2961 34592
rect -2881 35066 -2777 35079
rect -2881 34592 -2852 35066
rect -2806 34592 -2777 35066
rect -2881 34579 -2777 34592
rect -2697 35066 -2609 35079
rect -2697 34592 -2668 35066
rect -2622 34592 -2609 35066
rect -2697 34579 -2609 34592
rect 4753 35066 4841 35079
rect 4753 34592 4766 35066
rect 4812 34592 4841 35066
rect 4753 34579 4841 34592
rect 4921 35066 5025 35079
rect 4921 34592 4950 35066
rect 4996 34592 5025 35066
rect 4921 34579 5025 34592
rect 5105 35066 5209 35079
rect 5105 34592 5134 35066
rect 5180 34592 5209 35066
rect 5105 34579 5209 34592
rect 5289 35066 5377 35079
rect 5289 34592 5318 35066
rect 5364 34592 5377 35066
rect 5289 34579 5377 34592
rect 6239 35066 6327 35079
rect 6239 34592 6252 35066
rect 6298 34592 6327 35066
rect 6239 34579 6327 34592
rect 6407 35066 6511 35079
rect 6407 34592 6436 35066
rect 6482 34592 6511 35066
rect 6407 34579 6511 34592
rect 6591 35066 6695 35079
rect 6591 34592 6620 35066
rect 6666 34592 6695 35066
rect 6591 34579 6695 34592
rect 6775 35066 6863 35079
rect 6775 34592 6804 35066
rect 6850 34592 6863 35066
rect 6775 34579 6863 34592
rect 14225 35067 14313 35080
rect 14225 34593 14238 35067
rect 14284 34593 14313 35067
rect 14225 34580 14313 34593
rect 14393 35067 14497 35080
rect 14393 34593 14422 35067
rect 14468 34593 14497 35067
rect 14393 34580 14497 34593
rect 14577 35067 14681 35080
rect 14577 34593 14606 35067
rect 14652 34593 14681 35067
rect 14577 34580 14681 34593
rect 14761 35067 14849 35080
rect 14761 34593 14790 35067
rect 14836 34593 14849 35067
rect 14761 34580 14849 34593
rect 15711 35067 15799 35080
rect 15711 34593 15724 35067
rect 15770 34593 15799 35067
rect 15711 34580 15799 34593
rect 15879 35067 15983 35080
rect 15879 34593 15908 35067
rect 15954 34593 15983 35067
rect 15879 34580 15983 34593
rect 16063 35067 16167 35080
rect 16063 34593 16092 35067
rect 16138 34593 16167 35067
rect 16063 34580 16167 34593
rect 16247 35067 16335 35080
rect 16247 34593 16276 35067
rect 16322 34593 16335 35067
rect 16247 34580 16335 34593
rect 23697 35067 23785 35080
rect 23697 34593 23710 35067
rect 23756 34593 23785 35067
rect 23697 34580 23785 34593
rect 23865 35067 23969 35080
rect 23865 34593 23894 35067
rect 23940 34593 23969 35067
rect 23865 34580 23969 34593
rect 24049 35067 24153 35080
rect 24049 34593 24078 35067
rect 24124 34593 24153 35067
rect 24049 34580 24153 34593
rect 24233 35067 24321 35080
rect 24233 34593 24262 35067
rect 24308 34593 24321 35067
rect 24233 34580 24321 34593
rect 25183 35067 25271 35080
rect 25183 34593 25196 35067
rect 25242 34593 25271 35067
rect 25183 34580 25271 34593
rect 25351 35067 25455 35080
rect 25351 34593 25380 35067
rect 25426 34593 25455 35067
rect 25351 34580 25455 34593
rect 25535 35067 25639 35080
rect 25535 34593 25564 35067
rect 25610 34593 25639 35067
rect 25535 34580 25639 34593
rect 25719 35067 25807 35080
rect 25719 34593 25748 35067
rect 25794 34593 25807 35067
rect 25719 34580 25807 34593
rect 33169 35067 33257 35080
rect 33169 34593 33182 35067
rect 33228 34593 33257 35067
rect 33169 34580 33257 34593
rect 33337 35067 33441 35080
rect 33337 34593 33366 35067
rect 33412 34593 33441 35067
rect 33337 34580 33441 34593
rect 33521 35067 33625 35080
rect 33521 34593 33550 35067
rect 33596 34593 33625 35067
rect 33521 34580 33625 34593
rect 33705 35067 33793 35080
rect 33705 34593 33734 35067
rect 33780 34593 33793 35067
rect 33705 34580 33793 34593
rect 34655 35067 34743 35080
rect 34655 34593 34668 35067
rect 34714 34593 34743 35067
rect 34655 34580 34743 34593
rect 34823 35067 34927 35080
rect 34823 34593 34852 35067
rect 34898 34593 34927 35067
rect 34823 34580 34927 34593
rect 35007 35067 35111 35080
rect 35007 34593 35036 35067
rect 35082 34593 35111 35067
rect 35007 34580 35111 34593
rect 35191 35067 35279 35080
rect 35191 34593 35220 35067
rect 35266 34593 35279 35067
rect 35191 34580 35279 34593
rect 42641 35067 42729 35080
rect 42641 34593 42654 35067
rect 42700 34593 42729 35067
rect 42641 34580 42729 34593
rect 42809 35067 42913 35080
rect 42809 34593 42838 35067
rect 42884 34593 42913 35067
rect 42809 34580 42913 34593
rect 42993 35067 43097 35080
rect 42993 34593 43022 35067
rect 43068 34593 43097 35067
rect 42993 34580 43097 34593
rect 43177 35067 43265 35080
rect 43177 34593 43206 35067
rect 43252 34593 43265 35067
rect 43177 34580 43265 34593
rect 44127 35067 44215 35080
rect 44127 34593 44140 35067
rect 44186 34593 44215 35067
rect 44127 34580 44215 34593
rect 44295 35067 44399 35080
rect 44295 34593 44324 35067
rect 44370 34593 44399 35067
rect 44295 34580 44399 34593
rect 44479 35067 44583 35080
rect 44479 34593 44508 35067
rect 44554 34593 44583 35067
rect 44479 34580 44583 34593
rect 44663 35067 44751 35080
rect 44663 34593 44692 35067
rect 44738 34593 44751 35067
rect 44663 34580 44751 34593
rect -4719 32861 -4631 32874
rect -4719 32387 -4706 32861
rect -4660 32387 -4631 32861
rect -4719 32374 -4631 32387
rect -4551 32861 -4447 32874
rect -4551 32387 -4522 32861
rect -4476 32387 -4447 32861
rect -4551 32374 -4447 32387
rect -4367 32861 -4263 32874
rect -4367 32387 -4338 32861
rect -4292 32387 -4263 32861
rect -4367 32374 -4263 32387
rect -4183 32861 -4095 32874
rect -4183 32387 -4154 32861
rect -4108 32387 -4095 32861
rect -4183 32374 -4095 32387
rect -3233 32862 -3145 32875
rect -3233 32388 -3220 32862
rect -3174 32388 -3145 32862
rect -3233 32375 -3145 32388
rect -3065 32862 -2961 32875
rect -3065 32388 -3036 32862
rect -2990 32388 -2961 32862
rect -3065 32375 -2961 32388
rect -2881 32862 -2777 32875
rect -2881 32388 -2852 32862
rect -2806 32388 -2777 32862
rect -2881 32375 -2777 32388
rect -2697 32862 -2609 32875
rect -2697 32388 -2668 32862
rect -2622 32388 -2609 32862
rect -2697 32375 -2609 32388
rect 4753 32861 4841 32874
rect 4753 32387 4766 32861
rect 4812 32387 4841 32861
rect 4753 32374 4841 32387
rect 4921 32861 5025 32874
rect 4921 32387 4950 32861
rect 4996 32387 5025 32861
rect 4921 32374 5025 32387
rect 5105 32861 5209 32874
rect 5105 32387 5134 32861
rect 5180 32387 5209 32861
rect 5105 32374 5209 32387
rect 5289 32861 5377 32874
rect 5289 32387 5318 32861
rect 5364 32387 5377 32861
rect 5289 32374 5377 32387
rect 6239 32862 6327 32875
rect 6239 32388 6252 32862
rect 6298 32388 6327 32862
rect 6239 32375 6327 32388
rect 6407 32862 6511 32875
rect 6407 32388 6436 32862
rect 6482 32388 6511 32862
rect 6407 32375 6511 32388
rect 6591 32862 6695 32875
rect 6591 32388 6620 32862
rect 6666 32388 6695 32862
rect 6591 32375 6695 32388
rect 6775 32862 6863 32875
rect 6775 32388 6804 32862
rect 6850 32388 6863 32862
rect 6775 32375 6863 32388
rect 14225 32862 14313 32875
rect 14225 32388 14238 32862
rect 14284 32388 14313 32862
rect 14225 32375 14313 32388
rect 14393 32862 14497 32875
rect 14393 32388 14422 32862
rect 14468 32388 14497 32862
rect 14393 32375 14497 32388
rect 14577 32862 14681 32875
rect 14577 32388 14606 32862
rect 14652 32388 14681 32862
rect 14577 32375 14681 32388
rect 14761 32862 14849 32875
rect 14761 32388 14790 32862
rect 14836 32388 14849 32862
rect 14761 32375 14849 32388
rect 15711 32863 15799 32876
rect 15711 32389 15724 32863
rect 15770 32389 15799 32863
rect 15711 32376 15799 32389
rect 15879 32863 15983 32876
rect 15879 32389 15908 32863
rect 15954 32389 15983 32863
rect 15879 32376 15983 32389
rect 16063 32863 16167 32876
rect 16063 32389 16092 32863
rect 16138 32389 16167 32863
rect 16063 32376 16167 32389
rect 16247 32863 16335 32876
rect 16247 32389 16276 32863
rect 16322 32389 16335 32863
rect 16247 32376 16335 32389
rect 23697 32862 23785 32875
rect 23697 32388 23710 32862
rect 23756 32388 23785 32862
rect 23697 32375 23785 32388
rect 23865 32862 23969 32875
rect 23865 32388 23894 32862
rect 23940 32388 23969 32862
rect 23865 32375 23969 32388
rect 24049 32862 24153 32875
rect 24049 32388 24078 32862
rect 24124 32388 24153 32862
rect 24049 32375 24153 32388
rect 24233 32862 24321 32875
rect 24233 32388 24262 32862
rect 24308 32388 24321 32862
rect 24233 32375 24321 32388
rect 25183 32863 25271 32876
rect 25183 32389 25196 32863
rect 25242 32389 25271 32863
rect 25183 32376 25271 32389
rect 25351 32863 25455 32876
rect 25351 32389 25380 32863
rect 25426 32389 25455 32863
rect 25351 32376 25455 32389
rect 25535 32863 25639 32876
rect 25535 32389 25564 32863
rect 25610 32389 25639 32863
rect 25535 32376 25639 32389
rect 25719 32863 25807 32876
rect 25719 32389 25748 32863
rect 25794 32389 25807 32863
rect 25719 32376 25807 32389
rect 33169 32862 33257 32875
rect 33169 32388 33182 32862
rect 33228 32388 33257 32862
rect 33169 32375 33257 32388
rect 33337 32862 33441 32875
rect 33337 32388 33366 32862
rect 33412 32388 33441 32862
rect 33337 32375 33441 32388
rect 33521 32862 33625 32875
rect 33521 32388 33550 32862
rect 33596 32388 33625 32862
rect 33521 32375 33625 32388
rect 33705 32862 33793 32875
rect 33705 32388 33734 32862
rect 33780 32388 33793 32862
rect 33705 32375 33793 32388
rect 34655 32863 34743 32876
rect 34655 32389 34668 32863
rect 34714 32389 34743 32863
rect 34655 32376 34743 32389
rect 34823 32863 34927 32876
rect 34823 32389 34852 32863
rect 34898 32389 34927 32863
rect 34823 32376 34927 32389
rect 35007 32863 35111 32876
rect 35007 32389 35036 32863
rect 35082 32389 35111 32863
rect 35007 32376 35111 32389
rect 35191 32863 35279 32876
rect 35191 32389 35220 32863
rect 35266 32389 35279 32863
rect 35191 32376 35279 32389
rect 42641 32862 42729 32875
rect 42641 32388 42654 32862
rect 42700 32388 42729 32862
rect 42641 32375 42729 32388
rect 42809 32862 42913 32875
rect 42809 32388 42838 32862
rect 42884 32388 42913 32862
rect 42809 32375 42913 32388
rect 42993 32862 43097 32875
rect 42993 32388 43022 32862
rect 43068 32388 43097 32862
rect 42993 32375 43097 32388
rect 43177 32862 43265 32875
rect 43177 32388 43206 32862
rect 43252 32388 43265 32862
rect 43177 32375 43265 32388
rect 44127 32863 44215 32876
rect 44127 32389 44140 32863
rect 44186 32389 44215 32863
rect 44127 32376 44215 32389
rect 44295 32863 44399 32876
rect 44295 32389 44324 32863
rect 44370 32389 44399 32863
rect 44295 32376 44399 32389
rect 44479 32863 44583 32876
rect 44479 32389 44508 32863
rect 44554 32389 44583 32863
rect 44479 32376 44583 32389
rect 44663 32863 44751 32876
rect 44663 32389 44692 32863
rect 44738 32389 44751 32863
rect 44663 32376 44751 32389
rect -9861 31746 -9773 31759
rect -9861 31172 -9848 31746
rect -9802 31172 -9773 31746
rect -9861 31159 -9773 31172
rect -9673 31746 -9585 31759
rect -9673 31172 -9644 31746
rect -9598 31172 -9585 31746
rect -9673 31159 -9585 31172
rect -8973 31746 -8885 31759
rect -8973 31172 -8960 31746
rect -8914 31172 -8885 31746
rect -8973 31159 -8885 31172
rect -8785 31746 -8697 31759
rect -8785 31172 -8756 31746
rect -8710 31172 -8697 31746
rect -8785 31159 -8697 31172
rect -8493 31746 -8405 31759
rect -8493 31172 -8480 31746
rect -8434 31172 -8405 31746
rect -8493 31159 -8405 31172
rect -8305 31746 -8217 31759
rect -8305 31172 -8276 31746
rect -8230 31172 -8217 31746
rect -8305 31159 -8217 31172
rect -389 31746 -301 31759
rect -389 31172 -376 31746
rect -330 31172 -301 31746
rect -389 31159 -301 31172
rect -201 31746 -113 31759
rect -201 31172 -172 31746
rect -126 31172 -113 31746
rect -201 31159 -113 31172
rect 499 31746 587 31759
rect 499 31172 512 31746
rect 558 31172 587 31746
rect 499 31159 587 31172
rect 687 31746 775 31759
rect 687 31172 716 31746
rect 762 31172 775 31746
rect 687 31159 775 31172
rect 979 31746 1067 31759
rect 979 31172 992 31746
rect 1038 31172 1067 31746
rect 979 31159 1067 31172
rect 1167 31746 1255 31759
rect 1167 31172 1196 31746
rect 1242 31172 1255 31746
rect 1167 31159 1255 31172
rect 9083 31747 9171 31760
rect 9083 31173 9096 31747
rect 9142 31173 9171 31747
rect 9083 31160 9171 31173
rect 9271 31747 9359 31760
rect 9271 31173 9300 31747
rect 9346 31173 9359 31747
rect 9271 31160 9359 31173
rect 9971 31747 10059 31760
rect 9971 31173 9984 31747
rect 10030 31173 10059 31747
rect 9971 31160 10059 31173
rect 10159 31747 10247 31760
rect 10159 31173 10188 31747
rect 10234 31173 10247 31747
rect 10159 31160 10247 31173
rect 10451 31747 10539 31760
rect 10451 31173 10464 31747
rect 10510 31173 10539 31747
rect 10451 31160 10539 31173
rect 10639 31747 10727 31760
rect 10639 31173 10668 31747
rect 10714 31173 10727 31747
rect 10639 31160 10727 31173
rect 18555 31747 18643 31760
rect 18555 31173 18568 31747
rect 18614 31173 18643 31747
rect 18555 31160 18643 31173
rect 18743 31747 18831 31760
rect 18743 31173 18772 31747
rect 18818 31173 18831 31747
rect 18743 31160 18831 31173
rect 19443 31747 19531 31760
rect 19443 31173 19456 31747
rect 19502 31173 19531 31747
rect 19443 31160 19531 31173
rect 19631 31747 19719 31760
rect 19631 31173 19660 31747
rect 19706 31173 19719 31747
rect 19631 31160 19719 31173
rect 19923 31747 20011 31760
rect 19923 31173 19936 31747
rect 19982 31173 20011 31747
rect 19923 31160 20011 31173
rect 20111 31747 20199 31760
rect 20111 31173 20140 31747
rect 20186 31173 20199 31747
rect 20111 31160 20199 31173
rect 28027 31747 28115 31760
rect 28027 31173 28040 31747
rect 28086 31173 28115 31747
rect 28027 31160 28115 31173
rect 28215 31747 28303 31760
rect 28215 31173 28244 31747
rect 28290 31173 28303 31747
rect 28215 31160 28303 31173
rect 28915 31747 29003 31760
rect 28915 31173 28928 31747
rect 28974 31173 29003 31747
rect 28915 31160 29003 31173
rect 29103 31747 29191 31760
rect 29103 31173 29132 31747
rect 29178 31173 29191 31747
rect 29103 31160 29191 31173
rect 29395 31747 29483 31760
rect 29395 31173 29408 31747
rect 29454 31173 29483 31747
rect 29395 31160 29483 31173
rect 29583 31747 29671 31760
rect 29583 31173 29612 31747
rect 29658 31173 29671 31747
rect 29583 31160 29671 31173
rect 37499 31747 37587 31760
rect 37499 31173 37512 31747
rect 37558 31173 37587 31747
rect 37499 31160 37587 31173
rect 37687 31747 37775 31760
rect 37687 31173 37716 31747
rect 37762 31173 37775 31747
rect 37687 31160 37775 31173
rect 38387 31747 38475 31760
rect 38387 31173 38400 31747
rect 38446 31173 38475 31747
rect 38387 31160 38475 31173
rect 38575 31747 38663 31760
rect 38575 31173 38604 31747
rect 38650 31173 38663 31747
rect 38575 31160 38663 31173
rect 38867 31747 38955 31760
rect 38867 31173 38880 31747
rect 38926 31173 38955 31747
rect 38867 31160 38955 31173
rect 39055 31747 39143 31760
rect 39055 31173 39084 31747
rect 39130 31173 39143 31747
rect 39055 31160 39143 31173
rect -10755 30326 -10667 30339
rect -10755 29752 -10742 30326
rect -10696 29752 -10667 30326
rect -10755 29739 -10667 29752
rect -10567 30326 -10479 30339
rect -10567 29752 -10538 30326
rect -10492 29752 -10479 30326
rect -10567 29739 -10479 29752
rect -7633 30570 -7545 30583
rect -7633 29996 -7620 30570
rect -7574 29996 -7545 30570
rect -7633 29983 -7545 29996
rect -7445 30570 -7341 30583
rect -7445 29996 -7416 30570
rect -7370 29996 -7341 30570
rect -7445 29983 -7341 29996
rect -7241 30570 -7153 30583
rect -7241 29996 -7212 30570
rect -7166 29996 -7153 30570
rect -7241 29983 -7153 29996
rect -6949 30570 -6861 30583
rect -6949 29996 -6936 30570
rect -6890 29996 -6861 30570
rect -6949 29983 -6861 29996
rect -6761 30570 -6657 30583
rect -6761 29996 -6732 30570
rect -6686 29996 -6657 30570
rect -6761 29983 -6657 29996
rect -6557 30570 -6469 30583
rect -6557 29996 -6528 30570
rect -6482 29996 -6469 30570
rect -6557 29983 -6469 29996
rect -6265 30570 -6177 30583
rect -6265 29996 -6252 30570
rect -6206 29996 -6177 30570
rect -6265 29983 -6177 29996
rect -6077 30570 -5989 30583
rect -6077 29996 -6048 30570
rect -6002 29996 -5989 30570
rect -6077 29983 -5989 29996
rect -4719 30656 -4631 30669
rect -4719 30182 -4706 30656
rect -4660 30182 -4631 30656
rect -4719 30169 -4631 30182
rect -4551 30656 -4447 30669
rect -4551 30182 -4522 30656
rect -4476 30182 -4447 30656
rect -4551 30169 -4447 30182
rect -4367 30656 -4263 30669
rect -4367 30182 -4338 30656
rect -4292 30182 -4263 30656
rect -4367 30169 -4263 30182
rect -4183 30656 -4095 30669
rect -4183 30182 -4154 30656
rect -4108 30182 -4095 30656
rect -4183 30169 -4095 30182
rect -9861 29406 -9773 29419
rect -9861 28832 -9848 29406
rect -9802 28832 -9773 29406
rect -9861 28819 -9773 28832
rect -9673 29406 -9585 29419
rect -9673 28832 -9644 29406
rect -9598 28832 -9585 29406
rect -9673 28819 -9585 28832
rect -8973 29406 -8885 29419
rect -8973 28832 -8960 29406
rect -8914 28832 -8885 29406
rect -8973 28819 -8885 28832
rect -8785 29406 -8697 29419
rect -8785 28832 -8756 29406
rect -8710 28832 -8697 29406
rect -8785 28819 -8697 28832
rect -8493 29406 -8405 29419
rect -8493 28832 -8480 29406
rect -8434 28832 -8405 29406
rect -8493 28819 -8405 28832
rect -8305 29406 -8217 29419
rect -8305 28832 -8276 29406
rect -8230 28832 -8217 29406
rect -8305 28819 -8217 28832
rect -1283 30326 -1195 30339
rect -1283 29752 -1270 30326
rect -1224 29752 -1195 30326
rect -1283 29739 -1195 29752
rect -1095 30326 -1007 30339
rect -1095 29752 -1066 30326
rect -1020 29752 -1007 30326
rect -1095 29739 -1007 29752
rect 1839 30570 1927 30583
rect 1839 29996 1852 30570
rect 1898 29996 1927 30570
rect 1839 29983 1927 29996
rect 2027 30570 2131 30583
rect 2027 29996 2056 30570
rect 2102 29996 2131 30570
rect 2027 29983 2131 29996
rect 2231 30570 2319 30583
rect 2231 29996 2260 30570
rect 2306 29996 2319 30570
rect 2231 29983 2319 29996
rect 2523 30570 2611 30583
rect 2523 29996 2536 30570
rect 2582 29996 2611 30570
rect 2523 29983 2611 29996
rect 2711 30570 2815 30583
rect 2711 29996 2740 30570
rect 2786 29996 2815 30570
rect 2711 29983 2815 29996
rect 2915 30570 3003 30583
rect 2915 29996 2944 30570
rect 2990 29996 3003 30570
rect 2915 29983 3003 29996
rect 3207 30570 3295 30583
rect 3207 29996 3220 30570
rect 3266 29996 3295 30570
rect 3207 29983 3295 29996
rect 3395 30570 3483 30583
rect 3395 29996 3424 30570
rect 3470 29996 3483 30570
rect 3395 29983 3483 29996
rect 4753 30656 4841 30669
rect 4753 30182 4766 30656
rect 4812 30182 4841 30656
rect 4753 30169 4841 30182
rect 4921 30656 5025 30669
rect 4921 30182 4950 30656
rect 4996 30182 5025 30656
rect 4921 30169 5025 30182
rect 5105 30656 5209 30669
rect 5105 30182 5134 30656
rect 5180 30182 5209 30656
rect 5105 30169 5209 30182
rect 5289 30656 5377 30669
rect 5289 30182 5318 30656
rect 5364 30182 5377 30656
rect 5289 30169 5377 30182
rect -389 29406 -301 29419
rect -389 28832 -376 29406
rect -330 28832 -301 29406
rect -389 28819 -301 28832
rect -201 29406 -113 29419
rect -201 28832 -172 29406
rect -126 28832 -113 29406
rect -201 28819 -113 28832
rect 499 29406 587 29419
rect 499 28832 512 29406
rect 558 28832 587 29406
rect 499 28819 587 28832
rect 687 29406 775 29419
rect 687 28832 716 29406
rect 762 28832 775 29406
rect 687 28819 775 28832
rect 979 29406 1067 29419
rect 979 28832 992 29406
rect 1038 28832 1067 29406
rect 979 28819 1067 28832
rect 1167 29406 1255 29419
rect 1167 28832 1196 29406
rect 1242 28832 1255 29406
rect 1167 28819 1255 28832
rect 8189 30327 8277 30340
rect 8189 29753 8202 30327
rect 8248 29753 8277 30327
rect 8189 29740 8277 29753
rect 8377 30327 8465 30340
rect 8377 29753 8406 30327
rect 8452 29753 8465 30327
rect 8377 29740 8465 29753
rect 11311 30571 11399 30584
rect 11311 29997 11324 30571
rect 11370 29997 11399 30571
rect 11311 29984 11399 29997
rect 11499 30571 11603 30584
rect 11499 29997 11528 30571
rect 11574 29997 11603 30571
rect 11499 29984 11603 29997
rect 11703 30571 11791 30584
rect 11703 29997 11732 30571
rect 11778 29997 11791 30571
rect 11703 29984 11791 29997
rect 11995 30571 12083 30584
rect 11995 29997 12008 30571
rect 12054 29997 12083 30571
rect 11995 29984 12083 29997
rect 12183 30571 12287 30584
rect 12183 29997 12212 30571
rect 12258 29997 12287 30571
rect 12183 29984 12287 29997
rect 12387 30571 12475 30584
rect 12387 29997 12416 30571
rect 12462 29997 12475 30571
rect 12387 29984 12475 29997
rect 12679 30571 12767 30584
rect 12679 29997 12692 30571
rect 12738 29997 12767 30571
rect 12679 29984 12767 29997
rect 12867 30571 12955 30584
rect 12867 29997 12896 30571
rect 12942 29997 12955 30571
rect 12867 29984 12955 29997
rect 14225 30657 14313 30670
rect 14225 30183 14238 30657
rect 14284 30183 14313 30657
rect 14225 30170 14313 30183
rect 14393 30657 14497 30670
rect 14393 30183 14422 30657
rect 14468 30183 14497 30657
rect 14393 30170 14497 30183
rect 14577 30657 14681 30670
rect 14577 30183 14606 30657
rect 14652 30183 14681 30657
rect 14577 30170 14681 30183
rect 14761 30657 14849 30670
rect 14761 30183 14790 30657
rect 14836 30183 14849 30657
rect 14761 30170 14849 30183
rect 9083 29407 9171 29420
rect 9083 28833 9096 29407
rect 9142 28833 9171 29407
rect 9083 28820 9171 28833
rect 9271 29407 9359 29420
rect 9271 28833 9300 29407
rect 9346 28833 9359 29407
rect 9271 28820 9359 28833
rect 9971 29407 10059 29420
rect 9971 28833 9984 29407
rect 10030 28833 10059 29407
rect 9971 28820 10059 28833
rect 10159 29407 10247 29420
rect 10159 28833 10188 29407
rect 10234 28833 10247 29407
rect 10159 28820 10247 28833
rect 10451 29407 10539 29420
rect 10451 28833 10464 29407
rect 10510 28833 10539 29407
rect 10451 28820 10539 28833
rect 10639 29407 10727 29420
rect 10639 28833 10668 29407
rect 10714 28833 10727 29407
rect 10639 28820 10727 28833
rect 17661 30327 17749 30340
rect 17661 29753 17674 30327
rect 17720 29753 17749 30327
rect 17661 29740 17749 29753
rect 17849 30327 17937 30340
rect 17849 29753 17878 30327
rect 17924 29753 17937 30327
rect 17849 29740 17937 29753
rect 20783 30571 20871 30584
rect 20783 29997 20796 30571
rect 20842 29997 20871 30571
rect 20783 29984 20871 29997
rect 20971 30571 21075 30584
rect 20971 29997 21000 30571
rect 21046 29997 21075 30571
rect 20971 29984 21075 29997
rect 21175 30571 21263 30584
rect 21175 29997 21204 30571
rect 21250 29997 21263 30571
rect 21175 29984 21263 29997
rect 21467 30571 21555 30584
rect 21467 29997 21480 30571
rect 21526 29997 21555 30571
rect 21467 29984 21555 29997
rect 21655 30571 21759 30584
rect 21655 29997 21684 30571
rect 21730 29997 21759 30571
rect 21655 29984 21759 29997
rect 21859 30571 21947 30584
rect 21859 29997 21888 30571
rect 21934 29997 21947 30571
rect 21859 29984 21947 29997
rect 22151 30571 22239 30584
rect 22151 29997 22164 30571
rect 22210 29997 22239 30571
rect 22151 29984 22239 29997
rect 22339 30571 22427 30584
rect 22339 29997 22368 30571
rect 22414 29997 22427 30571
rect 22339 29984 22427 29997
rect 23697 30657 23785 30670
rect 23697 30183 23710 30657
rect 23756 30183 23785 30657
rect 23697 30170 23785 30183
rect 23865 30657 23969 30670
rect 23865 30183 23894 30657
rect 23940 30183 23969 30657
rect 23865 30170 23969 30183
rect 24049 30657 24153 30670
rect 24049 30183 24078 30657
rect 24124 30183 24153 30657
rect 24049 30170 24153 30183
rect 24233 30657 24321 30670
rect 24233 30183 24262 30657
rect 24308 30183 24321 30657
rect 24233 30170 24321 30183
rect 18555 29407 18643 29420
rect 18555 28833 18568 29407
rect 18614 28833 18643 29407
rect 18555 28820 18643 28833
rect 18743 29407 18831 29420
rect 18743 28833 18772 29407
rect 18818 28833 18831 29407
rect 18743 28820 18831 28833
rect 19443 29407 19531 29420
rect 19443 28833 19456 29407
rect 19502 28833 19531 29407
rect 19443 28820 19531 28833
rect 19631 29407 19719 29420
rect 19631 28833 19660 29407
rect 19706 28833 19719 29407
rect 19631 28820 19719 28833
rect 19923 29407 20011 29420
rect 19923 28833 19936 29407
rect 19982 28833 20011 29407
rect 19923 28820 20011 28833
rect 20111 29407 20199 29420
rect 20111 28833 20140 29407
rect 20186 28833 20199 29407
rect 20111 28820 20199 28833
rect 27133 30327 27221 30340
rect 27133 29753 27146 30327
rect 27192 29753 27221 30327
rect 27133 29740 27221 29753
rect 27321 30327 27409 30340
rect 27321 29753 27350 30327
rect 27396 29753 27409 30327
rect 27321 29740 27409 29753
rect 30255 30571 30343 30584
rect 30255 29997 30268 30571
rect 30314 29997 30343 30571
rect 30255 29984 30343 29997
rect 30443 30571 30547 30584
rect 30443 29997 30472 30571
rect 30518 29997 30547 30571
rect 30443 29984 30547 29997
rect 30647 30571 30735 30584
rect 30647 29997 30676 30571
rect 30722 29997 30735 30571
rect 30647 29984 30735 29997
rect 30939 30571 31027 30584
rect 30939 29997 30952 30571
rect 30998 29997 31027 30571
rect 30939 29984 31027 29997
rect 31127 30571 31231 30584
rect 31127 29997 31156 30571
rect 31202 29997 31231 30571
rect 31127 29984 31231 29997
rect 31331 30571 31419 30584
rect 31331 29997 31360 30571
rect 31406 29997 31419 30571
rect 31331 29984 31419 29997
rect 31623 30571 31711 30584
rect 31623 29997 31636 30571
rect 31682 29997 31711 30571
rect 31623 29984 31711 29997
rect 31811 30571 31899 30584
rect 31811 29997 31840 30571
rect 31886 29997 31899 30571
rect 31811 29984 31899 29997
rect 33169 30657 33257 30670
rect 33169 30183 33182 30657
rect 33228 30183 33257 30657
rect 33169 30170 33257 30183
rect 33337 30657 33441 30670
rect 33337 30183 33366 30657
rect 33412 30183 33441 30657
rect 33337 30170 33441 30183
rect 33521 30657 33625 30670
rect 33521 30183 33550 30657
rect 33596 30183 33625 30657
rect 33521 30170 33625 30183
rect 33705 30657 33793 30670
rect 33705 30183 33734 30657
rect 33780 30183 33793 30657
rect 33705 30170 33793 30183
rect 28027 29407 28115 29420
rect 28027 28833 28040 29407
rect 28086 28833 28115 29407
rect 28027 28820 28115 28833
rect 28215 29407 28303 29420
rect 28215 28833 28244 29407
rect 28290 28833 28303 29407
rect 28215 28820 28303 28833
rect 28915 29407 29003 29420
rect 28915 28833 28928 29407
rect 28974 28833 29003 29407
rect 28915 28820 29003 28833
rect 29103 29407 29191 29420
rect 29103 28833 29132 29407
rect 29178 28833 29191 29407
rect 29103 28820 29191 28833
rect 29395 29407 29483 29420
rect 29395 28833 29408 29407
rect 29454 28833 29483 29407
rect 29395 28820 29483 28833
rect 29583 29407 29671 29420
rect 29583 28833 29612 29407
rect 29658 28833 29671 29407
rect 29583 28820 29671 28833
rect 36605 30327 36693 30340
rect 36605 29753 36618 30327
rect 36664 29753 36693 30327
rect 36605 29740 36693 29753
rect 36793 30327 36881 30340
rect 36793 29753 36822 30327
rect 36868 29753 36881 30327
rect 36793 29740 36881 29753
rect 39727 30571 39815 30584
rect 39727 29997 39740 30571
rect 39786 29997 39815 30571
rect 39727 29984 39815 29997
rect 39915 30571 40019 30584
rect 39915 29997 39944 30571
rect 39990 29997 40019 30571
rect 39915 29984 40019 29997
rect 40119 30571 40207 30584
rect 40119 29997 40148 30571
rect 40194 29997 40207 30571
rect 40119 29984 40207 29997
rect 40411 30571 40499 30584
rect 40411 29997 40424 30571
rect 40470 29997 40499 30571
rect 40411 29984 40499 29997
rect 40599 30571 40703 30584
rect 40599 29997 40628 30571
rect 40674 29997 40703 30571
rect 40599 29984 40703 29997
rect 40803 30571 40891 30584
rect 40803 29997 40832 30571
rect 40878 29997 40891 30571
rect 40803 29984 40891 29997
rect 41095 30571 41183 30584
rect 41095 29997 41108 30571
rect 41154 29997 41183 30571
rect 41095 29984 41183 29997
rect 41283 30571 41371 30584
rect 41283 29997 41312 30571
rect 41358 29997 41371 30571
rect 41283 29984 41371 29997
rect 42641 30657 42729 30670
rect 42641 30183 42654 30657
rect 42700 30183 42729 30657
rect 42641 30170 42729 30183
rect 42809 30657 42913 30670
rect 42809 30183 42838 30657
rect 42884 30183 42913 30657
rect 42809 30170 42913 30183
rect 42993 30657 43097 30670
rect 42993 30183 43022 30657
rect 43068 30183 43097 30657
rect 42993 30170 43097 30183
rect 43177 30657 43265 30670
rect 43177 30183 43206 30657
rect 43252 30183 43265 30657
rect 43177 30170 43265 30183
rect 37499 29407 37587 29420
rect 37499 28833 37512 29407
rect 37558 28833 37587 29407
rect 37499 28820 37587 28833
rect 37687 29407 37775 29420
rect 37687 28833 37716 29407
rect 37762 28833 37775 29407
rect 37687 28820 37775 28833
rect 38387 29407 38475 29420
rect 38387 28833 38400 29407
rect 38446 28833 38475 29407
rect 38387 28820 38475 28833
rect 38575 29407 38663 29420
rect 38575 28833 38604 29407
rect 38650 28833 38663 29407
rect 38575 28820 38663 28833
rect 38867 29407 38955 29420
rect 38867 28833 38880 29407
rect 38926 28833 38955 29407
rect 38867 28820 38955 28833
rect 39055 29407 39143 29420
rect 39055 28833 39084 29407
rect 39130 28833 39143 29407
rect 39055 28820 39143 28833
rect -12468 28396 -12380 28409
rect -12468 27822 -12455 28396
rect -12409 27822 -12380 28396
rect -12468 27809 -12380 27822
rect -12280 28396 -12192 28409
rect -12280 27822 -12251 28396
rect -12205 27822 -12192 28396
rect -12280 27809 -12192 27822
rect -7977 24969 -7889 24982
rect -7977 24495 -7964 24969
rect -7918 24495 -7889 24969
rect -7977 24482 -7889 24495
rect -7809 24969 -7705 24982
rect -7809 24495 -7780 24969
rect -7734 24495 -7705 24969
rect -7809 24482 -7705 24495
rect -7625 24969 -7521 24982
rect -7625 24495 -7596 24969
rect -7550 24495 -7521 24969
rect -7625 24482 -7521 24495
rect -7441 24969 -7353 24982
rect -7441 24495 -7412 24969
rect -7366 24495 -7353 24969
rect -7441 24482 -7353 24495
rect -3935 24966 -3847 24979
rect -3935 24492 -3922 24966
rect -3876 24492 -3847 24966
rect -3935 24479 -3847 24492
rect -3767 24966 -3663 24979
rect -3767 24492 -3738 24966
rect -3692 24492 -3663 24966
rect -3767 24479 -3663 24492
rect -3583 24966 -3479 24979
rect -3583 24492 -3554 24966
rect -3508 24492 -3479 24966
rect -3583 24479 -3479 24492
rect -3399 24966 -3311 24979
rect -3399 24492 -3370 24966
rect -3324 24492 -3311 24966
rect -3399 24479 -3311 24492
rect 107 24966 195 24979
rect 107 24492 120 24966
rect 166 24492 195 24966
rect 107 24479 195 24492
rect 275 24966 379 24979
rect 275 24492 304 24966
rect 350 24492 379 24966
rect 275 24479 379 24492
rect 459 24966 563 24979
rect 459 24492 488 24966
rect 534 24492 563 24966
rect 459 24479 563 24492
rect 643 24966 731 24979
rect 643 24492 672 24966
rect 718 24492 731 24966
rect 643 24479 731 24492
rect 4149 24966 4237 24979
rect 4149 24492 4162 24966
rect 4208 24492 4237 24966
rect 4149 24479 4237 24492
rect 4317 24966 4421 24979
rect 4317 24492 4346 24966
rect 4392 24492 4421 24966
rect 4317 24479 4421 24492
rect 4501 24966 4605 24979
rect 4501 24492 4530 24966
rect 4576 24492 4605 24966
rect 4501 24479 4605 24492
rect 4685 24966 4773 24979
rect 4685 24492 4714 24966
rect 4760 24492 4773 24966
rect 4685 24479 4773 24492
rect 8191 24966 8279 24979
rect 8191 24492 8204 24966
rect 8250 24492 8279 24966
rect 8191 24479 8279 24492
rect 8359 24966 8463 24979
rect 8359 24492 8388 24966
rect 8434 24492 8463 24966
rect 8359 24479 8463 24492
rect 8543 24966 8647 24979
rect 8543 24492 8572 24966
rect 8618 24492 8647 24966
rect 8543 24479 8647 24492
rect 8727 24966 8815 24979
rect 8727 24492 8756 24966
rect 8802 24492 8815 24966
rect 8727 24479 8815 24492
rect 12233 24966 12321 24979
rect 12233 24492 12246 24966
rect 12292 24492 12321 24966
rect 12233 24479 12321 24492
rect 12401 24966 12505 24979
rect 12401 24492 12430 24966
rect 12476 24492 12505 24966
rect 12401 24479 12505 24492
rect 12585 24966 12689 24979
rect 12585 24492 12614 24966
rect 12660 24492 12689 24966
rect 12585 24479 12689 24492
rect 12769 24966 12857 24979
rect 12769 24492 12798 24966
rect 12844 24492 12857 24966
rect 12769 24479 12857 24492
rect 16275 24966 16363 24979
rect 16275 24492 16288 24966
rect 16334 24492 16363 24966
rect 16275 24479 16363 24492
rect 16443 24966 16547 24979
rect 16443 24492 16472 24966
rect 16518 24492 16547 24966
rect 16443 24479 16547 24492
rect 16627 24966 16731 24979
rect 16627 24492 16656 24966
rect 16702 24492 16731 24966
rect 16627 24479 16731 24492
rect 16811 24966 16899 24979
rect 16811 24492 16840 24966
rect 16886 24492 16899 24966
rect 16811 24479 16899 24492
rect -7977 22764 -7889 22777
rect -7977 22290 -7964 22764
rect -7918 22290 -7889 22764
rect -7977 22277 -7889 22290
rect -7809 22764 -7705 22777
rect -7809 22290 -7780 22764
rect -7734 22290 -7705 22764
rect -7809 22277 -7705 22290
rect -7625 22764 -7521 22777
rect -7625 22290 -7596 22764
rect -7550 22290 -7521 22764
rect -7625 22277 -7521 22290
rect -7441 22764 -7353 22777
rect -7441 22290 -7412 22764
rect -7366 22290 -7353 22764
rect -7441 22277 -7353 22290
rect -6491 22764 -6403 22777
rect -6491 22290 -6478 22764
rect -6432 22290 -6403 22764
rect -6491 22277 -6403 22290
rect -6323 22764 -6219 22777
rect -6323 22290 -6294 22764
rect -6248 22290 -6219 22764
rect -6323 22277 -6219 22290
rect -6139 22764 -6035 22777
rect -6139 22290 -6110 22764
rect -6064 22290 -6035 22764
rect -6139 22277 -6035 22290
rect -5955 22764 -5867 22777
rect -5955 22290 -5926 22764
rect -5880 22290 -5867 22764
rect -5955 22277 -5867 22290
rect -3935 22761 -3847 22774
rect -3935 22287 -3922 22761
rect -3876 22287 -3847 22761
rect -3935 22274 -3847 22287
rect -3767 22761 -3663 22774
rect -3767 22287 -3738 22761
rect -3692 22287 -3663 22761
rect -3767 22274 -3663 22287
rect -3583 22761 -3479 22774
rect -3583 22287 -3554 22761
rect -3508 22287 -3479 22761
rect -3583 22274 -3479 22287
rect -3399 22761 -3311 22774
rect -3399 22287 -3370 22761
rect -3324 22287 -3311 22761
rect -3399 22274 -3311 22287
rect -2449 22761 -2361 22774
rect -2449 22287 -2436 22761
rect -2390 22287 -2361 22761
rect -2449 22274 -2361 22287
rect -2281 22761 -2177 22774
rect -2281 22287 -2252 22761
rect -2206 22287 -2177 22761
rect -2281 22274 -2177 22287
rect -2097 22761 -1993 22774
rect -2097 22287 -2068 22761
rect -2022 22287 -1993 22761
rect -2097 22274 -1993 22287
rect -1913 22761 -1825 22774
rect -1913 22287 -1884 22761
rect -1838 22287 -1825 22761
rect -1913 22274 -1825 22287
rect 107 22761 195 22774
rect 107 22287 120 22761
rect 166 22287 195 22761
rect 107 22274 195 22287
rect 275 22761 379 22774
rect 275 22287 304 22761
rect 350 22287 379 22761
rect 275 22274 379 22287
rect 459 22761 563 22774
rect 459 22287 488 22761
rect 534 22287 563 22761
rect 459 22274 563 22287
rect 643 22761 731 22774
rect 643 22287 672 22761
rect 718 22287 731 22761
rect 643 22274 731 22287
rect 1593 22761 1681 22774
rect 1593 22287 1606 22761
rect 1652 22287 1681 22761
rect 1593 22274 1681 22287
rect 1761 22761 1865 22774
rect 1761 22287 1790 22761
rect 1836 22287 1865 22761
rect 1761 22274 1865 22287
rect 1945 22761 2049 22774
rect 1945 22287 1974 22761
rect 2020 22287 2049 22761
rect 1945 22274 2049 22287
rect 2129 22761 2217 22774
rect 2129 22287 2158 22761
rect 2204 22287 2217 22761
rect 2129 22274 2217 22287
rect 4149 22761 4237 22774
rect 4149 22287 4162 22761
rect 4208 22287 4237 22761
rect 4149 22274 4237 22287
rect 4317 22761 4421 22774
rect 4317 22287 4346 22761
rect 4392 22287 4421 22761
rect 4317 22274 4421 22287
rect 4501 22761 4605 22774
rect 4501 22287 4530 22761
rect 4576 22287 4605 22761
rect 4501 22274 4605 22287
rect 4685 22761 4773 22774
rect 4685 22287 4714 22761
rect 4760 22287 4773 22761
rect 4685 22274 4773 22287
rect 5635 22761 5723 22774
rect 5635 22287 5648 22761
rect 5694 22287 5723 22761
rect 5635 22274 5723 22287
rect 5803 22761 5907 22774
rect 5803 22287 5832 22761
rect 5878 22287 5907 22761
rect 5803 22274 5907 22287
rect 5987 22761 6091 22774
rect 5987 22287 6016 22761
rect 6062 22287 6091 22761
rect 5987 22274 6091 22287
rect 6171 22761 6259 22774
rect 6171 22287 6200 22761
rect 6246 22287 6259 22761
rect 6171 22274 6259 22287
rect 8191 22761 8279 22774
rect 8191 22287 8204 22761
rect 8250 22287 8279 22761
rect 8191 22274 8279 22287
rect 8359 22761 8463 22774
rect 8359 22287 8388 22761
rect 8434 22287 8463 22761
rect 8359 22274 8463 22287
rect 8543 22761 8647 22774
rect 8543 22287 8572 22761
rect 8618 22287 8647 22761
rect 8543 22274 8647 22287
rect 8727 22761 8815 22774
rect 8727 22287 8756 22761
rect 8802 22287 8815 22761
rect 8727 22274 8815 22287
rect 9677 22761 9765 22774
rect 9677 22287 9690 22761
rect 9736 22287 9765 22761
rect 9677 22274 9765 22287
rect 9845 22761 9949 22774
rect 9845 22287 9874 22761
rect 9920 22287 9949 22761
rect 9845 22274 9949 22287
rect 10029 22761 10133 22774
rect 10029 22287 10058 22761
rect 10104 22287 10133 22761
rect 10029 22274 10133 22287
rect 10213 22761 10301 22774
rect 10213 22287 10242 22761
rect 10288 22287 10301 22761
rect 10213 22274 10301 22287
rect 12233 22761 12321 22774
rect 12233 22287 12246 22761
rect 12292 22287 12321 22761
rect 12233 22274 12321 22287
rect 12401 22761 12505 22774
rect 12401 22287 12430 22761
rect 12476 22287 12505 22761
rect 12401 22274 12505 22287
rect 12585 22761 12689 22774
rect 12585 22287 12614 22761
rect 12660 22287 12689 22761
rect 12585 22274 12689 22287
rect 12769 22761 12857 22774
rect 12769 22287 12798 22761
rect 12844 22287 12857 22761
rect 12769 22274 12857 22287
rect 13719 22761 13807 22774
rect 13719 22287 13732 22761
rect 13778 22287 13807 22761
rect 13719 22274 13807 22287
rect 13887 22761 13991 22774
rect 13887 22287 13916 22761
rect 13962 22287 13991 22761
rect 13887 22274 13991 22287
rect 14071 22761 14175 22774
rect 14071 22287 14100 22761
rect 14146 22287 14175 22761
rect 14071 22274 14175 22287
rect 14255 22761 14343 22774
rect 14255 22287 14284 22761
rect 14330 22287 14343 22761
rect 14255 22274 14343 22287
rect 16275 22761 16363 22774
rect 16275 22287 16288 22761
rect 16334 22287 16363 22761
rect 16275 22274 16363 22287
rect 16443 22761 16547 22774
rect 16443 22287 16472 22761
rect 16518 22287 16547 22761
rect 16443 22274 16547 22287
rect 16627 22761 16731 22774
rect 16627 22287 16656 22761
rect 16702 22287 16731 22761
rect 16627 22274 16731 22287
rect 16811 22761 16899 22774
rect 16811 22287 16840 22761
rect 16886 22287 16899 22761
rect 16811 22274 16899 22287
rect 17761 22761 17849 22774
rect 17761 22287 17774 22761
rect 17820 22287 17849 22761
rect 17761 22274 17849 22287
rect 17929 22761 18033 22774
rect 17929 22287 17958 22761
rect 18004 22287 18033 22761
rect 17929 22274 18033 22287
rect 18113 22761 18217 22774
rect 18113 22287 18142 22761
rect 18188 22287 18217 22761
rect 18113 22274 18217 22287
rect 18297 22761 18385 22774
rect 18297 22287 18326 22761
rect 18372 22287 18385 22761
rect 18297 22274 18385 22287
rect -7977 20559 -7889 20572
rect -7977 20085 -7964 20559
rect -7918 20085 -7889 20559
rect -7977 20072 -7889 20085
rect -7809 20559 -7705 20572
rect -7809 20085 -7780 20559
rect -7734 20085 -7705 20559
rect -7809 20072 -7705 20085
rect -7625 20559 -7521 20572
rect -7625 20085 -7596 20559
rect -7550 20085 -7521 20559
rect -7625 20072 -7521 20085
rect -7441 20559 -7353 20572
rect -7441 20085 -7412 20559
rect -7366 20085 -7353 20559
rect -7441 20072 -7353 20085
rect -6491 20560 -6403 20573
rect -6491 20086 -6478 20560
rect -6432 20086 -6403 20560
rect -6491 20073 -6403 20086
rect -6323 20560 -6219 20573
rect -6323 20086 -6294 20560
rect -6248 20086 -6219 20560
rect -6323 20073 -6219 20086
rect -6139 20560 -6035 20573
rect -6139 20086 -6110 20560
rect -6064 20086 -6035 20560
rect -6139 20073 -6035 20086
rect -5955 20560 -5867 20573
rect -5955 20086 -5926 20560
rect -5880 20086 -5867 20560
rect -5955 20073 -5867 20086
rect -3935 20556 -3847 20569
rect -3935 20082 -3922 20556
rect -3876 20082 -3847 20556
rect -3935 20069 -3847 20082
rect -3767 20556 -3663 20569
rect -3767 20082 -3738 20556
rect -3692 20082 -3663 20556
rect -3767 20069 -3663 20082
rect -3583 20556 -3479 20569
rect -3583 20082 -3554 20556
rect -3508 20082 -3479 20556
rect -3583 20069 -3479 20082
rect -3399 20556 -3311 20569
rect -3399 20082 -3370 20556
rect -3324 20082 -3311 20556
rect -3399 20069 -3311 20082
rect -2449 20557 -2361 20570
rect -2449 20083 -2436 20557
rect -2390 20083 -2361 20557
rect -2449 20070 -2361 20083
rect -2281 20557 -2177 20570
rect -2281 20083 -2252 20557
rect -2206 20083 -2177 20557
rect -2281 20070 -2177 20083
rect -2097 20557 -1993 20570
rect -2097 20083 -2068 20557
rect -2022 20083 -1993 20557
rect -2097 20070 -1993 20083
rect -1913 20557 -1825 20570
rect -1913 20083 -1884 20557
rect -1838 20083 -1825 20557
rect -1913 20070 -1825 20083
rect 107 20556 195 20569
rect 107 20082 120 20556
rect 166 20082 195 20556
rect 107 20069 195 20082
rect 275 20556 379 20569
rect 275 20082 304 20556
rect 350 20082 379 20556
rect 275 20069 379 20082
rect 459 20556 563 20569
rect 459 20082 488 20556
rect 534 20082 563 20556
rect 459 20069 563 20082
rect 643 20556 731 20569
rect 643 20082 672 20556
rect 718 20082 731 20556
rect 643 20069 731 20082
rect 1593 20557 1681 20570
rect 1593 20083 1606 20557
rect 1652 20083 1681 20557
rect 1593 20070 1681 20083
rect 1761 20557 1865 20570
rect 1761 20083 1790 20557
rect 1836 20083 1865 20557
rect 1761 20070 1865 20083
rect 1945 20557 2049 20570
rect 1945 20083 1974 20557
rect 2020 20083 2049 20557
rect 1945 20070 2049 20083
rect 2129 20557 2217 20570
rect 2129 20083 2158 20557
rect 2204 20083 2217 20557
rect 2129 20070 2217 20083
rect 4149 20556 4237 20569
rect 4149 20082 4162 20556
rect 4208 20082 4237 20556
rect 4149 20069 4237 20082
rect 4317 20556 4421 20569
rect 4317 20082 4346 20556
rect 4392 20082 4421 20556
rect 4317 20069 4421 20082
rect 4501 20556 4605 20569
rect 4501 20082 4530 20556
rect 4576 20082 4605 20556
rect 4501 20069 4605 20082
rect 4685 20556 4773 20569
rect 4685 20082 4714 20556
rect 4760 20082 4773 20556
rect 4685 20069 4773 20082
rect 5635 20557 5723 20570
rect 5635 20083 5648 20557
rect 5694 20083 5723 20557
rect 5635 20070 5723 20083
rect 5803 20557 5907 20570
rect 5803 20083 5832 20557
rect 5878 20083 5907 20557
rect 5803 20070 5907 20083
rect 5987 20557 6091 20570
rect 5987 20083 6016 20557
rect 6062 20083 6091 20557
rect 5987 20070 6091 20083
rect 6171 20557 6259 20570
rect 6171 20083 6200 20557
rect 6246 20083 6259 20557
rect 6171 20070 6259 20083
rect 8191 20556 8279 20569
rect 8191 20082 8204 20556
rect 8250 20082 8279 20556
rect 8191 20069 8279 20082
rect 8359 20556 8463 20569
rect 8359 20082 8388 20556
rect 8434 20082 8463 20556
rect 8359 20069 8463 20082
rect 8543 20556 8647 20569
rect 8543 20082 8572 20556
rect 8618 20082 8647 20556
rect 8543 20069 8647 20082
rect 8727 20556 8815 20569
rect 8727 20082 8756 20556
rect 8802 20082 8815 20556
rect 8727 20069 8815 20082
rect 9677 20557 9765 20570
rect 9677 20083 9690 20557
rect 9736 20083 9765 20557
rect 9677 20070 9765 20083
rect 9845 20557 9949 20570
rect 9845 20083 9874 20557
rect 9920 20083 9949 20557
rect 9845 20070 9949 20083
rect 10029 20557 10133 20570
rect 10029 20083 10058 20557
rect 10104 20083 10133 20557
rect 10029 20070 10133 20083
rect 10213 20557 10301 20570
rect 10213 20083 10242 20557
rect 10288 20083 10301 20557
rect 10213 20070 10301 20083
rect 12233 20556 12321 20569
rect 12233 20082 12246 20556
rect 12292 20082 12321 20556
rect 12233 20069 12321 20082
rect 12401 20556 12505 20569
rect 12401 20082 12430 20556
rect 12476 20082 12505 20556
rect 12401 20069 12505 20082
rect 12585 20556 12689 20569
rect 12585 20082 12614 20556
rect 12660 20082 12689 20556
rect 12585 20069 12689 20082
rect 12769 20556 12857 20569
rect 12769 20082 12798 20556
rect 12844 20082 12857 20556
rect 12769 20069 12857 20082
rect 13719 20557 13807 20570
rect 13719 20083 13732 20557
rect 13778 20083 13807 20557
rect 13719 20070 13807 20083
rect 13887 20557 13991 20570
rect 13887 20083 13916 20557
rect 13962 20083 13991 20557
rect 13887 20070 13991 20083
rect 14071 20557 14175 20570
rect 14071 20083 14100 20557
rect 14146 20083 14175 20557
rect 14071 20070 14175 20083
rect 14255 20557 14343 20570
rect 14255 20083 14284 20557
rect 14330 20083 14343 20557
rect 14255 20070 14343 20083
rect 16275 20556 16363 20569
rect 16275 20082 16288 20556
rect 16334 20082 16363 20556
rect 16275 20069 16363 20082
rect 16443 20556 16547 20569
rect 16443 20082 16472 20556
rect 16518 20082 16547 20556
rect 16443 20069 16547 20082
rect 16627 20556 16731 20569
rect 16627 20082 16656 20556
rect 16702 20082 16731 20556
rect 16627 20069 16731 20082
rect 16811 20556 16899 20569
rect 16811 20082 16840 20556
rect 16886 20082 16899 20556
rect 16811 20069 16899 20082
rect 17761 20557 17849 20570
rect 17761 20083 17774 20557
rect 17820 20083 17849 20557
rect 17761 20070 17849 20083
rect 17929 20557 18033 20570
rect 17929 20083 17958 20557
rect 18004 20083 18033 20557
rect 17929 20070 18033 20083
rect 18113 20557 18217 20570
rect 18113 20083 18142 20557
rect 18188 20083 18217 20557
rect 18113 20070 18217 20083
rect 18297 20557 18385 20570
rect 18297 20083 18326 20557
rect 18372 20083 18385 20557
rect 18297 20070 18385 20083
rect -7977 18354 -7889 18367
rect -7977 17880 -7964 18354
rect -7918 17880 -7889 18354
rect -7977 17867 -7889 17880
rect -7809 18354 -7705 18367
rect -7809 17880 -7780 18354
rect -7734 17880 -7705 18354
rect -7809 17867 -7705 17880
rect -7625 18354 -7521 18367
rect -7625 17880 -7596 18354
rect -7550 17880 -7521 18354
rect -7625 17867 -7521 17880
rect -7441 18354 -7353 18367
rect -7441 17880 -7412 18354
rect -7366 17880 -7353 18354
rect -7441 17867 -7353 17880
rect -3935 18351 -3847 18364
rect -3935 17877 -3922 18351
rect -3876 17877 -3847 18351
rect -3935 17864 -3847 17877
rect -3767 18351 -3663 18364
rect -3767 17877 -3738 18351
rect -3692 17877 -3663 18351
rect -3767 17864 -3663 17877
rect -3583 18351 -3479 18364
rect -3583 17877 -3554 18351
rect -3508 17877 -3479 18351
rect -3583 17864 -3479 17877
rect -3399 18351 -3311 18364
rect -3399 17877 -3370 18351
rect -3324 17877 -3311 18351
rect -3399 17864 -3311 17877
rect 107 18351 195 18364
rect 107 17877 120 18351
rect 166 17877 195 18351
rect 107 17864 195 17877
rect 275 18351 379 18364
rect 275 17877 304 18351
rect 350 17877 379 18351
rect 275 17864 379 17877
rect 459 18351 563 18364
rect 459 17877 488 18351
rect 534 17877 563 18351
rect 459 17864 563 17877
rect 643 18351 731 18364
rect 643 17877 672 18351
rect 718 17877 731 18351
rect 643 17864 731 17877
rect 4149 18351 4237 18364
rect 4149 17877 4162 18351
rect 4208 17877 4237 18351
rect 4149 17864 4237 17877
rect 4317 18351 4421 18364
rect 4317 17877 4346 18351
rect 4392 17877 4421 18351
rect 4317 17864 4421 17877
rect 4501 18351 4605 18364
rect 4501 17877 4530 18351
rect 4576 17877 4605 18351
rect 4501 17864 4605 17877
rect 4685 18351 4773 18364
rect 4685 17877 4714 18351
rect 4760 17877 4773 18351
rect 4685 17864 4773 17877
rect 8191 18351 8279 18364
rect 8191 17877 8204 18351
rect 8250 17877 8279 18351
rect 8191 17864 8279 17877
rect 8359 18351 8463 18364
rect 8359 17877 8388 18351
rect 8434 17877 8463 18351
rect 8359 17864 8463 17877
rect 8543 18351 8647 18364
rect 8543 17877 8572 18351
rect 8618 17877 8647 18351
rect 8543 17864 8647 17877
rect 8727 18351 8815 18364
rect 8727 17877 8756 18351
rect 8802 17877 8815 18351
rect 8727 17864 8815 17877
rect 12233 18351 12321 18364
rect 12233 17877 12246 18351
rect 12292 17877 12321 18351
rect 12233 17864 12321 17877
rect 12401 18351 12505 18364
rect 12401 17877 12430 18351
rect 12476 17877 12505 18351
rect 12401 17864 12505 17877
rect 12585 18351 12689 18364
rect 12585 17877 12614 18351
rect 12660 17877 12689 18351
rect 12585 17864 12689 17877
rect 12769 18351 12857 18364
rect 12769 17877 12798 18351
rect 12844 17877 12857 18351
rect 12769 17864 12857 17877
rect 16275 18351 16363 18364
rect 16275 17877 16288 18351
rect 16334 17877 16363 18351
rect 16275 17864 16363 17877
rect 16443 18351 16547 18364
rect 16443 17877 16472 18351
rect 16518 17877 16547 18351
rect 16443 17864 16547 17877
rect 16627 18351 16731 18364
rect 16627 17877 16656 18351
rect 16702 17877 16731 18351
rect 16627 17864 16731 17877
rect 16811 18351 16899 18364
rect 16811 17877 16840 18351
rect 16886 17877 16899 18351
rect 16811 17864 16899 17877
rect -11989 15390 -11901 15403
rect -11989 14916 -11976 15390
rect -11930 14916 -11901 15390
rect -11989 14903 -11901 14916
rect -11821 15390 -11717 15403
rect -11821 14916 -11792 15390
rect -11746 14916 -11717 15390
rect -11821 14903 -11717 14916
rect -11637 15390 -11533 15403
rect -11637 14916 -11608 15390
rect -11562 14916 -11533 15390
rect -11637 14903 -11533 14916
rect -11453 15390 -11365 15403
rect -11453 14916 -11424 15390
rect -11378 14916 -11365 15390
rect -11453 14903 -11365 14916
rect -7977 15390 -7889 15403
rect -7977 14916 -7964 15390
rect -7918 14916 -7889 15390
rect -7977 14903 -7889 14916
rect -7809 15390 -7705 15403
rect -7809 14916 -7780 15390
rect -7734 14916 -7705 15390
rect -7809 14903 -7705 14916
rect -7625 15390 -7521 15403
rect -7625 14916 -7596 15390
rect -7550 14916 -7521 15390
rect -7625 14903 -7521 14916
rect -7441 15390 -7353 15403
rect -7441 14916 -7412 15390
rect -7366 14916 -7353 15390
rect -7441 14903 -7353 14916
rect -3935 15390 -3847 15403
rect -3935 14916 -3922 15390
rect -3876 14916 -3847 15390
rect -3935 14903 -3847 14916
rect -3767 15390 -3663 15403
rect -3767 14916 -3738 15390
rect -3692 14916 -3663 15390
rect -3767 14903 -3663 14916
rect -3583 15390 -3479 15403
rect -3583 14916 -3554 15390
rect -3508 14916 -3479 15390
rect -3583 14903 -3479 14916
rect -3399 15390 -3311 15403
rect -3399 14916 -3370 15390
rect -3324 14916 -3311 15390
rect -3399 14903 -3311 14916
rect 107 15390 195 15403
rect 107 14916 120 15390
rect 166 14916 195 15390
rect 107 14903 195 14916
rect 275 15390 379 15403
rect 275 14916 304 15390
rect 350 14916 379 15390
rect 275 14903 379 14916
rect 459 15390 563 15403
rect 459 14916 488 15390
rect 534 14916 563 15390
rect 459 14903 563 14916
rect 643 15390 731 15403
rect 643 14916 672 15390
rect 718 14916 731 15390
rect 643 14903 731 14916
rect 4149 15390 4237 15403
rect 4149 14916 4162 15390
rect 4208 14916 4237 15390
rect 4149 14903 4237 14916
rect 4317 15390 4421 15403
rect 4317 14916 4346 15390
rect 4392 14916 4421 15390
rect 4317 14903 4421 14916
rect 4501 15390 4605 15403
rect 4501 14916 4530 15390
rect 4576 14916 4605 15390
rect 4501 14903 4605 14916
rect 4685 15390 4773 15403
rect 4685 14916 4714 15390
rect 4760 14916 4773 15390
rect 4685 14903 4773 14916
rect 8191 15390 8279 15403
rect 8191 14916 8204 15390
rect 8250 14916 8279 15390
rect 8191 14903 8279 14916
rect 8359 15390 8463 15403
rect 8359 14916 8388 15390
rect 8434 14916 8463 15390
rect 8359 14903 8463 14916
rect 8543 15390 8647 15403
rect 8543 14916 8572 15390
rect 8618 14916 8647 15390
rect 8543 14903 8647 14916
rect 8727 15390 8815 15403
rect 8727 14916 8756 15390
rect 8802 14916 8815 15390
rect 8727 14903 8815 14916
rect 12233 15390 12321 15403
rect 12233 14916 12246 15390
rect 12292 14916 12321 15390
rect 12233 14903 12321 14916
rect 12401 15390 12505 15403
rect 12401 14916 12430 15390
rect 12476 14916 12505 15390
rect 12401 14903 12505 14916
rect 12585 15390 12689 15403
rect 12585 14916 12614 15390
rect 12660 14916 12689 15390
rect 12585 14903 12689 14916
rect 12769 15390 12857 15403
rect 12769 14916 12798 15390
rect 12844 14916 12857 15390
rect 12769 14903 12857 14916
rect -11989 13185 -11901 13198
rect -11989 12711 -11976 13185
rect -11930 12711 -11901 13185
rect -11989 12698 -11901 12711
rect -11821 13185 -11717 13198
rect -11821 12711 -11792 13185
rect -11746 12711 -11717 13185
rect -11821 12698 -11717 12711
rect -11637 13185 -11533 13198
rect -11637 12711 -11608 13185
rect -11562 12711 -11533 13185
rect -11637 12698 -11533 12711
rect -11453 13185 -11365 13198
rect -11453 12711 -11424 13185
rect -11378 12711 -11365 13185
rect -11453 12698 -11365 12711
rect -10503 13185 -10415 13198
rect -10503 12711 -10490 13185
rect -10444 12711 -10415 13185
rect -10503 12698 -10415 12711
rect -10335 13185 -10231 13198
rect -10335 12711 -10306 13185
rect -10260 12711 -10231 13185
rect -10335 12698 -10231 12711
rect -10151 13185 -10047 13198
rect -10151 12711 -10122 13185
rect -10076 12711 -10047 13185
rect -10151 12698 -10047 12711
rect -9967 13185 -9879 13198
rect -9967 12711 -9938 13185
rect -9892 12711 -9879 13185
rect -9967 12698 -9879 12711
rect -7977 13185 -7889 13198
rect -7977 12711 -7964 13185
rect -7918 12711 -7889 13185
rect -7977 12698 -7889 12711
rect -7809 13185 -7705 13198
rect -7809 12711 -7780 13185
rect -7734 12711 -7705 13185
rect -7809 12698 -7705 12711
rect -7625 13185 -7521 13198
rect -7625 12711 -7596 13185
rect -7550 12711 -7521 13185
rect -7625 12698 -7521 12711
rect -7441 13185 -7353 13198
rect -7441 12711 -7412 13185
rect -7366 12711 -7353 13185
rect -7441 12698 -7353 12711
rect -6491 13185 -6403 13198
rect -6491 12711 -6478 13185
rect -6432 12711 -6403 13185
rect -6491 12698 -6403 12711
rect -6323 13185 -6219 13198
rect -6323 12711 -6294 13185
rect -6248 12711 -6219 13185
rect -6323 12698 -6219 12711
rect -6139 13185 -6035 13198
rect -6139 12711 -6110 13185
rect -6064 12711 -6035 13185
rect -6139 12698 -6035 12711
rect -5955 13185 -5867 13198
rect -5955 12711 -5926 13185
rect -5880 12711 -5867 13185
rect -5955 12698 -5867 12711
rect -3935 13185 -3847 13198
rect -3935 12711 -3922 13185
rect -3876 12711 -3847 13185
rect -3935 12698 -3847 12711
rect -3767 13185 -3663 13198
rect -3767 12711 -3738 13185
rect -3692 12711 -3663 13185
rect -3767 12698 -3663 12711
rect -3583 13185 -3479 13198
rect -3583 12711 -3554 13185
rect -3508 12711 -3479 13185
rect -3583 12698 -3479 12711
rect -3399 13185 -3311 13198
rect -3399 12711 -3370 13185
rect -3324 12711 -3311 13185
rect -3399 12698 -3311 12711
rect -2449 13185 -2361 13198
rect -2449 12711 -2436 13185
rect -2390 12711 -2361 13185
rect -2449 12698 -2361 12711
rect -2281 13185 -2177 13198
rect -2281 12711 -2252 13185
rect -2206 12711 -2177 13185
rect -2281 12698 -2177 12711
rect -2097 13185 -1993 13198
rect -2097 12711 -2068 13185
rect -2022 12711 -1993 13185
rect -2097 12698 -1993 12711
rect -1913 13185 -1825 13198
rect -1913 12711 -1884 13185
rect -1838 12711 -1825 13185
rect -1913 12698 -1825 12711
rect 107 13185 195 13198
rect 107 12711 120 13185
rect 166 12711 195 13185
rect 107 12698 195 12711
rect 275 13185 379 13198
rect 275 12711 304 13185
rect 350 12711 379 13185
rect 275 12698 379 12711
rect 459 13185 563 13198
rect 459 12711 488 13185
rect 534 12711 563 13185
rect 459 12698 563 12711
rect 643 13185 731 13198
rect 643 12711 672 13185
rect 718 12711 731 13185
rect 643 12698 731 12711
rect 1593 13185 1681 13198
rect 1593 12711 1606 13185
rect 1652 12711 1681 13185
rect 1593 12698 1681 12711
rect 1761 13185 1865 13198
rect 1761 12711 1790 13185
rect 1836 12711 1865 13185
rect 1761 12698 1865 12711
rect 1945 13185 2049 13198
rect 1945 12711 1974 13185
rect 2020 12711 2049 13185
rect 1945 12698 2049 12711
rect 2129 13185 2217 13198
rect 2129 12711 2158 13185
rect 2204 12711 2217 13185
rect 2129 12698 2217 12711
rect 4149 13185 4237 13198
rect 4149 12711 4162 13185
rect 4208 12711 4237 13185
rect 4149 12698 4237 12711
rect 4317 13185 4421 13198
rect 4317 12711 4346 13185
rect 4392 12711 4421 13185
rect 4317 12698 4421 12711
rect 4501 13185 4605 13198
rect 4501 12711 4530 13185
rect 4576 12711 4605 13185
rect 4501 12698 4605 12711
rect 4685 13185 4773 13198
rect 4685 12711 4714 13185
rect 4760 12711 4773 13185
rect 4685 12698 4773 12711
rect 5635 13185 5723 13198
rect 5635 12711 5648 13185
rect 5694 12711 5723 13185
rect 5635 12698 5723 12711
rect 5803 13185 5907 13198
rect 5803 12711 5832 13185
rect 5878 12711 5907 13185
rect 5803 12698 5907 12711
rect 5987 13185 6091 13198
rect 5987 12711 6016 13185
rect 6062 12711 6091 13185
rect 5987 12698 6091 12711
rect 6171 13185 6259 13198
rect 6171 12711 6200 13185
rect 6246 12711 6259 13185
rect 6171 12698 6259 12711
rect 8191 13185 8279 13198
rect 8191 12711 8204 13185
rect 8250 12711 8279 13185
rect 8191 12698 8279 12711
rect 8359 13185 8463 13198
rect 8359 12711 8388 13185
rect 8434 12711 8463 13185
rect 8359 12698 8463 12711
rect 8543 13185 8647 13198
rect 8543 12711 8572 13185
rect 8618 12711 8647 13185
rect 8543 12698 8647 12711
rect 8727 13185 8815 13198
rect 8727 12711 8756 13185
rect 8802 12711 8815 13185
rect 8727 12698 8815 12711
rect 9677 13185 9765 13198
rect 9677 12711 9690 13185
rect 9736 12711 9765 13185
rect 9677 12698 9765 12711
rect 9845 13185 9949 13198
rect 9845 12711 9874 13185
rect 9920 12711 9949 13185
rect 9845 12698 9949 12711
rect 10029 13185 10133 13198
rect 10029 12711 10058 13185
rect 10104 12711 10133 13185
rect 10029 12698 10133 12711
rect 10213 13185 10301 13198
rect 10213 12711 10242 13185
rect 10288 12711 10301 13185
rect 10213 12698 10301 12711
rect 12233 13185 12321 13198
rect 12233 12711 12246 13185
rect 12292 12711 12321 13185
rect 12233 12698 12321 12711
rect 12401 13185 12505 13198
rect 12401 12711 12430 13185
rect 12476 12711 12505 13185
rect 12401 12698 12505 12711
rect 12585 13185 12689 13198
rect 12585 12711 12614 13185
rect 12660 12711 12689 13185
rect 12585 12698 12689 12711
rect 12769 13185 12857 13198
rect 12769 12711 12798 13185
rect 12844 12711 12857 13185
rect 12769 12698 12857 12711
rect 13719 13185 13807 13198
rect 13719 12711 13732 13185
rect 13778 12711 13807 13185
rect 13719 12698 13807 12711
rect 13887 13185 13991 13198
rect 13887 12711 13916 13185
rect 13962 12711 13991 13185
rect 13887 12698 13991 12711
rect 14071 13185 14175 13198
rect 14071 12711 14100 13185
rect 14146 12711 14175 13185
rect 14071 12698 14175 12711
rect 14255 13185 14343 13198
rect 14255 12711 14284 13185
rect 14330 12711 14343 13185
rect 14255 12698 14343 12711
rect -11989 10980 -11901 10993
rect -11989 10506 -11976 10980
rect -11930 10506 -11901 10980
rect -11989 10493 -11901 10506
rect -11821 10980 -11717 10993
rect -11821 10506 -11792 10980
rect -11746 10506 -11717 10980
rect -11821 10493 -11717 10506
rect -11637 10980 -11533 10993
rect -11637 10506 -11608 10980
rect -11562 10506 -11533 10980
rect -11637 10493 -11533 10506
rect -11453 10980 -11365 10993
rect -11453 10506 -11424 10980
rect -11378 10506 -11365 10980
rect -11453 10493 -11365 10506
rect -10503 10981 -10415 10994
rect -10503 10507 -10490 10981
rect -10444 10507 -10415 10981
rect -10503 10494 -10415 10507
rect -10335 10981 -10231 10994
rect -10335 10507 -10306 10981
rect -10260 10507 -10231 10981
rect -10335 10494 -10231 10507
rect -10151 10981 -10047 10994
rect -10151 10507 -10122 10981
rect -10076 10507 -10047 10981
rect -10151 10494 -10047 10507
rect -9967 10981 -9879 10994
rect -9967 10507 -9938 10981
rect -9892 10507 -9879 10981
rect -9967 10494 -9879 10507
rect -7977 10980 -7889 10993
rect -7977 10506 -7964 10980
rect -7918 10506 -7889 10980
rect -7977 10493 -7889 10506
rect -7809 10980 -7705 10993
rect -7809 10506 -7780 10980
rect -7734 10506 -7705 10980
rect -7809 10493 -7705 10506
rect -7625 10980 -7521 10993
rect -7625 10506 -7596 10980
rect -7550 10506 -7521 10980
rect -7625 10493 -7521 10506
rect -7441 10980 -7353 10993
rect -7441 10506 -7412 10980
rect -7366 10506 -7353 10980
rect -7441 10493 -7353 10506
rect -6491 10981 -6403 10994
rect -6491 10507 -6478 10981
rect -6432 10507 -6403 10981
rect -6491 10494 -6403 10507
rect -6323 10981 -6219 10994
rect -6323 10507 -6294 10981
rect -6248 10507 -6219 10981
rect -6323 10494 -6219 10507
rect -6139 10981 -6035 10994
rect -6139 10507 -6110 10981
rect -6064 10507 -6035 10981
rect -6139 10494 -6035 10507
rect -5955 10981 -5867 10994
rect -5955 10507 -5926 10981
rect -5880 10507 -5867 10981
rect -5955 10494 -5867 10507
rect -3935 10980 -3847 10993
rect -3935 10506 -3922 10980
rect -3876 10506 -3847 10980
rect -3935 10493 -3847 10506
rect -3767 10980 -3663 10993
rect -3767 10506 -3738 10980
rect -3692 10506 -3663 10980
rect -3767 10493 -3663 10506
rect -3583 10980 -3479 10993
rect -3583 10506 -3554 10980
rect -3508 10506 -3479 10980
rect -3583 10493 -3479 10506
rect -3399 10980 -3311 10993
rect -3399 10506 -3370 10980
rect -3324 10506 -3311 10980
rect -3399 10493 -3311 10506
rect -2449 10981 -2361 10994
rect -2449 10507 -2436 10981
rect -2390 10507 -2361 10981
rect -2449 10494 -2361 10507
rect -2281 10981 -2177 10994
rect -2281 10507 -2252 10981
rect -2206 10507 -2177 10981
rect -2281 10494 -2177 10507
rect -2097 10981 -1993 10994
rect -2097 10507 -2068 10981
rect -2022 10507 -1993 10981
rect -2097 10494 -1993 10507
rect -1913 10981 -1825 10994
rect -1913 10507 -1884 10981
rect -1838 10507 -1825 10981
rect -1913 10494 -1825 10507
rect 107 10980 195 10993
rect 107 10506 120 10980
rect 166 10506 195 10980
rect 107 10493 195 10506
rect 275 10980 379 10993
rect 275 10506 304 10980
rect 350 10506 379 10980
rect 275 10493 379 10506
rect 459 10980 563 10993
rect 459 10506 488 10980
rect 534 10506 563 10980
rect 459 10493 563 10506
rect 643 10980 731 10993
rect 643 10506 672 10980
rect 718 10506 731 10980
rect 643 10493 731 10506
rect 1593 10981 1681 10994
rect 1593 10507 1606 10981
rect 1652 10507 1681 10981
rect 1593 10494 1681 10507
rect 1761 10981 1865 10994
rect 1761 10507 1790 10981
rect 1836 10507 1865 10981
rect 1761 10494 1865 10507
rect 1945 10981 2049 10994
rect 1945 10507 1974 10981
rect 2020 10507 2049 10981
rect 1945 10494 2049 10507
rect 2129 10981 2217 10994
rect 2129 10507 2158 10981
rect 2204 10507 2217 10981
rect 2129 10494 2217 10507
rect 4149 10980 4237 10993
rect 4149 10506 4162 10980
rect 4208 10506 4237 10980
rect 4149 10493 4237 10506
rect 4317 10980 4421 10993
rect 4317 10506 4346 10980
rect 4392 10506 4421 10980
rect 4317 10493 4421 10506
rect 4501 10980 4605 10993
rect 4501 10506 4530 10980
rect 4576 10506 4605 10980
rect 4501 10493 4605 10506
rect 4685 10980 4773 10993
rect 4685 10506 4714 10980
rect 4760 10506 4773 10980
rect 4685 10493 4773 10506
rect 5635 10981 5723 10994
rect 5635 10507 5648 10981
rect 5694 10507 5723 10981
rect 5635 10494 5723 10507
rect 5803 10981 5907 10994
rect 5803 10507 5832 10981
rect 5878 10507 5907 10981
rect 5803 10494 5907 10507
rect 5987 10981 6091 10994
rect 5987 10507 6016 10981
rect 6062 10507 6091 10981
rect 5987 10494 6091 10507
rect 6171 10981 6259 10994
rect 6171 10507 6200 10981
rect 6246 10507 6259 10981
rect 6171 10494 6259 10507
rect 8191 10980 8279 10993
rect 8191 10506 8204 10980
rect 8250 10506 8279 10980
rect 8191 10493 8279 10506
rect 8359 10980 8463 10993
rect 8359 10506 8388 10980
rect 8434 10506 8463 10980
rect 8359 10493 8463 10506
rect 8543 10980 8647 10993
rect 8543 10506 8572 10980
rect 8618 10506 8647 10980
rect 8543 10493 8647 10506
rect 8727 10980 8815 10993
rect 8727 10506 8756 10980
rect 8802 10506 8815 10980
rect 8727 10493 8815 10506
rect 9677 10981 9765 10994
rect 9677 10507 9690 10981
rect 9736 10507 9765 10981
rect 9677 10494 9765 10507
rect 9845 10981 9949 10994
rect 9845 10507 9874 10981
rect 9920 10507 9949 10981
rect 9845 10494 9949 10507
rect 10029 10981 10133 10994
rect 10029 10507 10058 10981
rect 10104 10507 10133 10981
rect 10029 10494 10133 10507
rect 10213 10981 10301 10994
rect 10213 10507 10242 10981
rect 10288 10507 10301 10981
rect 10213 10494 10301 10507
rect 12233 10980 12321 10993
rect 12233 10506 12246 10980
rect 12292 10506 12321 10980
rect 12233 10493 12321 10506
rect 12401 10980 12505 10993
rect 12401 10506 12430 10980
rect 12476 10506 12505 10980
rect 12401 10493 12505 10506
rect 12585 10980 12689 10993
rect 12585 10506 12614 10980
rect 12660 10506 12689 10980
rect 12585 10493 12689 10506
rect 12769 10980 12857 10993
rect 12769 10506 12798 10980
rect 12844 10506 12857 10980
rect 12769 10493 12857 10506
rect 13719 10981 13807 10994
rect 13719 10507 13732 10981
rect 13778 10507 13807 10981
rect 13719 10494 13807 10507
rect 13887 10981 13991 10994
rect 13887 10507 13916 10981
rect 13962 10507 13991 10981
rect 13887 10494 13991 10507
rect 14071 10981 14175 10994
rect 14071 10507 14100 10981
rect 14146 10507 14175 10981
rect 14071 10494 14175 10507
rect 14255 10981 14343 10994
rect 14255 10507 14284 10981
rect 14330 10507 14343 10981
rect 14255 10494 14343 10507
rect -11989 8775 -11901 8788
rect -11989 8301 -11976 8775
rect -11930 8301 -11901 8775
rect -11989 8288 -11901 8301
rect -11821 8775 -11717 8788
rect -11821 8301 -11792 8775
rect -11746 8301 -11717 8775
rect -11821 8288 -11717 8301
rect -11637 8775 -11533 8788
rect -11637 8301 -11608 8775
rect -11562 8301 -11533 8775
rect -11637 8288 -11533 8301
rect -11453 8775 -11365 8788
rect -11453 8301 -11424 8775
rect -11378 8301 -11365 8775
rect -11453 8288 -11365 8301
rect -7977 8775 -7889 8788
rect -7977 8301 -7964 8775
rect -7918 8301 -7889 8775
rect -7977 8288 -7889 8301
rect -7809 8775 -7705 8788
rect -7809 8301 -7780 8775
rect -7734 8301 -7705 8775
rect -7809 8288 -7705 8301
rect -7625 8775 -7521 8788
rect -7625 8301 -7596 8775
rect -7550 8301 -7521 8775
rect -7625 8288 -7521 8301
rect -7441 8775 -7353 8788
rect -7441 8301 -7412 8775
rect -7366 8301 -7353 8775
rect -7441 8288 -7353 8301
rect -3935 8775 -3847 8788
rect -3935 8301 -3922 8775
rect -3876 8301 -3847 8775
rect -3935 8288 -3847 8301
rect -3767 8775 -3663 8788
rect -3767 8301 -3738 8775
rect -3692 8301 -3663 8775
rect -3767 8288 -3663 8301
rect -3583 8775 -3479 8788
rect -3583 8301 -3554 8775
rect -3508 8301 -3479 8775
rect -3583 8288 -3479 8301
rect -3399 8775 -3311 8788
rect -3399 8301 -3370 8775
rect -3324 8301 -3311 8775
rect -3399 8288 -3311 8301
rect 107 8775 195 8788
rect 107 8301 120 8775
rect 166 8301 195 8775
rect 107 8288 195 8301
rect 275 8775 379 8788
rect 275 8301 304 8775
rect 350 8301 379 8775
rect 275 8288 379 8301
rect 459 8775 563 8788
rect 459 8301 488 8775
rect 534 8301 563 8775
rect 459 8288 563 8301
rect 643 8775 731 8788
rect 643 8301 672 8775
rect 718 8301 731 8775
rect 643 8288 731 8301
rect 4149 8775 4237 8788
rect 4149 8301 4162 8775
rect 4208 8301 4237 8775
rect 4149 8288 4237 8301
rect 4317 8775 4421 8788
rect 4317 8301 4346 8775
rect 4392 8301 4421 8775
rect 4317 8288 4421 8301
rect 4501 8775 4605 8788
rect 4501 8301 4530 8775
rect 4576 8301 4605 8775
rect 4501 8288 4605 8301
rect 4685 8775 4773 8788
rect 4685 8301 4714 8775
rect 4760 8301 4773 8775
rect 4685 8288 4773 8301
rect 8191 8775 8279 8788
rect 8191 8301 8204 8775
rect 8250 8301 8279 8775
rect 8191 8288 8279 8301
rect 8359 8775 8463 8788
rect 8359 8301 8388 8775
rect 8434 8301 8463 8775
rect 8359 8288 8463 8301
rect 8543 8775 8647 8788
rect 8543 8301 8572 8775
rect 8618 8301 8647 8775
rect 8543 8288 8647 8301
rect 8727 8775 8815 8788
rect 8727 8301 8756 8775
rect 8802 8301 8815 8775
rect 8727 8288 8815 8301
rect 12233 8775 12321 8788
rect 12233 8301 12246 8775
rect 12292 8301 12321 8775
rect 12233 8288 12321 8301
rect 12401 8775 12505 8788
rect 12401 8301 12430 8775
rect 12476 8301 12505 8775
rect 12401 8288 12505 8301
rect 12585 8775 12689 8788
rect 12585 8301 12614 8775
rect 12660 8301 12689 8775
rect 12585 8288 12689 8301
rect 12769 8775 12857 8788
rect 12769 8301 12798 8775
rect 12844 8301 12857 8775
rect 12769 8288 12857 8301
rect -10931 5167 -10831 5220
rect -10931 4933 -10909 5167
rect -10863 4933 -10831 5167
rect -10931 4880 -10831 4933
rect -10771 5192 -10661 5220
rect -10771 4958 -10739 5192
rect -10693 4958 -10661 5192
rect -10771 4880 -10661 4958
rect -10601 5167 -10491 5220
rect -10601 4933 -10569 5167
rect -10523 4933 -10491 5167
rect -10601 4880 -10491 4933
rect -10431 5192 -10321 5220
rect -10431 4958 -10399 5192
rect -10353 4958 -10321 5192
rect -10431 4880 -10321 4958
rect -10261 5167 -10151 5220
rect -10261 4933 -10229 5167
rect -10183 4933 -10151 5167
rect -10261 4880 -10151 4933
rect -10091 5167 -9991 5220
rect -10091 4933 -10059 5167
rect -10013 4933 -9991 5167
rect -10091 4880 -9991 4933
rect -8519 4854 -8431 4867
rect -8519 4680 -8506 4854
rect -8460 4680 -8431 4854
rect -8519 4667 -8431 4680
rect -8351 4854 -8263 4867
rect -8351 4680 -8322 4854
rect -8276 4680 -8263 4854
rect -8351 4667 -8263 4680
rect -8059 4854 -7971 4867
rect -8059 4680 -8046 4854
rect -8000 4680 -7971 4854
rect -8059 4667 -7971 4680
rect -7891 4854 -7803 4867
rect -7891 4680 -7862 4854
rect -7816 4680 -7803 4854
rect -7891 4667 -7803 4680
rect -9489 4349 -9401 4362
rect -9489 3575 -9476 4349
rect -9430 3575 -9401 4349
rect -9489 3562 -9401 3575
rect -9321 4349 -9233 4362
rect -9321 3575 -9292 4349
rect -9246 3575 -9233 4349
rect -9321 3562 -9233 3575
rect -7089 4349 -7001 4362
rect -7089 3575 -7076 4349
rect -7030 3575 -7001 4349
rect -7089 3562 -7001 3575
rect -6921 4349 -6833 4362
rect -6921 3575 -6892 4349
rect -6846 3575 -6833 4349
rect -6921 3562 -6833 3575
rect -11037 1664 -10949 1677
rect -11037 1530 -11024 1664
rect -10978 1530 -10949 1664
rect -11037 1517 -10949 1530
rect -10869 1664 -10781 1677
rect -10869 1530 -10840 1664
rect -10794 1530 -10781 1664
rect -10869 1517 -10781 1530
rect -10177 1664 -10089 1677
rect -10177 1530 -10164 1664
rect -10118 1530 -10089 1664
rect -10177 1517 -10089 1530
rect -10009 1664 -9921 1677
rect -10009 1530 -9980 1664
rect -9934 1530 -9921 1664
rect -10009 1517 -9921 1530
rect -9717 1684 -9629 1697
rect -9717 1510 -9704 1684
rect -9658 1510 -9629 1684
rect -9717 1497 -9629 1510
rect -9429 1684 -9325 1697
rect -9429 1510 -9400 1684
rect -9354 1510 -9325 1684
rect -9429 1497 -9325 1510
rect -9125 1684 -9021 1697
rect -9125 1510 -9096 1684
rect -9050 1510 -9021 1684
rect -9125 1497 -9021 1510
rect -8821 1684 -8717 1697
rect -8821 1510 -8792 1684
rect -8746 1510 -8717 1684
rect -8821 1497 -8717 1510
rect -8517 1684 -8413 1697
rect -8517 1510 -8488 1684
rect -8442 1510 -8413 1684
rect -8517 1497 -8413 1510
rect -8213 1684 -8109 1697
rect -8213 1510 -8184 1684
rect -8138 1510 -8109 1684
rect -8213 1497 -8109 1510
rect -7909 1684 -7805 1697
rect -7909 1510 -7880 1684
rect -7834 1510 -7805 1684
rect -7909 1497 -7805 1510
rect -7605 1684 -7501 1697
rect -7605 1510 -7576 1684
rect -7530 1510 -7501 1684
rect -7605 1497 -7501 1510
rect -7301 1684 -7197 1697
rect -7301 1510 -7272 1684
rect -7226 1510 -7197 1684
rect -7301 1497 -7197 1510
rect -6997 1684 -6893 1697
rect -6997 1510 -6968 1684
rect -6922 1510 -6893 1684
rect -6997 1497 -6893 1510
rect -6693 1684 -6605 1697
rect -6693 1510 -6664 1684
rect -6618 1510 -6605 1684
rect -6693 1497 -6605 1510
rect -6401 1664 -6313 1677
rect -6401 1530 -6388 1664
rect -6342 1530 -6313 1664
rect -6401 1517 -6313 1530
rect -6233 1664 -6145 1677
rect -6233 1530 -6204 1664
rect -6158 1530 -6145 1664
rect -6233 1517 -6145 1530
rect -5541 1664 -5453 1677
rect -5541 1530 -5528 1664
rect -5482 1530 -5453 1664
rect -5541 1517 -5453 1530
rect -5373 1664 -5285 1677
rect -5373 1530 -5344 1664
rect -5298 1530 -5285 1664
rect -5373 1517 -5285 1530
<< ndiffc >>
rect 39973 38095 40019 38141
rect 40143 38095 40189 38141
rect 40313 38095 40359 38141
rect 40483 38095 40529 38141
rect 40653 38095 40699 38141
rect 40823 38095 40869 38141
rect -4706 35937 -4660 36111
rect -4522 35937 -4476 36111
rect -4338 35937 -4292 36111
rect -4154 35937 -4108 36111
rect 4766 35937 4812 36111
rect 4950 35937 4996 36111
rect 5134 35937 5180 36111
rect 5318 35937 5364 36111
rect 14238 35938 14284 36112
rect 14422 35938 14468 36112
rect 14606 35938 14652 36112
rect 14790 35938 14836 36112
rect 23710 35938 23756 36112
rect 23894 35938 23940 36112
rect 24078 35938 24124 36112
rect 24262 35938 24308 36112
rect 33182 35938 33228 36112
rect 33366 35938 33412 36112
rect 33550 35938 33596 36112
rect 33734 35938 33780 36112
rect 42654 35938 42700 36112
rect 42838 35938 42884 36112
rect 43022 35938 43068 36112
rect 43206 35938 43252 36112
rect -4706 33732 -4660 33906
rect -4522 33732 -4476 33906
rect -4338 33732 -4292 33906
rect -4154 33732 -4108 33906
rect -3220 33732 -3174 33906
rect -3036 33732 -2990 33906
rect -2852 33732 -2806 33906
rect -2668 33732 -2622 33906
rect 4766 33732 4812 33906
rect 4950 33732 4996 33906
rect 5134 33732 5180 33906
rect 5318 33732 5364 33906
rect 6252 33732 6298 33906
rect 6436 33732 6482 33906
rect 6620 33732 6666 33906
rect 6804 33732 6850 33906
rect 14238 33733 14284 33907
rect 14422 33733 14468 33907
rect 14606 33733 14652 33907
rect 14790 33733 14836 33907
rect 15724 33733 15770 33907
rect 15908 33733 15954 33907
rect 16092 33733 16138 33907
rect 16276 33733 16322 33907
rect 23710 33733 23756 33907
rect 23894 33733 23940 33907
rect 24078 33733 24124 33907
rect 24262 33733 24308 33907
rect 25196 33733 25242 33907
rect 25380 33733 25426 33907
rect 25564 33733 25610 33907
rect 25748 33733 25794 33907
rect 33182 33733 33228 33907
rect 33366 33733 33412 33907
rect 33550 33733 33596 33907
rect 33734 33733 33780 33907
rect 34668 33733 34714 33907
rect 34852 33733 34898 33907
rect 35036 33733 35082 33907
rect 35220 33733 35266 33907
rect 42654 33733 42700 33907
rect 42838 33733 42884 33907
rect 43022 33733 43068 33907
rect 43206 33733 43252 33907
rect 44140 33733 44186 33907
rect 44324 33733 44370 33907
rect 44508 33733 44554 33907
rect 44692 33733 44738 33907
rect -4706 31527 -4660 31701
rect -4522 31527 -4476 31701
rect -4338 31527 -4292 31701
rect -4154 31527 -4108 31701
rect -3220 31528 -3174 31702
rect -3036 31528 -2990 31702
rect -2852 31528 -2806 31702
rect -2668 31528 -2622 31702
rect 4766 31527 4812 31701
rect 4950 31527 4996 31701
rect 5134 31527 5180 31701
rect 5318 31527 5364 31701
rect 6252 31528 6298 31702
rect 6436 31528 6482 31702
rect 6620 31528 6666 31702
rect 6804 31528 6850 31702
rect 14238 31528 14284 31702
rect 14422 31528 14468 31702
rect 14606 31528 14652 31702
rect 14790 31528 14836 31702
rect 15724 31529 15770 31703
rect 15908 31529 15954 31703
rect 16092 31529 16138 31703
rect 16276 31529 16322 31703
rect 23710 31528 23756 31702
rect 23894 31528 23940 31702
rect 24078 31528 24124 31702
rect 24262 31528 24308 31702
rect 25196 31529 25242 31703
rect 25380 31529 25426 31703
rect 25564 31529 25610 31703
rect 25748 31529 25794 31703
rect 33182 31528 33228 31702
rect 33366 31528 33412 31702
rect 33550 31528 33596 31702
rect 33734 31528 33780 31702
rect 34668 31529 34714 31703
rect 34852 31529 34898 31703
rect 35036 31529 35082 31703
rect 35220 31529 35266 31703
rect 42654 31528 42700 31702
rect 42838 31528 42884 31702
rect 43022 31528 43068 31702
rect 43206 31528 43252 31702
rect 44140 31529 44186 31703
rect 44324 31529 44370 31703
rect 44508 31529 44554 31703
rect 44692 31529 44738 31703
rect -9848 30452 -9802 30626
rect -9644 30452 -9598 30626
rect -9440 30452 -9394 30626
rect -9164 30452 -9118 30626
rect -8960 30452 -8914 30626
rect -8756 30452 -8710 30626
rect -8480 30452 -8434 30626
rect -8276 30452 -8230 30626
rect -10742 29032 -10696 29206
rect -10538 29032 -10492 29206
rect -7620 29276 -7574 29450
rect -7416 29276 -7370 29450
rect -6936 29276 -6890 29450
rect -6732 29276 -6686 29450
rect -6252 29276 -6206 29450
rect -6048 29276 -6002 29450
rect -4706 29322 -4660 29496
rect -4522 29322 -4476 29496
rect -4338 29322 -4292 29496
rect -4154 29322 -4108 29496
rect -376 30452 -330 30626
rect -172 30452 -126 30626
rect 32 30452 78 30626
rect 308 30452 354 30626
rect 512 30452 558 30626
rect 716 30452 762 30626
rect 992 30452 1038 30626
rect 1196 30452 1242 30626
rect -1270 29032 -1224 29206
rect -1066 29032 -1020 29206
rect 1852 29276 1898 29450
rect 2056 29276 2102 29450
rect 2536 29276 2582 29450
rect 2740 29276 2786 29450
rect 3220 29276 3266 29450
rect 3424 29276 3470 29450
rect 4766 29322 4812 29496
rect 4950 29322 4996 29496
rect 5134 29322 5180 29496
rect 5318 29322 5364 29496
rect 9096 30453 9142 30627
rect 9300 30453 9346 30627
rect 9504 30453 9550 30627
rect 9780 30453 9826 30627
rect 9984 30453 10030 30627
rect 10188 30453 10234 30627
rect 10464 30453 10510 30627
rect 10668 30453 10714 30627
rect 8202 29033 8248 29207
rect 8406 29033 8452 29207
rect 11324 29277 11370 29451
rect 11528 29277 11574 29451
rect 12008 29277 12054 29451
rect 12212 29277 12258 29451
rect 12692 29277 12738 29451
rect 12896 29277 12942 29451
rect 14238 29323 14284 29497
rect 14422 29323 14468 29497
rect 14606 29323 14652 29497
rect 14790 29323 14836 29497
rect 18568 30453 18614 30627
rect 18772 30453 18818 30627
rect 18976 30453 19022 30627
rect 19252 30453 19298 30627
rect 19456 30453 19502 30627
rect 19660 30453 19706 30627
rect 19936 30453 19982 30627
rect 20140 30453 20186 30627
rect 17674 29033 17720 29207
rect 17878 29033 17924 29207
rect 20796 29277 20842 29451
rect 21000 29277 21046 29451
rect 21480 29277 21526 29451
rect 21684 29277 21730 29451
rect 22164 29277 22210 29451
rect 22368 29277 22414 29451
rect 23710 29323 23756 29497
rect 23894 29323 23940 29497
rect 24078 29323 24124 29497
rect 24262 29323 24308 29497
rect 28040 30453 28086 30627
rect 28244 30453 28290 30627
rect 28448 30453 28494 30627
rect 28724 30453 28770 30627
rect 28928 30453 28974 30627
rect 29132 30453 29178 30627
rect 29408 30453 29454 30627
rect 29612 30453 29658 30627
rect 27146 29033 27192 29207
rect 27350 29033 27396 29207
rect 30268 29277 30314 29451
rect 30472 29277 30518 29451
rect 30952 29277 30998 29451
rect 31156 29277 31202 29451
rect 31636 29277 31682 29451
rect 31840 29277 31886 29451
rect 33182 29323 33228 29497
rect 33366 29323 33412 29497
rect 33550 29323 33596 29497
rect 33734 29323 33780 29497
rect 37512 30453 37558 30627
rect 37716 30453 37762 30627
rect 37920 30453 37966 30627
rect 38196 30453 38242 30627
rect 38400 30453 38446 30627
rect 38604 30453 38650 30627
rect 38880 30453 38926 30627
rect 39084 30453 39130 30627
rect 36618 29033 36664 29207
rect 36822 29033 36868 29207
rect 39740 29277 39786 29451
rect 39944 29277 39990 29451
rect 40424 29277 40470 29451
rect 40628 29277 40674 29451
rect 41108 29277 41154 29451
rect 41312 29277 41358 29451
rect 42654 29323 42700 29497
rect 42838 29323 42884 29497
rect 43022 29323 43068 29497
rect 43206 29323 43252 29497
rect -9848 28112 -9802 28286
rect -9644 28112 -9598 28286
rect -9440 28112 -9394 28286
rect -9164 28112 -9118 28286
rect -8960 28112 -8914 28286
rect -8756 28112 -8710 28286
rect -8480 28112 -8434 28286
rect -8276 28112 -8230 28286
rect -376 28112 -330 28286
rect -172 28112 -126 28286
rect 32 28112 78 28286
rect 308 28112 354 28286
rect 512 28112 558 28286
rect 716 28112 762 28286
rect 992 28112 1038 28286
rect 1196 28112 1242 28286
rect 9096 28113 9142 28287
rect 9300 28113 9346 28287
rect 9504 28113 9550 28287
rect 9780 28113 9826 28287
rect 9984 28113 10030 28287
rect 10188 28113 10234 28287
rect 10464 28113 10510 28287
rect 10668 28113 10714 28287
rect 18568 28113 18614 28287
rect 18772 28113 18818 28287
rect 18976 28113 19022 28287
rect 19252 28113 19298 28287
rect 19456 28113 19502 28287
rect 19660 28113 19706 28287
rect 19936 28113 19982 28287
rect 20140 28113 20186 28287
rect 28040 28113 28086 28287
rect 28244 28113 28290 28287
rect 28448 28113 28494 28287
rect 28724 28113 28770 28287
rect 28928 28113 28974 28287
rect 29132 28113 29178 28287
rect 29408 28113 29454 28287
rect 29612 28113 29658 28287
rect 37512 28113 37558 28287
rect 37716 28113 37762 28287
rect 37920 28113 37966 28287
rect 38196 28113 38242 28287
rect 38400 28113 38446 28287
rect 38604 28113 38650 28287
rect 38880 28113 38926 28287
rect 39084 28113 39130 28287
rect -12455 27102 -12409 27276
rect -12251 27102 -12205 27276
rect -7964 23635 -7918 23809
rect -7780 23635 -7734 23809
rect -7596 23635 -7550 23809
rect -7412 23635 -7366 23809
rect -3922 23632 -3876 23806
rect -3738 23632 -3692 23806
rect -3554 23632 -3508 23806
rect -3370 23632 -3324 23806
rect 120 23632 166 23806
rect 304 23632 350 23806
rect 488 23632 534 23806
rect 672 23632 718 23806
rect 4162 23632 4208 23806
rect 4346 23632 4392 23806
rect 4530 23632 4576 23806
rect 4714 23632 4760 23806
rect 8204 23632 8250 23806
rect 8388 23632 8434 23806
rect 8572 23632 8618 23806
rect 8756 23632 8802 23806
rect 12246 23632 12292 23806
rect 12430 23632 12476 23806
rect 12614 23632 12660 23806
rect 12798 23632 12844 23806
rect 16288 23632 16334 23806
rect 16472 23632 16518 23806
rect 16656 23632 16702 23806
rect 16840 23632 16886 23806
rect -7964 21430 -7918 21604
rect -7780 21430 -7734 21604
rect -7596 21430 -7550 21604
rect -7412 21430 -7366 21604
rect -6478 21430 -6432 21604
rect -6294 21430 -6248 21604
rect -6110 21430 -6064 21604
rect -5926 21430 -5880 21604
rect -3922 21427 -3876 21601
rect -3738 21427 -3692 21601
rect -3554 21427 -3508 21601
rect -3370 21427 -3324 21601
rect -2436 21427 -2390 21601
rect -2252 21427 -2206 21601
rect -2068 21427 -2022 21601
rect -1884 21427 -1838 21601
rect 120 21427 166 21601
rect 304 21427 350 21601
rect 488 21427 534 21601
rect 672 21427 718 21601
rect 1606 21427 1652 21601
rect 1790 21427 1836 21601
rect 1974 21427 2020 21601
rect 2158 21427 2204 21601
rect 4162 21427 4208 21601
rect 4346 21427 4392 21601
rect 4530 21427 4576 21601
rect 4714 21427 4760 21601
rect 5648 21427 5694 21601
rect 5832 21427 5878 21601
rect 6016 21427 6062 21601
rect 6200 21427 6246 21601
rect 8204 21427 8250 21601
rect 8388 21427 8434 21601
rect 8572 21427 8618 21601
rect 8756 21427 8802 21601
rect 9690 21427 9736 21601
rect 9874 21427 9920 21601
rect 10058 21427 10104 21601
rect 10242 21427 10288 21601
rect 12246 21427 12292 21601
rect 12430 21427 12476 21601
rect 12614 21427 12660 21601
rect 12798 21427 12844 21601
rect 13732 21427 13778 21601
rect 13916 21427 13962 21601
rect 14100 21427 14146 21601
rect 14284 21427 14330 21601
rect 16288 21427 16334 21601
rect 16472 21427 16518 21601
rect 16656 21427 16702 21601
rect 16840 21427 16886 21601
rect 17774 21427 17820 21601
rect 17958 21427 18004 21601
rect 18142 21427 18188 21601
rect 18326 21427 18372 21601
rect -7964 19225 -7918 19399
rect -7780 19225 -7734 19399
rect -7596 19225 -7550 19399
rect -7412 19225 -7366 19399
rect -6478 19226 -6432 19400
rect -6294 19226 -6248 19400
rect -6110 19226 -6064 19400
rect -5926 19226 -5880 19400
rect -3922 19222 -3876 19396
rect -3738 19222 -3692 19396
rect -3554 19222 -3508 19396
rect -3370 19222 -3324 19396
rect -2436 19223 -2390 19397
rect -2252 19223 -2206 19397
rect -2068 19223 -2022 19397
rect -1884 19223 -1838 19397
rect 120 19222 166 19396
rect 304 19222 350 19396
rect 488 19222 534 19396
rect 672 19222 718 19396
rect 1606 19223 1652 19397
rect 1790 19223 1836 19397
rect 1974 19223 2020 19397
rect 2158 19223 2204 19397
rect 4162 19222 4208 19396
rect 4346 19222 4392 19396
rect 4530 19222 4576 19396
rect 4714 19222 4760 19396
rect 5648 19223 5694 19397
rect 5832 19223 5878 19397
rect 6016 19223 6062 19397
rect 6200 19223 6246 19397
rect 8204 19222 8250 19396
rect 8388 19222 8434 19396
rect 8572 19222 8618 19396
rect 8756 19222 8802 19396
rect 9690 19223 9736 19397
rect 9874 19223 9920 19397
rect 10058 19223 10104 19397
rect 10242 19223 10288 19397
rect 12246 19222 12292 19396
rect 12430 19222 12476 19396
rect 12614 19222 12660 19396
rect 12798 19222 12844 19396
rect 13732 19223 13778 19397
rect 13916 19223 13962 19397
rect 14100 19223 14146 19397
rect 14284 19223 14330 19397
rect 16288 19222 16334 19396
rect 16472 19222 16518 19396
rect 16656 19222 16702 19396
rect 16840 19222 16886 19396
rect 17774 19223 17820 19397
rect 17958 19223 18004 19397
rect 18142 19223 18188 19397
rect 18326 19223 18372 19397
rect -7964 17020 -7918 17194
rect -7780 17020 -7734 17194
rect -7596 17020 -7550 17194
rect -7412 17020 -7366 17194
rect -3922 17017 -3876 17191
rect -3738 17017 -3692 17191
rect -3554 17017 -3508 17191
rect -3370 17017 -3324 17191
rect 120 17017 166 17191
rect 304 17017 350 17191
rect 488 17017 534 17191
rect 672 17017 718 17191
rect 4162 17017 4208 17191
rect 4346 17017 4392 17191
rect 4530 17017 4576 17191
rect 4714 17017 4760 17191
rect 8204 17017 8250 17191
rect 8388 17017 8434 17191
rect 8572 17017 8618 17191
rect 8756 17017 8802 17191
rect 12246 17017 12292 17191
rect 12430 17017 12476 17191
rect 12614 17017 12660 17191
rect 12798 17017 12844 17191
rect 16288 17017 16334 17191
rect 16472 17017 16518 17191
rect 16656 17017 16702 17191
rect 16840 17017 16886 17191
rect -11976 14056 -11930 14230
rect -11792 14056 -11746 14230
rect -11608 14056 -11562 14230
rect -11424 14056 -11378 14230
rect -7964 14056 -7918 14230
rect -7780 14056 -7734 14230
rect -7596 14056 -7550 14230
rect -7412 14056 -7366 14230
rect -3922 14056 -3876 14230
rect -3738 14056 -3692 14230
rect -3554 14056 -3508 14230
rect -3370 14056 -3324 14230
rect 120 14056 166 14230
rect 304 14056 350 14230
rect 488 14056 534 14230
rect 672 14056 718 14230
rect 4162 14056 4208 14230
rect 4346 14056 4392 14230
rect 4530 14056 4576 14230
rect 4714 14056 4760 14230
rect 8204 14056 8250 14230
rect 8388 14056 8434 14230
rect 8572 14056 8618 14230
rect 8756 14056 8802 14230
rect 12246 14056 12292 14230
rect 12430 14056 12476 14230
rect 12614 14056 12660 14230
rect 12798 14056 12844 14230
rect -11976 11851 -11930 12025
rect -11792 11851 -11746 12025
rect -11608 11851 -11562 12025
rect -11424 11851 -11378 12025
rect -10490 11851 -10444 12025
rect -10306 11851 -10260 12025
rect -10122 11851 -10076 12025
rect -9938 11851 -9892 12025
rect -7964 11851 -7918 12025
rect -7780 11851 -7734 12025
rect -7596 11851 -7550 12025
rect -7412 11851 -7366 12025
rect -6478 11851 -6432 12025
rect -6294 11851 -6248 12025
rect -6110 11851 -6064 12025
rect -5926 11851 -5880 12025
rect -3922 11851 -3876 12025
rect -3738 11851 -3692 12025
rect -3554 11851 -3508 12025
rect -3370 11851 -3324 12025
rect -2436 11851 -2390 12025
rect -2252 11851 -2206 12025
rect -2068 11851 -2022 12025
rect -1884 11851 -1838 12025
rect 120 11851 166 12025
rect 304 11851 350 12025
rect 488 11851 534 12025
rect 672 11851 718 12025
rect 1606 11851 1652 12025
rect 1790 11851 1836 12025
rect 1974 11851 2020 12025
rect 2158 11851 2204 12025
rect 4162 11851 4208 12025
rect 4346 11851 4392 12025
rect 4530 11851 4576 12025
rect 4714 11851 4760 12025
rect 5648 11851 5694 12025
rect 5832 11851 5878 12025
rect 6016 11851 6062 12025
rect 6200 11851 6246 12025
rect 8204 11851 8250 12025
rect 8388 11851 8434 12025
rect 8572 11851 8618 12025
rect 8756 11851 8802 12025
rect 9690 11851 9736 12025
rect 9874 11851 9920 12025
rect 10058 11851 10104 12025
rect 10242 11851 10288 12025
rect 12246 11851 12292 12025
rect 12430 11851 12476 12025
rect 12614 11851 12660 12025
rect 12798 11851 12844 12025
rect 13732 11851 13778 12025
rect 13916 11851 13962 12025
rect 14100 11851 14146 12025
rect 14284 11851 14330 12025
rect -11976 9646 -11930 9820
rect -11792 9646 -11746 9820
rect -11608 9646 -11562 9820
rect -11424 9646 -11378 9820
rect -10490 9647 -10444 9821
rect -10306 9647 -10260 9821
rect -10122 9647 -10076 9821
rect -9938 9647 -9892 9821
rect -7964 9646 -7918 9820
rect -7780 9646 -7734 9820
rect -7596 9646 -7550 9820
rect -7412 9646 -7366 9820
rect -6478 9647 -6432 9821
rect -6294 9647 -6248 9821
rect -6110 9647 -6064 9821
rect -5926 9647 -5880 9821
rect -3922 9646 -3876 9820
rect -3738 9646 -3692 9820
rect -3554 9646 -3508 9820
rect -3370 9646 -3324 9820
rect -2436 9647 -2390 9821
rect -2252 9647 -2206 9821
rect -2068 9647 -2022 9821
rect -1884 9647 -1838 9821
rect 120 9646 166 9820
rect 304 9646 350 9820
rect 488 9646 534 9820
rect 672 9646 718 9820
rect 1606 9647 1652 9821
rect 1790 9647 1836 9821
rect 1974 9647 2020 9821
rect 2158 9647 2204 9821
rect 4162 9646 4208 9820
rect 4346 9646 4392 9820
rect 4530 9646 4576 9820
rect 4714 9646 4760 9820
rect 5648 9647 5694 9821
rect 5832 9647 5878 9821
rect 6016 9647 6062 9821
rect 6200 9647 6246 9821
rect 8204 9646 8250 9820
rect 8388 9646 8434 9820
rect 8572 9646 8618 9820
rect 8756 9646 8802 9820
rect 9690 9647 9736 9821
rect 9874 9647 9920 9821
rect 10058 9647 10104 9821
rect 10242 9647 10288 9821
rect 12246 9646 12292 9820
rect 12430 9646 12476 9820
rect 12614 9646 12660 9820
rect 12798 9646 12844 9820
rect 13732 9647 13778 9821
rect 13916 9647 13962 9821
rect 14100 9647 14146 9821
rect 14284 9647 14330 9821
rect -11976 7441 -11930 7615
rect -11792 7441 -11746 7615
rect -11608 7441 -11562 7615
rect -11424 7441 -11378 7615
rect -7964 7441 -7918 7615
rect -7780 7441 -7734 7615
rect -7596 7441 -7550 7615
rect -7412 7441 -7366 7615
rect -3922 7441 -3876 7615
rect -3738 7441 -3692 7615
rect -3554 7441 -3508 7615
rect -3370 7441 -3324 7615
rect 120 7441 166 7615
rect 304 7441 350 7615
rect 488 7441 534 7615
rect 672 7441 718 7615
rect 4162 7441 4208 7615
rect 4346 7441 4392 7615
rect 4530 7441 4576 7615
rect 4714 7441 4760 7615
rect 8204 7441 8250 7615
rect 8388 7441 8434 7615
rect 8572 7441 8618 7615
rect 8756 7441 8802 7615
rect 12246 7441 12292 7615
rect 12430 7441 12476 7615
rect 12614 7441 12660 7615
rect 12798 7441 12844 7615
rect -10909 4432 -10863 4478
rect -10739 4432 -10693 4478
rect -10569 4432 -10523 4478
rect -10399 4432 -10353 4478
rect -10229 4432 -10183 4478
rect -10059 4432 -10013 4478
rect -8506 3860 -8460 4034
rect -8322 3860 -8276 4034
rect -8046 3860 -8000 4034
rect -7862 3860 -7816 4034
rect -9476 2727 -9430 3101
rect -9292 2727 -9246 3101
rect -7076 2727 -7030 3101
rect -6892 2727 -6846 3101
rect -9842 354 -9796 728
rect -9538 354 -9492 728
rect -9234 354 -9188 728
rect -8930 354 -8884 728
rect -8626 354 -8580 728
rect -8322 354 -8276 728
rect -8046 354 -8000 728
rect -7742 354 -7696 728
rect -7438 354 -7392 728
rect -7134 354 -7088 728
rect -6830 354 -6784 728
rect -6526 354 -6480 728
rect -10008 -1031 -9962 -757
rect -9704 -1031 -9658 -757
rect -9400 -1031 -9354 -757
rect -9096 -1031 -9050 -757
rect -8792 -1031 -8746 -757
rect -8488 -1031 -8442 -757
rect -8184 -1031 -8138 -757
rect -7880 -1031 -7834 -757
rect -7576 -1031 -7530 -757
rect -7272 -1031 -7226 -757
rect -6968 -1031 -6922 -757
rect -6664 -1031 -6618 -757
rect -6360 -1031 -6314 -757
rect -10008 -1994 -9962 -1720
rect -9704 -1994 -9658 -1720
rect -9400 -1994 -9354 -1720
rect -9096 -1994 -9050 -1720
rect -8792 -1994 -8746 -1720
rect -8488 -1994 -8442 -1720
rect -8184 -1994 -8138 -1720
rect -7880 -1994 -7834 -1720
rect -7576 -1994 -7530 -1720
rect -7272 -1994 -7226 -1720
rect -6968 -1994 -6922 -1720
rect -6664 -1994 -6618 -1720
rect -6360 -1994 -6314 -1720
rect -8460 -2780 -8414 -2646
rect -8276 -2780 -8230 -2646
rect -8092 -2780 -8046 -2646
rect -7908 -2780 -7862 -2646
<< pdiffc >>
rect 39973 38596 40019 38830
rect 40143 38621 40189 38855
rect 40313 38596 40359 38830
rect 40483 38621 40529 38855
rect 40653 38596 40699 38830
rect 40823 38596 40869 38830
rect -4706 36797 -4660 37271
rect -4522 36797 -4476 37271
rect -4338 36797 -4292 37271
rect -4154 36797 -4108 37271
rect 4766 36797 4812 37271
rect 4950 36797 4996 37271
rect 5134 36797 5180 37271
rect 5318 36797 5364 37271
rect 14238 36798 14284 37272
rect 14422 36798 14468 37272
rect 14606 36798 14652 37272
rect 14790 36798 14836 37272
rect 23710 36798 23756 37272
rect 23894 36798 23940 37272
rect 24078 36798 24124 37272
rect 24262 36798 24308 37272
rect 33182 36798 33228 37272
rect 33366 36798 33412 37272
rect 33550 36798 33596 37272
rect 33734 36798 33780 37272
rect 42654 36798 42700 37272
rect 42838 36798 42884 37272
rect 43022 36798 43068 37272
rect 43206 36798 43252 37272
rect -4706 34592 -4660 35066
rect -4522 34592 -4476 35066
rect -4338 34592 -4292 35066
rect -4154 34592 -4108 35066
rect -3220 34592 -3174 35066
rect -3036 34592 -2990 35066
rect -2852 34592 -2806 35066
rect -2668 34592 -2622 35066
rect 4766 34592 4812 35066
rect 4950 34592 4996 35066
rect 5134 34592 5180 35066
rect 5318 34592 5364 35066
rect 6252 34592 6298 35066
rect 6436 34592 6482 35066
rect 6620 34592 6666 35066
rect 6804 34592 6850 35066
rect 14238 34593 14284 35067
rect 14422 34593 14468 35067
rect 14606 34593 14652 35067
rect 14790 34593 14836 35067
rect 15724 34593 15770 35067
rect 15908 34593 15954 35067
rect 16092 34593 16138 35067
rect 16276 34593 16322 35067
rect 23710 34593 23756 35067
rect 23894 34593 23940 35067
rect 24078 34593 24124 35067
rect 24262 34593 24308 35067
rect 25196 34593 25242 35067
rect 25380 34593 25426 35067
rect 25564 34593 25610 35067
rect 25748 34593 25794 35067
rect 33182 34593 33228 35067
rect 33366 34593 33412 35067
rect 33550 34593 33596 35067
rect 33734 34593 33780 35067
rect 34668 34593 34714 35067
rect 34852 34593 34898 35067
rect 35036 34593 35082 35067
rect 35220 34593 35266 35067
rect 42654 34593 42700 35067
rect 42838 34593 42884 35067
rect 43022 34593 43068 35067
rect 43206 34593 43252 35067
rect 44140 34593 44186 35067
rect 44324 34593 44370 35067
rect 44508 34593 44554 35067
rect 44692 34593 44738 35067
rect -4706 32387 -4660 32861
rect -4522 32387 -4476 32861
rect -4338 32387 -4292 32861
rect -4154 32387 -4108 32861
rect -3220 32388 -3174 32862
rect -3036 32388 -2990 32862
rect -2852 32388 -2806 32862
rect -2668 32388 -2622 32862
rect 4766 32387 4812 32861
rect 4950 32387 4996 32861
rect 5134 32387 5180 32861
rect 5318 32387 5364 32861
rect 6252 32388 6298 32862
rect 6436 32388 6482 32862
rect 6620 32388 6666 32862
rect 6804 32388 6850 32862
rect 14238 32388 14284 32862
rect 14422 32388 14468 32862
rect 14606 32388 14652 32862
rect 14790 32388 14836 32862
rect 15724 32389 15770 32863
rect 15908 32389 15954 32863
rect 16092 32389 16138 32863
rect 16276 32389 16322 32863
rect 23710 32388 23756 32862
rect 23894 32388 23940 32862
rect 24078 32388 24124 32862
rect 24262 32388 24308 32862
rect 25196 32389 25242 32863
rect 25380 32389 25426 32863
rect 25564 32389 25610 32863
rect 25748 32389 25794 32863
rect 33182 32388 33228 32862
rect 33366 32388 33412 32862
rect 33550 32388 33596 32862
rect 33734 32388 33780 32862
rect 34668 32389 34714 32863
rect 34852 32389 34898 32863
rect 35036 32389 35082 32863
rect 35220 32389 35266 32863
rect 42654 32388 42700 32862
rect 42838 32388 42884 32862
rect 43022 32388 43068 32862
rect 43206 32388 43252 32862
rect 44140 32389 44186 32863
rect 44324 32389 44370 32863
rect 44508 32389 44554 32863
rect 44692 32389 44738 32863
rect -9848 31172 -9802 31746
rect -9644 31172 -9598 31746
rect -8960 31172 -8914 31746
rect -8756 31172 -8710 31746
rect -8480 31172 -8434 31746
rect -8276 31172 -8230 31746
rect -376 31172 -330 31746
rect -172 31172 -126 31746
rect 512 31172 558 31746
rect 716 31172 762 31746
rect 992 31172 1038 31746
rect 1196 31172 1242 31746
rect 9096 31173 9142 31747
rect 9300 31173 9346 31747
rect 9984 31173 10030 31747
rect 10188 31173 10234 31747
rect 10464 31173 10510 31747
rect 10668 31173 10714 31747
rect 18568 31173 18614 31747
rect 18772 31173 18818 31747
rect 19456 31173 19502 31747
rect 19660 31173 19706 31747
rect 19936 31173 19982 31747
rect 20140 31173 20186 31747
rect 28040 31173 28086 31747
rect 28244 31173 28290 31747
rect 28928 31173 28974 31747
rect 29132 31173 29178 31747
rect 29408 31173 29454 31747
rect 29612 31173 29658 31747
rect 37512 31173 37558 31747
rect 37716 31173 37762 31747
rect 38400 31173 38446 31747
rect 38604 31173 38650 31747
rect 38880 31173 38926 31747
rect 39084 31173 39130 31747
rect -10742 29752 -10696 30326
rect -10538 29752 -10492 30326
rect -7620 29996 -7574 30570
rect -7416 29996 -7370 30570
rect -7212 29996 -7166 30570
rect -6936 29996 -6890 30570
rect -6732 29996 -6686 30570
rect -6528 29996 -6482 30570
rect -6252 29996 -6206 30570
rect -6048 29996 -6002 30570
rect -4706 30182 -4660 30656
rect -4522 30182 -4476 30656
rect -4338 30182 -4292 30656
rect -4154 30182 -4108 30656
rect -9848 28832 -9802 29406
rect -9644 28832 -9598 29406
rect -8960 28832 -8914 29406
rect -8756 28832 -8710 29406
rect -8480 28832 -8434 29406
rect -8276 28832 -8230 29406
rect -1270 29752 -1224 30326
rect -1066 29752 -1020 30326
rect 1852 29996 1898 30570
rect 2056 29996 2102 30570
rect 2260 29996 2306 30570
rect 2536 29996 2582 30570
rect 2740 29996 2786 30570
rect 2944 29996 2990 30570
rect 3220 29996 3266 30570
rect 3424 29996 3470 30570
rect 4766 30182 4812 30656
rect 4950 30182 4996 30656
rect 5134 30182 5180 30656
rect 5318 30182 5364 30656
rect -376 28832 -330 29406
rect -172 28832 -126 29406
rect 512 28832 558 29406
rect 716 28832 762 29406
rect 992 28832 1038 29406
rect 1196 28832 1242 29406
rect 8202 29753 8248 30327
rect 8406 29753 8452 30327
rect 11324 29997 11370 30571
rect 11528 29997 11574 30571
rect 11732 29997 11778 30571
rect 12008 29997 12054 30571
rect 12212 29997 12258 30571
rect 12416 29997 12462 30571
rect 12692 29997 12738 30571
rect 12896 29997 12942 30571
rect 14238 30183 14284 30657
rect 14422 30183 14468 30657
rect 14606 30183 14652 30657
rect 14790 30183 14836 30657
rect 9096 28833 9142 29407
rect 9300 28833 9346 29407
rect 9984 28833 10030 29407
rect 10188 28833 10234 29407
rect 10464 28833 10510 29407
rect 10668 28833 10714 29407
rect 17674 29753 17720 30327
rect 17878 29753 17924 30327
rect 20796 29997 20842 30571
rect 21000 29997 21046 30571
rect 21204 29997 21250 30571
rect 21480 29997 21526 30571
rect 21684 29997 21730 30571
rect 21888 29997 21934 30571
rect 22164 29997 22210 30571
rect 22368 29997 22414 30571
rect 23710 30183 23756 30657
rect 23894 30183 23940 30657
rect 24078 30183 24124 30657
rect 24262 30183 24308 30657
rect 18568 28833 18614 29407
rect 18772 28833 18818 29407
rect 19456 28833 19502 29407
rect 19660 28833 19706 29407
rect 19936 28833 19982 29407
rect 20140 28833 20186 29407
rect 27146 29753 27192 30327
rect 27350 29753 27396 30327
rect 30268 29997 30314 30571
rect 30472 29997 30518 30571
rect 30676 29997 30722 30571
rect 30952 29997 30998 30571
rect 31156 29997 31202 30571
rect 31360 29997 31406 30571
rect 31636 29997 31682 30571
rect 31840 29997 31886 30571
rect 33182 30183 33228 30657
rect 33366 30183 33412 30657
rect 33550 30183 33596 30657
rect 33734 30183 33780 30657
rect 28040 28833 28086 29407
rect 28244 28833 28290 29407
rect 28928 28833 28974 29407
rect 29132 28833 29178 29407
rect 29408 28833 29454 29407
rect 29612 28833 29658 29407
rect 36618 29753 36664 30327
rect 36822 29753 36868 30327
rect 39740 29997 39786 30571
rect 39944 29997 39990 30571
rect 40148 29997 40194 30571
rect 40424 29997 40470 30571
rect 40628 29997 40674 30571
rect 40832 29997 40878 30571
rect 41108 29997 41154 30571
rect 41312 29997 41358 30571
rect 42654 30183 42700 30657
rect 42838 30183 42884 30657
rect 43022 30183 43068 30657
rect 43206 30183 43252 30657
rect 37512 28833 37558 29407
rect 37716 28833 37762 29407
rect 38400 28833 38446 29407
rect 38604 28833 38650 29407
rect 38880 28833 38926 29407
rect 39084 28833 39130 29407
rect -12455 27822 -12409 28396
rect -12251 27822 -12205 28396
rect -7964 24495 -7918 24969
rect -7780 24495 -7734 24969
rect -7596 24495 -7550 24969
rect -7412 24495 -7366 24969
rect -3922 24492 -3876 24966
rect -3738 24492 -3692 24966
rect -3554 24492 -3508 24966
rect -3370 24492 -3324 24966
rect 120 24492 166 24966
rect 304 24492 350 24966
rect 488 24492 534 24966
rect 672 24492 718 24966
rect 4162 24492 4208 24966
rect 4346 24492 4392 24966
rect 4530 24492 4576 24966
rect 4714 24492 4760 24966
rect 8204 24492 8250 24966
rect 8388 24492 8434 24966
rect 8572 24492 8618 24966
rect 8756 24492 8802 24966
rect 12246 24492 12292 24966
rect 12430 24492 12476 24966
rect 12614 24492 12660 24966
rect 12798 24492 12844 24966
rect 16288 24492 16334 24966
rect 16472 24492 16518 24966
rect 16656 24492 16702 24966
rect 16840 24492 16886 24966
rect -7964 22290 -7918 22764
rect -7780 22290 -7734 22764
rect -7596 22290 -7550 22764
rect -7412 22290 -7366 22764
rect -6478 22290 -6432 22764
rect -6294 22290 -6248 22764
rect -6110 22290 -6064 22764
rect -5926 22290 -5880 22764
rect -3922 22287 -3876 22761
rect -3738 22287 -3692 22761
rect -3554 22287 -3508 22761
rect -3370 22287 -3324 22761
rect -2436 22287 -2390 22761
rect -2252 22287 -2206 22761
rect -2068 22287 -2022 22761
rect -1884 22287 -1838 22761
rect 120 22287 166 22761
rect 304 22287 350 22761
rect 488 22287 534 22761
rect 672 22287 718 22761
rect 1606 22287 1652 22761
rect 1790 22287 1836 22761
rect 1974 22287 2020 22761
rect 2158 22287 2204 22761
rect 4162 22287 4208 22761
rect 4346 22287 4392 22761
rect 4530 22287 4576 22761
rect 4714 22287 4760 22761
rect 5648 22287 5694 22761
rect 5832 22287 5878 22761
rect 6016 22287 6062 22761
rect 6200 22287 6246 22761
rect 8204 22287 8250 22761
rect 8388 22287 8434 22761
rect 8572 22287 8618 22761
rect 8756 22287 8802 22761
rect 9690 22287 9736 22761
rect 9874 22287 9920 22761
rect 10058 22287 10104 22761
rect 10242 22287 10288 22761
rect 12246 22287 12292 22761
rect 12430 22287 12476 22761
rect 12614 22287 12660 22761
rect 12798 22287 12844 22761
rect 13732 22287 13778 22761
rect 13916 22287 13962 22761
rect 14100 22287 14146 22761
rect 14284 22287 14330 22761
rect 16288 22287 16334 22761
rect 16472 22287 16518 22761
rect 16656 22287 16702 22761
rect 16840 22287 16886 22761
rect 17774 22287 17820 22761
rect 17958 22287 18004 22761
rect 18142 22287 18188 22761
rect 18326 22287 18372 22761
rect -7964 20085 -7918 20559
rect -7780 20085 -7734 20559
rect -7596 20085 -7550 20559
rect -7412 20085 -7366 20559
rect -6478 20086 -6432 20560
rect -6294 20086 -6248 20560
rect -6110 20086 -6064 20560
rect -5926 20086 -5880 20560
rect -3922 20082 -3876 20556
rect -3738 20082 -3692 20556
rect -3554 20082 -3508 20556
rect -3370 20082 -3324 20556
rect -2436 20083 -2390 20557
rect -2252 20083 -2206 20557
rect -2068 20083 -2022 20557
rect -1884 20083 -1838 20557
rect 120 20082 166 20556
rect 304 20082 350 20556
rect 488 20082 534 20556
rect 672 20082 718 20556
rect 1606 20083 1652 20557
rect 1790 20083 1836 20557
rect 1974 20083 2020 20557
rect 2158 20083 2204 20557
rect 4162 20082 4208 20556
rect 4346 20082 4392 20556
rect 4530 20082 4576 20556
rect 4714 20082 4760 20556
rect 5648 20083 5694 20557
rect 5832 20083 5878 20557
rect 6016 20083 6062 20557
rect 6200 20083 6246 20557
rect 8204 20082 8250 20556
rect 8388 20082 8434 20556
rect 8572 20082 8618 20556
rect 8756 20082 8802 20556
rect 9690 20083 9736 20557
rect 9874 20083 9920 20557
rect 10058 20083 10104 20557
rect 10242 20083 10288 20557
rect 12246 20082 12292 20556
rect 12430 20082 12476 20556
rect 12614 20082 12660 20556
rect 12798 20082 12844 20556
rect 13732 20083 13778 20557
rect 13916 20083 13962 20557
rect 14100 20083 14146 20557
rect 14284 20083 14330 20557
rect 16288 20082 16334 20556
rect 16472 20082 16518 20556
rect 16656 20082 16702 20556
rect 16840 20082 16886 20556
rect 17774 20083 17820 20557
rect 17958 20083 18004 20557
rect 18142 20083 18188 20557
rect 18326 20083 18372 20557
rect -7964 17880 -7918 18354
rect -7780 17880 -7734 18354
rect -7596 17880 -7550 18354
rect -7412 17880 -7366 18354
rect -3922 17877 -3876 18351
rect -3738 17877 -3692 18351
rect -3554 17877 -3508 18351
rect -3370 17877 -3324 18351
rect 120 17877 166 18351
rect 304 17877 350 18351
rect 488 17877 534 18351
rect 672 17877 718 18351
rect 4162 17877 4208 18351
rect 4346 17877 4392 18351
rect 4530 17877 4576 18351
rect 4714 17877 4760 18351
rect 8204 17877 8250 18351
rect 8388 17877 8434 18351
rect 8572 17877 8618 18351
rect 8756 17877 8802 18351
rect 12246 17877 12292 18351
rect 12430 17877 12476 18351
rect 12614 17877 12660 18351
rect 12798 17877 12844 18351
rect 16288 17877 16334 18351
rect 16472 17877 16518 18351
rect 16656 17877 16702 18351
rect 16840 17877 16886 18351
rect -11976 14916 -11930 15390
rect -11792 14916 -11746 15390
rect -11608 14916 -11562 15390
rect -11424 14916 -11378 15390
rect -7964 14916 -7918 15390
rect -7780 14916 -7734 15390
rect -7596 14916 -7550 15390
rect -7412 14916 -7366 15390
rect -3922 14916 -3876 15390
rect -3738 14916 -3692 15390
rect -3554 14916 -3508 15390
rect -3370 14916 -3324 15390
rect 120 14916 166 15390
rect 304 14916 350 15390
rect 488 14916 534 15390
rect 672 14916 718 15390
rect 4162 14916 4208 15390
rect 4346 14916 4392 15390
rect 4530 14916 4576 15390
rect 4714 14916 4760 15390
rect 8204 14916 8250 15390
rect 8388 14916 8434 15390
rect 8572 14916 8618 15390
rect 8756 14916 8802 15390
rect 12246 14916 12292 15390
rect 12430 14916 12476 15390
rect 12614 14916 12660 15390
rect 12798 14916 12844 15390
rect -11976 12711 -11930 13185
rect -11792 12711 -11746 13185
rect -11608 12711 -11562 13185
rect -11424 12711 -11378 13185
rect -10490 12711 -10444 13185
rect -10306 12711 -10260 13185
rect -10122 12711 -10076 13185
rect -9938 12711 -9892 13185
rect -7964 12711 -7918 13185
rect -7780 12711 -7734 13185
rect -7596 12711 -7550 13185
rect -7412 12711 -7366 13185
rect -6478 12711 -6432 13185
rect -6294 12711 -6248 13185
rect -6110 12711 -6064 13185
rect -5926 12711 -5880 13185
rect -3922 12711 -3876 13185
rect -3738 12711 -3692 13185
rect -3554 12711 -3508 13185
rect -3370 12711 -3324 13185
rect -2436 12711 -2390 13185
rect -2252 12711 -2206 13185
rect -2068 12711 -2022 13185
rect -1884 12711 -1838 13185
rect 120 12711 166 13185
rect 304 12711 350 13185
rect 488 12711 534 13185
rect 672 12711 718 13185
rect 1606 12711 1652 13185
rect 1790 12711 1836 13185
rect 1974 12711 2020 13185
rect 2158 12711 2204 13185
rect 4162 12711 4208 13185
rect 4346 12711 4392 13185
rect 4530 12711 4576 13185
rect 4714 12711 4760 13185
rect 5648 12711 5694 13185
rect 5832 12711 5878 13185
rect 6016 12711 6062 13185
rect 6200 12711 6246 13185
rect 8204 12711 8250 13185
rect 8388 12711 8434 13185
rect 8572 12711 8618 13185
rect 8756 12711 8802 13185
rect 9690 12711 9736 13185
rect 9874 12711 9920 13185
rect 10058 12711 10104 13185
rect 10242 12711 10288 13185
rect 12246 12711 12292 13185
rect 12430 12711 12476 13185
rect 12614 12711 12660 13185
rect 12798 12711 12844 13185
rect 13732 12711 13778 13185
rect 13916 12711 13962 13185
rect 14100 12711 14146 13185
rect 14284 12711 14330 13185
rect -11976 10506 -11930 10980
rect -11792 10506 -11746 10980
rect -11608 10506 -11562 10980
rect -11424 10506 -11378 10980
rect -10490 10507 -10444 10981
rect -10306 10507 -10260 10981
rect -10122 10507 -10076 10981
rect -9938 10507 -9892 10981
rect -7964 10506 -7918 10980
rect -7780 10506 -7734 10980
rect -7596 10506 -7550 10980
rect -7412 10506 -7366 10980
rect -6478 10507 -6432 10981
rect -6294 10507 -6248 10981
rect -6110 10507 -6064 10981
rect -5926 10507 -5880 10981
rect -3922 10506 -3876 10980
rect -3738 10506 -3692 10980
rect -3554 10506 -3508 10980
rect -3370 10506 -3324 10980
rect -2436 10507 -2390 10981
rect -2252 10507 -2206 10981
rect -2068 10507 -2022 10981
rect -1884 10507 -1838 10981
rect 120 10506 166 10980
rect 304 10506 350 10980
rect 488 10506 534 10980
rect 672 10506 718 10980
rect 1606 10507 1652 10981
rect 1790 10507 1836 10981
rect 1974 10507 2020 10981
rect 2158 10507 2204 10981
rect 4162 10506 4208 10980
rect 4346 10506 4392 10980
rect 4530 10506 4576 10980
rect 4714 10506 4760 10980
rect 5648 10507 5694 10981
rect 5832 10507 5878 10981
rect 6016 10507 6062 10981
rect 6200 10507 6246 10981
rect 8204 10506 8250 10980
rect 8388 10506 8434 10980
rect 8572 10506 8618 10980
rect 8756 10506 8802 10980
rect 9690 10507 9736 10981
rect 9874 10507 9920 10981
rect 10058 10507 10104 10981
rect 10242 10507 10288 10981
rect 12246 10506 12292 10980
rect 12430 10506 12476 10980
rect 12614 10506 12660 10980
rect 12798 10506 12844 10980
rect 13732 10507 13778 10981
rect 13916 10507 13962 10981
rect 14100 10507 14146 10981
rect 14284 10507 14330 10981
rect -11976 8301 -11930 8775
rect -11792 8301 -11746 8775
rect -11608 8301 -11562 8775
rect -11424 8301 -11378 8775
rect -7964 8301 -7918 8775
rect -7780 8301 -7734 8775
rect -7596 8301 -7550 8775
rect -7412 8301 -7366 8775
rect -3922 8301 -3876 8775
rect -3738 8301 -3692 8775
rect -3554 8301 -3508 8775
rect -3370 8301 -3324 8775
rect 120 8301 166 8775
rect 304 8301 350 8775
rect 488 8301 534 8775
rect 672 8301 718 8775
rect 4162 8301 4208 8775
rect 4346 8301 4392 8775
rect 4530 8301 4576 8775
rect 4714 8301 4760 8775
rect 8204 8301 8250 8775
rect 8388 8301 8434 8775
rect 8572 8301 8618 8775
rect 8756 8301 8802 8775
rect 12246 8301 12292 8775
rect 12430 8301 12476 8775
rect 12614 8301 12660 8775
rect 12798 8301 12844 8775
rect -10909 4933 -10863 5167
rect -10739 4958 -10693 5192
rect -10569 4933 -10523 5167
rect -10399 4958 -10353 5192
rect -10229 4933 -10183 5167
rect -10059 4933 -10013 5167
rect -8506 4680 -8460 4854
rect -8322 4680 -8276 4854
rect -8046 4680 -8000 4854
rect -7862 4680 -7816 4854
rect -9476 3575 -9430 4349
rect -9292 3575 -9246 4349
rect -7076 3575 -7030 4349
rect -6892 3575 -6846 4349
rect -11024 1530 -10978 1664
rect -10840 1530 -10794 1664
rect -10164 1530 -10118 1664
rect -9980 1530 -9934 1664
rect -9704 1510 -9658 1684
rect -9400 1510 -9354 1684
rect -9096 1510 -9050 1684
rect -8792 1510 -8746 1684
rect -8488 1510 -8442 1684
rect -8184 1510 -8138 1684
rect -7880 1510 -7834 1684
rect -7576 1510 -7530 1684
rect -7272 1510 -7226 1684
rect -6968 1510 -6922 1684
rect -6664 1510 -6618 1684
rect -6388 1530 -6342 1664
rect -6204 1530 -6158 1664
rect -5528 1530 -5482 1664
rect -5344 1530 -5298 1664
<< psubdiff >>
rect 40051 37941 40201 37963
rect 40051 37895 40103 37941
rect 40149 37895 40201 37941
rect 40051 37873 40201 37895
rect 40291 37941 40441 37963
rect 40291 37895 40343 37941
rect 40389 37895 40441 37941
rect 40291 37873 40441 37895
rect 40531 37941 40681 37963
rect 40531 37895 40583 37941
rect 40629 37895 40681 37941
rect 40531 37873 40681 37895
rect 40771 37941 40921 37963
rect 40771 37895 40823 37941
rect 40869 37895 40921 37941
rect 40771 37873 40921 37895
rect -4857 36238 -3957 36310
rect -4857 36194 -4785 36238
rect -4857 35854 -4844 36194
rect -4798 35854 -4785 36194
rect -4029 36194 -3957 36238
rect -4857 35810 -4785 35854
rect -4029 35854 -4016 36194
rect -3970 35854 -3957 36194
rect -4029 35810 -3957 35854
rect -4857 35738 -3957 35810
rect 4615 36238 5515 36310
rect 4615 36194 4687 36238
rect 4615 35854 4628 36194
rect 4674 35854 4687 36194
rect 5443 36194 5515 36238
rect 4615 35810 4687 35854
rect 5443 35854 5456 36194
rect 5502 35854 5515 36194
rect 5443 35810 5515 35854
rect 4615 35738 5515 35810
rect 14087 36239 14987 36311
rect 14087 36195 14159 36239
rect 14087 35855 14100 36195
rect 14146 35855 14159 36195
rect 14915 36195 14987 36239
rect 14087 35811 14159 35855
rect 14915 35855 14928 36195
rect 14974 35855 14987 36195
rect 14915 35811 14987 35855
rect 14087 35739 14987 35811
rect 23559 36239 24459 36311
rect 23559 36195 23631 36239
rect 23559 35855 23572 36195
rect 23618 35855 23631 36195
rect 24387 36195 24459 36239
rect 23559 35811 23631 35855
rect 24387 35855 24400 36195
rect 24446 35855 24459 36195
rect 24387 35811 24459 35855
rect 23559 35739 24459 35811
rect 33031 36239 33931 36311
rect 33031 36195 33103 36239
rect 33031 35855 33044 36195
rect 33090 35855 33103 36195
rect 33859 36195 33931 36239
rect 33031 35811 33103 35855
rect 33859 35855 33872 36195
rect 33918 35855 33931 36195
rect 33859 35811 33931 35855
rect 33031 35739 33931 35811
rect 42503 36239 43403 36311
rect 42503 36195 42575 36239
rect 42503 35855 42516 36195
rect 42562 35855 42575 36195
rect 43331 36195 43403 36239
rect 42503 35811 42575 35855
rect 43331 35855 43344 36195
rect 43390 35855 43403 36195
rect 43331 35811 43403 35855
rect 42503 35739 43403 35811
rect -4857 34033 -3957 34105
rect -4857 33989 -4785 34033
rect -4857 33649 -4844 33989
rect -4798 33649 -4785 33989
rect -4029 33989 -3957 34033
rect -4857 33605 -4785 33649
rect -4029 33649 -4016 33989
rect -3970 33649 -3957 33989
rect -4029 33605 -3957 33649
rect -4857 33533 -3957 33605
rect -3371 34033 -2471 34105
rect -3371 33989 -3299 34033
rect -3371 33649 -3358 33989
rect -3312 33649 -3299 33989
rect -2543 33989 -2471 34033
rect -3371 33605 -3299 33649
rect -2543 33649 -2530 33989
rect -2484 33649 -2471 33989
rect -2543 33605 -2471 33649
rect -3371 33533 -2471 33605
rect 4615 34033 5515 34105
rect 4615 33989 4687 34033
rect 4615 33649 4628 33989
rect 4674 33649 4687 33989
rect 5443 33989 5515 34033
rect 4615 33605 4687 33649
rect 5443 33649 5456 33989
rect 5502 33649 5515 33989
rect 5443 33605 5515 33649
rect 4615 33533 5515 33605
rect 6101 34033 7001 34105
rect 6101 33989 6173 34033
rect 6101 33649 6114 33989
rect 6160 33649 6173 33989
rect 6929 33989 7001 34033
rect 6101 33605 6173 33649
rect 6929 33649 6942 33989
rect 6988 33649 7001 33989
rect 6929 33605 7001 33649
rect 6101 33533 7001 33605
rect 14087 34034 14987 34106
rect 14087 33990 14159 34034
rect 14087 33650 14100 33990
rect 14146 33650 14159 33990
rect 14915 33990 14987 34034
rect 14087 33606 14159 33650
rect 14915 33650 14928 33990
rect 14974 33650 14987 33990
rect 14915 33606 14987 33650
rect 14087 33534 14987 33606
rect 15573 34034 16473 34106
rect 15573 33990 15645 34034
rect 15573 33650 15586 33990
rect 15632 33650 15645 33990
rect 16401 33990 16473 34034
rect 15573 33606 15645 33650
rect 16401 33650 16414 33990
rect 16460 33650 16473 33990
rect 16401 33606 16473 33650
rect 15573 33534 16473 33606
rect 23559 34034 24459 34106
rect 23559 33990 23631 34034
rect 23559 33650 23572 33990
rect 23618 33650 23631 33990
rect 24387 33990 24459 34034
rect 23559 33606 23631 33650
rect 24387 33650 24400 33990
rect 24446 33650 24459 33990
rect 24387 33606 24459 33650
rect 23559 33534 24459 33606
rect 25045 34034 25945 34106
rect 25045 33990 25117 34034
rect 25045 33650 25058 33990
rect 25104 33650 25117 33990
rect 25873 33990 25945 34034
rect 25045 33606 25117 33650
rect 25873 33650 25886 33990
rect 25932 33650 25945 33990
rect 25873 33606 25945 33650
rect 25045 33534 25945 33606
rect 33031 34034 33931 34106
rect 33031 33990 33103 34034
rect 33031 33650 33044 33990
rect 33090 33650 33103 33990
rect 33859 33990 33931 34034
rect 33031 33606 33103 33650
rect 33859 33650 33872 33990
rect 33918 33650 33931 33990
rect 33859 33606 33931 33650
rect 33031 33534 33931 33606
rect 34517 34034 35417 34106
rect 34517 33990 34589 34034
rect 34517 33650 34530 33990
rect 34576 33650 34589 33990
rect 35345 33990 35417 34034
rect 34517 33606 34589 33650
rect 35345 33650 35358 33990
rect 35404 33650 35417 33990
rect 35345 33606 35417 33650
rect 34517 33534 35417 33606
rect 42503 34034 43403 34106
rect 42503 33990 42575 34034
rect 42503 33650 42516 33990
rect 42562 33650 42575 33990
rect 43331 33990 43403 34034
rect 42503 33606 42575 33650
rect 43331 33650 43344 33990
rect 43390 33650 43403 33990
rect 43331 33606 43403 33650
rect 42503 33534 43403 33606
rect 43989 34034 44889 34106
rect 43989 33990 44061 34034
rect 43989 33650 44002 33990
rect 44048 33650 44061 33990
rect 44817 33990 44889 34034
rect 43989 33606 44061 33650
rect 44817 33650 44830 33990
rect 44876 33650 44889 33990
rect 44817 33606 44889 33650
rect 43989 33534 44889 33606
rect -4857 31828 -3957 31900
rect -4857 31784 -4785 31828
rect -4857 31444 -4844 31784
rect -4798 31444 -4785 31784
rect -4029 31784 -3957 31828
rect -4857 31400 -4785 31444
rect -4029 31444 -4016 31784
rect -3970 31444 -3957 31784
rect -4029 31400 -3957 31444
rect -4857 31328 -3957 31400
rect -3371 31829 -2471 31901
rect -3371 31785 -3299 31829
rect -3371 31445 -3358 31785
rect -3312 31445 -3299 31785
rect -2543 31785 -2471 31829
rect -3371 31401 -3299 31445
rect -2543 31445 -2530 31785
rect -2484 31445 -2471 31785
rect -2543 31401 -2471 31445
rect -3371 31329 -2471 31401
rect 4615 31828 5515 31900
rect 4615 31784 4687 31828
rect 4615 31444 4628 31784
rect 4674 31444 4687 31784
rect 5443 31784 5515 31828
rect 4615 31400 4687 31444
rect 5443 31444 5456 31784
rect 5502 31444 5515 31784
rect 5443 31400 5515 31444
rect 4615 31328 5515 31400
rect 6101 31829 7001 31901
rect 6101 31785 6173 31829
rect 6101 31445 6114 31785
rect 6160 31445 6173 31785
rect 6929 31785 7001 31829
rect 6101 31401 6173 31445
rect 6929 31445 6942 31785
rect 6988 31445 7001 31785
rect 6929 31401 7001 31445
rect 6101 31329 7001 31401
rect 14087 31829 14987 31901
rect 14087 31785 14159 31829
rect 14087 31445 14100 31785
rect 14146 31445 14159 31785
rect 14915 31785 14987 31829
rect 14087 31401 14159 31445
rect 14915 31445 14928 31785
rect 14974 31445 14987 31785
rect 14915 31401 14987 31445
rect 14087 31329 14987 31401
rect 15573 31830 16473 31902
rect 15573 31786 15645 31830
rect 15573 31446 15586 31786
rect 15632 31446 15645 31786
rect 16401 31786 16473 31830
rect 15573 31402 15645 31446
rect 16401 31446 16414 31786
rect 16460 31446 16473 31786
rect 16401 31402 16473 31446
rect 15573 31330 16473 31402
rect 23559 31829 24459 31901
rect 23559 31785 23631 31829
rect 23559 31445 23572 31785
rect 23618 31445 23631 31785
rect 24387 31785 24459 31829
rect 23559 31401 23631 31445
rect 24387 31445 24400 31785
rect 24446 31445 24459 31785
rect 24387 31401 24459 31445
rect 23559 31329 24459 31401
rect 25045 31830 25945 31902
rect 25045 31786 25117 31830
rect 25045 31446 25058 31786
rect 25104 31446 25117 31786
rect 25873 31786 25945 31830
rect 25045 31402 25117 31446
rect 25873 31446 25886 31786
rect 25932 31446 25945 31786
rect 25873 31402 25945 31446
rect 25045 31330 25945 31402
rect 33031 31829 33931 31901
rect 33031 31785 33103 31829
rect 33031 31445 33044 31785
rect 33090 31445 33103 31785
rect 33859 31785 33931 31829
rect 33031 31401 33103 31445
rect 33859 31445 33872 31785
rect 33918 31445 33931 31785
rect 33859 31401 33931 31445
rect 33031 31329 33931 31401
rect 34517 31830 35417 31902
rect 34517 31786 34589 31830
rect 34517 31446 34530 31786
rect 34576 31446 34589 31786
rect 35345 31786 35417 31830
rect 34517 31402 34589 31446
rect 35345 31446 35358 31786
rect 35404 31446 35417 31786
rect 35345 31402 35417 31446
rect 34517 31330 35417 31402
rect 42503 31829 43403 31901
rect 42503 31785 42575 31829
rect 42503 31445 42516 31785
rect 42562 31445 42575 31785
rect 43331 31785 43403 31829
rect 42503 31401 42575 31445
rect 43331 31445 43344 31785
rect 43390 31445 43403 31785
rect 43331 31401 43403 31445
rect 42503 31329 43403 31401
rect 43989 31830 44889 31902
rect 43989 31786 44061 31830
rect 43989 31446 44002 31786
rect 44048 31446 44061 31786
rect 44817 31786 44889 31830
rect 43989 31402 44061 31446
rect 44817 31446 44830 31786
rect 44876 31446 44889 31786
rect 44817 31402 44889 31446
rect 43989 31330 44889 31402
rect -9999 30753 -8079 30825
rect -9999 30709 -9927 30753
rect -9999 30369 -9986 30709
rect -9940 30369 -9927 30709
rect -9315 30709 -9243 30753
rect -9999 30325 -9927 30369
rect -9315 30369 -9302 30709
rect -9256 30369 -9243 30709
rect -8631 30709 -8559 30753
rect -9315 30325 -9243 30369
rect -8631 30369 -8618 30709
rect -8572 30369 -8559 30709
rect -8151 30709 -8079 30753
rect -8631 30325 -8559 30369
rect -8151 30369 -8138 30709
rect -8092 30369 -8079 30709
rect -8151 30325 -8079 30369
rect -9999 30253 -8079 30325
rect -527 30753 1393 30825
rect -527 30709 -455 30753
rect -10893 29333 -10341 29405
rect -10893 29289 -10821 29333
rect -10893 28949 -10880 29289
rect -10834 28949 -10821 29289
rect -10413 29289 -10341 29333
rect -10893 28905 -10821 28949
rect -10413 28949 -10400 29289
rect -10354 28949 -10341 29289
rect -10413 28905 -10341 28949
rect -10893 28833 -10341 28905
rect -7771 29577 -7219 29649
rect -7771 29533 -7699 29577
rect -7771 29193 -7758 29533
rect -7712 29193 -7699 29533
rect -7291 29533 -7219 29577
rect -7771 29149 -7699 29193
rect -7291 29193 -7278 29533
rect -7232 29193 -7219 29533
rect -7291 29149 -7219 29193
rect -7771 29077 -7219 29149
rect -7087 29577 -6535 29649
rect -7087 29533 -7015 29577
rect -7087 29193 -7074 29533
rect -7028 29193 -7015 29533
rect -6607 29533 -6535 29577
rect -7087 29149 -7015 29193
rect -6607 29193 -6594 29533
rect -6548 29193 -6535 29533
rect -6607 29149 -6535 29193
rect -7087 29077 -6535 29149
rect -6403 29577 -5851 29649
rect -6403 29533 -6331 29577
rect -6403 29193 -6390 29533
rect -6344 29193 -6331 29533
rect -5923 29533 -5851 29577
rect -6403 29149 -6331 29193
rect -5923 29193 -5910 29533
rect -5864 29193 -5851 29533
rect -5923 29149 -5851 29193
rect -6403 29077 -5851 29149
rect -4857 29623 -3957 29695
rect -4857 29579 -4785 29623
rect -4857 29239 -4844 29579
rect -4798 29239 -4785 29579
rect -4029 29579 -3957 29623
rect -4857 29195 -4785 29239
rect -4029 29239 -4016 29579
rect -3970 29239 -3957 29579
rect -527 30369 -514 30709
rect -468 30369 -455 30709
rect 157 30709 229 30753
rect -527 30325 -455 30369
rect 157 30369 170 30709
rect 216 30369 229 30709
rect 841 30709 913 30753
rect 157 30325 229 30369
rect 841 30369 854 30709
rect 900 30369 913 30709
rect 1321 30709 1393 30753
rect 841 30325 913 30369
rect 1321 30369 1334 30709
rect 1380 30369 1393 30709
rect 1321 30325 1393 30369
rect -527 30253 1393 30325
rect 8945 30754 10865 30826
rect 8945 30710 9017 30754
rect -4029 29195 -3957 29239
rect -4857 29123 -3957 29195
rect -1421 29333 -869 29405
rect -1421 29289 -1349 29333
rect -1421 28949 -1408 29289
rect -1362 28949 -1349 29289
rect -941 29289 -869 29333
rect -1421 28905 -1349 28949
rect -941 28949 -928 29289
rect -882 28949 -869 29289
rect -941 28905 -869 28949
rect -1421 28833 -869 28905
rect 1701 29577 2253 29649
rect 1701 29533 1773 29577
rect 1701 29193 1714 29533
rect 1760 29193 1773 29533
rect 2181 29533 2253 29577
rect 1701 29149 1773 29193
rect 2181 29193 2194 29533
rect 2240 29193 2253 29533
rect 2181 29149 2253 29193
rect 1701 29077 2253 29149
rect 2385 29577 2937 29649
rect 2385 29533 2457 29577
rect 2385 29193 2398 29533
rect 2444 29193 2457 29533
rect 2865 29533 2937 29577
rect 2385 29149 2457 29193
rect 2865 29193 2878 29533
rect 2924 29193 2937 29533
rect 2865 29149 2937 29193
rect 2385 29077 2937 29149
rect 3069 29577 3621 29649
rect 3069 29533 3141 29577
rect 3069 29193 3082 29533
rect 3128 29193 3141 29533
rect 3549 29533 3621 29577
rect 3069 29149 3141 29193
rect 3549 29193 3562 29533
rect 3608 29193 3621 29533
rect 3549 29149 3621 29193
rect 3069 29077 3621 29149
rect 4615 29623 5515 29695
rect 4615 29579 4687 29623
rect 4615 29239 4628 29579
rect 4674 29239 4687 29579
rect 5443 29579 5515 29623
rect 4615 29195 4687 29239
rect 5443 29239 5456 29579
rect 5502 29239 5515 29579
rect 8945 30370 8958 30710
rect 9004 30370 9017 30710
rect 9629 30710 9701 30754
rect 8945 30326 9017 30370
rect 9629 30370 9642 30710
rect 9688 30370 9701 30710
rect 10313 30710 10385 30754
rect 9629 30326 9701 30370
rect 10313 30370 10326 30710
rect 10372 30370 10385 30710
rect 10793 30710 10865 30754
rect 10313 30326 10385 30370
rect 10793 30370 10806 30710
rect 10852 30370 10865 30710
rect 10793 30326 10865 30370
rect 8945 30254 10865 30326
rect 18417 30754 20337 30826
rect 18417 30710 18489 30754
rect 5443 29195 5515 29239
rect 4615 29123 5515 29195
rect 8051 29334 8603 29406
rect 8051 29290 8123 29334
rect 8051 28950 8064 29290
rect 8110 28950 8123 29290
rect 8531 29290 8603 29334
rect 8051 28906 8123 28950
rect 8531 28950 8544 29290
rect 8590 28950 8603 29290
rect 8531 28906 8603 28950
rect 8051 28834 8603 28906
rect 11173 29578 11725 29650
rect 11173 29534 11245 29578
rect 11173 29194 11186 29534
rect 11232 29194 11245 29534
rect 11653 29534 11725 29578
rect 11173 29150 11245 29194
rect 11653 29194 11666 29534
rect 11712 29194 11725 29534
rect 11653 29150 11725 29194
rect 11173 29078 11725 29150
rect 11857 29578 12409 29650
rect 11857 29534 11929 29578
rect 11857 29194 11870 29534
rect 11916 29194 11929 29534
rect 12337 29534 12409 29578
rect 11857 29150 11929 29194
rect 12337 29194 12350 29534
rect 12396 29194 12409 29534
rect 12337 29150 12409 29194
rect 11857 29078 12409 29150
rect 12541 29578 13093 29650
rect 12541 29534 12613 29578
rect 12541 29194 12554 29534
rect 12600 29194 12613 29534
rect 13021 29534 13093 29578
rect 12541 29150 12613 29194
rect 13021 29194 13034 29534
rect 13080 29194 13093 29534
rect 13021 29150 13093 29194
rect 12541 29078 13093 29150
rect 14087 29624 14987 29696
rect 14087 29580 14159 29624
rect 14087 29240 14100 29580
rect 14146 29240 14159 29580
rect 14915 29580 14987 29624
rect 14087 29196 14159 29240
rect 14915 29240 14928 29580
rect 14974 29240 14987 29580
rect 18417 30370 18430 30710
rect 18476 30370 18489 30710
rect 19101 30710 19173 30754
rect 18417 30326 18489 30370
rect 19101 30370 19114 30710
rect 19160 30370 19173 30710
rect 19785 30710 19857 30754
rect 19101 30326 19173 30370
rect 19785 30370 19798 30710
rect 19844 30370 19857 30710
rect 20265 30710 20337 30754
rect 19785 30326 19857 30370
rect 20265 30370 20278 30710
rect 20324 30370 20337 30710
rect 20265 30326 20337 30370
rect 18417 30254 20337 30326
rect 27889 30754 29809 30826
rect 27889 30710 27961 30754
rect 14915 29196 14987 29240
rect 14087 29124 14987 29196
rect 17523 29334 18075 29406
rect 17523 29290 17595 29334
rect 17523 28950 17536 29290
rect 17582 28950 17595 29290
rect 18003 29290 18075 29334
rect 17523 28906 17595 28950
rect 18003 28950 18016 29290
rect 18062 28950 18075 29290
rect 18003 28906 18075 28950
rect 17523 28834 18075 28906
rect 20645 29578 21197 29650
rect 20645 29534 20717 29578
rect 20645 29194 20658 29534
rect 20704 29194 20717 29534
rect 21125 29534 21197 29578
rect 20645 29150 20717 29194
rect 21125 29194 21138 29534
rect 21184 29194 21197 29534
rect 21125 29150 21197 29194
rect 20645 29078 21197 29150
rect 21329 29578 21881 29650
rect 21329 29534 21401 29578
rect 21329 29194 21342 29534
rect 21388 29194 21401 29534
rect 21809 29534 21881 29578
rect 21329 29150 21401 29194
rect 21809 29194 21822 29534
rect 21868 29194 21881 29534
rect 21809 29150 21881 29194
rect 21329 29078 21881 29150
rect 22013 29578 22565 29650
rect 22013 29534 22085 29578
rect 22013 29194 22026 29534
rect 22072 29194 22085 29534
rect 22493 29534 22565 29578
rect 22013 29150 22085 29194
rect 22493 29194 22506 29534
rect 22552 29194 22565 29534
rect 22493 29150 22565 29194
rect 22013 29078 22565 29150
rect 23559 29624 24459 29696
rect 23559 29580 23631 29624
rect 23559 29240 23572 29580
rect 23618 29240 23631 29580
rect 24387 29580 24459 29624
rect 23559 29196 23631 29240
rect 24387 29240 24400 29580
rect 24446 29240 24459 29580
rect 27889 30370 27902 30710
rect 27948 30370 27961 30710
rect 28573 30710 28645 30754
rect 27889 30326 27961 30370
rect 28573 30370 28586 30710
rect 28632 30370 28645 30710
rect 29257 30710 29329 30754
rect 28573 30326 28645 30370
rect 29257 30370 29270 30710
rect 29316 30370 29329 30710
rect 29737 30710 29809 30754
rect 29257 30326 29329 30370
rect 29737 30370 29750 30710
rect 29796 30370 29809 30710
rect 29737 30326 29809 30370
rect 27889 30254 29809 30326
rect 37361 30754 39281 30826
rect 37361 30710 37433 30754
rect 24387 29196 24459 29240
rect 23559 29124 24459 29196
rect 26995 29334 27547 29406
rect 26995 29290 27067 29334
rect 26995 28950 27008 29290
rect 27054 28950 27067 29290
rect 27475 29290 27547 29334
rect 26995 28906 27067 28950
rect 27475 28950 27488 29290
rect 27534 28950 27547 29290
rect 27475 28906 27547 28950
rect 26995 28834 27547 28906
rect 30117 29578 30669 29650
rect 30117 29534 30189 29578
rect 30117 29194 30130 29534
rect 30176 29194 30189 29534
rect 30597 29534 30669 29578
rect 30117 29150 30189 29194
rect 30597 29194 30610 29534
rect 30656 29194 30669 29534
rect 30597 29150 30669 29194
rect 30117 29078 30669 29150
rect 30801 29578 31353 29650
rect 30801 29534 30873 29578
rect 30801 29194 30814 29534
rect 30860 29194 30873 29534
rect 31281 29534 31353 29578
rect 30801 29150 30873 29194
rect 31281 29194 31294 29534
rect 31340 29194 31353 29534
rect 31281 29150 31353 29194
rect 30801 29078 31353 29150
rect 31485 29578 32037 29650
rect 31485 29534 31557 29578
rect 31485 29194 31498 29534
rect 31544 29194 31557 29534
rect 31965 29534 32037 29578
rect 31485 29150 31557 29194
rect 31965 29194 31978 29534
rect 32024 29194 32037 29534
rect 31965 29150 32037 29194
rect 31485 29078 32037 29150
rect 33031 29624 33931 29696
rect 33031 29580 33103 29624
rect 33031 29240 33044 29580
rect 33090 29240 33103 29580
rect 33859 29580 33931 29624
rect 33031 29196 33103 29240
rect 33859 29240 33872 29580
rect 33918 29240 33931 29580
rect 37361 30370 37374 30710
rect 37420 30370 37433 30710
rect 38045 30710 38117 30754
rect 37361 30326 37433 30370
rect 38045 30370 38058 30710
rect 38104 30370 38117 30710
rect 38729 30710 38801 30754
rect 38045 30326 38117 30370
rect 38729 30370 38742 30710
rect 38788 30370 38801 30710
rect 39209 30710 39281 30754
rect 38729 30326 38801 30370
rect 39209 30370 39222 30710
rect 39268 30370 39281 30710
rect 39209 30326 39281 30370
rect 37361 30254 39281 30326
rect 33859 29196 33931 29240
rect 33031 29124 33931 29196
rect 36467 29334 37019 29406
rect 36467 29290 36539 29334
rect 36467 28950 36480 29290
rect 36526 28950 36539 29290
rect 36947 29290 37019 29334
rect 36467 28906 36539 28950
rect 36947 28950 36960 29290
rect 37006 28950 37019 29290
rect 36947 28906 37019 28950
rect 36467 28834 37019 28906
rect 39589 29578 40141 29650
rect 39589 29534 39661 29578
rect 39589 29194 39602 29534
rect 39648 29194 39661 29534
rect 40069 29534 40141 29578
rect 39589 29150 39661 29194
rect 40069 29194 40082 29534
rect 40128 29194 40141 29534
rect 40069 29150 40141 29194
rect 39589 29078 40141 29150
rect 40273 29578 40825 29650
rect 40273 29534 40345 29578
rect 40273 29194 40286 29534
rect 40332 29194 40345 29534
rect 40753 29534 40825 29578
rect 40273 29150 40345 29194
rect 40753 29194 40766 29534
rect 40812 29194 40825 29534
rect 40753 29150 40825 29194
rect 40273 29078 40825 29150
rect 40957 29578 41509 29650
rect 40957 29534 41029 29578
rect 40957 29194 40970 29534
rect 41016 29194 41029 29534
rect 41437 29534 41509 29578
rect 40957 29150 41029 29194
rect 41437 29194 41450 29534
rect 41496 29194 41509 29534
rect 41437 29150 41509 29194
rect 40957 29078 41509 29150
rect 42503 29624 43403 29696
rect 42503 29580 42575 29624
rect 42503 29240 42516 29580
rect 42562 29240 42575 29580
rect 43331 29580 43403 29624
rect 42503 29196 42575 29240
rect 43331 29240 43344 29580
rect 43390 29240 43403 29580
rect 43331 29196 43403 29240
rect 42503 29124 43403 29196
rect -9999 28413 -8079 28485
rect -9999 28369 -9927 28413
rect -9999 28029 -9986 28369
rect -9940 28029 -9927 28369
rect -9315 28369 -9243 28413
rect -9999 27985 -9927 28029
rect -9315 28029 -9302 28369
rect -9256 28029 -9243 28369
rect -8631 28369 -8559 28413
rect -9315 27985 -9243 28029
rect -8631 28029 -8618 28369
rect -8572 28029 -8559 28369
rect -8151 28369 -8079 28413
rect -8631 27985 -8559 28029
rect -8151 28029 -8138 28369
rect -8092 28029 -8079 28369
rect -8151 27985 -8079 28029
rect -9999 27913 -8079 27985
rect -527 28413 1393 28485
rect -527 28369 -455 28413
rect -527 28029 -514 28369
rect -468 28029 -455 28369
rect 157 28369 229 28413
rect -527 27985 -455 28029
rect 157 28029 170 28369
rect 216 28029 229 28369
rect 841 28369 913 28413
rect 157 27985 229 28029
rect 841 28029 854 28369
rect 900 28029 913 28369
rect 1321 28369 1393 28413
rect 841 27985 913 28029
rect 1321 28029 1334 28369
rect 1380 28029 1393 28369
rect 1321 27985 1393 28029
rect -527 27913 1393 27985
rect 8945 28414 10865 28486
rect 8945 28370 9017 28414
rect 8945 28030 8958 28370
rect 9004 28030 9017 28370
rect 9629 28370 9701 28414
rect 8945 27986 9017 28030
rect 9629 28030 9642 28370
rect 9688 28030 9701 28370
rect 10313 28370 10385 28414
rect 9629 27986 9701 28030
rect 10313 28030 10326 28370
rect 10372 28030 10385 28370
rect 10793 28370 10865 28414
rect 10313 27986 10385 28030
rect 10793 28030 10806 28370
rect 10852 28030 10865 28370
rect 10793 27986 10865 28030
rect 8945 27914 10865 27986
rect 18417 28414 20337 28486
rect 18417 28370 18489 28414
rect 18417 28030 18430 28370
rect 18476 28030 18489 28370
rect 19101 28370 19173 28414
rect 18417 27986 18489 28030
rect 19101 28030 19114 28370
rect 19160 28030 19173 28370
rect 19785 28370 19857 28414
rect 19101 27986 19173 28030
rect 19785 28030 19798 28370
rect 19844 28030 19857 28370
rect 20265 28370 20337 28414
rect 19785 27986 19857 28030
rect 20265 28030 20278 28370
rect 20324 28030 20337 28370
rect 20265 27986 20337 28030
rect 18417 27914 20337 27986
rect 27889 28414 29809 28486
rect 27889 28370 27961 28414
rect 27889 28030 27902 28370
rect 27948 28030 27961 28370
rect 28573 28370 28645 28414
rect 27889 27986 27961 28030
rect 28573 28030 28586 28370
rect 28632 28030 28645 28370
rect 29257 28370 29329 28414
rect 28573 27986 28645 28030
rect 29257 28030 29270 28370
rect 29316 28030 29329 28370
rect 29737 28370 29809 28414
rect 29257 27986 29329 28030
rect 29737 28030 29750 28370
rect 29796 28030 29809 28370
rect 29737 27986 29809 28030
rect 27889 27914 29809 27986
rect 37361 28414 39281 28486
rect 37361 28370 37433 28414
rect 37361 28030 37374 28370
rect 37420 28030 37433 28370
rect 38045 28370 38117 28414
rect 37361 27986 37433 28030
rect 38045 28030 38058 28370
rect 38104 28030 38117 28370
rect 38729 28370 38801 28414
rect 38045 27986 38117 28030
rect 38729 28030 38742 28370
rect 38788 28030 38801 28370
rect 39209 28370 39281 28414
rect 38729 27986 38801 28030
rect 39209 28030 39222 28370
rect 39268 28030 39281 28370
rect 39209 27986 39281 28030
rect 37361 27914 39281 27986
rect -12606 27403 -12054 27475
rect -12606 27359 -12534 27403
rect -12606 27019 -12593 27359
rect -12547 27019 -12534 27359
rect -12126 27359 -12054 27403
rect -12606 26975 -12534 27019
rect -12126 27019 -12113 27359
rect -12067 27019 -12054 27359
rect -12126 26975 -12054 27019
rect -12606 26903 -12054 26975
rect -8115 23936 -7215 24008
rect -8115 23892 -8043 23936
rect -8115 23552 -8102 23892
rect -8056 23552 -8043 23892
rect -7287 23892 -7215 23936
rect -8115 23508 -8043 23552
rect -7287 23552 -7274 23892
rect -7228 23552 -7215 23892
rect -7287 23508 -7215 23552
rect -8115 23436 -7215 23508
rect -4073 23933 -3173 24005
rect -4073 23889 -4001 23933
rect -4073 23549 -4060 23889
rect -4014 23549 -4001 23889
rect -3245 23889 -3173 23933
rect -4073 23505 -4001 23549
rect -3245 23549 -3232 23889
rect -3186 23549 -3173 23889
rect -3245 23505 -3173 23549
rect -4073 23433 -3173 23505
rect -31 23933 869 24005
rect -31 23889 41 23933
rect -31 23549 -18 23889
rect 28 23549 41 23889
rect 797 23889 869 23933
rect -31 23505 41 23549
rect 797 23549 810 23889
rect 856 23549 869 23889
rect 797 23505 869 23549
rect -31 23433 869 23505
rect 4011 23933 4911 24005
rect 4011 23889 4083 23933
rect 4011 23549 4024 23889
rect 4070 23549 4083 23889
rect 4839 23889 4911 23933
rect 4011 23505 4083 23549
rect 4839 23549 4852 23889
rect 4898 23549 4911 23889
rect 4839 23505 4911 23549
rect 4011 23433 4911 23505
rect 8053 23933 8953 24005
rect 8053 23889 8125 23933
rect 8053 23549 8066 23889
rect 8112 23549 8125 23889
rect 8881 23889 8953 23933
rect 8053 23505 8125 23549
rect 8881 23549 8894 23889
rect 8940 23549 8953 23889
rect 8881 23505 8953 23549
rect 8053 23433 8953 23505
rect 12095 23933 12995 24005
rect 12095 23889 12167 23933
rect 12095 23549 12108 23889
rect 12154 23549 12167 23889
rect 12923 23889 12995 23933
rect 12095 23505 12167 23549
rect 12923 23549 12936 23889
rect 12982 23549 12995 23889
rect 12923 23505 12995 23549
rect 12095 23433 12995 23505
rect 16137 23933 17037 24005
rect 16137 23889 16209 23933
rect 16137 23549 16150 23889
rect 16196 23549 16209 23889
rect 16965 23889 17037 23933
rect 16137 23505 16209 23549
rect 16965 23549 16978 23889
rect 17024 23549 17037 23889
rect 16965 23505 17037 23549
rect 16137 23433 17037 23505
rect -8115 21731 -7215 21803
rect -8115 21687 -8043 21731
rect -8115 21347 -8102 21687
rect -8056 21347 -8043 21687
rect -7287 21687 -7215 21731
rect -8115 21303 -8043 21347
rect -7287 21347 -7274 21687
rect -7228 21347 -7215 21687
rect -7287 21303 -7215 21347
rect -8115 21231 -7215 21303
rect -6629 21731 -5729 21803
rect -6629 21687 -6557 21731
rect -6629 21347 -6616 21687
rect -6570 21347 -6557 21687
rect -5801 21687 -5729 21731
rect -6629 21303 -6557 21347
rect -5801 21347 -5788 21687
rect -5742 21347 -5729 21687
rect -5801 21303 -5729 21347
rect -6629 21231 -5729 21303
rect -4073 21728 -3173 21800
rect -4073 21684 -4001 21728
rect -4073 21344 -4060 21684
rect -4014 21344 -4001 21684
rect -3245 21684 -3173 21728
rect -4073 21300 -4001 21344
rect -3245 21344 -3232 21684
rect -3186 21344 -3173 21684
rect -3245 21300 -3173 21344
rect -4073 21228 -3173 21300
rect -2587 21728 -1687 21800
rect -2587 21684 -2515 21728
rect -2587 21344 -2574 21684
rect -2528 21344 -2515 21684
rect -1759 21684 -1687 21728
rect -2587 21300 -2515 21344
rect -1759 21344 -1746 21684
rect -1700 21344 -1687 21684
rect -1759 21300 -1687 21344
rect -2587 21228 -1687 21300
rect -31 21728 869 21800
rect -31 21684 41 21728
rect -31 21344 -18 21684
rect 28 21344 41 21684
rect 797 21684 869 21728
rect -31 21300 41 21344
rect 797 21344 810 21684
rect 856 21344 869 21684
rect 797 21300 869 21344
rect -31 21228 869 21300
rect 1455 21728 2355 21800
rect 1455 21684 1527 21728
rect 1455 21344 1468 21684
rect 1514 21344 1527 21684
rect 2283 21684 2355 21728
rect 1455 21300 1527 21344
rect 2283 21344 2296 21684
rect 2342 21344 2355 21684
rect 2283 21300 2355 21344
rect 1455 21228 2355 21300
rect 4011 21728 4911 21800
rect 4011 21684 4083 21728
rect 4011 21344 4024 21684
rect 4070 21344 4083 21684
rect 4839 21684 4911 21728
rect 4011 21300 4083 21344
rect 4839 21344 4852 21684
rect 4898 21344 4911 21684
rect 4839 21300 4911 21344
rect 4011 21228 4911 21300
rect 5497 21728 6397 21800
rect 5497 21684 5569 21728
rect 5497 21344 5510 21684
rect 5556 21344 5569 21684
rect 6325 21684 6397 21728
rect 5497 21300 5569 21344
rect 6325 21344 6338 21684
rect 6384 21344 6397 21684
rect 6325 21300 6397 21344
rect 5497 21228 6397 21300
rect 8053 21728 8953 21800
rect 8053 21684 8125 21728
rect 8053 21344 8066 21684
rect 8112 21344 8125 21684
rect 8881 21684 8953 21728
rect 8053 21300 8125 21344
rect 8881 21344 8894 21684
rect 8940 21344 8953 21684
rect 8881 21300 8953 21344
rect 8053 21228 8953 21300
rect 9539 21728 10439 21800
rect 9539 21684 9611 21728
rect 9539 21344 9552 21684
rect 9598 21344 9611 21684
rect 10367 21684 10439 21728
rect 9539 21300 9611 21344
rect 10367 21344 10380 21684
rect 10426 21344 10439 21684
rect 10367 21300 10439 21344
rect 9539 21228 10439 21300
rect 12095 21728 12995 21800
rect 12095 21684 12167 21728
rect 12095 21344 12108 21684
rect 12154 21344 12167 21684
rect 12923 21684 12995 21728
rect 12095 21300 12167 21344
rect 12923 21344 12936 21684
rect 12982 21344 12995 21684
rect 12923 21300 12995 21344
rect 12095 21228 12995 21300
rect 13581 21728 14481 21800
rect 13581 21684 13653 21728
rect 13581 21344 13594 21684
rect 13640 21344 13653 21684
rect 14409 21684 14481 21728
rect 13581 21300 13653 21344
rect 14409 21344 14422 21684
rect 14468 21344 14481 21684
rect 14409 21300 14481 21344
rect 13581 21228 14481 21300
rect 16137 21728 17037 21800
rect 16137 21684 16209 21728
rect 16137 21344 16150 21684
rect 16196 21344 16209 21684
rect 16965 21684 17037 21728
rect 16137 21300 16209 21344
rect 16965 21344 16978 21684
rect 17024 21344 17037 21684
rect 16965 21300 17037 21344
rect 16137 21228 17037 21300
rect 17623 21728 18523 21800
rect 17623 21684 17695 21728
rect 17623 21344 17636 21684
rect 17682 21344 17695 21684
rect 18451 21684 18523 21728
rect 17623 21300 17695 21344
rect 18451 21344 18464 21684
rect 18510 21344 18523 21684
rect 18451 21300 18523 21344
rect 17623 21228 18523 21300
rect -8115 19526 -7215 19598
rect -8115 19482 -8043 19526
rect -8115 19142 -8102 19482
rect -8056 19142 -8043 19482
rect -7287 19482 -7215 19526
rect -8115 19098 -8043 19142
rect -7287 19142 -7274 19482
rect -7228 19142 -7215 19482
rect -7287 19098 -7215 19142
rect -8115 19026 -7215 19098
rect -6629 19527 -5729 19599
rect -6629 19483 -6557 19527
rect -6629 19143 -6616 19483
rect -6570 19143 -6557 19483
rect -5801 19483 -5729 19527
rect -6629 19099 -6557 19143
rect -5801 19143 -5788 19483
rect -5742 19143 -5729 19483
rect -5801 19099 -5729 19143
rect -6629 19027 -5729 19099
rect -4073 19523 -3173 19595
rect -4073 19479 -4001 19523
rect -4073 19139 -4060 19479
rect -4014 19139 -4001 19479
rect -3245 19479 -3173 19523
rect -4073 19095 -4001 19139
rect -3245 19139 -3232 19479
rect -3186 19139 -3173 19479
rect -3245 19095 -3173 19139
rect -4073 19023 -3173 19095
rect -2587 19524 -1687 19596
rect -2587 19480 -2515 19524
rect -2587 19140 -2574 19480
rect -2528 19140 -2515 19480
rect -1759 19480 -1687 19524
rect -2587 19096 -2515 19140
rect -1759 19140 -1746 19480
rect -1700 19140 -1687 19480
rect -1759 19096 -1687 19140
rect -2587 19024 -1687 19096
rect -31 19523 869 19595
rect -31 19479 41 19523
rect -31 19139 -18 19479
rect 28 19139 41 19479
rect 797 19479 869 19523
rect -31 19095 41 19139
rect 797 19139 810 19479
rect 856 19139 869 19479
rect 797 19095 869 19139
rect -31 19023 869 19095
rect 1455 19524 2355 19596
rect 1455 19480 1527 19524
rect 1455 19140 1468 19480
rect 1514 19140 1527 19480
rect 2283 19480 2355 19524
rect 1455 19096 1527 19140
rect 2283 19140 2296 19480
rect 2342 19140 2355 19480
rect 2283 19096 2355 19140
rect 1455 19024 2355 19096
rect 4011 19523 4911 19595
rect 4011 19479 4083 19523
rect 4011 19139 4024 19479
rect 4070 19139 4083 19479
rect 4839 19479 4911 19523
rect 4011 19095 4083 19139
rect 4839 19139 4852 19479
rect 4898 19139 4911 19479
rect 4839 19095 4911 19139
rect 4011 19023 4911 19095
rect 5497 19524 6397 19596
rect 5497 19480 5569 19524
rect 5497 19140 5510 19480
rect 5556 19140 5569 19480
rect 6325 19480 6397 19524
rect 5497 19096 5569 19140
rect 6325 19140 6338 19480
rect 6384 19140 6397 19480
rect 6325 19096 6397 19140
rect 5497 19024 6397 19096
rect 8053 19523 8953 19595
rect 8053 19479 8125 19523
rect 8053 19139 8066 19479
rect 8112 19139 8125 19479
rect 8881 19479 8953 19523
rect 8053 19095 8125 19139
rect 8881 19139 8894 19479
rect 8940 19139 8953 19479
rect 8881 19095 8953 19139
rect 8053 19023 8953 19095
rect 9539 19524 10439 19596
rect 9539 19480 9611 19524
rect 9539 19140 9552 19480
rect 9598 19140 9611 19480
rect 10367 19480 10439 19524
rect 9539 19096 9611 19140
rect 10367 19140 10380 19480
rect 10426 19140 10439 19480
rect 10367 19096 10439 19140
rect 9539 19024 10439 19096
rect 12095 19523 12995 19595
rect 12095 19479 12167 19523
rect 12095 19139 12108 19479
rect 12154 19139 12167 19479
rect 12923 19479 12995 19523
rect 12095 19095 12167 19139
rect 12923 19139 12936 19479
rect 12982 19139 12995 19479
rect 12923 19095 12995 19139
rect 12095 19023 12995 19095
rect 13581 19524 14481 19596
rect 13581 19480 13653 19524
rect 13581 19140 13594 19480
rect 13640 19140 13653 19480
rect 14409 19480 14481 19524
rect 13581 19096 13653 19140
rect 14409 19140 14422 19480
rect 14468 19140 14481 19480
rect 14409 19096 14481 19140
rect 13581 19024 14481 19096
rect 16137 19523 17037 19595
rect 16137 19479 16209 19523
rect 16137 19139 16150 19479
rect 16196 19139 16209 19479
rect 16965 19479 17037 19523
rect 16137 19095 16209 19139
rect 16965 19139 16978 19479
rect 17024 19139 17037 19479
rect 16965 19095 17037 19139
rect 16137 19023 17037 19095
rect 17623 19524 18523 19596
rect 17623 19480 17695 19524
rect 17623 19140 17636 19480
rect 17682 19140 17695 19480
rect 18451 19480 18523 19524
rect 17623 19096 17695 19140
rect 18451 19140 18464 19480
rect 18510 19140 18523 19480
rect 18451 19096 18523 19140
rect 17623 19024 18523 19096
rect -8115 17321 -7215 17393
rect -8115 17277 -8043 17321
rect -8115 16937 -8102 17277
rect -8056 16937 -8043 17277
rect -7287 17277 -7215 17321
rect -8115 16893 -8043 16937
rect -7287 16937 -7274 17277
rect -7228 16937 -7215 17277
rect -7287 16893 -7215 16937
rect -8115 16821 -7215 16893
rect -4073 17318 -3173 17390
rect -4073 17274 -4001 17318
rect -4073 16934 -4060 17274
rect -4014 16934 -4001 17274
rect -3245 17274 -3173 17318
rect -4073 16890 -4001 16934
rect -3245 16934 -3232 17274
rect -3186 16934 -3173 17274
rect -3245 16890 -3173 16934
rect -4073 16818 -3173 16890
rect -31 17318 869 17390
rect -31 17274 41 17318
rect -31 16934 -18 17274
rect 28 16934 41 17274
rect 797 17274 869 17318
rect -31 16890 41 16934
rect 797 16934 810 17274
rect 856 16934 869 17274
rect 797 16890 869 16934
rect -31 16818 869 16890
rect 4011 17318 4911 17390
rect 4011 17274 4083 17318
rect 4011 16934 4024 17274
rect 4070 16934 4083 17274
rect 4839 17274 4911 17318
rect 4011 16890 4083 16934
rect 4839 16934 4852 17274
rect 4898 16934 4911 17274
rect 4839 16890 4911 16934
rect 4011 16818 4911 16890
rect 8053 17318 8953 17390
rect 8053 17274 8125 17318
rect 8053 16934 8066 17274
rect 8112 16934 8125 17274
rect 8881 17274 8953 17318
rect 8053 16890 8125 16934
rect 8881 16934 8894 17274
rect 8940 16934 8953 17274
rect 8881 16890 8953 16934
rect 8053 16818 8953 16890
rect 12095 17318 12995 17390
rect 12095 17274 12167 17318
rect 12095 16934 12108 17274
rect 12154 16934 12167 17274
rect 12923 17274 12995 17318
rect 12095 16890 12167 16934
rect 12923 16934 12936 17274
rect 12982 16934 12995 17274
rect 12923 16890 12995 16934
rect 12095 16818 12995 16890
rect 16137 17318 17037 17390
rect 16137 17274 16209 17318
rect 16137 16934 16150 17274
rect 16196 16934 16209 17274
rect 16965 17274 17037 17318
rect 16137 16890 16209 16934
rect 16965 16934 16978 17274
rect 17024 16934 17037 17274
rect 16965 16890 17037 16934
rect 16137 16818 17037 16890
rect -12127 14357 -11227 14429
rect -12127 14313 -12055 14357
rect -12127 13973 -12114 14313
rect -12068 13973 -12055 14313
rect -11299 14313 -11227 14357
rect -12127 13929 -12055 13973
rect -11299 13973 -11286 14313
rect -11240 13973 -11227 14313
rect -11299 13929 -11227 13973
rect -12127 13857 -11227 13929
rect -8115 14357 -7215 14429
rect -8115 14313 -8043 14357
rect -8115 13973 -8102 14313
rect -8056 13973 -8043 14313
rect -7287 14313 -7215 14357
rect -8115 13929 -8043 13973
rect -7287 13973 -7274 14313
rect -7228 13973 -7215 14313
rect -7287 13929 -7215 13973
rect -8115 13857 -7215 13929
rect -4073 14357 -3173 14429
rect -4073 14313 -4001 14357
rect -4073 13973 -4060 14313
rect -4014 13973 -4001 14313
rect -3245 14313 -3173 14357
rect -4073 13929 -4001 13973
rect -3245 13973 -3232 14313
rect -3186 13973 -3173 14313
rect -3245 13929 -3173 13973
rect -4073 13857 -3173 13929
rect -31 14357 869 14429
rect -31 14313 41 14357
rect -31 13973 -18 14313
rect 28 13973 41 14313
rect 797 14313 869 14357
rect -31 13929 41 13973
rect 797 13973 810 14313
rect 856 13973 869 14313
rect 797 13929 869 13973
rect -31 13857 869 13929
rect 4011 14357 4911 14429
rect 4011 14313 4083 14357
rect 4011 13973 4024 14313
rect 4070 13973 4083 14313
rect 4839 14313 4911 14357
rect 4011 13929 4083 13973
rect 4839 13973 4852 14313
rect 4898 13973 4911 14313
rect 4839 13929 4911 13973
rect 4011 13857 4911 13929
rect 8053 14357 8953 14429
rect 8053 14313 8125 14357
rect 8053 13973 8066 14313
rect 8112 13973 8125 14313
rect 8881 14313 8953 14357
rect 8053 13929 8125 13973
rect 8881 13973 8894 14313
rect 8940 13973 8953 14313
rect 8881 13929 8953 13973
rect 8053 13857 8953 13929
rect 12095 14357 12995 14429
rect 12095 14313 12167 14357
rect 12095 13973 12108 14313
rect 12154 13973 12167 14313
rect 12923 14313 12995 14357
rect 12095 13929 12167 13973
rect 12923 13973 12936 14313
rect 12982 13973 12995 14313
rect 12923 13929 12995 13973
rect 12095 13857 12995 13929
rect -12127 12152 -11227 12224
rect -12127 12108 -12055 12152
rect -12127 11768 -12114 12108
rect -12068 11768 -12055 12108
rect -11299 12108 -11227 12152
rect -12127 11724 -12055 11768
rect -11299 11768 -11286 12108
rect -11240 11768 -11227 12108
rect -11299 11724 -11227 11768
rect -12127 11652 -11227 11724
rect -10641 12152 -9741 12224
rect -10641 12108 -10569 12152
rect -10641 11768 -10628 12108
rect -10582 11768 -10569 12108
rect -9813 12108 -9741 12152
rect -10641 11724 -10569 11768
rect -9813 11768 -9800 12108
rect -9754 11768 -9741 12108
rect -9813 11724 -9741 11768
rect -10641 11652 -9741 11724
rect -8115 12152 -7215 12224
rect -8115 12108 -8043 12152
rect -8115 11768 -8102 12108
rect -8056 11768 -8043 12108
rect -7287 12108 -7215 12152
rect -8115 11724 -8043 11768
rect -7287 11768 -7274 12108
rect -7228 11768 -7215 12108
rect -7287 11724 -7215 11768
rect -8115 11652 -7215 11724
rect -6629 12152 -5729 12224
rect -6629 12108 -6557 12152
rect -6629 11768 -6616 12108
rect -6570 11768 -6557 12108
rect -5801 12108 -5729 12152
rect -6629 11724 -6557 11768
rect -5801 11768 -5788 12108
rect -5742 11768 -5729 12108
rect -5801 11724 -5729 11768
rect -6629 11652 -5729 11724
rect -4073 12152 -3173 12224
rect -4073 12108 -4001 12152
rect -4073 11768 -4060 12108
rect -4014 11768 -4001 12108
rect -3245 12108 -3173 12152
rect -4073 11724 -4001 11768
rect -3245 11768 -3232 12108
rect -3186 11768 -3173 12108
rect -3245 11724 -3173 11768
rect -4073 11652 -3173 11724
rect -2587 12152 -1687 12224
rect -2587 12108 -2515 12152
rect -2587 11768 -2574 12108
rect -2528 11768 -2515 12108
rect -1759 12108 -1687 12152
rect -2587 11724 -2515 11768
rect -1759 11768 -1746 12108
rect -1700 11768 -1687 12108
rect -1759 11724 -1687 11768
rect -2587 11652 -1687 11724
rect -31 12152 869 12224
rect -31 12108 41 12152
rect -31 11768 -18 12108
rect 28 11768 41 12108
rect 797 12108 869 12152
rect -31 11724 41 11768
rect 797 11768 810 12108
rect 856 11768 869 12108
rect 797 11724 869 11768
rect -31 11652 869 11724
rect 1455 12152 2355 12224
rect 1455 12108 1527 12152
rect 1455 11768 1468 12108
rect 1514 11768 1527 12108
rect 2283 12108 2355 12152
rect 1455 11724 1527 11768
rect 2283 11768 2296 12108
rect 2342 11768 2355 12108
rect 2283 11724 2355 11768
rect 1455 11652 2355 11724
rect 4011 12152 4911 12224
rect 4011 12108 4083 12152
rect 4011 11768 4024 12108
rect 4070 11768 4083 12108
rect 4839 12108 4911 12152
rect 4011 11724 4083 11768
rect 4839 11768 4852 12108
rect 4898 11768 4911 12108
rect 4839 11724 4911 11768
rect 4011 11652 4911 11724
rect 5497 12152 6397 12224
rect 5497 12108 5569 12152
rect 5497 11768 5510 12108
rect 5556 11768 5569 12108
rect 6325 12108 6397 12152
rect 5497 11724 5569 11768
rect 6325 11768 6338 12108
rect 6384 11768 6397 12108
rect 6325 11724 6397 11768
rect 5497 11652 6397 11724
rect 8053 12152 8953 12224
rect 8053 12108 8125 12152
rect 8053 11768 8066 12108
rect 8112 11768 8125 12108
rect 8881 12108 8953 12152
rect 8053 11724 8125 11768
rect 8881 11768 8894 12108
rect 8940 11768 8953 12108
rect 8881 11724 8953 11768
rect 8053 11652 8953 11724
rect 9539 12152 10439 12224
rect 9539 12108 9611 12152
rect 9539 11768 9552 12108
rect 9598 11768 9611 12108
rect 10367 12108 10439 12152
rect 9539 11724 9611 11768
rect 10367 11768 10380 12108
rect 10426 11768 10439 12108
rect 10367 11724 10439 11768
rect 9539 11652 10439 11724
rect 12095 12152 12995 12224
rect 12095 12108 12167 12152
rect 12095 11768 12108 12108
rect 12154 11768 12167 12108
rect 12923 12108 12995 12152
rect 12095 11724 12167 11768
rect 12923 11768 12936 12108
rect 12982 11768 12995 12108
rect 12923 11724 12995 11768
rect 12095 11652 12995 11724
rect 13581 12152 14481 12224
rect 13581 12108 13653 12152
rect 13581 11768 13594 12108
rect 13640 11768 13653 12108
rect 14409 12108 14481 12152
rect 13581 11724 13653 11768
rect 14409 11768 14422 12108
rect 14468 11768 14481 12108
rect 14409 11724 14481 11768
rect 13581 11652 14481 11724
rect -12127 9947 -11227 10019
rect -12127 9903 -12055 9947
rect -12127 9563 -12114 9903
rect -12068 9563 -12055 9903
rect -11299 9903 -11227 9947
rect -12127 9519 -12055 9563
rect -11299 9563 -11286 9903
rect -11240 9563 -11227 9903
rect -11299 9519 -11227 9563
rect -12127 9447 -11227 9519
rect -10641 9948 -9741 10020
rect -10641 9904 -10569 9948
rect -10641 9564 -10628 9904
rect -10582 9564 -10569 9904
rect -9813 9904 -9741 9948
rect -10641 9520 -10569 9564
rect -9813 9564 -9800 9904
rect -9754 9564 -9741 9904
rect -9813 9520 -9741 9564
rect -10641 9448 -9741 9520
rect -8115 9947 -7215 10019
rect -8115 9903 -8043 9947
rect -8115 9563 -8102 9903
rect -8056 9563 -8043 9903
rect -7287 9903 -7215 9947
rect -8115 9519 -8043 9563
rect -7287 9563 -7274 9903
rect -7228 9563 -7215 9903
rect -7287 9519 -7215 9563
rect -8115 9447 -7215 9519
rect -6629 9948 -5729 10020
rect -6629 9904 -6557 9948
rect -6629 9564 -6616 9904
rect -6570 9564 -6557 9904
rect -5801 9904 -5729 9948
rect -6629 9520 -6557 9564
rect -5801 9564 -5788 9904
rect -5742 9564 -5729 9904
rect -5801 9520 -5729 9564
rect -6629 9448 -5729 9520
rect -4073 9947 -3173 10019
rect -4073 9903 -4001 9947
rect -4073 9563 -4060 9903
rect -4014 9563 -4001 9903
rect -3245 9903 -3173 9947
rect -4073 9519 -4001 9563
rect -3245 9563 -3232 9903
rect -3186 9563 -3173 9903
rect -3245 9519 -3173 9563
rect -4073 9447 -3173 9519
rect -2587 9948 -1687 10020
rect -2587 9904 -2515 9948
rect -2587 9564 -2574 9904
rect -2528 9564 -2515 9904
rect -1759 9904 -1687 9948
rect -2587 9520 -2515 9564
rect -1759 9564 -1746 9904
rect -1700 9564 -1687 9904
rect -1759 9520 -1687 9564
rect -2587 9448 -1687 9520
rect -31 9947 869 10019
rect -31 9903 41 9947
rect -31 9563 -18 9903
rect 28 9563 41 9903
rect 797 9903 869 9947
rect -31 9519 41 9563
rect 797 9563 810 9903
rect 856 9563 869 9903
rect 797 9519 869 9563
rect -31 9447 869 9519
rect 1455 9948 2355 10020
rect 1455 9904 1527 9948
rect 1455 9564 1468 9904
rect 1514 9564 1527 9904
rect 2283 9904 2355 9948
rect 1455 9520 1527 9564
rect 2283 9564 2296 9904
rect 2342 9564 2355 9904
rect 2283 9520 2355 9564
rect 1455 9448 2355 9520
rect 4011 9947 4911 10019
rect 4011 9903 4083 9947
rect 4011 9563 4024 9903
rect 4070 9563 4083 9903
rect 4839 9903 4911 9947
rect 4011 9519 4083 9563
rect 4839 9563 4852 9903
rect 4898 9563 4911 9903
rect 4839 9519 4911 9563
rect 4011 9447 4911 9519
rect 5497 9948 6397 10020
rect 5497 9904 5569 9948
rect 5497 9564 5510 9904
rect 5556 9564 5569 9904
rect 6325 9904 6397 9948
rect 5497 9520 5569 9564
rect 6325 9564 6338 9904
rect 6384 9564 6397 9904
rect 6325 9520 6397 9564
rect 5497 9448 6397 9520
rect 8053 9947 8953 10019
rect 8053 9903 8125 9947
rect 8053 9563 8066 9903
rect 8112 9563 8125 9903
rect 8881 9903 8953 9947
rect 8053 9519 8125 9563
rect 8881 9563 8894 9903
rect 8940 9563 8953 9903
rect 8881 9519 8953 9563
rect 8053 9447 8953 9519
rect 9539 9948 10439 10020
rect 9539 9904 9611 9948
rect 9539 9564 9552 9904
rect 9598 9564 9611 9904
rect 10367 9904 10439 9948
rect 9539 9520 9611 9564
rect 10367 9564 10380 9904
rect 10426 9564 10439 9904
rect 10367 9520 10439 9564
rect 9539 9448 10439 9520
rect 12095 9947 12995 10019
rect 12095 9903 12167 9947
rect 12095 9563 12108 9903
rect 12154 9563 12167 9903
rect 12923 9903 12995 9947
rect 12095 9519 12167 9563
rect 12923 9563 12936 9903
rect 12982 9563 12995 9903
rect 12923 9519 12995 9563
rect 12095 9447 12995 9519
rect 13581 9948 14481 10020
rect 13581 9904 13653 9948
rect 13581 9564 13594 9904
rect 13640 9564 13653 9904
rect 14409 9904 14481 9948
rect 13581 9520 13653 9564
rect 14409 9564 14422 9904
rect 14468 9564 14481 9904
rect 14409 9520 14481 9564
rect 13581 9448 14481 9520
rect -12127 7742 -11227 7814
rect -12127 7698 -12055 7742
rect -12127 7358 -12114 7698
rect -12068 7358 -12055 7698
rect -11299 7698 -11227 7742
rect -12127 7314 -12055 7358
rect -11299 7358 -11286 7698
rect -11240 7358 -11227 7698
rect -11299 7314 -11227 7358
rect -12127 7242 -11227 7314
rect -8115 7742 -7215 7814
rect -8115 7698 -8043 7742
rect -8115 7358 -8102 7698
rect -8056 7358 -8043 7698
rect -7287 7698 -7215 7742
rect -8115 7314 -8043 7358
rect -7287 7358 -7274 7698
rect -7228 7358 -7215 7698
rect -7287 7314 -7215 7358
rect -8115 7242 -7215 7314
rect -4073 7742 -3173 7814
rect -4073 7698 -4001 7742
rect -4073 7358 -4060 7698
rect -4014 7358 -4001 7698
rect -3245 7698 -3173 7742
rect -4073 7314 -4001 7358
rect -3245 7358 -3232 7698
rect -3186 7358 -3173 7698
rect -3245 7314 -3173 7358
rect -4073 7242 -3173 7314
rect -31 7742 869 7814
rect -31 7698 41 7742
rect -31 7358 -18 7698
rect 28 7358 41 7698
rect 797 7698 869 7742
rect -31 7314 41 7358
rect 797 7358 810 7698
rect 856 7358 869 7698
rect 797 7314 869 7358
rect -31 7242 869 7314
rect 4011 7742 4911 7814
rect 4011 7698 4083 7742
rect 4011 7358 4024 7698
rect 4070 7358 4083 7698
rect 4839 7698 4911 7742
rect 4011 7314 4083 7358
rect 4839 7358 4852 7698
rect 4898 7358 4911 7698
rect 4839 7314 4911 7358
rect 4011 7242 4911 7314
rect 8053 7742 8953 7814
rect 8053 7698 8125 7742
rect 8053 7358 8066 7698
rect 8112 7358 8125 7698
rect 8881 7698 8953 7742
rect 8053 7314 8125 7358
rect 8881 7358 8894 7698
rect 8940 7358 8953 7698
rect 8881 7314 8953 7358
rect 8053 7242 8953 7314
rect 12095 7742 12995 7814
rect 12095 7698 12167 7742
rect 12095 7358 12108 7698
rect 12154 7358 12167 7698
rect 12923 7698 12995 7742
rect 12095 7314 12167 7358
rect 12923 7358 12936 7698
rect 12982 7358 12995 7698
rect 12923 7314 12995 7358
rect 12095 7242 12995 7314
rect -10831 4278 -10681 4300
rect -10831 4232 -10779 4278
rect -10733 4232 -10681 4278
rect -10831 4210 -10681 4232
rect -10591 4278 -10441 4300
rect -10591 4232 -10539 4278
rect -10493 4232 -10441 4278
rect -10591 4210 -10441 4232
rect -10351 4278 -10201 4300
rect -10351 4232 -10299 4278
rect -10253 4232 -10201 4278
rect -10351 4210 -10201 4232
rect -10111 4278 -9961 4300
rect -10111 4232 -10059 4278
rect -10013 4232 -9961 4278
rect -10111 4210 -9961 4232
rect -8657 4161 -7665 4233
rect -8657 4117 -8585 4161
rect -8657 3777 -8644 4117
rect -8598 3777 -8585 4117
rect -8197 4117 -8125 4161
rect -8657 3733 -8585 3777
rect -8197 3777 -8184 4117
rect -8138 3777 -8125 4117
rect -7737 4117 -7665 4161
rect -8197 3733 -8125 3777
rect -7737 3777 -7724 4117
rect -7678 3777 -7665 4117
rect -7737 3733 -7665 3777
rect -8657 3661 -7665 3733
rect -9627 3228 -9095 3300
rect -9627 2648 -9555 3228
rect -9167 2648 -9095 3228
rect -9627 2635 -9095 2648
rect -9627 2589 -9511 2635
rect -9211 2589 -9095 2635
rect -9627 2576 -9095 2589
rect -7227 3228 -6695 3300
rect -7227 2648 -7155 3228
rect -6767 2648 -6695 3228
rect -7227 2635 -6695 2648
rect -7227 2589 -7111 2635
rect -6811 2589 -6695 2635
rect -7227 2576 -6695 2589
rect -9993 855 -6329 927
rect -9993 811 -9921 855
rect -9993 271 -9980 811
rect -9934 271 -9921 811
rect -8197 811 -8125 855
rect -9993 227 -9921 271
rect -8197 271 -8184 811
rect -8138 271 -8125 811
rect -6401 811 -6329 855
rect -8197 227 -8125 271
rect -6401 271 -6388 811
rect -6342 271 -6329 811
rect -6401 227 -6329 271
rect -9993 155 -6329 227
rect -10354 -304 -5968 -232
rect -10354 -403 -10154 -304
rect -10354 -903 -10304 -403
rect -10204 -903 -10154 -403
rect -6168 -403 -5968 -304
rect -10354 -1848 -10154 -903
rect -6168 -903 -6118 -403
rect -6018 -903 -5968 -403
rect -10354 -2348 -10304 -1848
rect -10204 -2348 -10154 -1848
rect -6168 -1848 -5968 -903
rect -10354 -2447 -10154 -2348
rect -6168 -2348 -6118 -1848
rect -6018 -2348 -5968 -1848
rect -6168 -2447 -5968 -2348
rect -10354 -2519 -5968 -2447
rect -8611 -2563 -8539 -2519
rect -8611 -2863 -8598 -2563
rect -8552 -2863 -8539 -2563
rect -7783 -2563 -7711 -2519
rect -8611 -2907 -8539 -2863
rect -7783 -2863 -7770 -2563
rect -7724 -2863 -7711 -2563
rect -7783 -2907 -7711 -2863
rect -8611 -2979 -7711 -2907
<< nsubdiff >>
rect 40051 39021 40201 39043
rect 40051 38975 40103 39021
rect 40149 38975 40201 39021
rect 40051 38953 40201 38975
rect 40291 39021 40441 39043
rect 40291 38975 40343 39021
rect 40389 38975 40441 39021
rect 40291 38953 40441 38975
rect 40531 39021 40681 39043
rect 40531 38975 40583 39021
rect 40629 38975 40681 39021
rect 40531 38953 40681 38975
rect 40771 39021 40921 39043
rect 40771 38975 40823 39021
rect 40869 38975 40921 39021
rect 40771 38953 40921 38975
rect -4857 37398 -3957 37470
rect -4857 37354 -4785 37398
rect -4857 36714 -4844 37354
rect -4798 36714 -4785 37354
rect -4029 37354 -3957 37398
rect -4857 36670 -4785 36714
rect -4029 36714 -4016 37354
rect -3970 36714 -3957 37354
rect -4029 36670 -3957 36714
rect -4857 36598 -3957 36670
rect 4615 37398 5515 37470
rect 4615 37354 4687 37398
rect 4615 36714 4628 37354
rect 4674 36714 4687 37354
rect 5443 37354 5515 37398
rect 4615 36670 4687 36714
rect 5443 36714 5456 37354
rect 5502 36714 5515 37354
rect 5443 36670 5515 36714
rect 4615 36598 5515 36670
rect 14087 37399 14987 37471
rect 14087 37355 14159 37399
rect 14087 36715 14100 37355
rect 14146 36715 14159 37355
rect 14915 37355 14987 37399
rect 14087 36671 14159 36715
rect 14915 36715 14928 37355
rect 14974 36715 14987 37355
rect 14915 36671 14987 36715
rect 14087 36599 14987 36671
rect 23559 37399 24459 37471
rect 23559 37355 23631 37399
rect 23559 36715 23572 37355
rect 23618 36715 23631 37355
rect 24387 37355 24459 37399
rect 23559 36671 23631 36715
rect 24387 36715 24400 37355
rect 24446 36715 24459 37355
rect 24387 36671 24459 36715
rect 23559 36599 24459 36671
rect 33031 37399 33931 37471
rect 33031 37355 33103 37399
rect 33031 36715 33044 37355
rect 33090 36715 33103 37355
rect 33859 37355 33931 37399
rect 33031 36671 33103 36715
rect 33859 36715 33872 37355
rect 33918 36715 33931 37355
rect 33859 36671 33931 36715
rect 33031 36599 33931 36671
rect 42503 37399 43403 37471
rect 42503 37355 42575 37399
rect 42503 36715 42516 37355
rect 42562 36715 42575 37355
rect 43331 37355 43403 37399
rect 42503 36671 42575 36715
rect 43331 36715 43344 37355
rect 43390 36715 43403 37355
rect 43331 36671 43403 36715
rect 42503 36599 43403 36671
rect -4857 35193 -3957 35265
rect -4857 35149 -4785 35193
rect -4857 34509 -4844 35149
rect -4798 34509 -4785 35149
rect -4029 35149 -3957 35193
rect -4857 34465 -4785 34509
rect -4029 34509 -4016 35149
rect -3970 34509 -3957 35149
rect -4029 34465 -3957 34509
rect -4857 34393 -3957 34465
rect -3371 35193 -2471 35265
rect -3371 35149 -3299 35193
rect -3371 34509 -3358 35149
rect -3312 34509 -3299 35149
rect -2543 35149 -2471 35193
rect -3371 34465 -3299 34509
rect -2543 34509 -2530 35149
rect -2484 34509 -2471 35149
rect -2543 34465 -2471 34509
rect -3371 34393 -2471 34465
rect 4615 35193 5515 35265
rect 4615 35149 4687 35193
rect 4615 34509 4628 35149
rect 4674 34509 4687 35149
rect 5443 35149 5515 35193
rect 4615 34465 4687 34509
rect 5443 34509 5456 35149
rect 5502 34509 5515 35149
rect 5443 34465 5515 34509
rect 4615 34393 5515 34465
rect 6101 35193 7001 35265
rect 6101 35149 6173 35193
rect 6101 34509 6114 35149
rect 6160 34509 6173 35149
rect 6929 35149 7001 35193
rect 6101 34465 6173 34509
rect 6929 34509 6942 35149
rect 6988 34509 7001 35149
rect 6929 34465 7001 34509
rect 6101 34393 7001 34465
rect 14087 35194 14987 35266
rect 14087 35150 14159 35194
rect 14087 34510 14100 35150
rect 14146 34510 14159 35150
rect 14915 35150 14987 35194
rect 14087 34466 14159 34510
rect 14915 34510 14928 35150
rect 14974 34510 14987 35150
rect 14915 34466 14987 34510
rect 14087 34394 14987 34466
rect 15573 35194 16473 35266
rect 15573 35150 15645 35194
rect 15573 34510 15586 35150
rect 15632 34510 15645 35150
rect 16401 35150 16473 35194
rect 15573 34466 15645 34510
rect 16401 34510 16414 35150
rect 16460 34510 16473 35150
rect 16401 34466 16473 34510
rect 15573 34394 16473 34466
rect 23559 35194 24459 35266
rect 23559 35150 23631 35194
rect 23559 34510 23572 35150
rect 23618 34510 23631 35150
rect 24387 35150 24459 35194
rect 23559 34466 23631 34510
rect 24387 34510 24400 35150
rect 24446 34510 24459 35150
rect 24387 34466 24459 34510
rect 23559 34394 24459 34466
rect 25045 35194 25945 35266
rect 25045 35150 25117 35194
rect 25045 34510 25058 35150
rect 25104 34510 25117 35150
rect 25873 35150 25945 35194
rect 25045 34466 25117 34510
rect 25873 34510 25886 35150
rect 25932 34510 25945 35150
rect 25873 34466 25945 34510
rect 25045 34394 25945 34466
rect 33031 35194 33931 35266
rect 33031 35150 33103 35194
rect 33031 34510 33044 35150
rect 33090 34510 33103 35150
rect 33859 35150 33931 35194
rect 33031 34466 33103 34510
rect 33859 34510 33872 35150
rect 33918 34510 33931 35150
rect 33859 34466 33931 34510
rect 33031 34394 33931 34466
rect 34517 35194 35417 35266
rect 34517 35150 34589 35194
rect 34517 34510 34530 35150
rect 34576 34510 34589 35150
rect 35345 35150 35417 35194
rect 34517 34466 34589 34510
rect 35345 34510 35358 35150
rect 35404 34510 35417 35150
rect 35345 34466 35417 34510
rect 34517 34394 35417 34466
rect 42503 35194 43403 35266
rect 42503 35150 42575 35194
rect 42503 34510 42516 35150
rect 42562 34510 42575 35150
rect 43331 35150 43403 35194
rect 42503 34466 42575 34510
rect 43331 34510 43344 35150
rect 43390 34510 43403 35150
rect 43331 34466 43403 34510
rect 42503 34394 43403 34466
rect 43989 35194 44889 35266
rect 43989 35150 44061 35194
rect 43989 34510 44002 35150
rect 44048 34510 44061 35150
rect 44817 35150 44889 35194
rect 43989 34466 44061 34510
rect 44817 34510 44830 35150
rect 44876 34510 44889 35150
rect 44817 34466 44889 34510
rect 43989 34394 44889 34466
rect -4857 32988 -3957 33060
rect -4857 32944 -4785 32988
rect -4857 32304 -4844 32944
rect -4798 32304 -4785 32944
rect -4029 32944 -3957 32988
rect -4857 32260 -4785 32304
rect -4029 32304 -4016 32944
rect -3970 32304 -3957 32944
rect -4029 32260 -3957 32304
rect -4857 32188 -3957 32260
rect -3371 32989 -2471 33061
rect -3371 32945 -3299 32989
rect -3371 32305 -3358 32945
rect -3312 32305 -3299 32945
rect -2543 32945 -2471 32989
rect -3371 32261 -3299 32305
rect -2543 32305 -2530 32945
rect -2484 32305 -2471 32945
rect -2543 32261 -2471 32305
rect -3371 32189 -2471 32261
rect 4615 32988 5515 33060
rect 4615 32944 4687 32988
rect 4615 32304 4628 32944
rect 4674 32304 4687 32944
rect 5443 32944 5515 32988
rect 4615 32260 4687 32304
rect 5443 32304 5456 32944
rect 5502 32304 5515 32944
rect 5443 32260 5515 32304
rect 4615 32188 5515 32260
rect 6101 32989 7001 33061
rect 6101 32945 6173 32989
rect 6101 32305 6114 32945
rect 6160 32305 6173 32945
rect 6929 32945 7001 32989
rect 6101 32261 6173 32305
rect 6929 32305 6942 32945
rect 6988 32305 7001 32945
rect 6929 32261 7001 32305
rect 6101 32189 7001 32261
rect 14087 32989 14987 33061
rect 14087 32945 14159 32989
rect 14087 32305 14100 32945
rect 14146 32305 14159 32945
rect 14915 32945 14987 32989
rect 14087 32261 14159 32305
rect 14915 32305 14928 32945
rect 14974 32305 14987 32945
rect 14915 32261 14987 32305
rect 14087 32189 14987 32261
rect 15573 32990 16473 33062
rect 15573 32946 15645 32990
rect 15573 32306 15586 32946
rect 15632 32306 15645 32946
rect 16401 32946 16473 32990
rect 15573 32262 15645 32306
rect 16401 32306 16414 32946
rect 16460 32306 16473 32946
rect 16401 32262 16473 32306
rect 15573 32190 16473 32262
rect 23559 32989 24459 33061
rect 23559 32945 23631 32989
rect 23559 32305 23572 32945
rect 23618 32305 23631 32945
rect 24387 32945 24459 32989
rect 23559 32261 23631 32305
rect 24387 32305 24400 32945
rect 24446 32305 24459 32945
rect 24387 32261 24459 32305
rect 23559 32189 24459 32261
rect 25045 32990 25945 33062
rect 25045 32946 25117 32990
rect 25045 32306 25058 32946
rect 25104 32306 25117 32946
rect 25873 32946 25945 32990
rect 25045 32262 25117 32306
rect 25873 32306 25886 32946
rect 25932 32306 25945 32946
rect 25873 32262 25945 32306
rect 25045 32190 25945 32262
rect 33031 32989 33931 33061
rect 33031 32945 33103 32989
rect 33031 32305 33044 32945
rect 33090 32305 33103 32945
rect 33859 32945 33931 32989
rect 33031 32261 33103 32305
rect 33859 32305 33872 32945
rect 33918 32305 33931 32945
rect 33859 32261 33931 32305
rect 33031 32189 33931 32261
rect 34517 32990 35417 33062
rect 34517 32946 34589 32990
rect 34517 32306 34530 32946
rect 34576 32306 34589 32946
rect 35345 32946 35417 32990
rect 34517 32262 34589 32306
rect 35345 32306 35358 32946
rect 35404 32306 35417 32946
rect 35345 32262 35417 32306
rect 34517 32190 35417 32262
rect 42503 32989 43403 33061
rect 42503 32945 42575 32989
rect 42503 32305 42516 32945
rect 42562 32305 42575 32945
rect 43331 32945 43403 32989
rect 42503 32261 42575 32305
rect 43331 32305 43344 32945
rect 43390 32305 43403 32945
rect 43331 32261 43403 32305
rect 42503 32189 43403 32261
rect 43989 32990 44889 33062
rect 43989 32946 44061 32990
rect 43989 32306 44002 32946
rect 44048 32306 44061 32946
rect 44817 32946 44889 32990
rect 43989 32262 44061 32306
rect 44817 32306 44830 32946
rect 44876 32306 44889 32946
rect 44817 32262 44889 32306
rect 43989 32190 44889 32262
rect -9999 31873 -9447 31945
rect -9999 31829 -9927 31873
rect -9999 31089 -9986 31829
rect -9940 31089 -9927 31829
rect -9519 31829 -9447 31873
rect -9999 31045 -9927 31089
rect -9519 31089 -9506 31829
rect -9460 31089 -9447 31829
rect -9519 31045 -9447 31089
rect -9999 30973 -9447 31045
rect -9111 31873 -8079 31945
rect -9111 31829 -9039 31873
rect -9111 31089 -9098 31829
rect -9052 31089 -9039 31829
rect -8631 31829 -8559 31873
rect -9111 31045 -9039 31089
rect -8631 31089 -8618 31829
rect -8572 31089 -8559 31829
rect -8151 31829 -8079 31873
rect -8631 31045 -8559 31089
rect -8151 31089 -8138 31829
rect -8092 31089 -8079 31829
rect -527 31873 25 31945
rect -527 31829 -455 31873
rect -8151 31045 -8079 31089
rect -9111 30973 -8079 31045
rect -527 31089 -514 31829
rect -468 31089 -455 31829
rect -47 31829 25 31873
rect -527 31045 -455 31089
rect -47 31089 -34 31829
rect 12 31089 25 31829
rect -47 31045 25 31089
rect -527 30973 25 31045
rect 361 31873 1393 31945
rect 361 31829 433 31873
rect 361 31089 374 31829
rect 420 31089 433 31829
rect 841 31829 913 31873
rect 361 31045 433 31089
rect 841 31089 854 31829
rect 900 31089 913 31829
rect 1321 31829 1393 31873
rect 841 31045 913 31089
rect 1321 31089 1334 31829
rect 1380 31089 1393 31829
rect 8945 31874 9497 31946
rect 8945 31830 9017 31874
rect 1321 31045 1393 31089
rect 361 30973 1393 31045
rect 8945 31090 8958 31830
rect 9004 31090 9017 31830
rect 9425 31830 9497 31874
rect 8945 31046 9017 31090
rect 9425 31090 9438 31830
rect 9484 31090 9497 31830
rect 9425 31046 9497 31090
rect 8945 30974 9497 31046
rect 9833 31874 10865 31946
rect 9833 31830 9905 31874
rect 9833 31090 9846 31830
rect 9892 31090 9905 31830
rect 10313 31830 10385 31874
rect 9833 31046 9905 31090
rect 10313 31090 10326 31830
rect 10372 31090 10385 31830
rect 10793 31830 10865 31874
rect 10313 31046 10385 31090
rect 10793 31090 10806 31830
rect 10852 31090 10865 31830
rect 18417 31874 18969 31946
rect 18417 31830 18489 31874
rect 10793 31046 10865 31090
rect 9833 30974 10865 31046
rect 18417 31090 18430 31830
rect 18476 31090 18489 31830
rect 18897 31830 18969 31874
rect 18417 31046 18489 31090
rect 18897 31090 18910 31830
rect 18956 31090 18969 31830
rect 18897 31046 18969 31090
rect 18417 30974 18969 31046
rect 19305 31874 20337 31946
rect 19305 31830 19377 31874
rect 19305 31090 19318 31830
rect 19364 31090 19377 31830
rect 19785 31830 19857 31874
rect 19305 31046 19377 31090
rect 19785 31090 19798 31830
rect 19844 31090 19857 31830
rect 20265 31830 20337 31874
rect 19785 31046 19857 31090
rect 20265 31090 20278 31830
rect 20324 31090 20337 31830
rect 27889 31874 28441 31946
rect 27889 31830 27961 31874
rect 20265 31046 20337 31090
rect 19305 30974 20337 31046
rect 27889 31090 27902 31830
rect 27948 31090 27961 31830
rect 28369 31830 28441 31874
rect 27889 31046 27961 31090
rect 28369 31090 28382 31830
rect 28428 31090 28441 31830
rect 28369 31046 28441 31090
rect 27889 30974 28441 31046
rect 28777 31874 29809 31946
rect 28777 31830 28849 31874
rect 28777 31090 28790 31830
rect 28836 31090 28849 31830
rect 29257 31830 29329 31874
rect 28777 31046 28849 31090
rect 29257 31090 29270 31830
rect 29316 31090 29329 31830
rect 29737 31830 29809 31874
rect 29257 31046 29329 31090
rect 29737 31090 29750 31830
rect 29796 31090 29809 31830
rect 37361 31874 37913 31946
rect 37361 31830 37433 31874
rect 29737 31046 29809 31090
rect 28777 30974 29809 31046
rect 37361 31090 37374 31830
rect 37420 31090 37433 31830
rect 37841 31830 37913 31874
rect 37361 31046 37433 31090
rect 37841 31090 37854 31830
rect 37900 31090 37913 31830
rect 37841 31046 37913 31090
rect 37361 30974 37913 31046
rect 38249 31874 39281 31946
rect 38249 31830 38321 31874
rect 38249 31090 38262 31830
rect 38308 31090 38321 31830
rect 38729 31830 38801 31874
rect 38249 31046 38321 31090
rect 38729 31090 38742 31830
rect 38788 31090 38801 31830
rect 39209 31830 39281 31874
rect 38729 31046 38801 31090
rect 39209 31090 39222 31830
rect 39268 31090 39281 31830
rect 39209 31046 39281 31090
rect 38249 30974 39281 31046
rect -4857 30783 -3957 30855
rect -10893 30453 -10341 30525
rect -10893 30409 -10821 30453
rect -10893 29669 -10880 30409
rect -10834 29669 -10821 30409
rect -10413 30409 -10341 30453
rect -10893 29625 -10821 29669
rect -10413 29669 -10400 30409
rect -10354 29669 -10341 30409
rect -7771 30697 -5851 30769
rect -7771 30653 -7699 30697
rect -7771 29913 -7758 30653
rect -7712 29913 -7699 30653
rect -7087 30653 -7015 30697
rect -7771 29869 -7699 29913
rect -7087 29913 -7074 30653
rect -7028 29913 -7015 30653
rect -6403 30653 -6331 30697
rect -7087 29869 -7015 29913
rect -6403 29913 -6390 30653
rect -6344 29913 -6331 30653
rect -5923 30653 -5851 30697
rect -6403 29869 -6331 29913
rect -5923 29913 -5910 30653
rect -5864 29913 -5851 30653
rect -4857 30739 -4785 30783
rect -4857 30099 -4844 30739
rect -4798 30099 -4785 30739
rect -4029 30739 -3957 30783
rect -4857 30055 -4785 30099
rect -4029 30099 -4016 30739
rect -3970 30099 -3957 30739
rect 4615 30783 5515 30855
rect -4029 30055 -3957 30099
rect -4857 29983 -3957 30055
rect -1421 30453 -869 30525
rect -1421 30409 -1349 30453
rect -5923 29869 -5851 29913
rect -7771 29797 -5851 29869
rect -10413 29625 -10341 29669
rect -10893 29553 -10341 29625
rect -9999 29533 -9447 29605
rect -9999 29489 -9927 29533
rect -9999 28749 -9986 29489
rect -9940 28749 -9927 29489
rect -9519 29489 -9447 29533
rect -9999 28705 -9927 28749
rect -9519 28749 -9506 29489
rect -9460 28749 -9447 29489
rect -9519 28705 -9447 28749
rect -9999 28633 -9447 28705
rect -9111 29533 -8079 29605
rect -9111 29489 -9039 29533
rect -9111 28749 -9098 29489
rect -9052 28749 -9039 29489
rect -8631 29489 -8559 29533
rect -9111 28705 -9039 28749
rect -8631 28749 -8618 29489
rect -8572 28749 -8559 29489
rect -8151 29489 -8079 29533
rect -8631 28705 -8559 28749
rect -8151 28749 -8138 29489
rect -8092 28749 -8079 29489
rect -1421 29669 -1408 30409
rect -1362 29669 -1349 30409
rect -941 30409 -869 30453
rect -1421 29625 -1349 29669
rect -941 29669 -928 30409
rect -882 29669 -869 30409
rect 1701 30697 3621 30769
rect 1701 30653 1773 30697
rect 1701 29913 1714 30653
rect 1760 29913 1773 30653
rect 2385 30653 2457 30697
rect 1701 29869 1773 29913
rect 2385 29913 2398 30653
rect 2444 29913 2457 30653
rect 3069 30653 3141 30697
rect 2385 29869 2457 29913
rect 3069 29913 3082 30653
rect 3128 29913 3141 30653
rect 3549 30653 3621 30697
rect 3069 29869 3141 29913
rect 3549 29913 3562 30653
rect 3608 29913 3621 30653
rect 4615 30739 4687 30783
rect 4615 30099 4628 30739
rect 4674 30099 4687 30739
rect 5443 30739 5515 30783
rect 4615 30055 4687 30099
rect 5443 30099 5456 30739
rect 5502 30099 5515 30739
rect 14087 30784 14987 30856
rect 5443 30055 5515 30099
rect 4615 29983 5515 30055
rect 8051 30454 8603 30526
rect 8051 30410 8123 30454
rect 3549 29869 3621 29913
rect 1701 29797 3621 29869
rect -941 29625 -869 29669
rect -1421 29553 -869 29625
rect -527 29533 25 29605
rect -527 29489 -455 29533
rect -8151 28705 -8079 28749
rect -9111 28633 -8079 28705
rect -527 28749 -514 29489
rect -468 28749 -455 29489
rect -47 29489 25 29533
rect -527 28705 -455 28749
rect -47 28749 -34 29489
rect 12 28749 25 29489
rect -47 28705 25 28749
rect -527 28633 25 28705
rect 361 29533 1393 29605
rect 361 29489 433 29533
rect 361 28749 374 29489
rect 420 28749 433 29489
rect 841 29489 913 29533
rect 361 28705 433 28749
rect 841 28749 854 29489
rect 900 28749 913 29489
rect 1321 29489 1393 29533
rect 841 28705 913 28749
rect 1321 28749 1334 29489
rect 1380 28749 1393 29489
rect 8051 29670 8064 30410
rect 8110 29670 8123 30410
rect 8531 30410 8603 30454
rect 8051 29626 8123 29670
rect 8531 29670 8544 30410
rect 8590 29670 8603 30410
rect 11173 30698 13093 30770
rect 11173 30654 11245 30698
rect 11173 29914 11186 30654
rect 11232 29914 11245 30654
rect 11857 30654 11929 30698
rect 11173 29870 11245 29914
rect 11857 29914 11870 30654
rect 11916 29914 11929 30654
rect 12541 30654 12613 30698
rect 11857 29870 11929 29914
rect 12541 29914 12554 30654
rect 12600 29914 12613 30654
rect 13021 30654 13093 30698
rect 12541 29870 12613 29914
rect 13021 29914 13034 30654
rect 13080 29914 13093 30654
rect 14087 30740 14159 30784
rect 14087 30100 14100 30740
rect 14146 30100 14159 30740
rect 14915 30740 14987 30784
rect 14087 30056 14159 30100
rect 14915 30100 14928 30740
rect 14974 30100 14987 30740
rect 23559 30784 24459 30856
rect 14915 30056 14987 30100
rect 14087 29984 14987 30056
rect 17523 30454 18075 30526
rect 17523 30410 17595 30454
rect 13021 29870 13093 29914
rect 11173 29798 13093 29870
rect 8531 29626 8603 29670
rect 8051 29554 8603 29626
rect 8945 29534 9497 29606
rect 8945 29490 9017 29534
rect 1321 28705 1393 28749
rect 361 28633 1393 28705
rect 8945 28750 8958 29490
rect 9004 28750 9017 29490
rect 9425 29490 9497 29534
rect 8945 28706 9017 28750
rect 9425 28750 9438 29490
rect 9484 28750 9497 29490
rect 9425 28706 9497 28750
rect 8945 28634 9497 28706
rect 9833 29534 10865 29606
rect 9833 29490 9905 29534
rect 9833 28750 9846 29490
rect 9892 28750 9905 29490
rect 10313 29490 10385 29534
rect 9833 28706 9905 28750
rect 10313 28750 10326 29490
rect 10372 28750 10385 29490
rect 10793 29490 10865 29534
rect 10313 28706 10385 28750
rect 10793 28750 10806 29490
rect 10852 28750 10865 29490
rect 17523 29670 17536 30410
rect 17582 29670 17595 30410
rect 18003 30410 18075 30454
rect 17523 29626 17595 29670
rect 18003 29670 18016 30410
rect 18062 29670 18075 30410
rect 20645 30698 22565 30770
rect 20645 30654 20717 30698
rect 20645 29914 20658 30654
rect 20704 29914 20717 30654
rect 21329 30654 21401 30698
rect 20645 29870 20717 29914
rect 21329 29914 21342 30654
rect 21388 29914 21401 30654
rect 22013 30654 22085 30698
rect 21329 29870 21401 29914
rect 22013 29914 22026 30654
rect 22072 29914 22085 30654
rect 22493 30654 22565 30698
rect 22013 29870 22085 29914
rect 22493 29914 22506 30654
rect 22552 29914 22565 30654
rect 23559 30740 23631 30784
rect 23559 30100 23572 30740
rect 23618 30100 23631 30740
rect 24387 30740 24459 30784
rect 23559 30056 23631 30100
rect 24387 30100 24400 30740
rect 24446 30100 24459 30740
rect 33031 30784 33931 30856
rect 24387 30056 24459 30100
rect 23559 29984 24459 30056
rect 26995 30454 27547 30526
rect 26995 30410 27067 30454
rect 22493 29870 22565 29914
rect 20645 29798 22565 29870
rect 18003 29626 18075 29670
rect 17523 29554 18075 29626
rect 18417 29534 18969 29606
rect 18417 29490 18489 29534
rect 10793 28706 10865 28750
rect 9833 28634 10865 28706
rect 18417 28750 18430 29490
rect 18476 28750 18489 29490
rect 18897 29490 18969 29534
rect 18417 28706 18489 28750
rect 18897 28750 18910 29490
rect 18956 28750 18969 29490
rect 18897 28706 18969 28750
rect 18417 28634 18969 28706
rect 19305 29534 20337 29606
rect 19305 29490 19377 29534
rect 19305 28750 19318 29490
rect 19364 28750 19377 29490
rect 19785 29490 19857 29534
rect 19305 28706 19377 28750
rect 19785 28750 19798 29490
rect 19844 28750 19857 29490
rect 20265 29490 20337 29534
rect 19785 28706 19857 28750
rect 20265 28750 20278 29490
rect 20324 28750 20337 29490
rect 26995 29670 27008 30410
rect 27054 29670 27067 30410
rect 27475 30410 27547 30454
rect 26995 29626 27067 29670
rect 27475 29670 27488 30410
rect 27534 29670 27547 30410
rect 30117 30698 32037 30770
rect 30117 30654 30189 30698
rect 30117 29914 30130 30654
rect 30176 29914 30189 30654
rect 30801 30654 30873 30698
rect 30117 29870 30189 29914
rect 30801 29914 30814 30654
rect 30860 29914 30873 30654
rect 31485 30654 31557 30698
rect 30801 29870 30873 29914
rect 31485 29914 31498 30654
rect 31544 29914 31557 30654
rect 31965 30654 32037 30698
rect 31485 29870 31557 29914
rect 31965 29914 31978 30654
rect 32024 29914 32037 30654
rect 33031 30740 33103 30784
rect 33031 30100 33044 30740
rect 33090 30100 33103 30740
rect 33859 30740 33931 30784
rect 33031 30056 33103 30100
rect 33859 30100 33872 30740
rect 33918 30100 33931 30740
rect 42503 30784 43403 30856
rect 33859 30056 33931 30100
rect 33031 29984 33931 30056
rect 36467 30454 37019 30526
rect 36467 30410 36539 30454
rect 31965 29870 32037 29914
rect 30117 29798 32037 29870
rect 27475 29626 27547 29670
rect 26995 29554 27547 29626
rect 27889 29534 28441 29606
rect 27889 29490 27961 29534
rect 20265 28706 20337 28750
rect 19305 28634 20337 28706
rect 27889 28750 27902 29490
rect 27948 28750 27961 29490
rect 28369 29490 28441 29534
rect 27889 28706 27961 28750
rect 28369 28750 28382 29490
rect 28428 28750 28441 29490
rect 28369 28706 28441 28750
rect 27889 28634 28441 28706
rect 28777 29534 29809 29606
rect 28777 29490 28849 29534
rect 28777 28750 28790 29490
rect 28836 28750 28849 29490
rect 29257 29490 29329 29534
rect 28777 28706 28849 28750
rect 29257 28750 29270 29490
rect 29316 28750 29329 29490
rect 29737 29490 29809 29534
rect 29257 28706 29329 28750
rect 29737 28750 29750 29490
rect 29796 28750 29809 29490
rect 36467 29670 36480 30410
rect 36526 29670 36539 30410
rect 36947 30410 37019 30454
rect 36467 29626 36539 29670
rect 36947 29670 36960 30410
rect 37006 29670 37019 30410
rect 39589 30698 41509 30770
rect 39589 30654 39661 30698
rect 39589 29914 39602 30654
rect 39648 29914 39661 30654
rect 40273 30654 40345 30698
rect 39589 29870 39661 29914
rect 40273 29914 40286 30654
rect 40332 29914 40345 30654
rect 40957 30654 41029 30698
rect 40273 29870 40345 29914
rect 40957 29914 40970 30654
rect 41016 29914 41029 30654
rect 41437 30654 41509 30698
rect 40957 29870 41029 29914
rect 41437 29914 41450 30654
rect 41496 29914 41509 30654
rect 42503 30740 42575 30784
rect 42503 30100 42516 30740
rect 42562 30100 42575 30740
rect 43331 30740 43403 30784
rect 42503 30056 42575 30100
rect 43331 30100 43344 30740
rect 43390 30100 43403 30740
rect 43331 30056 43403 30100
rect 42503 29984 43403 30056
rect 41437 29870 41509 29914
rect 39589 29798 41509 29870
rect 36947 29626 37019 29670
rect 36467 29554 37019 29626
rect 37361 29534 37913 29606
rect 37361 29490 37433 29534
rect 29737 28706 29809 28750
rect 28777 28634 29809 28706
rect 37361 28750 37374 29490
rect 37420 28750 37433 29490
rect 37841 29490 37913 29534
rect 37361 28706 37433 28750
rect 37841 28750 37854 29490
rect 37900 28750 37913 29490
rect 37841 28706 37913 28750
rect 37361 28634 37913 28706
rect 38249 29534 39281 29606
rect 38249 29490 38321 29534
rect 38249 28750 38262 29490
rect 38308 28750 38321 29490
rect 38729 29490 38801 29534
rect 38249 28706 38321 28750
rect 38729 28750 38742 29490
rect 38788 28750 38801 29490
rect 39209 29490 39281 29534
rect 38729 28706 38801 28750
rect 39209 28750 39222 29490
rect 39268 28750 39281 29490
rect 39209 28706 39281 28750
rect 38249 28634 39281 28706
rect -12606 28523 -12054 28595
rect -12606 28479 -12534 28523
rect -12606 27739 -12593 28479
rect -12547 27739 -12534 28479
rect -12126 28479 -12054 28523
rect -12606 27695 -12534 27739
rect -12126 27739 -12113 28479
rect -12067 27739 -12054 28479
rect -12126 27695 -12054 27739
rect -12606 27623 -12054 27695
rect -8115 25096 -7215 25168
rect -8115 25052 -8043 25096
rect -8115 24412 -8102 25052
rect -8056 24412 -8043 25052
rect -7287 25052 -7215 25096
rect -8115 24368 -8043 24412
rect -7287 24412 -7274 25052
rect -7228 24412 -7215 25052
rect -7287 24368 -7215 24412
rect -8115 24296 -7215 24368
rect -4073 25093 -3173 25165
rect -4073 25049 -4001 25093
rect -4073 24409 -4060 25049
rect -4014 24409 -4001 25049
rect -3245 25049 -3173 25093
rect -4073 24365 -4001 24409
rect -3245 24409 -3232 25049
rect -3186 24409 -3173 25049
rect -3245 24365 -3173 24409
rect -4073 24293 -3173 24365
rect -31 25093 869 25165
rect -31 25049 41 25093
rect -31 24409 -18 25049
rect 28 24409 41 25049
rect 797 25049 869 25093
rect -31 24365 41 24409
rect 797 24409 810 25049
rect 856 24409 869 25049
rect 797 24365 869 24409
rect -31 24293 869 24365
rect 4011 25093 4911 25165
rect 4011 25049 4083 25093
rect 4011 24409 4024 25049
rect 4070 24409 4083 25049
rect 4839 25049 4911 25093
rect 4011 24365 4083 24409
rect 4839 24409 4852 25049
rect 4898 24409 4911 25049
rect 4839 24365 4911 24409
rect 4011 24293 4911 24365
rect 8053 25093 8953 25165
rect 8053 25049 8125 25093
rect 8053 24409 8066 25049
rect 8112 24409 8125 25049
rect 8881 25049 8953 25093
rect 8053 24365 8125 24409
rect 8881 24409 8894 25049
rect 8940 24409 8953 25049
rect 8881 24365 8953 24409
rect 8053 24293 8953 24365
rect 12095 25093 12995 25165
rect 12095 25049 12167 25093
rect 12095 24409 12108 25049
rect 12154 24409 12167 25049
rect 12923 25049 12995 25093
rect 12095 24365 12167 24409
rect 12923 24409 12936 25049
rect 12982 24409 12995 25049
rect 12923 24365 12995 24409
rect 12095 24293 12995 24365
rect 16137 25093 17037 25165
rect 16137 25049 16209 25093
rect 16137 24409 16150 25049
rect 16196 24409 16209 25049
rect 16965 25049 17037 25093
rect 16137 24365 16209 24409
rect 16965 24409 16978 25049
rect 17024 24409 17037 25049
rect 16965 24365 17037 24409
rect 16137 24293 17037 24365
rect -8115 22891 -7215 22963
rect -8115 22847 -8043 22891
rect -8115 22207 -8102 22847
rect -8056 22207 -8043 22847
rect -7287 22847 -7215 22891
rect -8115 22163 -8043 22207
rect -7287 22207 -7274 22847
rect -7228 22207 -7215 22847
rect -7287 22163 -7215 22207
rect -8115 22091 -7215 22163
rect -6629 22891 -5729 22963
rect -6629 22847 -6557 22891
rect -6629 22207 -6616 22847
rect -6570 22207 -6557 22847
rect -5801 22847 -5729 22891
rect -6629 22163 -6557 22207
rect -5801 22207 -5788 22847
rect -5742 22207 -5729 22847
rect -5801 22163 -5729 22207
rect -6629 22091 -5729 22163
rect -4073 22888 -3173 22960
rect -4073 22844 -4001 22888
rect -4073 22204 -4060 22844
rect -4014 22204 -4001 22844
rect -3245 22844 -3173 22888
rect -4073 22160 -4001 22204
rect -3245 22204 -3232 22844
rect -3186 22204 -3173 22844
rect -3245 22160 -3173 22204
rect -4073 22088 -3173 22160
rect -2587 22888 -1687 22960
rect -2587 22844 -2515 22888
rect -2587 22204 -2574 22844
rect -2528 22204 -2515 22844
rect -1759 22844 -1687 22888
rect -2587 22160 -2515 22204
rect -1759 22204 -1746 22844
rect -1700 22204 -1687 22844
rect -1759 22160 -1687 22204
rect -2587 22088 -1687 22160
rect -31 22888 869 22960
rect -31 22844 41 22888
rect -31 22204 -18 22844
rect 28 22204 41 22844
rect 797 22844 869 22888
rect -31 22160 41 22204
rect 797 22204 810 22844
rect 856 22204 869 22844
rect 797 22160 869 22204
rect -31 22088 869 22160
rect 1455 22888 2355 22960
rect 1455 22844 1527 22888
rect 1455 22204 1468 22844
rect 1514 22204 1527 22844
rect 2283 22844 2355 22888
rect 1455 22160 1527 22204
rect 2283 22204 2296 22844
rect 2342 22204 2355 22844
rect 2283 22160 2355 22204
rect 1455 22088 2355 22160
rect 4011 22888 4911 22960
rect 4011 22844 4083 22888
rect 4011 22204 4024 22844
rect 4070 22204 4083 22844
rect 4839 22844 4911 22888
rect 4011 22160 4083 22204
rect 4839 22204 4852 22844
rect 4898 22204 4911 22844
rect 4839 22160 4911 22204
rect 4011 22088 4911 22160
rect 5497 22888 6397 22960
rect 5497 22844 5569 22888
rect 5497 22204 5510 22844
rect 5556 22204 5569 22844
rect 6325 22844 6397 22888
rect 5497 22160 5569 22204
rect 6325 22204 6338 22844
rect 6384 22204 6397 22844
rect 6325 22160 6397 22204
rect 5497 22088 6397 22160
rect 8053 22888 8953 22960
rect 8053 22844 8125 22888
rect 8053 22204 8066 22844
rect 8112 22204 8125 22844
rect 8881 22844 8953 22888
rect 8053 22160 8125 22204
rect 8881 22204 8894 22844
rect 8940 22204 8953 22844
rect 8881 22160 8953 22204
rect 8053 22088 8953 22160
rect 9539 22888 10439 22960
rect 9539 22844 9611 22888
rect 9539 22204 9552 22844
rect 9598 22204 9611 22844
rect 10367 22844 10439 22888
rect 9539 22160 9611 22204
rect 10367 22204 10380 22844
rect 10426 22204 10439 22844
rect 10367 22160 10439 22204
rect 9539 22088 10439 22160
rect 12095 22888 12995 22960
rect 12095 22844 12167 22888
rect 12095 22204 12108 22844
rect 12154 22204 12167 22844
rect 12923 22844 12995 22888
rect 12095 22160 12167 22204
rect 12923 22204 12936 22844
rect 12982 22204 12995 22844
rect 12923 22160 12995 22204
rect 12095 22088 12995 22160
rect 13581 22888 14481 22960
rect 13581 22844 13653 22888
rect 13581 22204 13594 22844
rect 13640 22204 13653 22844
rect 14409 22844 14481 22888
rect 13581 22160 13653 22204
rect 14409 22204 14422 22844
rect 14468 22204 14481 22844
rect 14409 22160 14481 22204
rect 13581 22088 14481 22160
rect 16137 22888 17037 22960
rect 16137 22844 16209 22888
rect 16137 22204 16150 22844
rect 16196 22204 16209 22844
rect 16965 22844 17037 22888
rect 16137 22160 16209 22204
rect 16965 22204 16978 22844
rect 17024 22204 17037 22844
rect 16965 22160 17037 22204
rect 16137 22088 17037 22160
rect 17623 22888 18523 22960
rect 17623 22844 17695 22888
rect 17623 22204 17636 22844
rect 17682 22204 17695 22844
rect 18451 22844 18523 22888
rect 17623 22160 17695 22204
rect 18451 22204 18464 22844
rect 18510 22204 18523 22844
rect 18451 22160 18523 22204
rect 17623 22088 18523 22160
rect -8115 20686 -7215 20758
rect -8115 20642 -8043 20686
rect -8115 20002 -8102 20642
rect -8056 20002 -8043 20642
rect -7287 20642 -7215 20686
rect -8115 19958 -8043 20002
rect -7287 20002 -7274 20642
rect -7228 20002 -7215 20642
rect -7287 19958 -7215 20002
rect -8115 19886 -7215 19958
rect -6629 20687 -5729 20759
rect -6629 20643 -6557 20687
rect -6629 20003 -6616 20643
rect -6570 20003 -6557 20643
rect -5801 20643 -5729 20687
rect -6629 19959 -6557 20003
rect -5801 20003 -5788 20643
rect -5742 20003 -5729 20643
rect -5801 19959 -5729 20003
rect -6629 19887 -5729 19959
rect -4073 20683 -3173 20755
rect -4073 20639 -4001 20683
rect -4073 19999 -4060 20639
rect -4014 19999 -4001 20639
rect -3245 20639 -3173 20683
rect -4073 19955 -4001 19999
rect -3245 19999 -3232 20639
rect -3186 19999 -3173 20639
rect -3245 19955 -3173 19999
rect -4073 19883 -3173 19955
rect -2587 20684 -1687 20756
rect -2587 20640 -2515 20684
rect -2587 20000 -2574 20640
rect -2528 20000 -2515 20640
rect -1759 20640 -1687 20684
rect -2587 19956 -2515 20000
rect -1759 20000 -1746 20640
rect -1700 20000 -1687 20640
rect -1759 19956 -1687 20000
rect -2587 19884 -1687 19956
rect -31 20683 869 20755
rect -31 20639 41 20683
rect -31 19999 -18 20639
rect 28 19999 41 20639
rect 797 20639 869 20683
rect -31 19955 41 19999
rect 797 19999 810 20639
rect 856 19999 869 20639
rect 797 19955 869 19999
rect -31 19883 869 19955
rect 1455 20684 2355 20756
rect 1455 20640 1527 20684
rect 1455 20000 1468 20640
rect 1514 20000 1527 20640
rect 2283 20640 2355 20684
rect 1455 19956 1527 20000
rect 2283 20000 2296 20640
rect 2342 20000 2355 20640
rect 2283 19956 2355 20000
rect 1455 19884 2355 19956
rect 4011 20683 4911 20755
rect 4011 20639 4083 20683
rect 4011 19999 4024 20639
rect 4070 19999 4083 20639
rect 4839 20639 4911 20683
rect 4011 19955 4083 19999
rect 4839 19999 4852 20639
rect 4898 19999 4911 20639
rect 4839 19955 4911 19999
rect 4011 19883 4911 19955
rect 5497 20684 6397 20756
rect 5497 20640 5569 20684
rect 5497 20000 5510 20640
rect 5556 20000 5569 20640
rect 6325 20640 6397 20684
rect 5497 19956 5569 20000
rect 6325 20000 6338 20640
rect 6384 20000 6397 20640
rect 6325 19956 6397 20000
rect 5497 19884 6397 19956
rect 8053 20683 8953 20755
rect 8053 20639 8125 20683
rect 8053 19999 8066 20639
rect 8112 19999 8125 20639
rect 8881 20639 8953 20683
rect 8053 19955 8125 19999
rect 8881 19999 8894 20639
rect 8940 19999 8953 20639
rect 8881 19955 8953 19999
rect 8053 19883 8953 19955
rect 9539 20684 10439 20756
rect 9539 20640 9611 20684
rect 9539 20000 9552 20640
rect 9598 20000 9611 20640
rect 10367 20640 10439 20684
rect 9539 19956 9611 20000
rect 10367 20000 10380 20640
rect 10426 20000 10439 20640
rect 10367 19956 10439 20000
rect 9539 19884 10439 19956
rect 12095 20683 12995 20755
rect 12095 20639 12167 20683
rect 12095 19999 12108 20639
rect 12154 19999 12167 20639
rect 12923 20639 12995 20683
rect 12095 19955 12167 19999
rect 12923 19999 12936 20639
rect 12982 19999 12995 20639
rect 12923 19955 12995 19999
rect 12095 19883 12995 19955
rect 13581 20684 14481 20756
rect 13581 20640 13653 20684
rect 13581 20000 13594 20640
rect 13640 20000 13653 20640
rect 14409 20640 14481 20684
rect 13581 19956 13653 20000
rect 14409 20000 14422 20640
rect 14468 20000 14481 20640
rect 14409 19956 14481 20000
rect 13581 19884 14481 19956
rect 16137 20683 17037 20755
rect 16137 20639 16209 20683
rect 16137 19999 16150 20639
rect 16196 19999 16209 20639
rect 16965 20639 17037 20683
rect 16137 19955 16209 19999
rect 16965 19999 16978 20639
rect 17024 19999 17037 20639
rect 16965 19955 17037 19999
rect 16137 19883 17037 19955
rect 17623 20684 18523 20756
rect 17623 20640 17695 20684
rect 17623 20000 17636 20640
rect 17682 20000 17695 20640
rect 18451 20640 18523 20684
rect 17623 19956 17695 20000
rect 18451 20000 18464 20640
rect 18510 20000 18523 20640
rect 18451 19956 18523 20000
rect 17623 19884 18523 19956
rect -8115 18481 -7215 18553
rect -8115 18437 -8043 18481
rect -8115 17797 -8102 18437
rect -8056 17797 -8043 18437
rect -7287 18437 -7215 18481
rect -8115 17753 -8043 17797
rect -7287 17797 -7274 18437
rect -7228 17797 -7215 18437
rect -7287 17753 -7215 17797
rect -8115 17681 -7215 17753
rect -4073 18478 -3173 18550
rect -4073 18434 -4001 18478
rect -4073 17794 -4060 18434
rect -4014 17794 -4001 18434
rect -3245 18434 -3173 18478
rect -4073 17750 -4001 17794
rect -3245 17794 -3232 18434
rect -3186 17794 -3173 18434
rect -3245 17750 -3173 17794
rect -4073 17678 -3173 17750
rect -31 18478 869 18550
rect -31 18434 41 18478
rect -31 17794 -18 18434
rect 28 17794 41 18434
rect 797 18434 869 18478
rect -31 17750 41 17794
rect 797 17794 810 18434
rect 856 17794 869 18434
rect 797 17750 869 17794
rect -31 17678 869 17750
rect 4011 18478 4911 18550
rect 4011 18434 4083 18478
rect 4011 17794 4024 18434
rect 4070 17794 4083 18434
rect 4839 18434 4911 18478
rect 4011 17750 4083 17794
rect 4839 17794 4852 18434
rect 4898 17794 4911 18434
rect 4839 17750 4911 17794
rect 4011 17678 4911 17750
rect 8053 18478 8953 18550
rect 8053 18434 8125 18478
rect 8053 17794 8066 18434
rect 8112 17794 8125 18434
rect 8881 18434 8953 18478
rect 8053 17750 8125 17794
rect 8881 17794 8894 18434
rect 8940 17794 8953 18434
rect 8881 17750 8953 17794
rect 8053 17678 8953 17750
rect 12095 18478 12995 18550
rect 12095 18434 12167 18478
rect 12095 17794 12108 18434
rect 12154 17794 12167 18434
rect 12923 18434 12995 18478
rect 12095 17750 12167 17794
rect 12923 17794 12936 18434
rect 12982 17794 12995 18434
rect 12923 17750 12995 17794
rect 12095 17678 12995 17750
rect 16137 18478 17037 18550
rect 16137 18434 16209 18478
rect 16137 17794 16150 18434
rect 16196 17794 16209 18434
rect 16965 18434 17037 18478
rect 16137 17750 16209 17794
rect 16965 17794 16978 18434
rect 17024 17794 17037 18434
rect 16965 17750 17037 17794
rect 16137 17678 17037 17750
rect -12127 15517 -11227 15589
rect -12127 15473 -12055 15517
rect -12127 14833 -12114 15473
rect -12068 14833 -12055 15473
rect -11299 15473 -11227 15517
rect -12127 14789 -12055 14833
rect -11299 14833 -11286 15473
rect -11240 14833 -11227 15473
rect -11299 14789 -11227 14833
rect -12127 14717 -11227 14789
rect -8115 15517 -7215 15589
rect -8115 15473 -8043 15517
rect -8115 14833 -8102 15473
rect -8056 14833 -8043 15473
rect -7287 15473 -7215 15517
rect -8115 14789 -8043 14833
rect -7287 14833 -7274 15473
rect -7228 14833 -7215 15473
rect -7287 14789 -7215 14833
rect -8115 14717 -7215 14789
rect -4073 15517 -3173 15589
rect -4073 15473 -4001 15517
rect -4073 14833 -4060 15473
rect -4014 14833 -4001 15473
rect -3245 15473 -3173 15517
rect -4073 14789 -4001 14833
rect -3245 14833 -3232 15473
rect -3186 14833 -3173 15473
rect -3245 14789 -3173 14833
rect -4073 14717 -3173 14789
rect -31 15517 869 15589
rect -31 15473 41 15517
rect -31 14833 -18 15473
rect 28 14833 41 15473
rect 797 15473 869 15517
rect -31 14789 41 14833
rect 797 14833 810 15473
rect 856 14833 869 15473
rect 797 14789 869 14833
rect -31 14717 869 14789
rect 4011 15517 4911 15589
rect 4011 15473 4083 15517
rect 4011 14833 4024 15473
rect 4070 14833 4083 15473
rect 4839 15473 4911 15517
rect 4011 14789 4083 14833
rect 4839 14833 4852 15473
rect 4898 14833 4911 15473
rect 4839 14789 4911 14833
rect 4011 14717 4911 14789
rect 8053 15517 8953 15589
rect 8053 15473 8125 15517
rect 8053 14833 8066 15473
rect 8112 14833 8125 15473
rect 8881 15473 8953 15517
rect 8053 14789 8125 14833
rect 8881 14833 8894 15473
rect 8940 14833 8953 15473
rect 8881 14789 8953 14833
rect 8053 14717 8953 14789
rect 12095 15517 12995 15589
rect 12095 15473 12167 15517
rect 12095 14833 12108 15473
rect 12154 14833 12167 15473
rect 12923 15473 12995 15517
rect 12095 14789 12167 14833
rect 12923 14833 12936 15473
rect 12982 14833 12995 15473
rect 12923 14789 12995 14833
rect 12095 14717 12995 14789
rect -12127 13312 -11227 13384
rect -12127 13268 -12055 13312
rect -12127 12628 -12114 13268
rect -12068 12628 -12055 13268
rect -11299 13268 -11227 13312
rect -12127 12584 -12055 12628
rect -11299 12628 -11286 13268
rect -11240 12628 -11227 13268
rect -11299 12584 -11227 12628
rect -12127 12512 -11227 12584
rect -10641 13312 -9741 13384
rect -10641 13268 -10569 13312
rect -10641 12628 -10628 13268
rect -10582 12628 -10569 13268
rect -9813 13268 -9741 13312
rect -10641 12584 -10569 12628
rect -9813 12628 -9800 13268
rect -9754 12628 -9741 13268
rect -9813 12584 -9741 12628
rect -10641 12512 -9741 12584
rect -8115 13312 -7215 13384
rect -8115 13268 -8043 13312
rect -8115 12628 -8102 13268
rect -8056 12628 -8043 13268
rect -7287 13268 -7215 13312
rect -8115 12584 -8043 12628
rect -7287 12628 -7274 13268
rect -7228 12628 -7215 13268
rect -7287 12584 -7215 12628
rect -8115 12512 -7215 12584
rect -6629 13312 -5729 13384
rect -6629 13268 -6557 13312
rect -6629 12628 -6616 13268
rect -6570 12628 -6557 13268
rect -5801 13268 -5729 13312
rect -6629 12584 -6557 12628
rect -5801 12628 -5788 13268
rect -5742 12628 -5729 13268
rect -5801 12584 -5729 12628
rect -6629 12512 -5729 12584
rect -4073 13312 -3173 13384
rect -4073 13268 -4001 13312
rect -4073 12628 -4060 13268
rect -4014 12628 -4001 13268
rect -3245 13268 -3173 13312
rect -4073 12584 -4001 12628
rect -3245 12628 -3232 13268
rect -3186 12628 -3173 13268
rect -3245 12584 -3173 12628
rect -4073 12512 -3173 12584
rect -2587 13312 -1687 13384
rect -2587 13268 -2515 13312
rect -2587 12628 -2574 13268
rect -2528 12628 -2515 13268
rect -1759 13268 -1687 13312
rect -2587 12584 -2515 12628
rect -1759 12628 -1746 13268
rect -1700 12628 -1687 13268
rect -1759 12584 -1687 12628
rect -2587 12512 -1687 12584
rect -31 13312 869 13384
rect -31 13268 41 13312
rect -31 12628 -18 13268
rect 28 12628 41 13268
rect 797 13268 869 13312
rect -31 12584 41 12628
rect 797 12628 810 13268
rect 856 12628 869 13268
rect 797 12584 869 12628
rect -31 12512 869 12584
rect 1455 13312 2355 13384
rect 1455 13268 1527 13312
rect 1455 12628 1468 13268
rect 1514 12628 1527 13268
rect 2283 13268 2355 13312
rect 1455 12584 1527 12628
rect 2283 12628 2296 13268
rect 2342 12628 2355 13268
rect 2283 12584 2355 12628
rect 1455 12512 2355 12584
rect 4011 13312 4911 13384
rect 4011 13268 4083 13312
rect 4011 12628 4024 13268
rect 4070 12628 4083 13268
rect 4839 13268 4911 13312
rect 4011 12584 4083 12628
rect 4839 12628 4852 13268
rect 4898 12628 4911 13268
rect 4839 12584 4911 12628
rect 4011 12512 4911 12584
rect 5497 13312 6397 13384
rect 5497 13268 5569 13312
rect 5497 12628 5510 13268
rect 5556 12628 5569 13268
rect 6325 13268 6397 13312
rect 5497 12584 5569 12628
rect 6325 12628 6338 13268
rect 6384 12628 6397 13268
rect 6325 12584 6397 12628
rect 5497 12512 6397 12584
rect 8053 13312 8953 13384
rect 8053 13268 8125 13312
rect 8053 12628 8066 13268
rect 8112 12628 8125 13268
rect 8881 13268 8953 13312
rect 8053 12584 8125 12628
rect 8881 12628 8894 13268
rect 8940 12628 8953 13268
rect 8881 12584 8953 12628
rect 8053 12512 8953 12584
rect 9539 13312 10439 13384
rect 9539 13268 9611 13312
rect 9539 12628 9552 13268
rect 9598 12628 9611 13268
rect 10367 13268 10439 13312
rect 9539 12584 9611 12628
rect 10367 12628 10380 13268
rect 10426 12628 10439 13268
rect 10367 12584 10439 12628
rect 9539 12512 10439 12584
rect 12095 13312 12995 13384
rect 12095 13268 12167 13312
rect 12095 12628 12108 13268
rect 12154 12628 12167 13268
rect 12923 13268 12995 13312
rect 12095 12584 12167 12628
rect 12923 12628 12936 13268
rect 12982 12628 12995 13268
rect 12923 12584 12995 12628
rect 12095 12512 12995 12584
rect 13581 13312 14481 13384
rect 13581 13268 13653 13312
rect 13581 12628 13594 13268
rect 13640 12628 13653 13268
rect 14409 13268 14481 13312
rect 13581 12584 13653 12628
rect 14409 12628 14422 13268
rect 14468 12628 14481 13268
rect 14409 12584 14481 12628
rect 13581 12512 14481 12584
rect -12127 11107 -11227 11179
rect -12127 11063 -12055 11107
rect -12127 10423 -12114 11063
rect -12068 10423 -12055 11063
rect -11299 11063 -11227 11107
rect -12127 10379 -12055 10423
rect -11299 10423 -11286 11063
rect -11240 10423 -11227 11063
rect -11299 10379 -11227 10423
rect -12127 10307 -11227 10379
rect -10641 11108 -9741 11180
rect -10641 11064 -10569 11108
rect -10641 10424 -10628 11064
rect -10582 10424 -10569 11064
rect -9813 11064 -9741 11108
rect -10641 10380 -10569 10424
rect -9813 10424 -9800 11064
rect -9754 10424 -9741 11064
rect -9813 10380 -9741 10424
rect -10641 10308 -9741 10380
rect -8115 11107 -7215 11179
rect -8115 11063 -8043 11107
rect -8115 10423 -8102 11063
rect -8056 10423 -8043 11063
rect -7287 11063 -7215 11107
rect -8115 10379 -8043 10423
rect -7287 10423 -7274 11063
rect -7228 10423 -7215 11063
rect -7287 10379 -7215 10423
rect -8115 10307 -7215 10379
rect -6629 11108 -5729 11180
rect -6629 11064 -6557 11108
rect -6629 10424 -6616 11064
rect -6570 10424 -6557 11064
rect -5801 11064 -5729 11108
rect -6629 10380 -6557 10424
rect -5801 10424 -5788 11064
rect -5742 10424 -5729 11064
rect -5801 10380 -5729 10424
rect -6629 10308 -5729 10380
rect -4073 11107 -3173 11179
rect -4073 11063 -4001 11107
rect -4073 10423 -4060 11063
rect -4014 10423 -4001 11063
rect -3245 11063 -3173 11107
rect -4073 10379 -4001 10423
rect -3245 10423 -3232 11063
rect -3186 10423 -3173 11063
rect -3245 10379 -3173 10423
rect -4073 10307 -3173 10379
rect -2587 11108 -1687 11180
rect -2587 11064 -2515 11108
rect -2587 10424 -2574 11064
rect -2528 10424 -2515 11064
rect -1759 11064 -1687 11108
rect -2587 10380 -2515 10424
rect -1759 10424 -1746 11064
rect -1700 10424 -1687 11064
rect -1759 10380 -1687 10424
rect -2587 10308 -1687 10380
rect -31 11107 869 11179
rect -31 11063 41 11107
rect -31 10423 -18 11063
rect 28 10423 41 11063
rect 797 11063 869 11107
rect -31 10379 41 10423
rect 797 10423 810 11063
rect 856 10423 869 11063
rect 797 10379 869 10423
rect -31 10307 869 10379
rect 1455 11108 2355 11180
rect 1455 11064 1527 11108
rect 1455 10424 1468 11064
rect 1514 10424 1527 11064
rect 2283 11064 2355 11108
rect 1455 10380 1527 10424
rect 2283 10424 2296 11064
rect 2342 10424 2355 11064
rect 2283 10380 2355 10424
rect 1455 10308 2355 10380
rect 4011 11107 4911 11179
rect 4011 11063 4083 11107
rect 4011 10423 4024 11063
rect 4070 10423 4083 11063
rect 4839 11063 4911 11107
rect 4011 10379 4083 10423
rect 4839 10423 4852 11063
rect 4898 10423 4911 11063
rect 4839 10379 4911 10423
rect 4011 10307 4911 10379
rect 5497 11108 6397 11180
rect 5497 11064 5569 11108
rect 5497 10424 5510 11064
rect 5556 10424 5569 11064
rect 6325 11064 6397 11108
rect 5497 10380 5569 10424
rect 6325 10424 6338 11064
rect 6384 10424 6397 11064
rect 6325 10380 6397 10424
rect 5497 10308 6397 10380
rect 8053 11107 8953 11179
rect 8053 11063 8125 11107
rect 8053 10423 8066 11063
rect 8112 10423 8125 11063
rect 8881 11063 8953 11107
rect 8053 10379 8125 10423
rect 8881 10423 8894 11063
rect 8940 10423 8953 11063
rect 8881 10379 8953 10423
rect 8053 10307 8953 10379
rect 9539 11108 10439 11180
rect 9539 11064 9611 11108
rect 9539 10424 9552 11064
rect 9598 10424 9611 11064
rect 10367 11064 10439 11108
rect 9539 10380 9611 10424
rect 10367 10424 10380 11064
rect 10426 10424 10439 11064
rect 10367 10380 10439 10424
rect 9539 10308 10439 10380
rect 12095 11107 12995 11179
rect 12095 11063 12167 11107
rect 12095 10423 12108 11063
rect 12154 10423 12167 11063
rect 12923 11063 12995 11107
rect 12095 10379 12167 10423
rect 12923 10423 12936 11063
rect 12982 10423 12995 11063
rect 12923 10379 12995 10423
rect 12095 10307 12995 10379
rect 13581 11108 14481 11180
rect 13581 11064 13653 11108
rect 13581 10424 13594 11064
rect 13640 10424 13653 11064
rect 14409 11064 14481 11108
rect 13581 10380 13653 10424
rect 14409 10424 14422 11064
rect 14468 10424 14481 11064
rect 14409 10380 14481 10424
rect 13581 10308 14481 10380
rect -12127 8902 -11227 8974
rect -12127 8858 -12055 8902
rect -12127 8218 -12114 8858
rect -12068 8218 -12055 8858
rect -11299 8858 -11227 8902
rect -12127 8174 -12055 8218
rect -11299 8218 -11286 8858
rect -11240 8218 -11227 8858
rect -11299 8174 -11227 8218
rect -12127 8102 -11227 8174
rect -8115 8902 -7215 8974
rect -8115 8858 -8043 8902
rect -8115 8218 -8102 8858
rect -8056 8218 -8043 8858
rect -7287 8858 -7215 8902
rect -8115 8174 -8043 8218
rect -7287 8218 -7274 8858
rect -7228 8218 -7215 8858
rect -7287 8174 -7215 8218
rect -8115 8102 -7215 8174
rect -4073 8902 -3173 8974
rect -4073 8858 -4001 8902
rect -4073 8218 -4060 8858
rect -4014 8218 -4001 8858
rect -3245 8858 -3173 8902
rect -4073 8174 -4001 8218
rect -3245 8218 -3232 8858
rect -3186 8218 -3173 8858
rect -3245 8174 -3173 8218
rect -4073 8102 -3173 8174
rect -31 8902 869 8974
rect -31 8858 41 8902
rect -31 8218 -18 8858
rect 28 8218 41 8858
rect 797 8858 869 8902
rect -31 8174 41 8218
rect 797 8218 810 8858
rect 856 8218 869 8858
rect 797 8174 869 8218
rect -31 8102 869 8174
rect 4011 8902 4911 8974
rect 4011 8858 4083 8902
rect 4011 8218 4024 8858
rect 4070 8218 4083 8858
rect 4839 8858 4911 8902
rect 4011 8174 4083 8218
rect 4839 8218 4852 8858
rect 4898 8218 4911 8858
rect 4839 8174 4911 8218
rect 4011 8102 4911 8174
rect 8053 8902 8953 8974
rect 8053 8858 8125 8902
rect 8053 8218 8066 8858
rect 8112 8218 8125 8858
rect 8881 8858 8953 8902
rect 8053 8174 8125 8218
rect 8881 8218 8894 8858
rect 8940 8218 8953 8858
rect 8881 8174 8953 8218
rect 8053 8102 8953 8174
rect 12095 8902 12995 8974
rect 12095 8858 12167 8902
rect 12095 8218 12108 8858
rect 12154 8218 12167 8858
rect 12923 8858 12995 8902
rect 12095 8174 12167 8218
rect 12923 8218 12936 8858
rect 12982 8218 12995 8858
rect 12923 8174 12995 8218
rect 12095 8102 12995 8174
rect -10831 5358 -10681 5380
rect -10831 5312 -10779 5358
rect -10733 5312 -10681 5358
rect -10831 5290 -10681 5312
rect -10591 5358 -10441 5380
rect -10591 5312 -10539 5358
rect -10493 5312 -10441 5358
rect -10591 5290 -10441 5312
rect -10351 5358 -10201 5380
rect -10351 5312 -10299 5358
rect -10253 5312 -10201 5358
rect -10351 5290 -10201 5312
rect -10111 5358 -9961 5380
rect -10111 5312 -10059 5358
rect -10013 5312 -9961 5358
rect -10111 5290 -9961 5312
rect -8657 4981 -7665 5053
rect -8657 4937 -8585 4981
rect -8657 4597 -8644 4937
rect -8598 4597 -8585 4937
rect -8197 4937 -8125 4981
rect -8657 4553 -8585 4597
rect -8197 4597 -8184 4937
rect -8138 4597 -8125 4937
rect -7737 4937 -7665 4981
rect -8197 4553 -8125 4597
rect -7737 4597 -7724 4937
rect -7678 4597 -7665 4937
rect -7737 4553 -7665 4597
rect -9627 4487 -9095 4500
rect -9627 4441 -9511 4487
rect -9211 4441 -9095 4487
rect -8657 4481 -7665 4553
rect -7227 4487 -6695 4500
rect -9627 4428 -9095 4441
rect -9627 3448 -9555 4428
rect -9167 3448 -9095 4428
rect -7227 4441 -7111 4487
rect -6811 4441 -6695 4487
rect -7227 4428 -6695 4441
rect -9627 3376 -9095 3448
rect -7227 3448 -7155 4428
rect -6767 3448 -6695 4428
rect -7227 3376 -6695 3448
rect -9855 1863 -6467 1883
rect -11175 1791 -10643 1863
rect -11175 1747 -11103 1791
rect -11175 1447 -11162 1747
rect -11116 1447 -11103 1747
rect -10715 1747 -10643 1791
rect -11175 1403 -11103 1447
rect -10715 1447 -10702 1747
rect -10656 1447 -10643 1747
rect -10715 1403 -10643 1447
rect -11175 1331 -10643 1403
rect -10315 1811 -6007 1863
rect -10315 1791 -9783 1811
rect -10315 1747 -10243 1791
rect -10315 1447 -10302 1747
rect -10256 1447 -10243 1747
rect -9855 1767 -9783 1791
rect -6539 1791 -6007 1811
rect -10315 1403 -10243 1447
rect -9855 1427 -9842 1767
rect -9796 1427 -9783 1767
rect -6539 1767 -6467 1791
rect -9855 1403 -9783 1427
rect -6539 1427 -6526 1767
rect -6480 1427 -6467 1767
rect -6079 1747 -6007 1791
rect -10315 1383 -9783 1403
rect -6539 1403 -6467 1427
rect -6079 1447 -6066 1747
rect -6020 1447 -6007 1747
rect -6079 1403 -6007 1447
rect -6539 1383 -6007 1403
rect -10315 1331 -6007 1383
rect -5679 1791 -5147 1863
rect -5679 1747 -5607 1791
rect -5679 1447 -5666 1747
rect -5620 1447 -5607 1747
rect -5219 1747 -5147 1791
rect -5679 1403 -5607 1447
rect -5219 1447 -5206 1747
rect -5160 1447 -5147 1747
rect -5219 1403 -5147 1447
rect -5679 1331 -5147 1403
rect -9855 1311 -6467 1331
<< psubdiffcont >>
rect 40103 37895 40149 37941
rect 40343 37895 40389 37941
rect 40583 37895 40629 37941
rect 40823 37895 40869 37941
rect -4844 35854 -4798 36194
rect -4016 35854 -3970 36194
rect 4628 35854 4674 36194
rect 5456 35854 5502 36194
rect 14100 35855 14146 36195
rect 14928 35855 14974 36195
rect 23572 35855 23618 36195
rect 24400 35855 24446 36195
rect 33044 35855 33090 36195
rect 33872 35855 33918 36195
rect 42516 35855 42562 36195
rect 43344 35855 43390 36195
rect -4844 33649 -4798 33989
rect -4016 33649 -3970 33989
rect -3358 33649 -3312 33989
rect -2530 33649 -2484 33989
rect 4628 33649 4674 33989
rect 5456 33649 5502 33989
rect 6114 33649 6160 33989
rect 6942 33649 6988 33989
rect 14100 33650 14146 33990
rect 14928 33650 14974 33990
rect 15586 33650 15632 33990
rect 16414 33650 16460 33990
rect 23572 33650 23618 33990
rect 24400 33650 24446 33990
rect 25058 33650 25104 33990
rect 25886 33650 25932 33990
rect 33044 33650 33090 33990
rect 33872 33650 33918 33990
rect 34530 33650 34576 33990
rect 35358 33650 35404 33990
rect 42516 33650 42562 33990
rect 43344 33650 43390 33990
rect 44002 33650 44048 33990
rect 44830 33650 44876 33990
rect -4844 31444 -4798 31784
rect -4016 31444 -3970 31784
rect -3358 31445 -3312 31785
rect -2530 31445 -2484 31785
rect 4628 31444 4674 31784
rect 5456 31444 5502 31784
rect 6114 31445 6160 31785
rect 6942 31445 6988 31785
rect 14100 31445 14146 31785
rect 14928 31445 14974 31785
rect 15586 31446 15632 31786
rect 16414 31446 16460 31786
rect 23572 31445 23618 31785
rect 24400 31445 24446 31785
rect 25058 31446 25104 31786
rect 25886 31446 25932 31786
rect 33044 31445 33090 31785
rect 33872 31445 33918 31785
rect 34530 31446 34576 31786
rect 35358 31446 35404 31786
rect 42516 31445 42562 31785
rect 43344 31445 43390 31785
rect 44002 31446 44048 31786
rect 44830 31446 44876 31786
rect -9986 30369 -9940 30709
rect -9302 30369 -9256 30709
rect -8618 30369 -8572 30709
rect -8138 30369 -8092 30709
rect -10880 28949 -10834 29289
rect -10400 28949 -10354 29289
rect -7758 29193 -7712 29533
rect -7278 29193 -7232 29533
rect -7074 29193 -7028 29533
rect -6594 29193 -6548 29533
rect -6390 29193 -6344 29533
rect -5910 29193 -5864 29533
rect -4844 29239 -4798 29579
rect -4016 29239 -3970 29579
rect -514 30369 -468 30709
rect 170 30369 216 30709
rect 854 30369 900 30709
rect 1334 30369 1380 30709
rect -1408 28949 -1362 29289
rect -928 28949 -882 29289
rect 1714 29193 1760 29533
rect 2194 29193 2240 29533
rect 2398 29193 2444 29533
rect 2878 29193 2924 29533
rect 3082 29193 3128 29533
rect 3562 29193 3608 29533
rect 4628 29239 4674 29579
rect 5456 29239 5502 29579
rect 8958 30370 9004 30710
rect 9642 30370 9688 30710
rect 10326 30370 10372 30710
rect 10806 30370 10852 30710
rect 8064 28950 8110 29290
rect 8544 28950 8590 29290
rect 11186 29194 11232 29534
rect 11666 29194 11712 29534
rect 11870 29194 11916 29534
rect 12350 29194 12396 29534
rect 12554 29194 12600 29534
rect 13034 29194 13080 29534
rect 14100 29240 14146 29580
rect 14928 29240 14974 29580
rect 18430 30370 18476 30710
rect 19114 30370 19160 30710
rect 19798 30370 19844 30710
rect 20278 30370 20324 30710
rect 17536 28950 17582 29290
rect 18016 28950 18062 29290
rect 20658 29194 20704 29534
rect 21138 29194 21184 29534
rect 21342 29194 21388 29534
rect 21822 29194 21868 29534
rect 22026 29194 22072 29534
rect 22506 29194 22552 29534
rect 23572 29240 23618 29580
rect 24400 29240 24446 29580
rect 27902 30370 27948 30710
rect 28586 30370 28632 30710
rect 29270 30370 29316 30710
rect 29750 30370 29796 30710
rect 27008 28950 27054 29290
rect 27488 28950 27534 29290
rect 30130 29194 30176 29534
rect 30610 29194 30656 29534
rect 30814 29194 30860 29534
rect 31294 29194 31340 29534
rect 31498 29194 31544 29534
rect 31978 29194 32024 29534
rect 33044 29240 33090 29580
rect 33872 29240 33918 29580
rect 37374 30370 37420 30710
rect 38058 30370 38104 30710
rect 38742 30370 38788 30710
rect 39222 30370 39268 30710
rect 36480 28950 36526 29290
rect 36960 28950 37006 29290
rect 39602 29194 39648 29534
rect 40082 29194 40128 29534
rect 40286 29194 40332 29534
rect 40766 29194 40812 29534
rect 40970 29194 41016 29534
rect 41450 29194 41496 29534
rect 42516 29240 42562 29580
rect 43344 29240 43390 29580
rect -9986 28029 -9940 28369
rect -9302 28029 -9256 28369
rect -8618 28029 -8572 28369
rect -8138 28029 -8092 28369
rect -514 28029 -468 28369
rect 170 28029 216 28369
rect 854 28029 900 28369
rect 1334 28029 1380 28369
rect 8958 28030 9004 28370
rect 9642 28030 9688 28370
rect 10326 28030 10372 28370
rect 10806 28030 10852 28370
rect 18430 28030 18476 28370
rect 19114 28030 19160 28370
rect 19798 28030 19844 28370
rect 20278 28030 20324 28370
rect 27902 28030 27948 28370
rect 28586 28030 28632 28370
rect 29270 28030 29316 28370
rect 29750 28030 29796 28370
rect 37374 28030 37420 28370
rect 38058 28030 38104 28370
rect 38742 28030 38788 28370
rect 39222 28030 39268 28370
rect -12593 27019 -12547 27359
rect -12113 27019 -12067 27359
rect -8102 23552 -8056 23892
rect -7274 23552 -7228 23892
rect -4060 23549 -4014 23889
rect -3232 23549 -3186 23889
rect -18 23549 28 23889
rect 810 23549 856 23889
rect 4024 23549 4070 23889
rect 4852 23549 4898 23889
rect 8066 23549 8112 23889
rect 8894 23549 8940 23889
rect 12108 23549 12154 23889
rect 12936 23549 12982 23889
rect 16150 23549 16196 23889
rect 16978 23549 17024 23889
rect -8102 21347 -8056 21687
rect -7274 21347 -7228 21687
rect -6616 21347 -6570 21687
rect -5788 21347 -5742 21687
rect -4060 21344 -4014 21684
rect -3232 21344 -3186 21684
rect -2574 21344 -2528 21684
rect -1746 21344 -1700 21684
rect -18 21344 28 21684
rect 810 21344 856 21684
rect 1468 21344 1514 21684
rect 2296 21344 2342 21684
rect 4024 21344 4070 21684
rect 4852 21344 4898 21684
rect 5510 21344 5556 21684
rect 6338 21344 6384 21684
rect 8066 21344 8112 21684
rect 8894 21344 8940 21684
rect 9552 21344 9598 21684
rect 10380 21344 10426 21684
rect 12108 21344 12154 21684
rect 12936 21344 12982 21684
rect 13594 21344 13640 21684
rect 14422 21344 14468 21684
rect 16150 21344 16196 21684
rect 16978 21344 17024 21684
rect 17636 21344 17682 21684
rect 18464 21344 18510 21684
rect -8102 19142 -8056 19482
rect -7274 19142 -7228 19482
rect -6616 19143 -6570 19483
rect -5788 19143 -5742 19483
rect -4060 19139 -4014 19479
rect -3232 19139 -3186 19479
rect -2574 19140 -2528 19480
rect -1746 19140 -1700 19480
rect -18 19139 28 19479
rect 810 19139 856 19479
rect 1468 19140 1514 19480
rect 2296 19140 2342 19480
rect 4024 19139 4070 19479
rect 4852 19139 4898 19479
rect 5510 19140 5556 19480
rect 6338 19140 6384 19480
rect 8066 19139 8112 19479
rect 8894 19139 8940 19479
rect 9552 19140 9598 19480
rect 10380 19140 10426 19480
rect 12108 19139 12154 19479
rect 12936 19139 12982 19479
rect 13594 19140 13640 19480
rect 14422 19140 14468 19480
rect 16150 19139 16196 19479
rect 16978 19139 17024 19479
rect 17636 19140 17682 19480
rect 18464 19140 18510 19480
rect -8102 16937 -8056 17277
rect -7274 16937 -7228 17277
rect -4060 16934 -4014 17274
rect -3232 16934 -3186 17274
rect -18 16934 28 17274
rect 810 16934 856 17274
rect 4024 16934 4070 17274
rect 4852 16934 4898 17274
rect 8066 16934 8112 17274
rect 8894 16934 8940 17274
rect 12108 16934 12154 17274
rect 12936 16934 12982 17274
rect 16150 16934 16196 17274
rect 16978 16934 17024 17274
rect -12114 13973 -12068 14313
rect -11286 13973 -11240 14313
rect -8102 13973 -8056 14313
rect -7274 13973 -7228 14313
rect -4060 13973 -4014 14313
rect -3232 13973 -3186 14313
rect -18 13973 28 14313
rect 810 13973 856 14313
rect 4024 13973 4070 14313
rect 4852 13973 4898 14313
rect 8066 13973 8112 14313
rect 8894 13973 8940 14313
rect 12108 13973 12154 14313
rect 12936 13973 12982 14313
rect -12114 11768 -12068 12108
rect -11286 11768 -11240 12108
rect -10628 11768 -10582 12108
rect -9800 11768 -9754 12108
rect -8102 11768 -8056 12108
rect -7274 11768 -7228 12108
rect -6616 11768 -6570 12108
rect -5788 11768 -5742 12108
rect -4060 11768 -4014 12108
rect -3232 11768 -3186 12108
rect -2574 11768 -2528 12108
rect -1746 11768 -1700 12108
rect -18 11768 28 12108
rect 810 11768 856 12108
rect 1468 11768 1514 12108
rect 2296 11768 2342 12108
rect 4024 11768 4070 12108
rect 4852 11768 4898 12108
rect 5510 11768 5556 12108
rect 6338 11768 6384 12108
rect 8066 11768 8112 12108
rect 8894 11768 8940 12108
rect 9552 11768 9598 12108
rect 10380 11768 10426 12108
rect 12108 11768 12154 12108
rect 12936 11768 12982 12108
rect 13594 11768 13640 12108
rect 14422 11768 14468 12108
rect -12114 9563 -12068 9903
rect -11286 9563 -11240 9903
rect -10628 9564 -10582 9904
rect -9800 9564 -9754 9904
rect -8102 9563 -8056 9903
rect -7274 9563 -7228 9903
rect -6616 9564 -6570 9904
rect -5788 9564 -5742 9904
rect -4060 9563 -4014 9903
rect -3232 9563 -3186 9903
rect -2574 9564 -2528 9904
rect -1746 9564 -1700 9904
rect -18 9563 28 9903
rect 810 9563 856 9903
rect 1468 9564 1514 9904
rect 2296 9564 2342 9904
rect 4024 9563 4070 9903
rect 4852 9563 4898 9903
rect 5510 9564 5556 9904
rect 6338 9564 6384 9904
rect 8066 9563 8112 9903
rect 8894 9563 8940 9903
rect 9552 9564 9598 9904
rect 10380 9564 10426 9904
rect 12108 9563 12154 9903
rect 12936 9563 12982 9903
rect 13594 9564 13640 9904
rect 14422 9564 14468 9904
rect -12114 7358 -12068 7698
rect -11286 7358 -11240 7698
rect -8102 7358 -8056 7698
rect -7274 7358 -7228 7698
rect -4060 7358 -4014 7698
rect -3232 7358 -3186 7698
rect -18 7358 28 7698
rect 810 7358 856 7698
rect 4024 7358 4070 7698
rect 4852 7358 4898 7698
rect 8066 7358 8112 7698
rect 8894 7358 8940 7698
rect 12108 7358 12154 7698
rect 12936 7358 12982 7698
rect -10779 4232 -10733 4278
rect -10539 4232 -10493 4278
rect -10299 4232 -10253 4278
rect -10059 4232 -10013 4278
rect -8644 3777 -8598 4117
rect -8184 3777 -8138 4117
rect -7724 3777 -7678 4117
rect -9511 2589 -9211 2635
rect -7111 2589 -6811 2635
rect -9980 271 -9934 811
rect -8184 271 -8138 811
rect -6388 271 -6342 811
rect -10304 -903 -10204 -403
rect -6118 -903 -6018 -403
rect -10304 -2348 -10204 -1848
rect -6118 -2348 -6018 -1848
rect -8598 -2863 -8552 -2563
rect -7770 -2863 -7724 -2563
<< nsubdiffcont >>
rect 40103 38975 40149 39021
rect 40343 38975 40389 39021
rect 40583 38975 40629 39021
rect 40823 38975 40869 39021
rect -4844 36714 -4798 37354
rect -4016 36714 -3970 37354
rect 4628 36714 4674 37354
rect 5456 36714 5502 37354
rect 14100 36715 14146 37355
rect 14928 36715 14974 37355
rect 23572 36715 23618 37355
rect 24400 36715 24446 37355
rect 33044 36715 33090 37355
rect 33872 36715 33918 37355
rect 42516 36715 42562 37355
rect 43344 36715 43390 37355
rect -4844 34509 -4798 35149
rect -4016 34509 -3970 35149
rect -3358 34509 -3312 35149
rect -2530 34509 -2484 35149
rect 4628 34509 4674 35149
rect 5456 34509 5502 35149
rect 6114 34509 6160 35149
rect 6942 34509 6988 35149
rect 14100 34510 14146 35150
rect 14928 34510 14974 35150
rect 15586 34510 15632 35150
rect 16414 34510 16460 35150
rect 23572 34510 23618 35150
rect 24400 34510 24446 35150
rect 25058 34510 25104 35150
rect 25886 34510 25932 35150
rect 33044 34510 33090 35150
rect 33872 34510 33918 35150
rect 34530 34510 34576 35150
rect 35358 34510 35404 35150
rect 42516 34510 42562 35150
rect 43344 34510 43390 35150
rect 44002 34510 44048 35150
rect 44830 34510 44876 35150
rect -4844 32304 -4798 32944
rect -4016 32304 -3970 32944
rect -3358 32305 -3312 32945
rect -2530 32305 -2484 32945
rect 4628 32304 4674 32944
rect 5456 32304 5502 32944
rect 6114 32305 6160 32945
rect 6942 32305 6988 32945
rect 14100 32305 14146 32945
rect 14928 32305 14974 32945
rect 15586 32306 15632 32946
rect 16414 32306 16460 32946
rect 23572 32305 23618 32945
rect 24400 32305 24446 32945
rect 25058 32306 25104 32946
rect 25886 32306 25932 32946
rect 33044 32305 33090 32945
rect 33872 32305 33918 32945
rect 34530 32306 34576 32946
rect 35358 32306 35404 32946
rect 42516 32305 42562 32945
rect 43344 32305 43390 32945
rect 44002 32306 44048 32946
rect 44830 32306 44876 32946
rect -9986 31089 -9940 31829
rect -9506 31089 -9460 31829
rect -9098 31089 -9052 31829
rect -8618 31089 -8572 31829
rect -8138 31089 -8092 31829
rect -514 31089 -468 31829
rect -34 31089 12 31829
rect 374 31089 420 31829
rect 854 31089 900 31829
rect 1334 31089 1380 31829
rect 8958 31090 9004 31830
rect 9438 31090 9484 31830
rect 9846 31090 9892 31830
rect 10326 31090 10372 31830
rect 10806 31090 10852 31830
rect 18430 31090 18476 31830
rect 18910 31090 18956 31830
rect 19318 31090 19364 31830
rect 19798 31090 19844 31830
rect 20278 31090 20324 31830
rect 27902 31090 27948 31830
rect 28382 31090 28428 31830
rect 28790 31090 28836 31830
rect 29270 31090 29316 31830
rect 29750 31090 29796 31830
rect 37374 31090 37420 31830
rect 37854 31090 37900 31830
rect 38262 31090 38308 31830
rect 38742 31090 38788 31830
rect 39222 31090 39268 31830
rect -10880 29669 -10834 30409
rect -10400 29669 -10354 30409
rect -7758 29913 -7712 30653
rect -7074 29913 -7028 30653
rect -6390 29913 -6344 30653
rect -5910 29913 -5864 30653
rect -4844 30099 -4798 30739
rect -4016 30099 -3970 30739
rect -9986 28749 -9940 29489
rect -9506 28749 -9460 29489
rect -9098 28749 -9052 29489
rect -8618 28749 -8572 29489
rect -8138 28749 -8092 29489
rect -1408 29669 -1362 30409
rect -928 29669 -882 30409
rect 1714 29913 1760 30653
rect 2398 29913 2444 30653
rect 3082 29913 3128 30653
rect 3562 29913 3608 30653
rect 4628 30099 4674 30739
rect 5456 30099 5502 30739
rect -514 28749 -468 29489
rect -34 28749 12 29489
rect 374 28749 420 29489
rect 854 28749 900 29489
rect 1334 28749 1380 29489
rect 8064 29670 8110 30410
rect 8544 29670 8590 30410
rect 11186 29914 11232 30654
rect 11870 29914 11916 30654
rect 12554 29914 12600 30654
rect 13034 29914 13080 30654
rect 14100 30100 14146 30740
rect 14928 30100 14974 30740
rect 8958 28750 9004 29490
rect 9438 28750 9484 29490
rect 9846 28750 9892 29490
rect 10326 28750 10372 29490
rect 10806 28750 10852 29490
rect 17536 29670 17582 30410
rect 18016 29670 18062 30410
rect 20658 29914 20704 30654
rect 21342 29914 21388 30654
rect 22026 29914 22072 30654
rect 22506 29914 22552 30654
rect 23572 30100 23618 30740
rect 24400 30100 24446 30740
rect 18430 28750 18476 29490
rect 18910 28750 18956 29490
rect 19318 28750 19364 29490
rect 19798 28750 19844 29490
rect 20278 28750 20324 29490
rect 27008 29670 27054 30410
rect 27488 29670 27534 30410
rect 30130 29914 30176 30654
rect 30814 29914 30860 30654
rect 31498 29914 31544 30654
rect 31978 29914 32024 30654
rect 33044 30100 33090 30740
rect 33872 30100 33918 30740
rect 27902 28750 27948 29490
rect 28382 28750 28428 29490
rect 28790 28750 28836 29490
rect 29270 28750 29316 29490
rect 29750 28750 29796 29490
rect 36480 29670 36526 30410
rect 36960 29670 37006 30410
rect 39602 29914 39648 30654
rect 40286 29914 40332 30654
rect 40970 29914 41016 30654
rect 41450 29914 41496 30654
rect 42516 30100 42562 30740
rect 43344 30100 43390 30740
rect 37374 28750 37420 29490
rect 37854 28750 37900 29490
rect 38262 28750 38308 29490
rect 38742 28750 38788 29490
rect 39222 28750 39268 29490
rect -12593 27739 -12547 28479
rect -12113 27739 -12067 28479
rect -8102 24412 -8056 25052
rect -7274 24412 -7228 25052
rect -4060 24409 -4014 25049
rect -3232 24409 -3186 25049
rect -18 24409 28 25049
rect 810 24409 856 25049
rect 4024 24409 4070 25049
rect 4852 24409 4898 25049
rect 8066 24409 8112 25049
rect 8894 24409 8940 25049
rect 12108 24409 12154 25049
rect 12936 24409 12982 25049
rect 16150 24409 16196 25049
rect 16978 24409 17024 25049
rect -8102 22207 -8056 22847
rect -7274 22207 -7228 22847
rect -6616 22207 -6570 22847
rect -5788 22207 -5742 22847
rect -4060 22204 -4014 22844
rect -3232 22204 -3186 22844
rect -2574 22204 -2528 22844
rect -1746 22204 -1700 22844
rect -18 22204 28 22844
rect 810 22204 856 22844
rect 1468 22204 1514 22844
rect 2296 22204 2342 22844
rect 4024 22204 4070 22844
rect 4852 22204 4898 22844
rect 5510 22204 5556 22844
rect 6338 22204 6384 22844
rect 8066 22204 8112 22844
rect 8894 22204 8940 22844
rect 9552 22204 9598 22844
rect 10380 22204 10426 22844
rect 12108 22204 12154 22844
rect 12936 22204 12982 22844
rect 13594 22204 13640 22844
rect 14422 22204 14468 22844
rect 16150 22204 16196 22844
rect 16978 22204 17024 22844
rect 17636 22204 17682 22844
rect 18464 22204 18510 22844
rect -8102 20002 -8056 20642
rect -7274 20002 -7228 20642
rect -6616 20003 -6570 20643
rect -5788 20003 -5742 20643
rect -4060 19999 -4014 20639
rect -3232 19999 -3186 20639
rect -2574 20000 -2528 20640
rect -1746 20000 -1700 20640
rect -18 19999 28 20639
rect 810 19999 856 20639
rect 1468 20000 1514 20640
rect 2296 20000 2342 20640
rect 4024 19999 4070 20639
rect 4852 19999 4898 20639
rect 5510 20000 5556 20640
rect 6338 20000 6384 20640
rect 8066 19999 8112 20639
rect 8894 19999 8940 20639
rect 9552 20000 9598 20640
rect 10380 20000 10426 20640
rect 12108 19999 12154 20639
rect 12936 19999 12982 20639
rect 13594 20000 13640 20640
rect 14422 20000 14468 20640
rect 16150 19999 16196 20639
rect 16978 19999 17024 20639
rect 17636 20000 17682 20640
rect 18464 20000 18510 20640
rect -8102 17797 -8056 18437
rect -7274 17797 -7228 18437
rect -4060 17794 -4014 18434
rect -3232 17794 -3186 18434
rect -18 17794 28 18434
rect 810 17794 856 18434
rect 4024 17794 4070 18434
rect 4852 17794 4898 18434
rect 8066 17794 8112 18434
rect 8894 17794 8940 18434
rect 12108 17794 12154 18434
rect 12936 17794 12982 18434
rect 16150 17794 16196 18434
rect 16978 17794 17024 18434
rect -12114 14833 -12068 15473
rect -11286 14833 -11240 15473
rect -8102 14833 -8056 15473
rect -7274 14833 -7228 15473
rect -4060 14833 -4014 15473
rect -3232 14833 -3186 15473
rect -18 14833 28 15473
rect 810 14833 856 15473
rect 4024 14833 4070 15473
rect 4852 14833 4898 15473
rect 8066 14833 8112 15473
rect 8894 14833 8940 15473
rect 12108 14833 12154 15473
rect 12936 14833 12982 15473
rect -12114 12628 -12068 13268
rect -11286 12628 -11240 13268
rect -10628 12628 -10582 13268
rect -9800 12628 -9754 13268
rect -8102 12628 -8056 13268
rect -7274 12628 -7228 13268
rect -6616 12628 -6570 13268
rect -5788 12628 -5742 13268
rect -4060 12628 -4014 13268
rect -3232 12628 -3186 13268
rect -2574 12628 -2528 13268
rect -1746 12628 -1700 13268
rect -18 12628 28 13268
rect 810 12628 856 13268
rect 1468 12628 1514 13268
rect 2296 12628 2342 13268
rect 4024 12628 4070 13268
rect 4852 12628 4898 13268
rect 5510 12628 5556 13268
rect 6338 12628 6384 13268
rect 8066 12628 8112 13268
rect 8894 12628 8940 13268
rect 9552 12628 9598 13268
rect 10380 12628 10426 13268
rect 12108 12628 12154 13268
rect 12936 12628 12982 13268
rect 13594 12628 13640 13268
rect 14422 12628 14468 13268
rect -12114 10423 -12068 11063
rect -11286 10423 -11240 11063
rect -10628 10424 -10582 11064
rect -9800 10424 -9754 11064
rect -8102 10423 -8056 11063
rect -7274 10423 -7228 11063
rect -6616 10424 -6570 11064
rect -5788 10424 -5742 11064
rect -4060 10423 -4014 11063
rect -3232 10423 -3186 11063
rect -2574 10424 -2528 11064
rect -1746 10424 -1700 11064
rect -18 10423 28 11063
rect 810 10423 856 11063
rect 1468 10424 1514 11064
rect 2296 10424 2342 11064
rect 4024 10423 4070 11063
rect 4852 10423 4898 11063
rect 5510 10424 5556 11064
rect 6338 10424 6384 11064
rect 8066 10423 8112 11063
rect 8894 10423 8940 11063
rect 9552 10424 9598 11064
rect 10380 10424 10426 11064
rect 12108 10423 12154 11063
rect 12936 10423 12982 11063
rect 13594 10424 13640 11064
rect 14422 10424 14468 11064
rect -12114 8218 -12068 8858
rect -11286 8218 -11240 8858
rect -8102 8218 -8056 8858
rect -7274 8218 -7228 8858
rect -4060 8218 -4014 8858
rect -3232 8218 -3186 8858
rect -18 8218 28 8858
rect 810 8218 856 8858
rect 4024 8218 4070 8858
rect 4852 8218 4898 8858
rect 8066 8218 8112 8858
rect 8894 8218 8940 8858
rect 12108 8218 12154 8858
rect 12936 8218 12982 8858
rect -10779 5312 -10733 5358
rect -10539 5312 -10493 5358
rect -10299 5312 -10253 5358
rect -10059 5312 -10013 5358
rect -8644 4597 -8598 4937
rect -8184 4597 -8138 4937
rect -7724 4597 -7678 4937
rect -9511 4441 -9211 4487
rect -7111 4441 -6811 4487
rect -11162 1447 -11116 1747
rect -10702 1447 -10656 1747
rect -10302 1447 -10256 1747
rect -9842 1427 -9796 1767
rect -6526 1427 -6480 1767
rect -6066 1447 -6020 1747
rect -5666 1447 -5620 1747
rect -5206 1447 -5160 1747
<< polysilicon >>
rect 40051 38883 40111 38933
rect 40221 38883 40281 38933
rect 40391 38883 40451 38933
rect 40561 38883 40621 38933
rect 40731 38883 40791 38933
rect 40051 38523 40111 38543
rect 40221 38523 40281 38543
rect 40391 38523 40451 38543
rect 40561 38523 40621 38543
rect 40051 38513 40621 38523
rect 40051 38486 40681 38513
rect 40051 38463 40608 38486
rect 40221 38283 40281 38463
rect 40561 38440 40608 38463
rect 40654 38440 40681 38486
rect 40561 38413 40681 38440
rect 40561 38283 40621 38413
rect 40731 38363 40791 38543
rect 40051 38223 40621 38283
rect 40671 38336 40791 38363
rect 40671 38290 40698 38336
rect 40744 38290 40791 38336
rect 40671 38263 40791 38290
rect 40051 38203 40111 38223
rect 40221 38203 40281 38223
rect 40391 38203 40451 38223
rect 40561 38203 40621 38223
rect 40731 38203 40791 38263
rect 40051 37983 40111 38033
rect 40221 37983 40281 38033
rect 40391 37983 40451 38033
rect 40561 37983 40621 38033
rect 40731 37983 40791 38033
rect -4631 37363 -4551 37376
rect -4631 37317 -4618 37363
rect -4564 37317 -4551 37363
rect -4631 37284 -4551 37317
rect -4447 37363 -4367 37376
rect -4447 37317 -4434 37363
rect -4380 37317 -4367 37363
rect -4447 37284 -4367 37317
rect -4263 37363 -4183 37376
rect -4263 37317 -4250 37363
rect -4196 37317 -4183 37363
rect -4263 37284 -4183 37317
rect -4631 36751 -4551 36784
rect -4631 36705 -4618 36751
rect -4564 36705 -4551 36751
rect -4631 36692 -4551 36705
rect -4447 36751 -4367 36784
rect -4447 36705 -4434 36751
rect -4380 36705 -4367 36751
rect -4447 36692 -4367 36705
rect -4263 36751 -4183 36784
rect -4263 36705 -4250 36751
rect -4196 36705 -4183 36751
rect -4263 36692 -4183 36705
rect 4841 37363 4921 37376
rect 4841 37317 4854 37363
rect 4908 37317 4921 37363
rect 4841 37284 4921 37317
rect 5025 37363 5105 37376
rect 5025 37317 5038 37363
rect 5092 37317 5105 37363
rect 5025 37284 5105 37317
rect 5209 37363 5289 37376
rect 5209 37317 5222 37363
rect 5276 37317 5289 37363
rect 5209 37284 5289 37317
rect 4841 36751 4921 36784
rect 4841 36705 4854 36751
rect 4908 36705 4921 36751
rect 4841 36692 4921 36705
rect 5025 36751 5105 36784
rect 5025 36705 5038 36751
rect 5092 36705 5105 36751
rect 5025 36692 5105 36705
rect 5209 36751 5289 36784
rect 5209 36705 5222 36751
rect 5276 36705 5289 36751
rect 5209 36692 5289 36705
rect 14313 37364 14393 37377
rect 14313 37318 14326 37364
rect 14380 37318 14393 37364
rect 14313 37285 14393 37318
rect 14497 37364 14577 37377
rect 14497 37318 14510 37364
rect 14564 37318 14577 37364
rect 14497 37285 14577 37318
rect 14681 37364 14761 37377
rect 14681 37318 14694 37364
rect 14748 37318 14761 37364
rect 14681 37285 14761 37318
rect 14313 36752 14393 36785
rect 14313 36706 14326 36752
rect 14380 36706 14393 36752
rect 14313 36693 14393 36706
rect 14497 36752 14577 36785
rect 14497 36706 14510 36752
rect 14564 36706 14577 36752
rect 14497 36693 14577 36706
rect 14681 36752 14761 36785
rect 14681 36706 14694 36752
rect 14748 36706 14761 36752
rect 14681 36693 14761 36706
rect 23785 37364 23865 37377
rect 23785 37318 23798 37364
rect 23852 37318 23865 37364
rect 23785 37285 23865 37318
rect 23969 37364 24049 37377
rect 23969 37318 23982 37364
rect 24036 37318 24049 37364
rect 23969 37285 24049 37318
rect 24153 37364 24233 37377
rect 24153 37318 24166 37364
rect 24220 37318 24233 37364
rect 24153 37285 24233 37318
rect 23785 36752 23865 36785
rect 23785 36706 23798 36752
rect 23852 36706 23865 36752
rect 23785 36693 23865 36706
rect 23969 36752 24049 36785
rect 23969 36706 23982 36752
rect 24036 36706 24049 36752
rect 23969 36693 24049 36706
rect 24153 36752 24233 36785
rect 24153 36706 24166 36752
rect 24220 36706 24233 36752
rect 24153 36693 24233 36706
rect 33257 37364 33337 37377
rect 33257 37318 33270 37364
rect 33324 37318 33337 37364
rect 33257 37285 33337 37318
rect 33441 37364 33521 37377
rect 33441 37318 33454 37364
rect 33508 37318 33521 37364
rect 33441 37285 33521 37318
rect 33625 37364 33705 37377
rect 33625 37318 33638 37364
rect 33692 37318 33705 37364
rect 33625 37285 33705 37318
rect 33257 36752 33337 36785
rect 33257 36706 33270 36752
rect 33324 36706 33337 36752
rect 33257 36693 33337 36706
rect 33441 36752 33521 36785
rect 33441 36706 33454 36752
rect 33508 36706 33521 36752
rect 33441 36693 33521 36706
rect 33625 36752 33705 36785
rect 33625 36706 33638 36752
rect 33692 36706 33705 36752
rect 33625 36693 33705 36706
rect 42729 37364 42809 37377
rect 42729 37318 42742 37364
rect 42796 37318 42809 37364
rect 42729 37285 42809 37318
rect 42913 37364 42993 37377
rect 42913 37318 42926 37364
rect 42980 37318 42993 37364
rect 42913 37285 42993 37318
rect 43097 37364 43177 37377
rect 43097 37318 43110 37364
rect 43164 37318 43177 37364
rect 43097 37285 43177 37318
rect 42729 36752 42809 36785
rect 42729 36706 42742 36752
rect 42796 36706 42809 36752
rect 42729 36693 42809 36706
rect 42913 36752 42993 36785
rect 42913 36706 42926 36752
rect 42980 36706 42993 36752
rect 42913 36693 42993 36706
rect 43097 36752 43177 36785
rect 43097 36706 43110 36752
rect 43164 36706 43177 36752
rect 43097 36693 43177 36706
rect -4631 36203 -4551 36216
rect -4631 36157 -4618 36203
rect -4564 36157 -4551 36203
rect -4631 36124 -4551 36157
rect -4447 36203 -4367 36216
rect -4447 36157 -4434 36203
rect -4380 36157 -4367 36203
rect -4447 36124 -4367 36157
rect -4263 36203 -4183 36216
rect -4263 36157 -4250 36203
rect -4196 36157 -4183 36203
rect -4263 36124 -4183 36157
rect -4631 35891 -4551 35924
rect -4631 35845 -4618 35891
rect -4564 35845 -4551 35891
rect -4631 35832 -4551 35845
rect -4447 35891 -4367 35924
rect -4447 35845 -4434 35891
rect -4380 35845 -4367 35891
rect -4447 35832 -4367 35845
rect -4263 35891 -4183 35924
rect -4263 35845 -4250 35891
rect -4196 35845 -4183 35891
rect -4263 35832 -4183 35845
rect 4841 36203 4921 36216
rect 4841 36157 4854 36203
rect 4908 36157 4921 36203
rect 4841 36124 4921 36157
rect 5025 36203 5105 36216
rect 5025 36157 5038 36203
rect 5092 36157 5105 36203
rect 5025 36124 5105 36157
rect 5209 36203 5289 36216
rect 5209 36157 5222 36203
rect 5276 36157 5289 36203
rect 5209 36124 5289 36157
rect 4841 35891 4921 35924
rect 4841 35845 4854 35891
rect 4908 35845 4921 35891
rect 4841 35832 4921 35845
rect 5025 35891 5105 35924
rect 5025 35845 5038 35891
rect 5092 35845 5105 35891
rect 5025 35832 5105 35845
rect 5209 35891 5289 35924
rect 5209 35845 5222 35891
rect 5276 35845 5289 35891
rect 5209 35832 5289 35845
rect 14313 36204 14393 36217
rect 14313 36158 14326 36204
rect 14380 36158 14393 36204
rect 14313 36125 14393 36158
rect 14497 36204 14577 36217
rect 14497 36158 14510 36204
rect 14564 36158 14577 36204
rect 14497 36125 14577 36158
rect 14681 36204 14761 36217
rect 14681 36158 14694 36204
rect 14748 36158 14761 36204
rect 14681 36125 14761 36158
rect 14313 35892 14393 35925
rect 14313 35846 14326 35892
rect 14380 35846 14393 35892
rect 14313 35833 14393 35846
rect 14497 35892 14577 35925
rect 14497 35846 14510 35892
rect 14564 35846 14577 35892
rect 14497 35833 14577 35846
rect 14681 35892 14761 35925
rect 14681 35846 14694 35892
rect 14748 35846 14761 35892
rect 14681 35833 14761 35846
rect 23785 36204 23865 36217
rect 23785 36158 23798 36204
rect 23852 36158 23865 36204
rect 23785 36125 23865 36158
rect 23969 36204 24049 36217
rect 23969 36158 23982 36204
rect 24036 36158 24049 36204
rect 23969 36125 24049 36158
rect 24153 36204 24233 36217
rect 24153 36158 24166 36204
rect 24220 36158 24233 36204
rect 24153 36125 24233 36158
rect 23785 35892 23865 35925
rect 23785 35846 23798 35892
rect 23852 35846 23865 35892
rect 23785 35833 23865 35846
rect 23969 35892 24049 35925
rect 23969 35846 23982 35892
rect 24036 35846 24049 35892
rect 23969 35833 24049 35846
rect 24153 35892 24233 35925
rect 24153 35846 24166 35892
rect 24220 35846 24233 35892
rect 24153 35833 24233 35846
rect 33257 36204 33337 36217
rect 33257 36158 33270 36204
rect 33324 36158 33337 36204
rect 33257 36125 33337 36158
rect 33441 36204 33521 36217
rect 33441 36158 33454 36204
rect 33508 36158 33521 36204
rect 33441 36125 33521 36158
rect 33625 36204 33705 36217
rect 33625 36158 33638 36204
rect 33692 36158 33705 36204
rect 33625 36125 33705 36158
rect 33257 35892 33337 35925
rect 33257 35846 33270 35892
rect 33324 35846 33337 35892
rect 33257 35833 33337 35846
rect 33441 35892 33521 35925
rect 33441 35846 33454 35892
rect 33508 35846 33521 35892
rect 33441 35833 33521 35846
rect 33625 35892 33705 35925
rect 33625 35846 33638 35892
rect 33692 35846 33705 35892
rect 33625 35833 33705 35846
rect 42729 36204 42809 36217
rect 42729 36158 42742 36204
rect 42796 36158 42809 36204
rect 42729 36125 42809 36158
rect 42913 36204 42993 36217
rect 42913 36158 42926 36204
rect 42980 36158 42993 36204
rect 42913 36125 42993 36158
rect 43097 36204 43177 36217
rect 43097 36158 43110 36204
rect 43164 36158 43177 36204
rect 43097 36125 43177 36158
rect 42729 35892 42809 35925
rect 42729 35846 42742 35892
rect 42796 35846 42809 35892
rect 42729 35833 42809 35846
rect 42913 35892 42993 35925
rect 42913 35846 42926 35892
rect 42980 35846 42993 35892
rect 42913 35833 42993 35846
rect 43097 35892 43177 35925
rect 43097 35846 43110 35892
rect 43164 35846 43177 35892
rect 43097 35833 43177 35846
rect -4631 35158 -4551 35171
rect -4631 35112 -4618 35158
rect -4564 35112 -4551 35158
rect -4631 35079 -4551 35112
rect -4447 35158 -4367 35171
rect -4447 35112 -4434 35158
rect -4380 35112 -4367 35158
rect -4447 35079 -4367 35112
rect -4263 35158 -4183 35171
rect -4263 35112 -4250 35158
rect -4196 35112 -4183 35158
rect -4263 35079 -4183 35112
rect -4631 34546 -4551 34579
rect -4631 34500 -4618 34546
rect -4564 34500 -4551 34546
rect -4631 34487 -4551 34500
rect -4447 34546 -4367 34579
rect -4447 34500 -4434 34546
rect -4380 34500 -4367 34546
rect -4447 34487 -4367 34500
rect -4263 34546 -4183 34579
rect -4263 34500 -4250 34546
rect -4196 34500 -4183 34546
rect -4263 34487 -4183 34500
rect -3145 35158 -3065 35171
rect -3145 35112 -3132 35158
rect -3078 35112 -3065 35158
rect -3145 35079 -3065 35112
rect -2961 35158 -2881 35171
rect -2961 35112 -2948 35158
rect -2894 35112 -2881 35158
rect -2961 35079 -2881 35112
rect -2777 35158 -2697 35171
rect -2777 35112 -2764 35158
rect -2710 35112 -2697 35158
rect -2777 35079 -2697 35112
rect -3145 34546 -3065 34579
rect -3145 34500 -3132 34546
rect -3078 34500 -3065 34546
rect -3145 34487 -3065 34500
rect -2961 34546 -2881 34579
rect -2961 34500 -2948 34546
rect -2894 34500 -2881 34546
rect -2961 34487 -2881 34500
rect -2777 34546 -2697 34579
rect -2777 34500 -2764 34546
rect -2710 34500 -2697 34546
rect -2777 34487 -2697 34500
rect 4841 35158 4921 35171
rect 4841 35112 4854 35158
rect 4908 35112 4921 35158
rect 4841 35079 4921 35112
rect 5025 35158 5105 35171
rect 5025 35112 5038 35158
rect 5092 35112 5105 35158
rect 5025 35079 5105 35112
rect 5209 35158 5289 35171
rect 5209 35112 5222 35158
rect 5276 35112 5289 35158
rect 5209 35079 5289 35112
rect 4841 34546 4921 34579
rect 4841 34500 4854 34546
rect 4908 34500 4921 34546
rect 4841 34487 4921 34500
rect 5025 34546 5105 34579
rect 5025 34500 5038 34546
rect 5092 34500 5105 34546
rect 5025 34487 5105 34500
rect 5209 34546 5289 34579
rect 5209 34500 5222 34546
rect 5276 34500 5289 34546
rect 5209 34487 5289 34500
rect 6327 35158 6407 35171
rect 6327 35112 6340 35158
rect 6394 35112 6407 35158
rect 6327 35079 6407 35112
rect 6511 35158 6591 35171
rect 6511 35112 6524 35158
rect 6578 35112 6591 35158
rect 6511 35079 6591 35112
rect 6695 35158 6775 35171
rect 6695 35112 6708 35158
rect 6762 35112 6775 35158
rect 6695 35079 6775 35112
rect 6327 34546 6407 34579
rect 6327 34500 6340 34546
rect 6394 34500 6407 34546
rect 6327 34487 6407 34500
rect 6511 34546 6591 34579
rect 6511 34500 6524 34546
rect 6578 34500 6591 34546
rect 6511 34487 6591 34500
rect 6695 34546 6775 34579
rect 6695 34500 6708 34546
rect 6762 34500 6775 34546
rect 6695 34487 6775 34500
rect 14313 35159 14393 35172
rect 14313 35113 14326 35159
rect 14380 35113 14393 35159
rect 14313 35080 14393 35113
rect 14497 35159 14577 35172
rect 14497 35113 14510 35159
rect 14564 35113 14577 35159
rect 14497 35080 14577 35113
rect 14681 35159 14761 35172
rect 14681 35113 14694 35159
rect 14748 35113 14761 35159
rect 14681 35080 14761 35113
rect 14313 34547 14393 34580
rect 14313 34501 14326 34547
rect 14380 34501 14393 34547
rect 14313 34488 14393 34501
rect 14497 34547 14577 34580
rect 14497 34501 14510 34547
rect 14564 34501 14577 34547
rect 14497 34488 14577 34501
rect 14681 34547 14761 34580
rect 14681 34501 14694 34547
rect 14748 34501 14761 34547
rect 14681 34488 14761 34501
rect 15799 35159 15879 35172
rect 15799 35113 15812 35159
rect 15866 35113 15879 35159
rect 15799 35080 15879 35113
rect 15983 35159 16063 35172
rect 15983 35113 15996 35159
rect 16050 35113 16063 35159
rect 15983 35080 16063 35113
rect 16167 35159 16247 35172
rect 16167 35113 16180 35159
rect 16234 35113 16247 35159
rect 16167 35080 16247 35113
rect 15799 34547 15879 34580
rect 15799 34501 15812 34547
rect 15866 34501 15879 34547
rect 15799 34488 15879 34501
rect 15983 34547 16063 34580
rect 15983 34501 15996 34547
rect 16050 34501 16063 34547
rect 15983 34488 16063 34501
rect 16167 34547 16247 34580
rect 16167 34501 16180 34547
rect 16234 34501 16247 34547
rect 16167 34488 16247 34501
rect 23785 35159 23865 35172
rect 23785 35113 23798 35159
rect 23852 35113 23865 35159
rect 23785 35080 23865 35113
rect 23969 35159 24049 35172
rect 23969 35113 23982 35159
rect 24036 35113 24049 35159
rect 23969 35080 24049 35113
rect 24153 35159 24233 35172
rect 24153 35113 24166 35159
rect 24220 35113 24233 35159
rect 24153 35080 24233 35113
rect 23785 34547 23865 34580
rect 23785 34501 23798 34547
rect 23852 34501 23865 34547
rect 23785 34488 23865 34501
rect 23969 34547 24049 34580
rect 23969 34501 23982 34547
rect 24036 34501 24049 34547
rect 23969 34488 24049 34501
rect 24153 34547 24233 34580
rect 24153 34501 24166 34547
rect 24220 34501 24233 34547
rect 24153 34488 24233 34501
rect 25271 35159 25351 35172
rect 25271 35113 25284 35159
rect 25338 35113 25351 35159
rect 25271 35080 25351 35113
rect 25455 35159 25535 35172
rect 25455 35113 25468 35159
rect 25522 35113 25535 35159
rect 25455 35080 25535 35113
rect 25639 35159 25719 35172
rect 25639 35113 25652 35159
rect 25706 35113 25719 35159
rect 25639 35080 25719 35113
rect 25271 34547 25351 34580
rect 25271 34501 25284 34547
rect 25338 34501 25351 34547
rect 25271 34488 25351 34501
rect 25455 34547 25535 34580
rect 25455 34501 25468 34547
rect 25522 34501 25535 34547
rect 25455 34488 25535 34501
rect 25639 34547 25719 34580
rect 25639 34501 25652 34547
rect 25706 34501 25719 34547
rect 25639 34488 25719 34501
rect 33257 35159 33337 35172
rect 33257 35113 33270 35159
rect 33324 35113 33337 35159
rect 33257 35080 33337 35113
rect 33441 35159 33521 35172
rect 33441 35113 33454 35159
rect 33508 35113 33521 35159
rect 33441 35080 33521 35113
rect 33625 35159 33705 35172
rect 33625 35113 33638 35159
rect 33692 35113 33705 35159
rect 33625 35080 33705 35113
rect 33257 34547 33337 34580
rect 33257 34501 33270 34547
rect 33324 34501 33337 34547
rect 33257 34488 33337 34501
rect 33441 34547 33521 34580
rect 33441 34501 33454 34547
rect 33508 34501 33521 34547
rect 33441 34488 33521 34501
rect 33625 34547 33705 34580
rect 33625 34501 33638 34547
rect 33692 34501 33705 34547
rect 33625 34488 33705 34501
rect 34743 35159 34823 35172
rect 34743 35113 34756 35159
rect 34810 35113 34823 35159
rect 34743 35080 34823 35113
rect 34927 35159 35007 35172
rect 34927 35113 34940 35159
rect 34994 35113 35007 35159
rect 34927 35080 35007 35113
rect 35111 35159 35191 35172
rect 35111 35113 35124 35159
rect 35178 35113 35191 35159
rect 35111 35080 35191 35113
rect 34743 34547 34823 34580
rect 34743 34501 34756 34547
rect 34810 34501 34823 34547
rect 34743 34488 34823 34501
rect 34927 34547 35007 34580
rect 34927 34501 34940 34547
rect 34994 34501 35007 34547
rect 34927 34488 35007 34501
rect 35111 34547 35191 34580
rect 35111 34501 35124 34547
rect 35178 34501 35191 34547
rect 35111 34488 35191 34501
rect 42729 35159 42809 35172
rect 42729 35113 42742 35159
rect 42796 35113 42809 35159
rect 42729 35080 42809 35113
rect 42913 35159 42993 35172
rect 42913 35113 42926 35159
rect 42980 35113 42993 35159
rect 42913 35080 42993 35113
rect 43097 35159 43177 35172
rect 43097 35113 43110 35159
rect 43164 35113 43177 35159
rect 43097 35080 43177 35113
rect 42729 34547 42809 34580
rect 42729 34501 42742 34547
rect 42796 34501 42809 34547
rect 42729 34488 42809 34501
rect 42913 34547 42993 34580
rect 42913 34501 42926 34547
rect 42980 34501 42993 34547
rect 42913 34488 42993 34501
rect 43097 34547 43177 34580
rect 43097 34501 43110 34547
rect 43164 34501 43177 34547
rect 43097 34488 43177 34501
rect 44215 35159 44295 35172
rect 44215 35113 44228 35159
rect 44282 35113 44295 35159
rect 44215 35080 44295 35113
rect 44399 35159 44479 35172
rect 44399 35113 44412 35159
rect 44466 35113 44479 35159
rect 44399 35080 44479 35113
rect 44583 35159 44663 35172
rect 44583 35113 44596 35159
rect 44650 35113 44663 35159
rect 44583 35080 44663 35113
rect 44215 34547 44295 34580
rect 44215 34501 44228 34547
rect 44282 34501 44295 34547
rect 44215 34488 44295 34501
rect 44399 34547 44479 34580
rect 44399 34501 44412 34547
rect 44466 34501 44479 34547
rect 44399 34488 44479 34501
rect 44583 34547 44663 34580
rect 44583 34501 44596 34547
rect 44650 34501 44663 34547
rect 44583 34488 44663 34501
rect -4631 33998 -4551 34011
rect -4631 33952 -4618 33998
rect -4564 33952 -4551 33998
rect -4631 33919 -4551 33952
rect -4447 33998 -4367 34011
rect -4447 33952 -4434 33998
rect -4380 33952 -4367 33998
rect -4447 33919 -4367 33952
rect -4263 33998 -4183 34011
rect -4263 33952 -4250 33998
rect -4196 33952 -4183 33998
rect -4263 33919 -4183 33952
rect -4631 33686 -4551 33719
rect -4631 33640 -4618 33686
rect -4564 33640 -4551 33686
rect -4631 33627 -4551 33640
rect -4447 33686 -4367 33719
rect -4447 33640 -4434 33686
rect -4380 33640 -4367 33686
rect -4447 33627 -4367 33640
rect -4263 33686 -4183 33719
rect -4263 33640 -4250 33686
rect -4196 33640 -4183 33686
rect -4263 33627 -4183 33640
rect -3145 33998 -3065 34011
rect -3145 33952 -3132 33998
rect -3078 33952 -3065 33998
rect -3145 33919 -3065 33952
rect -2961 33998 -2881 34011
rect -2961 33952 -2948 33998
rect -2894 33952 -2881 33998
rect -2961 33919 -2881 33952
rect -2777 33998 -2697 34011
rect -2777 33952 -2764 33998
rect -2710 33952 -2697 33998
rect -2777 33919 -2697 33952
rect -3145 33686 -3065 33719
rect -3145 33640 -3132 33686
rect -3078 33640 -3065 33686
rect -3145 33627 -3065 33640
rect -2961 33686 -2881 33719
rect -2961 33640 -2948 33686
rect -2894 33640 -2881 33686
rect -2961 33627 -2881 33640
rect -2777 33686 -2697 33719
rect -2777 33640 -2764 33686
rect -2710 33640 -2697 33686
rect -2777 33627 -2697 33640
rect 4841 33998 4921 34011
rect 4841 33952 4854 33998
rect 4908 33952 4921 33998
rect 4841 33919 4921 33952
rect 5025 33998 5105 34011
rect 5025 33952 5038 33998
rect 5092 33952 5105 33998
rect 5025 33919 5105 33952
rect 5209 33998 5289 34011
rect 5209 33952 5222 33998
rect 5276 33952 5289 33998
rect 5209 33919 5289 33952
rect 4841 33686 4921 33719
rect 4841 33640 4854 33686
rect 4908 33640 4921 33686
rect 4841 33627 4921 33640
rect 5025 33686 5105 33719
rect 5025 33640 5038 33686
rect 5092 33640 5105 33686
rect 5025 33627 5105 33640
rect 5209 33686 5289 33719
rect 5209 33640 5222 33686
rect 5276 33640 5289 33686
rect 5209 33627 5289 33640
rect 6327 33998 6407 34011
rect 6327 33952 6340 33998
rect 6394 33952 6407 33998
rect 6327 33919 6407 33952
rect 6511 33998 6591 34011
rect 6511 33952 6524 33998
rect 6578 33952 6591 33998
rect 6511 33919 6591 33952
rect 6695 33998 6775 34011
rect 6695 33952 6708 33998
rect 6762 33952 6775 33998
rect 6695 33919 6775 33952
rect 6327 33686 6407 33719
rect 6327 33640 6340 33686
rect 6394 33640 6407 33686
rect 6327 33627 6407 33640
rect 6511 33686 6591 33719
rect 6511 33640 6524 33686
rect 6578 33640 6591 33686
rect 6511 33627 6591 33640
rect 6695 33686 6775 33719
rect 6695 33640 6708 33686
rect 6762 33640 6775 33686
rect 6695 33627 6775 33640
rect 14313 33999 14393 34012
rect 14313 33953 14326 33999
rect 14380 33953 14393 33999
rect 14313 33920 14393 33953
rect 14497 33999 14577 34012
rect 14497 33953 14510 33999
rect 14564 33953 14577 33999
rect 14497 33920 14577 33953
rect 14681 33999 14761 34012
rect 14681 33953 14694 33999
rect 14748 33953 14761 33999
rect 14681 33920 14761 33953
rect 14313 33687 14393 33720
rect 14313 33641 14326 33687
rect 14380 33641 14393 33687
rect 14313 33628 14393 33641
rect 14497 33687 14577 33720
rect 14497 33641 14510 33687
rect 14564 33641 14577 33687
rect 14497 33628 14577 33641
rect 14681 33687 14761 33720
rect 14681 33641 14694 33687
rect 14748 33641 14761 33687
rect 14681 33628 14761 33641
rect 15799 33999 15879 34012
rect 15799 33953 15812 33999
rect 15866 33953 15879 33999
rect 15799 33920 15879 33953
rect 15983 33999 16063 34012
rect 15983 33953 15996 33999
rect 16050 33953 16063 33999
rect 15983 33920 16063 33953
rect 16167 33999 16247 34012
rect 16167 33953 16180 33999
rect 16234 33953 16247 33999
rect 16167 33920 16247 33953
rect 15799 33687 15879 33720
rect 15799 33641 15812 33687
rect 15866 33641 15879 33687
rect 15799 33628 15879 33641
rect 15983 33687 16063 33720
rect 15983 33641 15996 33687
rect 16050 33641 16063 33687
rect 15983 33628 16063 33641
rect 16167 33687 16247 33720
rect 16167 33641 16180 33687
rect 16234 33641 16247 33687
rect 16167 33628 16247 33641
rect 23785 33999 23865 34012
rect 23785 33953 23798 33999
rect 23852 33953 23865 33999
rect 23785 33920 23865 33953
rect 23969 33999 24049 34012
rect 23969 33953 23982 33999
rect 24036 33953 24049 33999
rect 23969 33920 24049 33953
rect 24153 33999 24233 34012
rect 24153 33953 24166 33999
rect 24220 33953 24233 33999
rect 24153 33920 24233 33953
rect 23785 33687 23865 33720
rect 23785 33641 23798 33687
rect 23852 33641 23865 33687
rect 23785 33628 23865 33641
rect 23969 33687 24049 33720
rect 23969 33641 23982 33687
rect 24036 33641 24049 33687
rect 23969 33628 24049 33641
rect 24153 33687 24233 33720
rect 24153 33641 24166 33687
rect 24220 33641 24233 33687
rect 24153 33628 24233 33641
rect 25271 33999 25351 34012
rect 25271 33953 25284 33999
rect 25338 33953 25351 33999
rect 25271 33920 25351 33953
rect 25455 33999 25535 34012
rect 25455 33953 25468 33999
rect 25522 33953 25535 33999
rect 25455 33920 25535 33953
rect 25639 33999 25719 34012
rect 25639 33953 25652 33999
rect 25706 33953 25719 33999
rect 25639 33920 25719 33953
rect 25271 33687 25351 33720
rect 25271 33641 25284 33687
rect 25338 33641 25351 33687
rect 25271 33628 25351 33641
rect 25455 33687 25535 33720
rect 25455 33641 25468 33687
rect 25522 33641 25535 33687
rect 25455 33628 25535 33641
rect 25639 33687 25719 33720
rect 25639 33641 25652 33687
rect 25706 33641 25719 33687
rect 25639 33628 25719 33641
rect 33257 33999 33337 34012
rect 33257 33953 33270 33999
rect 33324 33953 33337 33999
rect 33257 33920 33337 33953
rect 33441 33999 33521 34012
rect 33441 33953 33454 33999
rect 33508 33953 33521 33999
rect 33441 33920 33521 33953
rect 33625 33999 33705 34012
rect 33625 33953 33638 33999
rect 33692 33953 33705 33999
rect 33625 33920 33705 33953
rect 33257 33687 33337 33720
rect 33257 33641 33270 33687
rect 33324 33641 33337 33687
rect 33257 33628 33337 33641
rect 33441 33687 33521 33720
rect 33441 33641 33454 33687
rect 33508 33641 33521 33687
rect 33441 33628 33521 33641
rect 33625 33687 33705 33720
rect 33625 33641 33638 33687
rect 33692 33641 33705 33687
rect 33625 33628 33705 33641
rect 34743 33999 34823 34012
rect 34743 33953 34756 33999
rect 34810 33953 34823 33999
rect 34743 33920 34823 33953
rect 34927 33999 35007 34012
rect 34927 33953 34940 33999
rect 34994 33953 35007 33999
rect 34927 33920 35007 33953
rect 35111 33999 35191 34012
rect 35111 33953 35124 33999
rect 35178 33953 35191 33999
rect 35111 33920 35191 33953
rect 34743 33687 34823 33720
rect 34743 33641 34756 33687
rect 34810 33641 34823 33687
rect 34743 33628 34823 33641
rect 34927 33687 35007 33720
rect 34927 33641 34940 33687
rect 34994 33641 35007 33687
rect 34927 33628 35007 33641
rect 35111 33687 35191 33720
rect 35111 33641 35124 33687
rect 35178 33641 35191 33687
rect 35111 33628 35191 33641
rect 42729 33999 42809 34012
rect 42729 33953 42742 33999
rect 42796 33953 42809 33999
rect 42729 33920 42809 33953
rect 42913 33999 42993 34012
rect 42913 33953 42926 33999
rect 42980 33953 42993 33999
rect 42913 33920 42993 33953
rect 43097 33999 43177 34012
rect 43097 33953 43110 33999
rect 43164 33953 43177 33999
rect 43097 33920 43177 33953
rect 42729 33687 42809 33720
rect 42729 33641 42742 33687
rect 42796 33641 42809 33687
rect 42729 33628 42809 33641
rect 42913 33687 42993 33720
rect 42913 33641 42926 33687
rect 42980 33641 42993 33687
rect 42913 33628 42993 33641
rect 43097 33687 43177 33720
rect 43097 33641 43110 33687
rect 43164 33641 43177 33687
rect 43097 33628 43177 33641
rect 44215 33999 44295 34012
rect 44215 33953 44228 33999
rect 44282 33953 44295 33999
rect 44215 33920 44295 33953
rect 44399 33999 44479 34012
rect 44399 33953 44412 33999
rect 44466 33953 44479 33999
rect 44399 33920 44479 33953
rect 44583 33999 44663 34012
rect 44583 33953 44596 33999
rect 44650 33953 44663 33999
rect 44583 33920 44663 33953
rect 44215 33687 44295 33720
rect 44215 33641 44228 33687
rect 44282 33641 44295 33687
rect 44215 33628 44295 33641
rect 44399 33687 44479 33720
rect 44399 33641 44412 33687
rect 44466 33641 44479 33687
rect 44399 33628 44479 33641
rect 44583 33687 44663 33720
rect 44583 33641 44596 33687
rect 44650 33641 44663 33687
rect 44583 33628 44663 33641
rect -4631 32953 -4551 32966
rect -4631 32907 -4618 32953
rect -4564 32907 -4551 32953
rect -4631 32874 -4551 32907
rect -4447 32953 -4367 32966
rect -4447 32907 -4434 32953
rect -4380 32907 -4367 32953
rect -4447 32874 -4367 32907
rect -4263 32953 -4183 32966
rect -4263 32907 -4250 32953
rect -4196 32907 -4183 32953
rect -4263 32874 -4183 32907
rect -4631 32341 -4551 32374
rect -4631 32295 -4618 32341
rect -4564 32295 -4551 32341
rect -4631 32282 -4551 32295
rect -4447 32341 -4367 32374
rect -4447 32295 -4434 32341
rect -4380 32295 -4367 32341
rect -4447 32282 -4367 32295
rect -4263 32341 -4183 32374
rect -4263 32295 -4250 32341
rect -4196 32295 -4183 32341
rect -4263 32282 -4183 32295
rect -3145 32954 -3065 32967
rect -3145 32908 -3132 32954
rect -3078 32908 -3065 32954
rect -3145 32875 -3065 32908
rect -2961 32954 -2881 32967
rect -2961 32908 -2948 32954
rect -2894 32908 -2881 32954
rect -2961 32875 -2881 32908
rect -2777 32954 -2697 32967
rect -2777 32908 -2764 32954
rect -2710 32908 -2697 32954
rect -2777 32875 -2697 32908
rect -3145 32342 -3065 32375
rect -3145 32296 -3132 32342
rect -3078 32296 -3065 32342
rect -3145 32283 -3065 32296
rect -2961 32342 -2881 32375
rect -2961 32296 -2948 32342
rect -2894 32296 -2881 32342
rect -2961 32283 -2881 32296
rect -2777 32342 -2697 32375
rect -2777 32296 -2764 32342
rect -2710 32296 -2697 32342
rect -2777 32283 -2697 32296
rect 4841 32953 4921 32966
rect 4841 32907 4854 32953
rect 4908 32907 4921 32953
rect 4841 32874 4921 32907
rect 5025 32953 5105 32966
rect 5025 32907 5038 32953
rect 5092 32907 5105 32953
rect 5025 32874 5105 32907
rect 5209 32953 5289 32966
rect 5209 32907 5222 32953
rect 5276 32907 5289 32953
rect 5209 32874 5289 32907
rect 4841 32341 4921 32374
rect 4841 32295 4854 32341
rect 4908 32295 4921 32341
rect 4841 32282 4921 32295
rect 5025 32341 5105 32374
rect 5025 32295 5038 32341
rect 5092 32295 5105 32341
rect 5025 32282 5105 32295
rect 5209 32341 5289 32374
rect 5209 32295 5222 32341
rect 5276 32295 5289 32341
rect 5209 32282 5289 32295
rect 6327 32954 6407 32967
rect 6327 32908 6340 32954
rect 6394 32908 6407 32954
rect 6327 32875 6407 32908
rect 6511 32954 6591 32967
rect 6511 32908 6524 32954
rect 6578 32908 6591 32954
rect 6511 32875 6591 32908
rect 6695 32954 6775 32967
rect 6695 32908 6708 32954
rect 6762 32908 6775 32954
rect 6695 32875 6775 32908
rect 6327 32342 6407 32375
rect 6327 32296 6340 32342
rect 6394 32296 6407 32342
rect 6327 32283 6407 32296
rect 6511 32342 6591 32375
rect 6511 32296 6524 32342
rect 6578 32296 6591 32342
rect 6511 32283 6591 32296
rect 6695 32342 6775 32375
rect 6695 32296 6708 32342
rect 6762 32296 6775 32342
rect 6695 32283 6775 32296
rect 14313 32954 14393 32967
rect 14313 32908 14326 32954
rect 14380 32908 14393 32954
rect 14313 32875 14393 32908
rect 14497 32954 14577 32967
rect 14497 32908 14510 32954
rect 14564 32908 14577 32954
rect 14497 32875 14577 32908
rect 14681 32954 14761 32967
rect 14681 32908 14694 32954
rect 14748 32908 14761 32954
rect 14681 32875 14761 32908
rect 14313 32342 14393 32375
rect 14313 32296 14326 32342
rect 14380 32296 14393 32342
rect 14313 32283 14393 32296
rect 14497 32342 14577 32375
rect 14497 32296 14510 32342
rect 14564 32296 14577 32342
rect 14497 32283 14577 32296
rect 14681 32342 14761 32375
rect 14681 32296 14694 32342
rect 14748 32296 14761 32342
rect 14681 32283 14761 32296
rect 15799 32955 15879 32968
rect 15799 32909 15812 32955
rect 15866 32909 15879 32955
rect 15799 32876 15879 32909
rect 15983 32955 16063 32968
rect 15983 32909 15996 32955
rect 16050 32909 16063 32955
rect 15983 32876 16063 32909
rect 16167 32955 16247 32968
rect 16167 32909 16180 32955
rect 16234 32909 16247 32955
rect 16167 32876 16247 32909
rect 15799 32343 15879 32376
rect 15799 32297 15812 32343
rect 15866 32297 15879 32343
rect 15799 32284 15879 32297
rect 15983 32343 16063 32376
rect 15983 32297 15996 32343
rect 16050 32297 16063 32343
rect 15983 32284 16063 32297
rect 16167 32343 16247 32376
rect 16167 32297 16180 32343
rect 16234 32297 16247 32343
rect 16167 32284 16247 32297
rect 23785 32954 23865 32967
rect 23785 32908 23798 32954
rect 23852 32908 23865 32954
rect 23785 32875 23865 32908
rect 23969 32954 24049 32967
rect 23969 32908 23982 32954
rect 24036 32908 24049 32954
rect 23969 32875 24049 32908
rect 24153 32954 24233 32967
rect 24153 32908 24166 32954
rect 24220 32908 24233 32954
rect 24153 32875 24233 32908
rect 23785 32342 23865 32375
rect 23785 32296 23798 32342
rect 23852 32296 23865 32342
rect 23785 32283 23865 32296
rect 23969 32342 24049 32375
rect 23969 32296 23982 32342
rect 24036 32296 24049 32342
rect 23969 32283 24049 32296
rect 24153 32342 24233 32375
rect 24153 32296 24166 32342
rect 24220 32296 24233 32342
rect 24153 32283 24233 32296
rect 25271 32955 25351 32968
rect 25271 32909 25284 32955
rect 25338 32909 25351 32955
rect 25271 32876 25351 32909
rect 25455 32955 25535 32968
rect 25455 32909 25468 32955
rect 25522 32909 25535 32955
rect 25455 32876 25535 32909
rect 25639 32955 25719 32968
rect 25639 32909 25652 32955
rect 25706 32909 25719 32955
rect 25639 32876 25719 32909
rect 25271 32343 25351 32376
rect 25271 32297 25284 32343
rect 25338 32297 25351 32343
rect 25271 32284 25351 32297
rect 25455 32343 25535 32376
rect 25455 32297 25468 32343
rect 25522 32297 25535 32343
rect 25455 32284 25535 32297
rect 25639 32343 25719 32376
rect 25639 32297 25652 32343
rect 25706 32297 25719 32343
rect 25639 32284 25719 32297
rect 33257 32954 33337 32967
rect 33257 32908 33270 32954
rect 33324 32908 33337 32954
rect 33257 32875 33337 32908
rect 33441 32954 33521 32967
rect 33441 32908 33454 32954
rect 33508 32908 33521 32954
rect 33441 32875 33521 32908
rect 33625 32954 33705 32967
rect 33625 32908 33638 32954
rect 33692 32908 33705 32954
rect 33625 32875 33705 32908
rect 33257 32342 33337 32375
rect 33257 32296 33270 32342
rect 33324 32296 33337 32342
rect 33257 32283 33337 32296
rect 33441 32342 33521 32375
rect 33441 32296 33454 32342
rect 33508 32296 33521 32342
rect 33441 32283 33521 32296
rect 33625 32342 33705 32375
rect 33625 32296 33638 32342
rect 33692 32296 33705 32342
rect 33625 32283 33705 32296
rect 34743 32955 34823 32968
rect 34743 32909 34756 32955
rect 34810 32909 34823 32955
rect 34743 32876 34823 32909
rect 34927 32955 35007 32968
rect 34927 32909 34940 32955
rect 34994 32909 35007 32955
rect 34927 32876 35007 32909
rect 35111 32955 35191 32968
rect 35111 32909 35124 32955
rect 35178 32909 35191 32955
rect 35111 32876 35191 32909
rect 34743 32343 34823 32376
rect 34743 32297 34756 32343
rect 34810 32297 34823 32343
rect 34743 32284 34823 32297
rect 34927 32343 35007 32376
rect 34927 32297 34940 32343
rect 34994 32297 35007 32343
rect 34927 32284 35007 32297
rect 35111 32343 35191 32376
rect 35111 32297 35124 32343
rect 35178 32297 35191 32343
rect 35111 32284 35191 32297
rect 42729 32954 42809 32967
rect 42729 32908 42742 32954
rect 42796 32908 42809 32954
rect 42729 32875 42809 32908
rect 42913 32954 42993 32967
rect 42913 32908 42926 32954
rect 42980 32908 42993 32954
rect 42913 32875 42993 32908
rect 43097 32954 43177 32967
rect 43097 32908 43110 32954
rect 43164 32908 43177 32954
rect 43097 32875 43177 32908
rect 42729 32342 42809 32375
rect 42729 32296 42742 32342
rect 42796 32296 42809 32342
rect 42729 32283 42809 32296
rect 42913 32342 42993 32375
rect 42913 32296 42926 32342
rect 42980 32296 42993 32342
rect 42913 32283 42993 32296
rect 43097 32342 43177 32375
rect 43097 32296 43110 32342
rect 43164 32296 43177 32342
rect 43097 32283 43177 32296
rect 44215 32955 44295 32968
rect 44215 32909 44228 32955
rect 44282 32909 44295 32955
rect 44215 32876 44295 32909
rect 44399 32955 44479 32968
rect 44399 32909 44412 32955
rect 44466 32909 44479 32955
rect 44399 32876 44479 32909
rect 44583 32955 44663 32968
rect 44583 32909 44596 32955
rect 44650 32909 44663 32955
rect 44583 32876 44663 32909
rect 44215 32343 44295 32376
rect 44215 32297 44228 32343
rect 44282 32297 44295 32343
rect 44215 32284 44295 32297
rect 44399 32343 44479 32376
rect 44399 32297 44412 32343
rect 44466 32297 44479 32343
rect 44399 32284 44479 32297
rect 44583 32343 44663 32376
rect 44583 32297 44596 32343
rect 44650 32297 44663 32343
rect 44583 32284 44663 32297
rect -9773 31838 -9673 31851
rect -9773 31792 -9760 31838
rect -9686 31792 -9673 31838
rect -9773 31759 -9673 31792
rect -9773 31126 -9673 31159
rect -9773 31080 -9760 31126
rect -9686 31080 -9673 31126
rect -9773 31067 -9673 31080
rect -8885 31838 -8785 31851
rect -8885 31792 -8872 31838
rect -8798 31792 -8785 31838
rect -8885 31759 -8785 31792
rect -8885 31126 -8785 31159
rect -8885 31080 -8872 31126
rect -8798 31080 -8785 31126
rect -8885 31067 -8785 31080
rect -8405 31838 -8305 31851
rect -8405 31792 -8392 31838
rect -8318 31792 -8305 31838
rect -8405 31759 -8305 31792
rect -8405 31126 -8305 31159
rect -8405 31080 -8392 31126
rect -8318 31080 -8305 31126
rect -8405 31067 -8305 31080
rect -4631 31793 -4551 31806
rect -4631 31747 -4618 31793
rect -4564 31747 -4551 31793
rect -4631 31714 -4551 31747
rect -4447 31793 -4367 31806
rect -4447 31747 -4434 31793
rect -4380 31747 -4367 31793
rect -4447 31714 -4367 31747
rect -4263 31793 -4183 31806
rect -4263 31747 -4250 31793
rect -4196 31747 -4183 31793
rect -4263 31714 -4183 31747
rect -4631 31481 -4551 31514
rect -4631 31435 -4618 31481
rect -4564 31435 -4551 31481
rect -4631 31422 -4551 31435
rect -4447 31481 -4367 31514
rect -4447 31435 -4434 31481
rect -4380 31435 -4367 31481
rect -4447 31422 -4367 31435
rect -4263 31481 -4183 31514
rect -4263 31435 -4250 31481
rect -4196 31435 -4183 31481
rect -4263 31422 -4183 31435
rect -3145 31794 -3065 31807
rect -3145 31748 -3132 31794
rect -3078 31748 -3065 31794
rect -3145 31715 -3065 31748
rect -2961 31794 -2881 31807
rect -2961 31748 -2948 31794
rect -2894 31748 -2881 31794
rect -2961 31715 -2881 31748
rect -2777 31794 -2697 31807
rect -2777 31748 -2764 31794
rect -2710 31748 -2697 31794
rect -2777 31715 -2697 31748
rect -3145 31482 -3065 31515
rect -3145 31436 -3132 31482
rect -3078 31436 -3065 31482
rect -3145 31423 -3065 31436
rect -2961 31482 -2881 31515
rect -2961 31436 -2948 31482
rect -2894 31436 -2881 31482
rect -2961 31423 -2881 31436
rect -2777 31482 -2697 31515
rect -2777 31436 -2764 31482
rect -2710 31436 -2697 31482
rect -2777 31423 -2697 31436
rect -301 31838 -201 31851
rect -301 31792 -288 31838
rect -214 31792 -201 31838
rect -301 31759 -201 31792
rect -301 31126 -201 31159
rect -301 31080 -288 31126
rect -214 31080 -201 31126
rect -301 31067 -201 31080
rect 587 31838 687 31851
rect 587 31792 600 31838
rect 674 31792 687 31838
rect 587 31759 687 31792
rect 587 31126 687 31159
rect 587 31080 600 31126
rect 674 31080 687 31126
rect 587 31067 687 31080
rect 1067 31838 1167 31851
rect 1067 31792 1080 31838
rect 1154 31792 1167 31838
rect 1067 31759 1167 31792
rect 1067 31126 1167 31159
rect 1067 31080 1080 31126
rect 1154 31080 1167 31126
rect 1067 31067 1167 31080
rect 4841 31793 4921 31806
rect 4841 31747 4854 31793
rect 4908 31747 4921 31793
rect 4841 31714 4921 31747
rect 5025 31793 5105 31806
rect 5025 31747 5038 31793
rect 5092 31747 5105 31793
rect 5025 31714 5105 31747
rect 5209 31793 5289 31806
rect 5209 31747 5222 31793
rect 5276 31747 5289 31793
rect 5209 31714 5289 31747
rect 4841 31481 4921 31514
rect 4841 31435 4854 31481
rect 4908 31435 4921 31481
rect 4841 31422 4921 31435
rect 5025 31481 5105 31514
rect 5025 31435 5038 31481
rect 5092 31435 5105 31481
rect 5025 31422 5105 31435
rect 5209 31481 5289 31514
rect 5209 31435 5222 31481
rect 5276 31435 5289 31481
rect 5209 31422 5289 31435
rect 6327 31794 6407 31807
rect 6327 31748 6340 31794
rect 6394 31748 6407 31794
rect 6327 31715 6407 31748
rect 6511 31794 6591 31807
rect 6511 31748 6524 31794
rect 6578 31748 6591 31794
rect 6511 31715 6591 31748
rect 6695 31794 6775 31807
rect 6695 31748 6708 31794
rect 6762 31748 6775 31794
rect 6695 31715 6775 31748
rect 6327 31482 6407 31515
rect 6327 31436 6340 31482
rect 6394 31436 6407 31482
rect 6327 31423 6407 31436
rect 6511 31482 6591 31515
rect 6511 31436 6524 31482
rect 6578 31436 6591 31482
rect 6511 31423 6591 31436
rect 6695 31482 6775 31515
rect 6695 31436 6708 31482
rect 6762 31436 6775 31482
rect 6695 31423 6775 31436
rect 9171 31839 9271 31852
rect 9171 31793 9184 31839
rect 9258 31793 9271 31839
rect 9171 31760 9271 31793
rect 9171 31127 9271 31160
rect 9171 31081 9184 31127
rect 9258 31081 9271 31127
rect 9171 31068 9271 31081
rect 10059 31839 10159 31852
rect 10059 31793 10072 31839
rect 10146 31793 10159 31839
rect 10059 31760 10159 31793
rect 10059 31127 10159 31160
rect 10059 31081 10072 31127
rect 10146 31081 10159 31127
rect 10059 31068 10159 31081
rect 10539 31839 10639 31852
rect 10539 31793 10552 31839
rect 10626 31793 10639 31839
rect 10539 31760 10639 31793
rect 10539 31127 10639 31160
rect 10539 31081 10552 31127
rect 10626 31081 10639 31127
rect 10539 31068 10639 31081
rect 14313 31794 14393 31807
rect 14313 31748 14326 31794
rect 14380 31748 14393 31794
rect 14313 31715 14393 31748
rect 14497 31794 14577 31807
rect 14497 31748 14510 31794
rect 14564 31748 14577 31794
rect 14497 31715 14577 31748
rect 14681 31794 14761 31807
rect 14681 31748 14694 31794
rect 14748 31748 14761 31794
rect 14681 31715 14761 31748
rect 14313 31482 14393 31515
rect 14313 31436 14326 31482
rect 14380 31436 14393 31482
rect 14313 31423 14393 31436
rect 14497 31482 14577 31515
rect 14497 31436 14510 31482
rect 14564 31436 14577 31482
rect 14497 31423 14577 31436
rect 14681 31482 14761 31515
rect 14681 31436 14694 31482
rect 14748 31436 14761 31482
rect 14681 31423 14761 31436
rect 15799 31795 15879 31808
rect 15799 31749 15812 31795
rect 15866 31749 15879 31795
rect 15799 31716 15879 31749
rect 15983 31795 16063 31808
rect 15983 31749 15996 31795
rect 16050 31749 16063 31795
rect 15983 31716 16063 31749
rect 16167 31795 16247 31808
rect 16167 31749 16180 31795
rect 16234 31749 16247 31795
rect 16167 31716 16247 31749
rect 15799 31483 15879 31516
rect 15799 31437 15812 31483
rect 15866 31437 15879 31483
rect 15799 31424 15879 31437
rect 15983 31483 16063 31516
rect 15983 31437 15996 31483
rect 16050 31437 16063 31483
rect 15983 31424 16063 31437
rect 16167 31483 16247 31516
rect 16167 31437 16180 31483
rect 16234 31437 16247 31483
rect 16167 31424 16247 31437
rect 18643 31839 18743 31852
rect 18643 31793 18656 31839
rect 18730 31793 18743 31839
rect 18643 31760 18743 31793
rect 18643 31127 18743 31160
rect 18643 31081 18656 31127
rect 18730 31081 18743 31127
rect 18643 31068 18743 31081
rect 19531 31839 19631 31852
rect 19531 31793 19544 31839
rect 19618 31793 19631 31839
rect 19531 31760 19631 31793
rect 19531 31127 19631 31160
rect 19531 31081 19544 31127
rect 19618 31081 19631 31127
rect 19531 31068 19631 31081
rect 20011 31839 20111 31852
rect 20011 31793 20024 31839
rect 20098 31793 20111 31839
rect 20011 31760 20111 31793
rect 20011 31127 20111 31160
rect 20011 31081 20024 31127
rect 20098 31081 20111 31127
rect 20011 31068 20111 31081
rect 23785 31794 23865 31807
rect 23785 31748 23798 31794
rect 23852 31748 23865 31794
rect 23785 31715 23865 31748
rect 23969 31794 24049 31807
rect 23969 31748 23982 31794
rect 24036 31748 24049 31794
rect 23969 31715 24049 31748
rect 24153 31794 24233 31807
rect 24153 31748 24166 31794
rect 24220 31748 24233 31794
rect 24153 31715 24233 31748
rect 23785 31482 23865 31515
rect 23785 31436 23798 31482
rect 23852 31436 23865 31482
rect 23785 31423 23865 31436
rect 23969 31482 24049 31515
rect 23969 31436 23982 31482
rect 24036 31436 24049 31482
rect 23969 31423 24049 31436
rect 24153 31482 24233 31515
rect 24153 31436 24166 31482
rect 24220 31436 24233 31482
rect 24153 31423 24233 31436
rect 25271 31795 25351 31808
rect 25271 31749 25284 31795
rect 25338 31749 25351 31795
rect 25271 31716 25351 31749
rect 25455 31795 25535 31808
rect 25455 31749 25468 31795
rect 25522 31749 25535 31795
rect 25455 31716 25535 31749
rect 25639 31795 25719 31808
rect 25639 31749 25652 31795
rect 25706 31749 25719 31795
rect 25639 31716 25719 31749
rect 25271 31483 25351 31516
rect 25271 31437 25284 31483
rect 25338 31437 25351 31483
rect 25271 31424 25351 31437
rect 25455 31483 25535 31516
rect 25455 31437 25468 31483
rect 25522 31437 25535 31483
rect 25455 31424 25535 31437
rect 25639 31483 25719 31516
rect 25639 31437 25652 31483
rect 25706 31437 25719 31483
rect 25639 31424 25719 31437
rect 28115 31839 28215 31852
rect 28115 31793 28128 31839
rect 28202 31793 28215 31839
rect 28115 31760 28215 31793
rect 28115 31127 28215 31160
rect 28115 31081 28128 31127
rect 28202 31081 28215 31127
rect 28115 31068 28215 31081
rect 29003 31839 29103 31852
rect 29003 31793 29016 31839
rect 29090 31793 29103 31839
rect 29003 31760 29103 31793
rect 29003 31127 29103 31160
rect 29003 31081 29016 31127
rect 29090 31081 29103 31127
rect 29003 31068 29103 31081
rect 29483 31839 29583 31852
rect 29483 31793 29496 31839
rect 29570 31793 29583 31839
rect 29483 31760 29583 31793
rect 29483 31127 29583 31160
rect 29483 31081 29496 31127
rect 29570 31081 29583 31127
rect 29483 31068 29583 31081
rect 33257 31794 33337 31807
rect 33257 31748 33270 31794
rect 33324 31748 33337 31794
rect 33257 31715 33337 31748
rect 33441 31794 33521 31807
rect 33441 31748 33454 31794
rect 33508 31748 33521 31794
rect 33441 31715 33521 31748
rect 33625 31794 33705 31807
rect 33625 31748 33638 31794
rect 33692 31748 33705 31794
rect 33625 31715 33705 31748
rect 33257 31482 33337 31515
rect 33257 31436 33270 31482
rect 33324 31436 33337 31482
rect 33257 31423 33337 31436
rect 33441 31482 33521 31515
rect 33441 31436 33454 31482
rect 33508 31436 33521 31482
rect 33441 31423 33521 31436
rect 33625 31482 33705 31515
rect 33625 31436 33638 31482
rect 33692 31436 33705 31482
rect 33625 31423 33705 31436
rect 34743 31795 34823 31808
rect 34743 31749 34756 31795
rect 34810 31749 34823 31795
rect 34743 31716 34823 31749
rect 34927 31795 35007 31808
rect 34927 31749 34940 31795
rect 34994 31749 35007 31795
rect 34927 31716 35007 31749
rect 35111 31795 35191 31808
rect 35111 31749 35124 31795
rect 35178 31749 35191 31795
rect 35111 31716 35191 31749
rect 34743 31483 34823 31516
rect 34743 31437 34756 31483
rect 34810 31437 34823 31483
rect 34743 31424 34823 31437
rect 34927 31483 35007 31516
rect 34927 31437 34940 31483
rect 34994 31437 35007 31483
rect 34927 31424 35007 31437
rect 35111 31483 35191 31516
rect 35111 31437 35124 31483
rect 35178 31437 35191 31483
rect 35111 31424 35191 31437
rect 37587 31839 37687 31852
rect 37587 31793 37600 31839
rect 37674 31793 37687 31839
rect 37587 31760 37687 31793
rect 37587 31127 37687 31160
rect 37587 31081 37600 31127
rect 37674 31081 37687 31127
rect 37587 31068 37687 31081
rect 38475 31839 38575 31852
rect 38475 31793 38488 31839
rect 38562 31793 38575 31839
rect 38475 31760 38575 31793
rect 38475 31127 38575 31160
rect 38475 31081 38488 31127
rect 38562 31081 38575 31127
rect 38475 31068 38575 31081
rect 38955 31839 39055 31852
rect 38955 31793 38968 31839
rect 39042 31793 39055 31839
rect 38955 31760 39055 31793
rect 38955 31127 39055 31160
rect 38955 31081 38968 31127
rect 39042 31081 39055 31127
rect 38955 31068 39055 31081
rect 42729 31794 42809 31807
rect 42729 31748 42742 31794
rect 42796 31748 42809 31794
rect 42729 31715 42809 31748
rect 42913 31794 42993 31807
rect 42913 31748 42926 31794
rect 42980 31748 42993 31794
rect 42913 31715 42993 31748
rect 43097 31794 43177 31807
rect 43097 31748 43110 31794
rect 43164 31748 43177 31794
rect 43097 31715 43177 31748
rect 42729 31482 42809 31515
rect 42729 31436 42742 31482
rect 42796 31436 42809 31482
rect 42729 31423 42809 31436
rect 42913 31482 42993 31515
rect 42913 31436 42926 31482
rect 42980 31436 42993 31482
rect 42913 31423 42993 31436
rect 43097 31482 43177 31515
rect 43097 31436 43110 31482
rect 43164 31436 43177 31482
rect 43097 31423 43177 31436
rect 44215 31795 44295 31808
rect 44215 31749 44228 31795
rect 44282 31749 44295 31795
rect 44215 31716 44295 31749
rect 44399 31795 44479 31808
rect 44399 31749 44412 31795
rect 44466 31749 44479 31795
rect 44399 31716 44479 31749
rect 44583 31795 44663 31808
rect 44583 31749 44596 31795
rect 44650 31749 44663 31795
rect 44583 31716 44663 31749
rect 44215 31483 44295 31516
rect 44215 31437 44228 31483
rect 44282 31437 44295 31483
rect 44215 31424 44295 31437
rect 44399 31483 44479 31516
rect 44399 31437 44412 31483
rect 44466 31437 44479 31483
rect 44399 31424 44479 31437
rect 44583 31483 44663 31516
rect 44583 31437 44596 31483
rect 44650 31437 44663 31483
rect 44583 31424 44663 31437
rect -10667 30418 -10567 30431
rect -10667 30372 -10654 30418
rect -10580 30372 -10567 30418
rect -10667 30339 -10567 30372
rect -10667 29706 -10567 29739
rect -10667 29660 -10654 29706
rect -10580 29660 -10567 29706
rect -10667 29647 -10567 29660
rect -9773 30718 -9673 30731
rect -9773 30672 -9760 30718
rect -9686 30672 -9673 30718
rect -9773 30639 -9673 30672
rect -9569 30718 -9469 30731
rect -9569 30672 -9556 30718
rect -9482 30672 -9469 30718
rect -9569 30639 -9469 30672
rect -9773 30406 -9673 30439
rect -9773 30360 -9760 30406
rect -9686 30360 -9673 30406
rect -9773 30347 -9673 30360
rect -9569 30406 -9469 30439
rect -9569 30360 -9556 30406
rect -9482 30360 -9469 30406
rect -9569 30347 -9469 30360
rect -9089 30718 -8989 30731
rect -9089 30672 -9076 30718
rect -9002 30672 -8989 30718
rect -9089 30639 -8989 30672
rect -8885 30718 -8785 30731
rect -8885 30672 -8872 30718
rect -8798 30672 -8785 30718
rect -8885 30639 -8785 30672
rect -9089 30406 -8989 30439
rect -9089 30360 -9076 30406
rect -9002 30360 -8989 30406
rect -9089 30347 -8989 30360
rect -8885 30406 -8785 30439
rect -8885 30360 -8872 30406
rect -8798 30360 -8785 30406
rect -8885 30347 -8785 30360
rect -8405 30718 -8305 30731
rect -8405 30672 -8392 30718
rect -8318 30672 -8305 30718
rect -8405 30639 -8305 30672
rect -8405 30406 -8305 30439
rect -8405 30360 -8392 30406
rect -8318 30360 -8305 30406
rect -8405 30347 -8305 30360
rect -7545 30662 -7445 30675
rect -7545 30616 -7532 30662
rect -7458 30616 -7445 30662
rect -7545 30583 -7445 30616
rect -7341 30662 -7241 30675
rect -7341 30616 -7328 30662
rect -7254 30616 -7241 30662
rect -7341 30583 -7241 30616
rect -7545 29950 -7445 29983
rect -7545 29904 -7532 29950
rect -7458 29904 -7445 29950
rect -7545 29891 -7445 29904
rect -7341 29950 -7241 29983
rect -7341 29904 -7328 29950
rect -7254 29904 -7241 29950
rect -7341 29891 -7241 29904
rect -6861 30662 -6761 30675
rect -6861 30616 -6848 30662
rect -6774 30616 -6761 30662
rect -6861 30583 -6761 30616
rect -6657 30662 -6557 30675
rect -6657 30616 -6644 30662
rect -6570 30616 -6557 30662
rect -6657 30583 -6557 30616
rect -6861 29950 -6761 29983
rect -6861 29904 -6848 29950
rect -6774 29904 -6761 29950
rect -6861 29891 -6761 29904
rect -6657 29950 -6557 29983
rect -6657 29904 -6644 29950
rect -6570 29904 -6557 29950
rect -6657 29891 -6557 29904
rect -6177 30662 -6077 30675
rect -6177 30616 -6164 30662
rect -6090 30616 -6077 30662
rect -6177 30583 -6077 30616
rect -6177 29950 -6077 29983
rect -6177 29904 -6164 29950
rect -6090 29904 -6077 29950
rect -6177 29891 -6077 29904
rect -4631 30748 -4551 30761
rect -4631 30702 -4618 30748
rect -4564 30702 -4551 30748
rect -4631 30669 -4551 30702
rect -4447 30748 -4367 30761
rect -4447 30702 -4434 30748
rect -4380 30702 -4367 30748
rect -4447 30669 -4367 30702
rect -4263 30748 -4183 30761
rect -4263 30702 -4250 30748
rect -4196 30702 -4183 30748
rect -4263 30669 -4183 30702
rect -4631 30136 -4551 30169
rect -4631 30090 -4618 30136
rect -4564 30090 -4551 30136
rect -4631 30077 -4551 30090
rect -4447 30136 -4367 30169
rect -4447 30090 -4434 30136
rect -4380 30090 -4367 30136
rect -4447 30077 -4367 30090
rect -4263 30136 -4183 30169
rect -4263 30090 -4250 30136
rect -4196 30090 -4183 30136
rect -4263 30077 -4183 30090
rect -10667 29298 -10567 29311
rect -10667 29252 -10654 29298
rect -10580 29252 -10567 29298
rect -10667 29219 -10567 29252
rect -10667 28986 -10567 29019
rect -10667 28940 -10654 28986
rect -10580 28940 -10567 28986
rect -10667 28927 -10567 28940
rect -9773 29498 -9673 29511
rect -9773 29452 -9760 29498
rect -9686 29452 -9673 29498
rect -9773 29419 -9673 29452
rect -9773 28786 -9673 28819
rect -9773 28740 -9760 28786
rect -9686 28740 -9673 28786
rect -9773 28727 -9673 28740
rect -8885 29498 -8785 29511
rect -8885 29452 -8872 29498
rect -8798 29452 -8785 29498
rect -8885 29419 -8785 29452
rect -8885 28786 -8785 28819
rect -8885 28740 -8872 28786
rect -8798 28740 -8785 28786
rect -8885 28727 -8785 28740
rect -8405 29498 -8305 29511
rect -8405 29452 -8392 29498
rect -8318 29452 -8305 29498
rect -8405 29419 -8305 29452
rect -8405 28786 -8305 28819
rect -8405 28740 -8392 28786
rect -8318 28740 -8305 28786
rect -8405 28727 -8305 28740
rect -7545 29542 -7445 29555
rect -7545 29496 -7532 29542
rect -7458 29496 -7445 29542
rect -7545 29463 -7445 29496
rect -7545 29230 -7445 29263
rect -7545 29184 -7532 29230
rect -7458 29184 -7445 29230
rect -7545 29171 -7445 29184
rect -6861 29542 -6761 29555
rect -6861 29496 -6848 29542
rect -6774 29496 -6761 29542
rect -6861 29463 -6761 29496
rect -6861 29230 -6761 29263
rect -6861 29184 -6848 29230
rect -6774 29184 -6761 29230
rect -6861 29171 -6761 29184
rect -6177 29542 -6077 29555
rect -6177 29496 -6164 29542
rect -6090 29496 -6077 29542
rect -6177 29463 -6077 29496
rect -6177 29230 -6077 29263
rect -6177 29184 -6164 29230
rect -6090 29184 -6077 29230
rect -6177 29171 -6077 29184
rect -4631 29588 -4551 29601
rect -4631 29542 -4618 29588
rect -4564 29542 -4551 29588
rect -4631 29509 -4551 29542
rect -4447 29588 -4367 29601
rect -4447 29542 -4434 29588
rect -4380 29542 -4367 29588
rect -4447 29509 -4367 29542
rect -4263 29588 -4183 29601
rect -4263 29542 -4250 29588
rect -4196 29542 -4183 29588
rect -4263 29509 -4183 29542
rect -4631 29276 -4551 29309
rect -4631 29230 -4618 29276
rect -4564 29230 -4551 29276
rect -4631 29217 -4551 29230
rect -4447 29276 -4367 29309
rect -4447 29230 -4434 29276
rect -4380 29230 -4367 29276
rect -4447 29217 -4367 29230
rect -4263 29276 -4183 29309
rect -4263 29230 -4250 29276
rect -4196 29230 -4183 29276
rect -4263 29217 -4183 29230
rect -1195 30418 -1095 30431
rect -1195 30372 -1182 30418
rect -1108 30372 -1095 30418
rect -1195 30339 -1095 30372
rect -1195 29706 -1095 29739
rect -1195 29660 -1182 29706
rect -1108 29660 -1095 29706
rect -1195 29647 -1095 29660
rect -301 30718 -201 30731
rect -301 30672 -288 30718
rect -214 30672 -201 30718
rect -301 30639 -201 30672
rect -97 30718 3 30731
rect -97 30672 -84 30718
rect -10 30672 3 30718
rect -97 30639 3 30672
rect -301 30406 -201 30439
rect -301 30360 -288 30406
rect -214 30360 -201 30406
rect -301 30347 -201 30360
rect -97 30406 3 30439
rect -97 30360 -84 30406
rect -10 30360 3 30406
rect -97 30347 3 30360
rect 383 30718 483 30731
rect 383 30672 396 30718
rect 470 30672 483 30718
rect 383 30639 483 30672
rect 587 30718 687 30731
rect 587 30672 600 30718
rect 674 30672 687 30718
rect 587 30639 687 30672
rect 383 30406 483 30439
rect 383 30360 396 30406
rect 470 30360 483 30406
rect 383 30347 483 30360
rect 587 30406 687 30439
rect 587 30360 600 30406
rect 674 30360 687 30406
rect 587 30347 687 30360
rect 1067 30718 1167 30731
rect 1067 30672 1080 30718
rect 1154 30672 1167 30718
rect 1067 30639 1167 30672
rect 1067 30406 1167 30439
rect 1067 30360 1080 30406
rect 1154 30360 1167 30406
rect 1067 30347 1167 30360
rect 1927 30662 2027 30675
rect 1927 30616 1940 30662
rect 2014 30616 2027 30662
rect 1927 30583 2027 30616
rect 2131 30662 2231 30675
rect 2131 30616 2144 30662
rect 2218 30616 2231 30662
rect 2131 30583 2231 30616
rect 1927 29950 2027 29983
rect 1927 29904 1940 29950
rect 2014 29904 2027 29950
rect 1927 29891 2027 29904
rect 2131 29950 2231 29983
rect 2131 29904 2144 29950
rect 2218 29904 2231 29950
rect 2131 29891 2231 29904
rect 2611 30662 2711 30675
rect 2611 30616 2624 30662
rect 2698 30616 2711 30662
rect 2611 30583 2711 30616
rect 2815 30662 2915 30675
rect 2815 30616 2828 30662
rect 2902 30616 2915 30662
rect 2815 30583 2915 30616
rect 2611 29950 2711 29983
rect 2611 29904 2624 29950
rect 2698 29904 2711 29950
rect 2611 29891 2711 29904
rect 2815 29950 2915 29983
rect 2815 29904 2828 29950
rect 2902 29904 2915 29950
rect 2815 29891 2915 29904
rect 3295 30662 3395 30675
rect 3295 30616 3308 30662
rect 3382 30616 3395 30662
rect 3295 30583 3395 30616
rect 3295 29950 3395 29983
rect 3295 29904 3308 29950
rect 3382 29904 3395 29950
rect 3295 29891 3395 29904
rect 4841 30748 4921 30761
rect 4841 30702 4854 30748
rect 4908 30702 4921 30748
rect 4841 30669 4921 30702
rect 5025 30748 5105 30761
rect 5025 30702 5038 30748
rect 5092 30702 5105 30748
rect 5025 30669 5105 30702
rect 5209 30748 5289 30761
rect 5209 30702 5222 30748
rect 5276 30702 5289 30748
rect 5209 30669 5289 30702
rect 4841 30136 4921 30169
rect 4841 30090 4854 30136
rect 4908 30090 4921 30136
rect 4841 30077 4921 30090
rect 5025 30136 5105 30169
rect 5025 30090 5038 30136
rect 5092 30090 5105 30136
rect 5025 30077 5105 30090
rect 5209 30136 5289 30169
rect 5209 30090 5222 30136
rect 5276 30090 5289 30136
rect 5209 30077 5289 30090
rect -1195 29298 -1095 29311
rect -1195 29252 -1182 29298
rect -1108 29252 -1095 29298
rect -1195 29219 -1095 29252
rect -1195 28986 -1095 29019
rect -1195 28940 -1182 28986
rect -1108 28940 -1095 28986
rect -1195 28927 -1095 28940
rect -301 29498 -201 29511
rect -301 29452 -288 29498
rect -214 29452 -201 29498
rect -301 29419 -201 29452
rect -301 28786 -201 28819
rect -301 28740 -288 28786
rect -214 28740 -201 28786
rect -301 28727 -201 28740
rect 587 29498 687 29511
rect 587 29452 600 29498
rect 674 29452 687 29498
rect 587 29419 687 29452
rect 587 28786 687 28819
rect 587 28740 600 28786
rect 674 28740 687 28786
rect 587 28727 687 28740
rect 1067 29498 1167 29511
rect 1067 29452 1080 29498
rect 1154 29452 1167 29498
rect 1067 29419 1167 29452
rect 1067 28786 1167 28819
rect 1067 28740 1080 28786
rect 1154 28740 1167 28786
rect 1067 28727 1167 28740
rect 1927 29542 2027 29555
rect 1927 29496 1940 29542
rect 2014 29496 2027 29542
rect 1927 29463 2027 29496
rect 1927 29230 2027 29263
rect 1927 29184 1940 29230
rect 2014 29184 2027 29230
rect 1927 29171 2027 29184
rect 2611 29542 2711 29555
rect 2611 29496 2624 29542
rect 2698 29496 2711 29542
rect 2611 29463 2711 29496
rect 2611 29230 2711 29263
rect 2611 29184 2624 29230
rect 2698 29184 2711 29230
rect 2611 29171 2711 29184
rect 3295 29542 3395 29555
rect 3295 29496 3308 29542
rect 3382 29496 3395 29542
rect 3295 29463 3395 29496
rect 3295 29230 3395 29263
rect 3295 29184 3308 29230
rect 3382 29184 3395 29230
rect 3295 29171 3395 29184
rect 4841 29588 4921 29601
rect 4841 29542 4854 29588
rect 4908 29542 4921 29588
rect 4841 29509 4921 29542
rect 5025 29588 5105 29601
rect 5025 29542 5038 29588
rect 5092 29542 5105 29588
rect 5025 29509 5105 29542
rect 5209 29588 5289 29601
rect 5209 29542 5222 29588
rect 5276 29542 5289 29588
rect 5209 29509 5289 29542
rect 4841 29276 4921 29309
rect 4841 29230 4854 29276
rect 4908 29230 4921 29276
rect 4841 29217 4921 29230
rect 5025 29276 5105 29309
rect 5025 29230 5038 29276
rect 5092 29230 5105 29276
rect 5025 29217 5105 29230
rect 5209 29276 5289 29309
rect 5209 29230 5222 29276
rect 5276 29230 5289 29276
rect 5209 29217 5289 29230
rect 8277 30419 8377 30432
rect 8277 30373 8290 30419
rect 8364 30373 8377 30419
rect 8277 30340 8377 30373
rect 8277 29707 8377 29740
rect 8277 29661 8290 29707
rect 8364 29661 8377 29707
rect 8277 29648 8377 29661
rect 9171 30719 9271 30732
rect 9171 30673 9184 30719
rect 9258 30673 9271 30719
rect 9171 30640 9271 30673
rect 9375 30719 9475 30732
rect 9375 30673 9388 30719
rect 9462 30673 9475 30719
rect 9375 30640 9475 30673
rect 9171 30407 9271 30440
rect 9171 30361 9184 30407
rect 9258 30361 9271 30407
rect 9171 30348 9271 30361
rect 9375 30407 9475 30440
rect 9375 30361 9388 30407
rect 9462 30361 9475 30407
rect 9375 30348 9475 30361
rect 9855 30719 9955 30732
rect 9855 30673 9868 30719
rect 9942 30673 9955 30719
rect 9855 30640 9955 30673
rect 10059 30719 10159 30732
rect 10059 30673 10072 30719
rect 10146 30673 10159 30719
rect 10059 30640 10159 30673
rect 9855 30407 9955 30440
rect 9855 30361 9868 30407
rect 9942 30361 9955 30407
rect 9855 30348 9955 30361
rect 10059 30407 10159 30440
rect 10059 30361 10072 30407
rect 10146 30361 10159 30407
rect 10059 30348 10159 30361
rect 10539 30719 10639 30732
rect 10539 30673 10552 30719
rect 10626 30673 10639 30719
rect 10539 30640 10639 30673
rect 10539 30407 10639 30440
rect 10539 30361 10552 30407
rect 10626 30361 10639 30407
rect 10539 30348 10639 30361
rect 11399 30663 11499 30676
rect 11399 30617 11412 30663
rect 11486 30617 11499 30663
rect 11399 30584 11499 30617
rect 11603 30663 11703 30676
rect 11603 30617 11616 30663
rect 11690 30617 11703 30663
rect 11603 30584 11703 30617
rect 11399 29951 11499 29984
rect 11399 29905 11412 29951
rect 11486 29905 11499 29951
rect 11399 29892 11499 29905
rect 11603 29951 11703 29984
rect 11603 29905 11616 29951
rect 11690 29905 11703 29951
rect 11603 29892 11703 29905
rect 12083 30663 12183 30676
rect 12083 30617 12096 30663
rect 12170 30617 12183 30663
rect 12083 30584 12183 30617
rect 12287 30663 12387 30676
rect 12287 30617 12300 30663
rect 12374 30617 12387 30663
rect 12287 30584 12387 30617
rect 12083 29951 12183 29984
rect 12083 29905 12096 29951
rect 12170 29905 12183 29951
rect 12083 29892 12183 29905
rect 12287 29951 12387 29984
rect 12287 29905 12300 29951
rect 12374 29905 12387 29951
rect 12287 29892 12387 29905
rect 12767 30663 12867 30676
rect 12767 30617 12780 30663
rect 12854 30617 12867 30663
rect 12767 30584 12867 30617
rect 12767 29951 12867 29984
rect 12767 29905 12780 29951
rect 12854 29905 12867 29951
rect 12767 29892 12867 29905
rect 14313 30749 14393 30762
rect 14313 30703 14326 30749
rect 14380 30703 14393 30749
rect 14313 30670 14393 30703
rect 14497 30749 14577 30762
rect 14497 30703 14510 30749
rect 14564 30703 14577 30749
rect 14497 30670 14577 30703
rect 14681 30749 14761 30762
rect 14681 30703 14694 30749
rect 14748 30703 14761 30749
rect 14681 30670 14761 30703
rect 14313 30137 14393 30170
rect 14313 30091 14326 30137
rect 14380 30091 14393 30137
rect 14313 30078 14393 30091
rect 14497 30137 14577 30170
rect 14497 30091 14510 30137
rect 14564 30091 14577 30137
rect 14497 30078 14577 30091
rect 14681 30137 14761 30170
rect 14681 30091 14694 30137
rect 14748 30091 14761 30137
rect 14681 30078 14761 30091
rect 8277 29299 8377 29312
rect 8277 29253 8290 29299
rect 8364 29253 8377 29299
rect 8277 29220 8377 29253
rect 8277 28987 8377 29020
rect 8277 28941 8290 28987
rect 8364 28941 8377 28987
rect 8277 28928 8377 28941
rect 9171 29499 9271 29512
rect 9171 29453 9184 29499
rect 9258 29453 9271 29499
rect 9171 29420 9271 29453
rect 9171 28787 9271 28820
rect 9171 28741 9184 28787
rect 9258 28741 9271 28787
rect 9171 28728 9271 28741
rect 10059 29499 10159 29512
rect 10059 29453 10072 29499
rect 10146 29453 10159 29499
rect 10059 29420 10159 29453
rect 10059 28787 10159 28820
rect 10059 28741 10072 28787
rect 10146 28741 10159 28787
rect 10059 28728 10159 28741
rect 10539 29499 10639 29512
rect 10539 29453 10552 29499
rect 10626 29453 10639 29499
rect 10539 29420 10639 29453
rect 10539 28787 10639 28820
rect 10539 28741 10552 28787
rect 10626 28741 10639 28787
rect 10539 28728 10639 28741
rect 11399 29543 11499 29556
rect 11399 29497 11412 29543
rect 11486 29497 11499 29543
rect 11399 29464 11499 29497
rect 11399 29231 11499 29264
rect 11399 29185 11412 29231
rect 11486 29185 11499 29231
rect 11399 29172 11499 29185
rect 12083 29543 12183 29556
rect 12083 29497 12096 29543
rect 12170 29497 12183 29543
rect 12083 29464 12183 29497
rect 12083 29231 12183 29264
rect 12083 29185 12096 29231
rect 12170 29185 12183 29231
rect 12083 29172 12183 29185
rect 12767 29543 12867 29556
rect 12767 29497 12780 29543
rect 12854 29497 12867 29543
rect 12767 29464 12867 29497
rect 12767 29231 12867 29264
rect 12767 29185 12780 29231
rect 12854 29185 12867 29231
rect 12767 29172 12867 29185
rect 14313 29589 14393 29602
rect 14313 29543 14326 29589
rect 14380 29543 14393 29589
rect 14313 29510 14393 29543
rect 14497 29589 14577 29602
rect 14497 29543 14510 29589
rect 14564 29543 14577 29589
rect 14497 29510 14577 29543
rect 14681 29589 14761 29602
rect 14681 29543 14694 29589
rect 14748 29543 14761 29589
rect 14681 29510 14761 29543
rect 14313 29277 14393 29310
rect 14313 29231 14326 29277
rect 14380 29231 14393 29277
rect 14313 29218 14393 29231
rect 14497 29277 14577 29310
rect 14497 29231 14510 29277
rect 14564 29231 14577 29277
rect 14497 29218 14577 29231
rect 14681 29277 14761 29310
rect 14681 29231 14694 29277
rect 14748 29231 14761 29277
rect 14681 29218 14761 29231
rect 17749 30419 17849 30432
rect 17749 30373 17762 30419
rect 17836 30373 17849 30419
rect 17749 30340 17849 30373
rect 17749 29707 17849 29740
rect 17749 29661 17762 29707
rect 17836 29661 17849 29707
rect 17749 29648 17849 29661
rect 18643 30719 18743 30732
rect 18643 30673 18656 30719
rect 18730 30673 18743 30719
rect 18643 30640 18743 30673
rect 18847 30719 18947 30732
rect 18847 30673 18860 30719
rect 18934 30673 18947 30719
rect 18847 30640 18947 30673
rect 18643 30407 18743 30440
rect 18643 30361 18656 30407
rect 18730 30361 18743 30407
rect 18643 30348 18743 30361
rect 18847 30407 18947 30440
rect 18847 30361 18860 30407
rect 18934 30361 18947 30407
rect 18847 30348 18947 30361
rect 19327 30719 19427 30732
rect 19327 30673 19340 30719
rect 19414 30673 19427 30719
rect 19327 30640 19427 30673
rect 19531 30719 19631 30732
rect 19531 30673 19544 30719
rect 19618 30673 19631 30719
rect 19531 30640 19631 30673
rect 19327 30407 19427 30440
rect 19327 30361 19340 30407
rect 19414 30361 19427 30407
rect 19327 30348 19427 30361
rect 19531 30407 19631 30440
rect 19531 30361 19544 30407
rect 19618 30361 19631 30407
rect 19531 30348 19631 30361
rect 20011 30719 20111 30732
rect 20011 30673 20024 30719
rect 20098 30673 20111 30719
rect 20011 30640 20111 30673
rect 20011 30407 20111 30440
rect 20011 30361 20024 30407
rect 20098 30361 20111 30407
rect 20011 30348 20111 30361
rect 20871 30663 20971 30676
rect 20871 30617 20884 30663
rect 20958 30617 20971 30663
rect 20871 30584 20971 30617
rect 21075 30663 21175 30676
rect 21075 30617 21088 30663
rect 21162 30617 21175 30663
rect 21075 30584 21175 30617
rect 20871 29951 20971 29984
rect 20871 29905 20884 29951
rect 20958 29905 20971 29951
rect 20871 29892 20971 29905
rect 21075 29951 21175 29984
rect 21075 29905 21088 29951
rect 21162 29905 21175 29951
rect 21075 29892 21175 29905
rect 21555 30663 21655 30676
rect 21555 30617 21568 30663
rect 21642 30617 21655 30663
rect 21555 30584 21655 30617
rect 21759 30663 21859 30676
rect 21759 30617 21772 30663
rect 21846 30617 21859 30663
rect 21759 30584 21859 30617
rect 21555 29951 21655 29984
rect 21555 29905 21568 29951
rect 21642 29905 21655 29951
rect 21555 29892 21655 29905
rect 21759 29951 21859 29984
rect 21759 29905 21772 29951
rect 21846 29905 21859 29951
rect 21759 29892 21859 29905
rect 22239 30663 22339 30676
rect 22239 30617 22252 30663
rect 22326 30617 22339 30663
rect 22239 30584 22339 30617
rect 22239 29951 22339 29984
rect 22239 29905 22252 29951
rect 22326 29905 22339 29951
rect 22239 29892 22339 29905
rect 23785 30749 23865 30762
rect 23785 30703 23798 30749
rect 23852 30703 23865 30749
rect 23785 30670 23865 30703
rect 23969 30749 24049 30762
rect 23969 30703 23982 30749
rect 24036 30703 24049 30749
rect 23969 30670 24049 30703
rect 24153 30749 24233 30762
rect 24153 30703 24166 30749
rect 24220 30703 24233 30749
rect 24153 30670 24233 30703
rect 23785 30137 23865 30170
rect 23785 30091 23798 30137
rect 23852 30091 23865 30137
rect 23785 30078 23865 30091
rect 23969 30137 24049 30170
rect 23969 30091 23982 30137
rect 24036 30091 24049 30137
rect 23969 30078 24049 30091
rect 24153 30137 24233 30170
rect 24153 30091 24166 30137
rect 24220 30091 24233 30137
rect 24153 30078 24233 30091
rect 17749 29299 17849 29312
rect 17749 29253 17762 29299
rect 17836 29253 17849 29299
rect 17749 29220 17849 29253
rect 17749 28987 17849 29020
rect 17749 28941 17762 28987
rect 17836 28941 17849 28987
rect 17749 28928 17849 28941
rect 18643 29499 18743 29512
rect 18643 29453 18656 29499
rect 18730 29453 18743 29499
rect 18643 29420 18743 29453
rect 18643 28787 18743 28820
rect 18643 28741 18656 28787
rect 18730 28741 18743 28787
rect 18643 28728 18743 28741
rect 19531 29499 19631 29512
rect 19531 29453 19544 29499
rect 19618 29453 19631 29499
rect 19531 29420 19631 29453
rect 19531 28787 19631 28820
rect 19531 28741 19544 28787
rect 19618 28741 19631 28787
rect 19531 28728 19631 28741
rect 20011 29499 20111 29512
rect 20011 29453 20024 29499
rect 20098 29453 20111 29499
rect 20011 29420 20111 29453
rect 20011 28787 20111 28820
rect 20011 28741 20024 28787
rect 20098 28741 20111 28787
rect 20011 28728 20111 28741
rect 20871 29543 20971 29556
rect 20871 29497 20884 29543
rect 20958 29497 20971 29543
rect 20871 29464 20971 29497
rect 20871 29231 20971 29264
rect 20871 29185 20884 29231
rect 20958 29185 20971 29231
rect 20871 29172 20971 29185
rect 21555 29543 21655 29556
rect 21555 29497 21568 29543
rect 21642 29497 21655 29543
rect 21555 29464 21655 29497
rect 21555 29231 21655 29264
rect 21555 29185 21568 29231
rect 21642 29185 21655 29231
rect 21555 29172 21655 29185
rect 22239 29543 22339 29556
rect 22239 29497 22252 29543
rect 22326 29497 22339 29543
rect 22239 29464 22339 29497
rect 22239 29231 22339 29264
rect 22239 29185 22252 29231
rect 22326 29185 22339 29231
rect 22239 29172 22339 29185
rect 23785 29589 23865 29602
rect 23785 29543 23798 29589
rect 23852 29543 23865 29589
rect 23785 29510 23865 29543
rect 23969 29589 24049 29602
rect 23969 29543 23982 29589
rect 24036 29543 24049 29589
rect 23969 29510 24049 29543
rect 24153 29589 24233 29602
rect 24153 29543 24166 29589
rect 24220 29543 24233 29589
rect 24153 29510 24233 29543
rect 23785 29277 23865 29310
rect 23785 29231 23798 29277
rect 23852 29231 23865 29277
rect 23785 29218 23865 29231
rect 23969 29277 24049 29310
rect 23969 29231 23982 29277
rect 24036 29231 24049 29277
rect 23969 29218 24049 29231
rect 24153 29277 24233 29310
rect 24153 29231 24166 29277
rect 24220 29231 24233 29277
rect 24153 29218 24233 29231
rect 27221 30419 27321 30432
rect 27221 30373 27234 30419
rect 27308 30373 27321 30419
rect 27221 30340 27321 30373
rect 27221 29707 27321 29740
rect 27221 29661 27234 29707
rect 27308 29661 27321 29707
rect 27221 29648 27321 29661
rect 28115 30719 28215 30732
rect 28115 30673 28128 30719
rect 28202 30673 28215 30719
rect 28115 30640 28215 30673
rect 28319 30719 28419 30732
rect 28319 30673 28332 30719
rect 28406 30673 28419 30719
rect 28319 30640 28419 30673
rect 28115 30407 28215 30440
rect 28115 30361 28128 30407
rect 28202 30361 28215 30407
rect 28115 30348 28215 30361
rect 28319 30407 28419 30440
rect 28319 30361 28332 30407
rect 28406 30361 28419 30407
rect 28319 30348 28419 30361
rect 28799 30719 28899 30732
rect 28799 30673 28812 30719
rect 28886 30673 28899 30719
rect 28799 30640 28899 30673
rect 29003 30719 29103 30732
rect 29003 30673 29016 30719
rect 29090 30673 29103 30719
rect 29003 30640 29103 30673
rect 28799 30407 28899 30440
rect 28799 30361 28812 30407
rect 28886 30361 28899 30407
rect 28799 30348 28899 30361
rect 29003 30407 29103 30440
rect 29003 30361 29016 30407
rect 29090 30361 29103 30407
rect 29003 30348 29103 30361
rect 29483 30719 29583 30732
rect 29483 30673 29496 30719
rect 29570 30673 29583 30719
rect 29483 30640 29583 30673
rect 29483 30407 29583 30440
rect 29483 30361 29496 30407
rect 29570 30361 29583 30407
rect 29483 30348 29583 30361
rect 30343 30663 30443 30676
rect 30343 30617 30356 30663
rect 30430 30617 30443 30663
rect 30343 30584 30443 30617
rect 30547 30663 30647 30676
rect 30547 30617 30560 30663
rect 30634 30617 30647 30663
rect 30547 30584 30647 30617
rect 30343 29951 30443 29984
rect 30343 29905 30356 29951
rect 30430 29905 30443 29951
rect 30343 29892 30443 29905
rect 30547 29951 30647 29984
rect 30547 29905 30560 29951
rect 30634 29905 30647 29951
rect 30547 29892 30647 29905
rect 31027 30663 31127 30676
rect 31027 30617 31040 30663
rect 31114 30617 31127 30663
rect 31027 30584 31127 30617
rect 31231 30663 31331 30676
rect 31231 30617 31244 30663
rect 31318 30617 31331 30663
rect 31231 30584 31331 30617
rect 31027 29951 31127 29984
rect 31027 29905 31040 29951
rect 31114 29905 31127 29951
rect 31027 29892 31127 29905
rect 31231 29951 31331 29984
rect 31231 29905 31244 29951
rect 31318 29905 31331 29951
rect 31231 29892 31331 29905
rect 31711 30663 31811 30676
rect 31711 30617 31724 30663
rect 31798 30617 31811 30663
rect 31711 30584 31811 30617
rect 31711 29951 31811 29984
rect 31711 29905 31724 29951
rect 31798 29905 31811 29951
rect 31711 29892 31811 29905
rect 33257 30749 33337 30762
rect 33257 30703 33270 30749
rect 33324 30703 33337 30749
rect 33257 30670 33337 30703
rect 33441 30749 33521 30762
rect 33441 30703 33454 30749
rect 33508 30703 33521 30749
rect 33441 30670 33521 30703
rect 33625 30749 33705 30762
rect 33625 30703 33638 30749
rect 33692 30703 33705 30749
rect 33625 30670 33705 30703
rect 33257 30137 33337 30170
rect 33257 30091 33270 30137
rect 33324 30091 33337 30137
rect 33257 30078 33337 30091
rect 33441 30137 33521 30170
rect 33441 30091 33454 30137
rect 33508 30091 33521 30137
rect 33441 30078 33521 30091
rect 33625 30137 33705 30170
rect 33625 30091 33638 30137
rect 33692 30091 33705 30137
rect 33625 30078 33705 30091
rect 27221 29299 27321 29312
rect 27221 29253 27234 29299
rect 27308 29253 27321 29299
rect 27221 29220 27321 29253
rect 27221 28987 27321 29020
rect 27221 28941 27234 28987
rect 27308 28941 27321 28987
rect 27221 28928 27321 28941
rect 28115 29499 28215 29512
rect 28115 29453 28128 29499
rect 28202 29453 28215 29499
rect 28115 29420 28215 29453
rect 28115 28787 28215 28820
rect 28115 28741 28128 28787
rect 28202 28741 28215 28787
rect 28115 28728 28215 28741
rect 29003 29499 29103 29512
rect 29003 29453 29016 29499
rect 29090 29453 29103 29499
rect 29003 29420 29103 29453
rect 29003 28787 29103 28820
rect 29003 28741 29016 28787
rect 29090 28741 29103 28787
rect 29003 28728 29103 28741
rect 29483 29499 29583 29512
rect 29483 29453 29496 29499
rect 29570 29453 29583 29499
rect 29483 29420 29583 29453
rect 29483 28787 29583 28820
rect 29483 28741 29496 28787
rect 29570 28741 29583 28787
rect 29483 28728 29583 28741
rect 30343 29543 30443 29556
rect 30343 29497 30356 29543
rect 30430 29497 30443 29543
rect 30343 29464 30443 29497
rect 30343 29231 30443 29264
rect 30343 29185 30356 29231
rect 30430 29185 30443 29231
rect 30343 29172 30443 29185
rect 31027 29543 31127 29556
rect 31027 29497 31040 29543
rect 31114 29497 31127 29543
rect 31027 29464 31127 29497
rect 31027 29231 31127 29264
rect 31027 29185 31040 29231
rect 31114 29185 31127 29231
rect 31027 29172 31127 29185
rect 31711 29543 31811 29556
rect 31711 29497 31724 29543
rect 31798 29497 31811 29543
rect 31711 29464 31811 29497
rect 31711 29231 31811 29264
rect 31711 29185 31724 29231
rect 31798 29185 31811 29231
rect 31711 29172 31811 29185
rect 33257 29589 33337 29602
rect 33257 29543 33270 29589
rect 33324 29543 33337 29589
rect 33257 29510 33337 29543
rect 33441 29589 33521 29602
rect 33441 29543 33454 29589
rect 33508 29543 33521 29589
rect 33441 29510 33521 29543
rect 33625 29589 33705 29602
rect 33625 29543 33638 29589
rect 33692 29543 33705 29589
rect 33625 29510 33705 29543
rect 33257 29277 33337 29310
rect 33257 29231 33270 29277
rect 33324 29231 33337 29277
rect 33257 29218 33337 29231
rect 33441 29277 33521 29310
rect 33441 29231 33454 29277
rect 33508 29231 33521 29277
rect 33441 29218 33521 29231
rect 33625 29277 33705 29310
rect 33625 29231 33638 29277
rect 33692 29231 33705 29277
rect 33625 29218 33705 29231
rect 36693 30419 36793 30432
rect 36693 30373 36706 30419
rect 36780 30373 36793 30419
rect 36693 30340 36793 30373
rect 36693 29707 36793 29740
rect 36693 29661 36706 29707
rect 36780 29661 36793 29707
rect 36693 29648 36793 29661
rect 37587 30719 37687 30732
rect 37587 30673 37600 30719
rect 37674 30673 37687 30719
rect 37587 30640 37687 30673
rect 37791 30719 37891 30732
rect 37791 30673 37804 30719
rect 37878 30673 37891 30719
rect 37791 30640 37891 30673
rect 37587 30407 37687 30440
rect 37587 30361 37600 30407
rect 37674 30361 37687 30407
rect 37587 30348 37687 30361
rect 37791 30407 37891 30440
rect 37791 30361 37804 30407
rect 37878 30361 37891 30407
rect 37791 30348 37891 30361
rect 38271 30719 38371 30732
rect 38271 30673 38284 30719
rect 38358 30673 38371 30719
rect 38271 30640 38371 30673
rect 38475 30719 38575 30732
rect 38475 30673 38488 30719
rect 38562 30673 38575 30719
rect 38475 30640 38575 30673
rect 38271 30407 38371 30440
rect 38271 30361 38284 30407
rect 38358 30361 38371 30407
rect 38271 30348 38371 30361
rect 38475 30407 38575 30440
rect 38475 30361 38488 30407
rect 38562 30361 38575 30407
rect 38475 30348 38575 30361
rect 38955 30719 39055 30732
rect 38955 30673 38968 30719
rect 39042 30673 39055 30719
rect 38955 30640 39055 30673
rect 38955 30407 39055 30440
rect 38955 30361 38968 30407
rect 39042 30361 39055 30407
rect 38955 30348 39055 30361
rect 39815 30663 39915 30676
rect 39815 30617 39828 30663
rect 39902 30617 39915 30663
rect 39815 30584 39915 30617
rect 40019 30663 40119 30676
rect 40019 30617 40032 30663
rect 40106 30617 40119 30663
rect 40019 30584 40119 30617
rect 39815 29951 39915 29984
rect 39815 29905 39828 29951
rect 39902 29905 39915 29951
rect 39815 29892 39915 29905
rect 40019 29951 40119 29984
rect 40019 29905 40032 29951
rect 40106 29905 40119 29951
rect 40019 29892 40119 29905
rect 40499 30663 40599 30676
rect 40499 30617 40512 30663
rect 40586 30617 40599 30663
rect 40499 30584 40599 30617
rect 40703 30663 40803 30676
rect 40703 30617 40716 30663
rect 40790 30617 40803 30663
rect 40703 30584 40803 30617
rect 40499 29951 40599 29984
rect 40499 29905 40512 29951
rect 40586 29905 40599 29951
rect 40499 29892 40599 29905
rect 40703 29951 40803 29984
rect 40703 29905 40716 29951
rect 40790 29905 40803 29951
rect 40703 29892 40803 29905
rect 41183 30663 41283 30676
rect 41183 30617 41196 30663
rect 41270 30617 41283 30663
rect 41183 30584 41283 30617
rect 41183 29951 41283 29984
rect 41183 29905 41196 29951
rect 41270 29905 41283 29951
rect 41183 29892 41283 29905
rect 42729 30749 42809 30762
rect 42729 30703 42742 30749
rect 42796 30703 42809 30749
rect 42729 30670 42809 30703
rect 42913 30749 42993 30762
rect 42913 30703 42926 30749
rect 42980 30703 42993 30749
rect 42913 30670 42993 30703
rect 43097 30749 43177 30762
rect 43097 30703 43110 30749
rect 43164 30703 43177 30749
rect 43097 30670 43177 30703
rect 42729 30137 42809 30170
rect 42729 30091 42742 30137
rect 42796 30091 42809 30137
rect 42729 30078 42809 30091
rect 42913 30137 42993 30170
rect 42913 30091 42926 30137
rect 42980 30091 42993 30137
rect 42913 30078 42993 30091
rect 43097 30137 43177 30170
rect 43097 30091 43110 30137
rect 43164 30091 43177 30137
rect 43097 30078 43177 30091
rect 36693 29299 36793 29312
rect 36693 29253 36706 29299
rect 36780 29253 36793 29299
rect 36693 29220 36793 29253
rect 36693 28987 36793 29020
rect 36693 28941 36706 28987
rect 36780 28941 36793 28987
rect 36693 28928 36793 28941
rect 37587 29499 37687 29512
rect 37587 29453 37600 29499
rect 37674 29453 37687 29499
rect 37587 29420 37687 29453
rect 37587 28787 37687 28820
rect 37587 28741 37600 28787
rect 37674 28741 37687 28787
rect 37587 28728 37687 28741
rect 38475 29499 38575 29512
rect 38475 29453 38488 29499
rect 38562 29453 38575 29499
rect 38475 29420 38575 29453
rect 38475 28787 38575 28820
rect 38475 28741 38488 28787
rect 38562 28741 38575 28787
rect 38475 28728 38575 28741
rect 38955 29499 39055 29512
rect 38955 29453 38968 29499
rect 39042 29453 39055 29499
rect 38955 29420 39055 29453
rect 38955 28787 39055 28820
rect 38955 28741 38968 28787
rect 39042 28741 39055 28787
rect 38955 28728 39055 28741
rect 39815 29543 39915 29556
rect 39815 29497 39828 29543
rect 39902 29497 39915 29543
rect 39815 29464 39915 29497
rect 39815 29231 39915 29264
rect 39815 29185 39828 29231
rect 39902 29185 39915 29231
rect 39815 29172 39915 29185
rect 40499 29543 40599 29556
rect 40499 29497 40512 29543
rect 40586 29497 40599 29543
rect 40499 29464 40599 29497
rect 40499 29231 40599 29264
rect 40499 29185 40512 29231
rect 40586 29185 40599 29231
rect 40499 29172 40599 29185
rect 41183 29543 41283 29556
rect 41183 29497 41196 29543
rect 41270 29497 41283 29543
rect 41183 29464 41283 29497
rect 41183 29231 41283 29264
rect 41183 29185 41196 29231
rect 41270 29185 41283 29231
rect 41183 29172 41283 29185
rect 42729 29589 42809 29602
rect 42729 29543 42742 29589
rect 42796 29543 42809 29589
rect 42729 29510 42809 29543
rect 42913 29589 42993 29602
rect 42913 29543 42926 29589
rect 42980 29543 42993 29589
rect 42913 29510 42993 29543
rect 43097 29589 43177 29602
rect 43097 29543 43110 29589
rect 43164 29543 43177 29589
rect 43097 29510 43177 29543
rect 42729 29277 42809 29310
rect 42729 29231 42742 29277
rect 42796 29231 42809 29277
rect 42729 29218 42809 29231
rect 42913 29277 42993 29310
rect 42913 29231 42926 29277
rect 42980 29231 42993 29277
rect 42913 29218 42993 29231
rect 43097 29277 43177 29310
rect 43097 29231 43110 29277
rect 43164 29231 43177 29277
rect 43097 29218 43177 29231
rect -12380 28488 -12280 28501
rect -12380 28442 -12367 28488
rect -12293 28442 -12280 28488
rect -12380 28409 -12280 28442
rect -12380 27776 -12280 27809
rect -12380 27730 -12367 27776
rect -12293 27730 -12280 27776
rect -12380 27717 -12280 27730
rect -9773 28378 -9673 28391
rect -9773 28332 -9760 28378
rect -9686 28332 -9673 28378
rect -9773 28299 -9673 28332
rect -9569 28378 -9469 28391
rect -9569 28332 -9556 28378
rect -9482 28332 -9469 28378
rect -9569 28299 -9469 28332
rect -9773 28066 -9673 28099
rect -9773 28020 -9760 28066
rect -9686 28020 -9673 28066
rect -9773 28007 -9673 28020
rect -9569 28066 -9469 28099
rect -9569 28020 -9556 28066
rect -9482 28020 -9469 28066
rect -9569 28007 -9469 28020
rect -9089 28378 -8989 28391
rect -9089 28332 -9076 28378
rect -9002 28332 -8989 28378
rect -9089 28299 -8989 28332
rect -8885 28378 -8785 28391
rect -8885 28332 -8872 28378
rect -8798 28332 -8785 28378
rect -8885 28299 -8785 28332
rect -9089 28066 -8989 28099
rect -9089 28020 -9076 28066
rect -9002 28020 -8989 28066
rect -9089 28007 -8989 28020
rect -8885 28066 -8785 28099
rect -8885 28020 -8872 28066
rect -8798 28020 -8785 28066
rect -8885 28007 -8785 28020
rect -8405 28378 -8305 28391
rect -8405 28332 -8392 28378
rect -8318 28332 -8305 28378
rect -8405 28299 -8305 28332
rect -8405 28066 -8305 28099
rect -8405 28020 -8392 28066
rect -8318 28020 -8305 28066
rect -8405 28007 -8305 28020
rect -301 28378 -201 28391
rect -301 28332 -288 28378
rect -214 28332 -201 28378
rect -301 28299 -201 28332
rect -97 28378 3 28391
rect -97 28332 -84 28378
rect -10 28332 3 28378
rect -97 28299 3 28332
rect -301 28066 -201 28099
rect -301 28020 -288 28066
rect -214 28020 -201 28066
rect -301 28007 -201 28020
rect -97 28066 3 28099
rect -97 28020 -84 28066
rect -10 28020 3 28066
rect -97 28007 3 28020
rect 383 28378 483 28391
rect 383 28332 396 28378
rect 470 28332 483 28378
rect 383 28299 483 28332
rect 587 28378 687 28391
rect 587 28332 600 28378
rect 674 28332 687 28378
rect 587 28299 687 28332
rect 383 28066 483 28099
rect 383 28020 396 28066
rect 470 28020 483 28066
rect 383 28007 483 28020
rect 587 28066 687 28099
rect 587 28020 600 28066
rect 674 28020 687 28066
rect 587 28007 687 28020
rect 1067 28378 1167 28391
rect 1067 28332 1080 28378
rect 1154 28332 1167 28378
rect 1067 28299 1167 28332
rect 1067 28066 1167 28099
rect 1067 28020 1080 28066
rect 1154 28020 1167 28066
rect 1067 28007 1167 28020
rect 9171 28379 9271 28392
rect 9171 28333 9184 28379
rect 9258 28333 9271 28379
rect 9171 28300 9271 28333
rect 9375 28379 9475 28392
rect 9375 28333 9388 28379
rect 9462 28333 9475 28379
rect 9375 28300 9475 28333
rect 9171 28067 9271 28100
rect 9171 28021 9184 28067
rect 9258 28021 9271 28067
rect 9171 28008 9271 28021
rect 9375 28067 9475 28100
rect 9375 28021 9388 28067
rect 9462 28021 9475 28067
rect 9375 28008 9475 28021
rect 9855 28379 9955 28392
rect 9855 28333 9868 28379
rect 9942 28333 9955 28379
rect 9855 28300 9955 28333
rect 10059 28379 10159 28392
rect 10059 28333 10072 28379
rect 10146 28333 10159 28379
rect 10059 28300 10159 28333
rect 9855 28067 9955 28100
rect 9855 28021 9868 28067
rect 9942 28021 9955 28067
rect 9855 28008 9955 28021
rect 10059 28067 10159 28100
rect 10059 28021 10072 28067
rect 10146 28021 10159 28067
rect 10059 28008 10159 28021
rect 10539 28379 10639 28392
rect 10539 28333 10552 28379
rect 10626 28333 10639 28379
rect 10539 28300 10639 28333
rect 10539 28067 10639 28100
rect 10539 28021 10552 28067
rect 10626 28021 10639 28067
rect 10539 28008 10639 28021
rect 18643 28379 18743 28392
rect 18643 28333 18656 28379
rect 18730 28333 18743 28379
rect 18643 28300 18743 28333
rect 18847 28379 18947 28392
rect 18847 28333 18860 28379
rect 18934 28333 18947 28379
rect 18847 28300 18947 28333
rect 18643 28067 18743 28100
rect 18643 28021 18656 28067
rect 18730 28021 18743 28067
rect 18643 28008 18743 28021
rect 18847 28067 18947 28100
rect 18847 28021 18860 28067
rect 18934 28021 18947 28067
rect 18847 28008 18947 28021
rect 19327 28379 19427 28392
rect 19327 28333 19340 28379
rect 19414 28333 19427 28379
rect 19327 28300 19427 28333
rect 19531 28379 19631 28392
rect 19531 28333 19544 28379
rect 19618 28333 19631 28379
rect 19531 28300 19631 28333
rect 19327 28067 19427 28100
rect 19327 28021 19340 28067
rect 19414 28021 19427 28067
rect 19327 28008 19427 28021
rect 19531 28067 19631 28100
rect 19531 28021 19544 28067
rect 19618 28021 19631 28067
rect 19531 28008 19631 28021
rect 20011 28379 20111 28392
rect 20011 28333 20024 28379
rect 20098 28333 20111 28379
rect 20011 28300 20111 28333
rect 20011 28067 20111 28100
rect 20011 28021 20024 28067
rect 20098 28021 20111 28067
rect 20011 28008 20111 28021
rect 28115 28379 28215 28392
rect 28115 28333 28128 28379
rect 28202 28333 28215 28379
rect 28115 28300 28215 28333
rect 28319 28379 28419 28392
rect 28319 28333 28332 28379
rect 28406 28333 28419 28379
rect 28319 28300 28419 28333
rect 28115 28067 28215 28100
rect 28115 28021 28128 28067
rect 28202 28021 28215 28067
rect 28115 28008 28215 28021
rect 28319 28067 28419 28100
rect 28319 28021 28332 28067
rect 28406 28021 28419 28067
rect 28319 28008 28419 28021
rect 28799 28379 28899 28392
rect 28799 28333 28812 28379
rect 28886 28333 28899 28379
rect 28799 28300 28899 28333
rect 29003 28379 29103 28392
rect 29003 28333 29016 28379
rect 29090 28333 29103 28379
rect 29003 28300 29103 28333
rect 28799 28067 28899 28100
rect 28799 28021 28812 28067
rect 28886 28021 28899 28067
rect 28799 28008 28899 28021
rect 29003 28067 29103 28100
rect 29003 28021 29016 28067
rect 29090 28021 29103 28067
rect 29003 28008 29103 28021
rect 29483 28379 29583 28392
rect 29483 28333 29496 28379
rect 29570 28333 29583 28379
rect 29483 28300 29583 28333
rect 29483 28067 29583 28100
rect 29483 28021 29496 28067
rect 29570 28021 29583 28067
rect 29483 28008 29583 28021
rect 37587 28379 37687 28392
rect 37587 28333 37600 28379
rect 37674 28333 37687 28379
rect 37587 28300 37687 28333
rect 37791 28379 37891 28392
rect 37791 28333 37804 28379
rect 37878 28333 37891 28379
rect 37791 28300 37891 28333
rect 37587 28067 37687 28100
rect 37587 28021 37600 28067
rect 37674 28021 37687 28067
rect 37587 28008 37687 28021
rect 37791 28067 37891 28100
rect 37791 28021 37804 28067
rect 37878 28021 37891 28067
rect 37791 28008 37891 28021
rect 38271 28379 38371 28392
rect 38271 28333 38284 28379
rect 38358 28333 38371 28379
rect 38271 28300 38371 28333
rect 38475 28379 38575 28392
rect 38475 28333 38488 28379
rect 38562 28333 38575 28379
rect 38475 28300 38575 28333
rect 38271 28067 38371 28100
rect 38271 28021 38284 28067
rect 38358 28021 38371 28067
rect 38271 28008 38371 28021
rect 38475 28067 38575 28100
rect 38475 28021 38488 28067
rect 38562 28021 38575 28067
rect 38475 28008 38575 28021
rect 38955 28379 39055 28392
rect 38955 28333 38968 28379
rect 39042 28333 39055 28379
rect 38955 28300 39055 28333
rect 38955 28067 39055 28100
rect 38955 28021 38968 28067
rect 39042 28021 39055 28067
rect 38955 28008 39055 28021
rect -12380 27368 -12280 27381
rect -12380 27322 -12367 27368
rect -12293 27322 -12280 27368
rect -12380 27289 -12280 27322
rect -12380 27056 -12280 27089
rect -12380 27010 -12367 27056
rect -12293 27010 -12280 27056
rect -12380 26997 -12280 27010
rect -7889 25061 -7809 25074
rect -7889 25015 -7876 25061
rect -7822 25015 -7809 25061
rect -7889 24982 -7809 25015
rect -7705 25061 -7625 25074
rect -7705 25015 -7692 25061
rect -7638 25015 -7625 25061
rect -7705 24982 -7625 25015
rect -7521 25061 -7441 25074
rect -7521 25015 -7508 25061
rect -7454 25015 -7441 25061
rect -7521 24982 -7441 25015
rect -7889 24449 -7809 24482
rect -7889 24403 -7876 24449
rect -7822 24403 -7809 24449
rect -7889 24390 -7809 24403
rect -7705 24449 -7625 24482
rect -7705 24403 -7692 24449
rect -7638 24403 -7625 24449
rect -7705 24390 -7625 24403
rect -7521 24449 -7441 24482
rect -7521 24403 -7508 24449
rect -7454 24403 -7441 24449
rect -7521 24390 -7441 24403
rect -3847 25058 -3767 25071
rect -3847 25012 -3834 25058
rect -3780 25012 -3767 25058
rect -3847 24979 -3767 25012
rect -3663 25058 -3583 25071
rect -3663 25012 -3650 25058
rect -3596 25012 -3583 25058
rect -3663 24979 -3583 25012
rect -3479 25058 -3399 25071
rect -3479 25012 -3466 25058
rect -3412 25012 -3399 25058
rect -3479 24979 -3399 25012
rect -3847 24446 -3767 24479
rect -3847 24400 -3834 24446
rect -3780 24400 -3767 24446
rect -3847 24387 -3767 24400
rect -3663 24446 -3583 24479
rect -3663 24400 -3650 24446
rect -3596 24400 -3583 24446
rect -3663 24387 -3583 24400
rect -3479 24446 -3399 24479
rect -3479 24400 -3466 24446
rect -3412 24400 -3399 24446
rect -3479 24387 -3399 24400
rect 195 25058 275 25071
rect 195 25012 208 25058
rect 262 25012 275 25058
rect 195 24979 275 25012
rect 379 25058 459 25071
rect 379 25012 392 25058
rect 446 25012 459 25058
rect 379 24979 459 25012
rect 563 25058 643 25071
rect 563 25012 576 25058
rect 630 25012 643 25058
rect 563 24979 643 25012
rect 195 24446 275 24479
rect 195 24400 208 24446
rect 262 24400 275 24446
rect 195 24387 275 24400
rect 379 24446 459 24479
rect 379 24400 392 24446
rect 446 24400 459 24446
rect 379 24387 459 24400
rect 563 24446 643 24479
rect 563 24400 576 24446
rect 630 24400 643 24446
rect 563 24387 643 24400
rect 4237 25058 4317 25071
rect 4237 25012 4250 25058
rect 4304 25012 4317 25058
rect 4237 24979 4317 25012
rect 4421 25058 4501 25071
rect 4421 25012 4434 25058
rect 4488 25012 4501 25058
rect 4421 24979 4501 25012
rect 4605 25058 4685 25071
rect 4605 25012 4618 25058
rect 4672 25012 4685 25058
rect 4605 24979 4685 25012
rect 4237 24446 4317 24479
rect 4237 24400 4250 24446
rect 4304 24400 4317 24446
rect 4237 24387 4317 24400
rect 4421 24446 4501 24479
rect 4421 24400 4434 24446
rect 4488 24400 4501 24446
rect 4421 24387 4501 24400
rect 4605 24446 4685 24479
rect 4605 24400 4618 24446
rect 4672 24400 4685 24446
rect 4605 24387 4685 24400
rect 8279 25058 8359 25071
rect 8279 25012 8292 25058
rect 8346 25012 8359 25058
rect 8279 24979 8359 25012
rect 8463 25058 8543 25071
rect 8463 25012 8476 25058
rect 8530 25012 8543 25058
rect 8463 24979 8543 25012
rect 8647 25058 8727 25071
rect 8647 25012 8660 25058
rect 8714 25012 8727 25058
rect 8647 24979 8727 25012
rect 8279 24446 8359 24479
rect 8279 24400 8292 24446
rect 8346 24400 8359 24446
rect 8279 24387 8359 24400
rect 8463 24446 8543 24479
rect 8463 24400 8476 24446
rect 8530 24400 8543 24446
rect 8463 24387 8543 24400
rect 8647 24446 8727 24479
rect 8647 24400 8660 24446
rect 8714 24400 8727 24446
rect 8647 24387 8727 24400
rect 12321 25058 12401 25071
rect 12321 25012 12334 25058
rect 12388 25012 12401 25058
rect 12321 24979 12401 25012
rect 12505 25058 12585 25071
rect 12505 25012 12518 25058
rect 12572 25012 12585 25058
rect 12505 24979 12585 25012
rect 12689 25058 12769 25071
rect 12689 25012 12702 25058
rect 12756 25012 12769 25058
rect 12689 24979 12769 25012
rect 12321 24446 12401 24479
rect 12321 24400 12334 24446
rect 12388 24400 12401 24446
rect 12321 24387 12401 24400
rect 12505 24446 12585 24479
rect 12505 24400 12518 24446
rect 12572 24400 12585 24446
rect 12505 24387 12585 24400
rect 12689 24446 12769 24479
rect 12689 24400 12702 24446
rect 12756 24400 12769 24446
rect 12689 24387 12769 24400
rect 16363 25058 16443 25071
rect 16363 25012 16376 25058
rect 16430 25012 16443 25058
rect 16363 24979 16443 25012
rect 16547 25058 16627 25071
rect 16547 25012 16560 25058
rect 16614 25012 16627 25058
rect 16547 24979 16627 25012
rect 16731 25058 16811 25071
rect 16731 25012 16744 25058
rect 16798 25012 16811 25058
rect 16731 24979 16811 25012
rect 16363 24446 16443 24479
rect 16363 24400 16376 24446
rect 16430 24400 16443 24446
rect 16363 24387 16443 24400
rect 16547 24446 16627 24479
rect 16547 24400 16560 24446
rect 16614 24400 16627 24446
rect 16547 24387 16627 24400
rect 16731 24446 16811 24479
rect 16731 24400 16744 24446
rect 16798 24400 16811 24446
rect 16731 24387 16811 24400
rect -7889 23901 -7809 23914
rect -7889 23855 -7876 23901
rect -7822 23855 -7809 23901
rect -7889 23822 -7809 23855
rect -7705 23901 -7625 23914
rect -7705 23855 -7692 23901
rect -7638 23855 -7625 23901
rect -7705 23822 -7625 23855
rect -7521 23901 -7441 23914
rect -7521 23855 -7508 23901
rect -7454 23855 -7441 23901
rect -7521 23822 -7441 23855
rect -7889 23589 -7809 23622
rect -7889 23543 -7876 23589
rect -7822 23543 -7809 23589
rect -7889 23530 -7809 23543
rect -7705 23589 -7625 23622
rect -7705 23543 -7692 23589
rect -7638 23543 -7625 23589
rect -7705 23530 -7625 23543
rect -7521 23589 -7441 23622
rect -7521 23543 -7508 23589
rect -7454 23543 -7441 23589
rect -7521 23530 -7441 23543
rect -3847 23898 -3767 23911
rect -3847 23852 -3834 23898
rect -3780 23852 -3767 23898
rect -3847 23819 -3767 23852
rect -3663 23898 -3583 23911
rect -3663 23852 -3650 23898
rect -3596 23852 -3583 23898
rect -3663 23819 -3583 23852
rect -3479 23898 -3399 23911
rect -3479 23852 -3466 23898
rect -3412 23852 -3399 23898
rect -3479 23819 -3399 23852
rect -3847 23586 -3767 23619
rect -3847 23540 -3834 23586
rect -3780 23540 -3767 23586
rect -3847 23527 -3767 23540
rect -3663 23586 -3583 23619
rect -3663 23540 -3650 23586
rect -3596 23540 -3583 23586
rect -3663 23527 -3583 23540
rect -3479 23586 -3399 23619
rect -3479 23540 -3466 23586
rect -3412 23540 -3399 23586
rect -3479 23527 -3399 23540
rect 195 23898 275 23911
rect 195 23852 208 23898
rect 262 23852 275 23898
rect 195 23819 275 23852
rect 379 23898 459 23911
rect 379 23852 392 23898
rect 446 23852 459 23898
rect 379 23819 459 23852
rect 563 23898 643 23911
rect 563 23852 576 23898
rect 630 23852 643 23898
rect 563 23819 643 23852
rect 195 23586 275 23619
rect 195 23540 208 23586
rect 262 23540 275 23586
rect 195 23527 275 23540
rect 379 23586 459 23619
rect 379 23540 392 23586
rect 446 23540 459 23586
rect 379 23527 459 23540
rect 563 23586 643 23619
rect 563 23540 576 23586
rect 630 23540 643 23586
rect 563 23527 643 23540
rect 4237 23898 4317 23911
rect 4237 23852 4250 23898
rect 4304 23852 4317 23898
rect 4237 23819 4317 23852
rect 4421 23898 4501 23911
rect 4421 23852 4434 23898
rect 4488 23852 4501 23898
rect 4421 23819 4501 23852
rect 4605 23898 4685 23911
rect 4605 23852 4618 23898
rect 4672 23852 4685 23898
rect 4605 23819 4685 23852
rect 4237 23586 4317 23619
rect 4237 23540 4250 23586
rect 4304 23540 4317 23586
rect 4237 23527 4317 23540
rect 4421 23586 4501 23619
rect 4421 23540 4434 23586
rect 4488 23540 4501 23586
rect 4421 23527 4501 23540
rect 4605 23586 4685 23619
rect 4605 23540 4618 23586
rect 4672 23540 4685 23586
rect 4605 23527 4685 23540
rect 8279 23898 8359 23911
rect 8279 23852 8292 23898
rect 8346 23852 8359 23898
rect 8279 23819 8359 23852
rect 8463 23898 8543 23911
rect 8463 23852 8476 23898
rect 8530 23852 8543 23898
rect 8463 23819 8543 23852
rect 8647 23898 8727 23911
rect 8647 23852 8660 23898
rect 8714 23852 8727 23898
rect 8647 23819 8727 23852
rect 8279 23586 8359 23619
rect 8279 23540 8292 23586
rect 8346 23540 8359 23586
rect 8279 23527 8359 23540
rect 8463 23586 8543 23619
rect 8463 23540 8476 23586
rect 8530 23540 8543 23586
rect 8463 23527 8543 23540
rect 8647 23586 8727 23619
rect 8647 23540 8660 23586
rect 8714 23540 8727 23586
rect 8647 23527 8727 23540
rect 12321 23898 12401 23911
rect 12321 23852 12334 23898
rect 12388 23852 12401 23898
rect 12321 23819 12401 23852
rect 12505 23898 12585 23911
rect 12505 23852 12518 23898
rect 12572 23852 12585 23898
rect 12505 23819 12585 23852
rect 12689 23898 12769 23911
rect 12689 23852 12702 23898
rect 12756 23852 12769 23898
rect 12689 23819 12769 23852
rect 12321 23586 12401 23619
rect 12321 23540 12334 23586
rect 12388 23540 12401 23586
rect 12321 23527 12401 23540
rect 12505 23586 12585 23619
rect 12505 23540 12518 23586
rect 12572 23540 12585 23586
rect 12505 23527 12585 23540
rect 12689 23586 12769 23619
rect 12689 23540 12702 23586
rect 12756 23540 12769 23586
rect 12689 23527 12769 23540
rect 16363 23898 16443 23911
rect 16363 23852 16376 23898
rect 16430 23852 16443 23898
rect 16363 23819 16443 23852
rect 16547 23898 16627 23911
rect 16547 23852 16560 23898
rect 16614 23852 16627 23898
rect 16547 23819 16627 23852
rect 16731 23898 16811 23911
rect 16731 23852 16744 23898
rect 16798 23852 16811 23898
rect 16731 23819 16811 23852
rect 16363 23586 16443 23619
rect 16363 23540 16376 23586
rect 16430 23540 16443 23586
rect 16363 23527 16443 23540
rect 16547 23586 16627 23619
rect 16547 23540 16560 23586
rect 16614 23540 16627 23586
rect 16547 23527 16627 23540
rect 16731 23586 16811 23619
rect 16731 23540 16744 23586
rect 16798 23540 16811 23586
rect 16731 23527 16811 23540
rect -7889 22856 -7809 22869
rect -7889 22810 -7876 22856
rect -7822 22810 -7809 22856
rect -7889 22777 -7809 22810
rect -7705 22856 -7625 22869
rect -7705 22810 -7692 22856
rect -7638 22810 -7625 22856
rect -7705 22777 -7625 22810
rect -7521 22856 -7441 22869
rect -7521 22810 -7508 22856
rect -7454 22810 -7441 22856
rect -7521 22777 -7441 22810
rect -7889 22244 -7809 22277
rect -7889 22198 -7876 22244
rect -7822 22198 -7809 22244
rect -7889 22185 -7809 22198
rect -7705 22244 -7625 22277
rect -7705 22198 -7692 22244
rect -7638 22198 -7625 22244
rect -7705 22185 -7625 22198
rect -7521 22244 -7441 22277
rect -7521 22198 -7508 22244
rect -7454 22198 -7441 22244
rect -7521 22185 -7441 22198
rect -6403 22856 -6323 22869
rect -6403 22810 -6390 22856
rect -6336 22810 -6323 22856
rect -6403 22777 -6323 22810
rect -6219 22856 -6139 22869
rect -6219 22810 -6206 22856
rect -6152 22810 -6139 22856
rect -6219 22777 -6139 22810
rect -6035 22856 -5955 22869
rect -6035 22810 -6022 22856
rect -5968 22810 -5955 22856
rect -6035 22777 -5955 22810
rect -6403 22244 -6323 22277
rect -6403 22198 -6390 22244
rect -6336 22198 -6323 22244
rect -6403 22185 -6323 22198
rect -6219 22244 -6139 22277
rect -6219 22198 -6206 22244
rect -6152 22198 -6139 22244
rect -6219 22185 -6139 22198
rect -6035 22244 -5955 22277
rect -6035 22198 -6022 22244
rect -5968 22198 -5955 22244
rect -6035 22185 -5955 22198
rect -3847 22853 -3767 22866
rect -3847 22807 -3834 22853
rect -3780 22807 -3767 22853
rect -3847 22774 -3767 22807
rect -3663 22853 -3583 22866
rect -3663 22807 -3650 22853
rect -3596 22807 -3583 22853
rect -3663 22774 -3583 22807
rect -3479 22853 -3399 22866
rect -3479 22807 -3466 22853
rect -3412 22807 -3399 22853
rect -3479 22774 -3399 22807
rect -3847 22241 -3767 22274
rect -3847 22195 -3834 22241
rect -3780 22195 -3767 22241
rect -3847 22182 -3767 22195
rect -3663 22241 -3583 22274
rect -3663 22195 -3650 22241
rect -3596 22195 -3583 22241
rect -3663 22182 -3583 22195
rect -3479 22241 -3399 22274
rect -3479 22195 -3466 22241
rect -3412 22195 -3399 22241
rect -3479 22182 -3399 22195
rect -2361 22853 -2281 22866
rect -2361 22807 -2348 22853
rect -2294 22807 -2281 22853
rect -2361 22774 -2281 22807
rect -2177 22853 -2097 22866
rect -2177 22807 -2164 22853
rect -2110 22807 -2097 22853
rect -2177 22774 -2097 22807
rect -1993 22853 -1913 22866
rect -1993 22807 -1980 22853
rect -1926 22807 -1913 22853
rect -1993 22774 -1913 22807
rect -2361 22241 -2281 22274
rect -2361 22195 -2348 22241
rect -2294 22195 -2281 22241
rect -2361 22182 -2281 22195
rect -2177 22241 -2097 22274
rect -2177 22195 -2164 22241
rect -2110 22195 -2097 22241
rect -2177 22182 -2097 22195
rect -1993 22241 -1913 22274
rect -1993 22195 -1980 22241
rect -1926 22195 -1913 22241
rect -1993 22182 -1913 22195
rect 195 22853 275 22866
rect 195 22807 208 22853
rect 262 22807 275 22853
rect 195 22774 275 22807
rect 379 22853 459 22866
rect 379 22807 392 22853
rect 446 22807 459 22853
rect 379 22774 459 22807
rect 563 22853 643 22866
rect 563 22807 576 22853
rect 630 22807 643 22853
rect 563 22774 643 22807
rect 195 22241 275 22274
rect 195 22195 208 22241
rect 262 22195 275 22241
rect 195 22182 275 22195
rect 379 22241 459 22274
rect 379 22195 392 22241
rect 446 22195 459 22241
rect 379 22182 459 22195
rect 563 22241 643 22274
rect 563 22195 576 22241
rect 630 22195 643 22241
rect 563 22182 643 22195
rect 1681 22853 1761 22866
rect 1681 22807 1694 22853
rect 1748 22807 1761 22853
rect 1681 22774 1761 22807
rect 1865 22853 1945 22866
rect 1865 22807 1878 22853
rect 1932 22807 1945 22853
rect 1865 22774 1945 22807
rect 2049 22853 2129 22866
rect 2049 22807 2062 22853
rect 2116 22807 2129 22853
rect 2049 22774 2129 22807
rect 1681 22241 1761 22274
rect 1681 22195 1694 22241
rect 1748 22195 1761 22241
rect 1681 22182 1761 22195
rect 1865 22241 1945 22274
rect 1865 22195 1878 22241
rect 1932 22195 1945 22241
rect 1865 22182 1945 22195
rect 2049 22241 2129 22274
rect 2049 22195 2062 22241
rect 2116 22195 2129 22241
rect 2049 22182 2129 22195
rect 4237 22853 4317 22866
rect 4237 22807 4250 22853
rect 4304 22807 4317 22853
rect 4237 22774 4317 22807
rect 4421 22853 4501 22866
rect 4421 22807 4434 22853
rect 4488 22807 4501 22853
rect 4421 22774 4501 22807
rect 4605 22853 4685 22866
rect 4605 22807 4618 22853
rect 4672 22807 4685 22853
rect 4605 22774 4685 22807
rect 4237 22241 4317 22274
rect 4237 22195 4250 22241
rect 4304 22195 4317 22241
rect 4237 22182 4317 22195
rect 4421 22241 4501 22274
rect 4421 22195 4434 22241
rect 4488 22195 4501 22241
rect 4421 22182 4501 22195
rect 4605 22241 4685 22274
rect 4605 22195 4618 22241
rect 4672 22195 4685 22241
rect 4605 22182 4685 22195
rect 5723 22853 5803 22866
rect 5723 22807 5736 22853
rect 5790 22807 5803 22853
rect 5723 22774 5803 22807
rect 5907 22853 5987 22866
rect 5907 22807 5920 22853
rect 5974 22807 5987 22853
rect 5907 22774 5987 22807
rect 6091 22853 6171 22866
rect 6091 22807 6104 22853
rect 6158 22807 6171 22853
rect 6091 22774 6171 22807
rect 5723 22241 5803 22274
rect 5723 22195 5736 22241
rect 5790 22195 5803 22241
rect 5723 22182 5803 22195
rect 5907 22241 5987 22274
rect 5907 22195 5920 22241
rect 5974 22195 5987 22241
rect 5907 22182 5987 22195
rect 6091 22241 6171 22274
rect 6091 22195 6104 22241
rect 6158 22195 6171 22241
rect 6091 22182 6171 22195
rect 8279 22853 8359 22866
rect 8279 22807 8292 22853
rect 8346 22807 8359 22853
rect 8279 22774 8359 22807
rect 8463 22853 8543 22866
rect 8463 22807 8476 22853
rect 8530 22807 8543 22853
rect 8463 22774 8543 22807
rect 8647 22853 8727 22866
rect 8647 22807 8660 22853
rect 8714 22807 8727 22853
rect 8647 22774 8727 22807
rect 8279 22241 8359 22274
rect 8279 22195 8292 22241
rect 8346 22195 8359 22241
rect 8279 22182 8359 22195
rect 8463 22241 8543 22274
rect 8463 22195 8476 22241
rect 8530 22195 8543 22241
rect 8463 22182 8543 22195
rect 8647 22241 8727 22274
rect 8647 22195 8660 22241
rect 8714 22195 8727 22241
rect 8647 22182 8727 22195
rect 9765 22853 9845 22866
rect 9765 22807 9778 22853
rect 9832 22807 9845 22853
rect 9765 22774 9845 22807
rect 9949 22853 10029 22866
rect 9949 22807 9962 22853
rect 10016 22807 10029 22853
rect 9949 22774 10029 22807
rect 10133 22853 10213 22866
rect 10133 22807 10146 22853
rect 10200 22807 10213 22853
rect 10133 22774 10213 22807
rect 9765 22241 9845 22274
rect 9765 22195 9778 22241
rect 9832 22195 9845 22241
rect 9765 22182 9845 22195
rect 9949 22241 10029 22274
rect 9949 22195 9962 22241
rect 10016 22195 10029 22241
rect 9949 22182 10029 22195
rect 10133 22241 10213 22274
rect 10133 22195 10146 22241
rect 10200 22195 10213 22241
rect 10133 22182 10213 22195
rect 12321 22853 12401 22866
rect 12321 22807 12334 22853
rect 12388 22807 12401 22853
rect 12321 22774 12401 22807
rect 12505 22853 12585 22866
rect 12505 22807 12518 22853
rect 12572 22807 12585 22853
rect 12505 22774 12585 22807
rect 12689 22853 12769 22866
rect 12689 22807 12702 22853
rect 12756 22807 12769 22853
rect 12689 22774 12769 22807
rect 12321 22241 12401 22274
rect 12321 22195 12334 22241
rect 12388 22195 12401 22241
rect 12321 22182 12401 22195
rect 12505 22241 12585 22274
rect 12505 22195 12518 22241
rect 12572 22195 12585 22241
rect 12505 22182 12585 22195
rect 12689 22241 12769 22274
rect 12689 22195 12702 22241
rect 12756 22195 12769 22241
rect 12689 22182 12769 22195
rect 13807 22853 13887 22866
rect 13807 22807 13820 22853
rect 13874 22807 13887 22853
rect 13807 22774 13887 22807
rect 13991 22853 14071 22866
rect 13991 22807 14004 22853
rect 14058 22807 14071 22853
rect 13991 22774 14071 22807
rect 14175 22853 14255 22866
rect 14175 22807 14188 22853
rect 14242 22807 14255 22853
rect 14175 22774 14255 22807
rect 13807 22241 13887 22274
rect 13807 22195 13820 22241
rect 13874 22195 13887 22241
rect 13807 22182 13887 22195
rect 13991 22241 14071 22274
rect 13991 22195 14004 22241
rect 14058 22195 14071 22241
rect 13991 22182 14071 22195
rect 14175 22241 14255 22274
rect 14175 22195 14188 22241
rect 14242 22195 14255 22241
rect 14175 22182 14255 22195
rect 16363 22853 16443 22866
rect 16363 22807 16376 22853
rect 16430 22807 16443 22853
rect 16363 22774 16443 22807
rect 16547 22853 16627 22866
rect 16547 22807 16560 22853
rect 16614 22807 16627 22853
rect 16547 22774 16627 22807
rect 16731 22853 16811 22866
rect 16731 22807 16744 22853
rect 16798 22807 16811 22853
rect 16731 22774 16811 22807
rect 16363 22241 16443 22274
rect 16363 22195 16376 22241
rect 16430 22195 16443 22241
rect 16363 22182 16443 22195
rect 16547 22241 16627 22274
rect 16547 22195 16560 22241
rect 16614 22195 16627 22241
rect 16547 22182 16627 22195
rect 16731 22241 16811 22274
rect 16731 22195 16744 22241
rect 16798 22195 16811 22241
rect 16731 22182 16811 22195
rect 17849 22853 17929 22866
rect 17849 22807 17862 22853
rect 17916 22807 17929 22853
rect 17849 22774 17929 22807
rect 18033 22853 18113 22866
rect 18033 22807 18046 22853
rect 18100 22807 18113 22853
rect 18033 22774 18113 22807
rect 18217 22853 18297 22866
rect 18217 22807 18230 22853
rect 18284 22807 18297 22853
rect 18217 22774 18297 22807
rect 17849 22241 17929 22274
rect 17849 22195 17862 22241
rect 17916 22195 17929 22241
rect 17849 22182 17929 22195
rect 18033 22241 18113 22274
rect 18033 22195 18046 22241
rect 18100 22195 18113 22241
rect 18033 22182 18113 22195
rect 18217 22241 18297 22274
rect 18217 22195 18230 22241
rect 18284 22195 18297 22241
rect 18217 22182 18297 22195
rect -7889 21696 -7809 21709
rect -7889 21650 -7876 21696
rect -7822 21650 -7809 21696
rect -7889 21617 -7809 21650
rect -7705 21696 -7625 21709
rect -7705 21650 -7692 21696
rect -7638 21650 -7625 21696
rect -7705 21617 -7625 21650
rect -7521 21696 -7441 21709
rect -7521 21650 -7508 21696
rect -7454 21650 -7441 21696
rect -7521 21617 -7441 21650
rect -7889 21384 -7809 21417
rect -7889 21338 -7876 21384
rect -7822 21338 -7809 21384
rect -7889 21325 -7809 21338
rect -7705 21384 -7625 21417
rect -7705 21338 -7692 21384
rect -7638 21338 -7625 21384
rect -7705 21325 -7625 21338
rect -7521 21384 -7441 21417
rect -7521 21338 -7508 21384
rect -7454 21338 -7441 21384
rect -7521 21325 -7441 21338
rect -6403 21696 -6323 21709
rect -6403 21650 -6390 21696
rect -6336 21650 -6323 21696
rect -6403 21617 -6323 21650
rect -6219 21696 -6139 21709
rect -6219 21650 -6206 21696
rect -6152 21650 -6139 21696
rect -6219 21617 -6139 21650
rect -6035 21696 -5955 21709
rect -6035 21650 -6022 21696
rect -5968 21650 -5955 21696
rect -6035 21617 -5955 21650
rect -6403 21384 -6323 21417
rect -6403 21338 -6390 21384
rect -6336 21338 -6323 21384
rect -6403 21325 -6323 21338
rect -6219 21384 -6139 21417
rect -6219 21338 -6206 21384
rect -6152 21338 -6139 21384
rect -6219 21325 -6139 21338
rect -6035 21384 -5955 21417
rect -6035 21338 -6022 21384
rect -5968 21338 -5955 21384
rect -6035 21325 -5955 21338
rect -3847 21693 -3767 21706
rect -3847 21647 -3834 21693
rect -3780 21647 -3767 21693
rect -3847 21614 -3767 21647
rect -3663 21693 -3583 21706
rect -3663 21647 -3650 21693
rect -3596 21647 -3583 21693
rect -3663 21614 -3583 21647
rect -3479 21693 -3399 21706
rect -3479 21647 -3466 21693
rect -3412 21647 -3399 21693
rect -3479 21614 -3399 21647
rect -3847 21381 -3767 21414
rect -3847 21335 -3834 21381
rect -3780 21335 -3767 21381
rect -3847 21322 -3767 21335
rect -3663 21381 -3583 21414
rect -3663 21335 -3650 21381
rect -3596 21335 -3583 21381
rect -3663 21322 -3583 21335
rect -3479 21381 -3399 21414
rect -3479 21335 -3466 21381
rect -3412 21335 -3399 21381
rect -3479 21322 -3399 21335
rect -2361 21693 -2281 21706
rect -2361 21647 -2348 21693
rect -2294 21647 -2281 21693
rect -2361 21614 -2281 21647
rect -2177 21693 -2097 21706
rect -2177 21647 -2164 21693
rect -2110 21647 -2097 21693
rect -2177 21614 -2097 21647
rect -1993 21693 -1913 21706
rect -1993 21647 -1980 21693
rect -1926 21647 -1913 21693
rect -1993 21614 -1913 21647
rect -2361 21381 -2281 21414
rect -2361 21335 -2348 21381
rect -2294 21335 -2281 21381
rect -2361 21322 -2281 21335
rect -2177 21381 -2097 21414
rect -2177 21335 -2164 21381
rect -2110 21335 -2097 21381
rect -2177 21322 -2097 21335
rect -1993 21381 -1913 21414
rect -1993 21335 -1980 21381
rect -1926 21335 -1913 21381
rect -1993 21322 -1913 21335
rect 195 21693 275 21706
rect 195 21647 208 21693
rect 262 21647 275 21693
rect 195 21614 275 21647
rect 379 21693 459 21706
rect 379 21647 392 21693
rect 446 21647 459 21693
rect 379 21614 459 21647
rect 563 21693 643 21706
rect 563 21647 576 21693
rect 630 21647 643 21693
rect 563 21614 643 21647
rect 195 21381 275 21414
rect 195 21335 208 21381
rect 262 21335 275 21381
rect 195 21322 275 21335
rect 379 21381 459 21414
rect 379 21335 392 21381
rect 446 21335 459 21381
rect 379 21322 459 21335
rect 563 21381 643 21414
rect 563 21335 576 21381
rect 630 21335 643 21381
rect 563 21322 643 21335
rect 1681 21693 1761 21706
rect 1681 21647 1694 21693
rect 1748 21647 1761 21693
rect 1681 21614 1761 21647
rect 1865 21693 1945 21706
rect 1865 21647 1878 21693
rect 1932 21647 1945 21693
rect 1865 21614 1945 21647
rect 2049 21693 2129 21706
rect 2049 21647 2062 21693
rect 2116 21647 2129 21693
rect 2049 21614 2129 21647
rect 1681 21381 1761 21414
rect 1681 21335 1694 21381
rect 1748 21335 1761 21381
rect 1681 21322 1761 21335
rect 1865 21381 1945 21414
rect 1865 21335 1878 21381
rect 1932 21335 1945 21381
rect 1865 21322 1945 21335
rect 2049 21381 2129 21414
rect 2049 21335 2062 21381
rect 2116 21335 2129 21381
rect 2049 21322 2129 21335
rect 4237 21693 4317 21706
rect 4237 21647 4250 21693
rect 4304 21647 4317 21693
rect 4237 21614 4317 21647
rect 4421 21693 4501 21706
rect 4421 21647 4434 21693
rect 4488 21647 4501 21693
rect 4421 21614 4501 21647
rect 4605 21693 4685 21706
rect 4605 21647 4618 21693
rect 4672 21647 4685 21693
rect 4605 21614 4685 21647
rect 4237 21381 4317 21414
rect 4237 21335 4250 21381
rect 4304 21335 4317 21381
rect 4237 21322 4317 21335
rect 4421 21381 4501 21414
rect 4421 21335 4434 21381
rect 4488 21335 4501 21381
rect 4421 21322 4501 21335
rect 4605 21381 4685 21414
rect 4605 21335 4618 21381
rect 4672 21335 4685 21381
rect 4605 21322 4685 21335
rect 5723 21693 5803 21706
rect 5723 21647 5736 21693
rect 5790 21647 5803 21693
rect 5723 21614 5803 21647
rect 5907 21693 5987 21706
rect 5907 21647 5920 21693
rect 5974 21647 5987 21693
rect 5907 21614 5987 21647
rect 6091 21693 6171 21706
rect 6091 21647 6104 21693
rect 6158 21647 6171 21693
rect 6091 21614 6171 21647
rect 5723 21381 5803 21414
rect 5723 21335 5736 21381
rect 5790 21335 5803 21381
rect 5723 21322 5803 21335
rect 5907 21381 5987 21414
rect 5907 21335 5920 21381
rect 5974 21335 5987 21381
rect 5907 21322 5987 21335
rect 6091 21381 6171 21414
rect 6091 21335 6104 21381
rect 6158 21335 6171 21381
rect 6091 21322 6171 21335
rect 8279 21693 8359 21706
rect 8279 21647 8292 21693
rect 8346 21647 8359 21693
rect 8279 21614 8359 21647
rect 8463 21693 8543 21706
rect 8463 21647 8476 21693
rect 8530 21647 8543 21693
rect 8463 21614 8543 21647
rect 8647 21693 8727 21706
rect 8647 21647 8660 21693
rect 8714 21647 8727 21693
rect 8647 21614 8727 21647
rect 8279 21381 8359 21414
rect 8279 21335 8292 21381
rect 8346 21335 8359 21381
rect 8279 21322 8359 21335
rect 8463 21381 8543 21414
rect 8463 21335 8476 21381
rect 8530 21335 8543 21381
rect 8463 21322 8543 21335
rect 8647 21381 8727 21414
rect 8647 21335 8660 21381
rect 8714 21335 8727 21381
rect 8647 21322 8727 21335
rect 9765 21693 9845 21706
rect 9765 21647 9778 21693
rect 9832 21647 9845 21693
rect 9765 21614 9845 21647
rect 9949 21693 10029 21706
rect 9949 21647 9962 21693
rect 10016 21647 10029 21693
rect 9949 21614 10029 21647
rect 10133 21693 10213 21706
rect 10133 21647 10146 21693
rect 10200 21647 10213 21693
rect 10133 21614 10213 21647
rect 9765 21381 9845 21414
rect 9765 21335 9778 21381
rect 9832 21335 9845 21381
rect 9765 21322 9845 21335
rect 9949 21381 10029 21414
rect 9949 21335 9962 21381
rect 10016 21335 10029 21381
rect 9949 21322 10029 21335
rect 10133 21381 10213 21414
rect 10133 21335 10146 21381
rect 10200 21335 10213 21381
rect 10133 21322 10213 21335
rect 12321 21693 12401 21706
rect 12321 21647 12334 21693
rect 12388 21647 12401 21693
rect 12321 21614 12401 21647
rect 12505 21693 12585 21706
rect 12505 21647 12518 21693
rect 12572 21647 12585 21693
rect 12505 21614 12585 21647
rect 12689 21693 12769 21706
rect 12689 21647 12702 21693
rect 12756 21647 12769 21693
rect 12689 21614 12769 21647
rect 12321 21381 12401 21414
rect 12321 21335 12334 21381
rect 12388 21335 12401 21381
rect 12321 21322 12401 21335
rect 12505 21381 12585 21414
rect 12505 21335 12518 21381
rect 12572 21335 12585 21381
rect 12505 21322 12585 21335
rect 12689 21381 12769 21414
rect 12689 21335 12702 21381
rect 12756 21335 12769 21381
rect 12689 21322 12769 21335
rect 13807 21693 13887 21706
rect 13807 21647 13820 21693
rect 13874 21647 13887 21693
rect 13807 21614 13887 21647
rect 13991 21693 14071 21706
rect 13991 21647 14004 21693
rect 14058 21647 14071 21693
rect 13991 21614 14071 21647
rect 14175 21693 14255 21706
rect 14175 21647 14188 21693
rect 14242 21647 14255 21693
rect 14175 21614 14255 21647
rect 13807 21381 13887 21414
rect 13807 21335 13820 21381
rect 13874 21335 13887 21381
rect 13807 21322 13887 21335
rect 13991 21381 14071 21414
rect 13991 21335 14004 21381
rect 14058 21335 14071 21381
rect 13991 21322 14071 21335
rect 14175 21381 14255 21414
rect 14175 21335 14188 21381
rect 14242 21335 14255 21381
rect 14175 21322 14255 21335
rect 16363 21693 16443 21706
rect 16363 21647 16376 21693
rect 16430 21647 16443 21693
rect 16363 21614 16443 21647
rect 16547 21693 16627 21706
rect 16547 21647 16560 21693
rect 16614 21647 16627 21693
rect 16547 21614 16627 21647
rect 16731 21693 16811 21706
rect 16731 21647 16744 21693
rect 16798 21647 16811 21693
rect 16731 21614 16811 21647
rect 16363 21381 16443 21414
rect 16363 21335 16376 21381
rect 16430 21335 16443 21381
rect 16363 21322 16443 21335
rect 16547 21381 16627 21414
rect 16547 21335 16560 21381
rect 16614 21335 16627 21381
rect 16547 21322 16627 21335
rect 16731 21381 16811 21414
rect 16731 21335 16744 21381
rect 16798 21335 16811 21381
rect 16731 21322 16811 21335
rect 17849 21693 17929 21706
rect 17849 21647 17862 21693
rect 17916 21647 17929 21693
rect 17849 21614 17929 21647
rect 18033 21693 18113 21706
rect 18033 21647 18046 21693
rect 18100 21647 18113 21693
rect 18033 21614 18113 21647
rect 18217 21693 18297 21706
rect 18217 21647 18230 21693
rect 18284 21647 18297 21693
rect 18217 21614 18297 21647
rect 17849 21381 17929 21414
rect 17849 21335 17862 21381
rect 17916 21335 17929 21381
rect 17849 21322 17929 21335
rect 18033 21381 18113 21414
rect 18033 21335 18046 21381
rect 18100 21335 18113 21381
rect 18033 21322 18113 21335
rect 18217 21381 18297 21414
rect 18217 21335 18230 21381
rect 18284 21335 18297 21381
rect 18217 21322 18297 21335
rect -7889 20651 -7809 20664
rect -7889 20605 -7876 20651
rect -7822 20605 -7809 20651
rect -7889 20572 -7809 20605
rect -7705 20651 -7625 20664
rect -7705 20605 -7692 20651
rect -7638 20605 -7625 20651
rect -7705 20572 -7625 20605
rect -7521 20651 -7441 20664
rect -7521 20605 -7508 20651
rect -7454 20605 -7441 20651
rect -7521 20572 -7441 20605
rect -7889 20039 -7809 20072
rect -7889 19993 -7876 20039
rect -7822 19993 -7809 20039
rect -7889 19980 -7809 19993
rect -7705 20039 -7625 20072
rect -7705 19993 -7692 20039
rect -7638 19993 -7625 20039
rect -7705 19980 -7625 19993
rect -7521 20039 -7441 20072
rect -7521 19993 -7508 20039
rect -7454 19993 -7441 20039
rect -7521 19980 -7441 19993
rect -6403 20652 -6323 20665
rect -6403 20606 -6390 20652
rect -6336 20606 -6323 20652
rect -6403 20573 -6323 20606
rect -6219 20652 -6139 20665
rect -6219 20606 -6206 20652
rect -6152 20606 -6139 20652
rect -6219 20573 -6139 20606
rect -6035 20652 -5955 20665
rect -6035 20606 -6022 20652
rect -5968 20606 -5955 20652
rect -6035 20573 -5955 20606
rect -6403 20040 -6323 20073
rect -6403 19994 -6390 20040
rect -6336 19994 -6323 20040
rect -6403 19981 -6323 19994
rect -6219 20040 -6139 20073
rect -6219 19994 -6206 20040
rect -6152 19994 -6139 20040
rect -6219 19981 -6139 19994
rect -6035 20040 -5955 20073
rect -6035 19994 -6022 20040
rect -5968 19994 -5955 20040
rect -6035 19981 -5955 19994
rect -3847 20648 -3767 20661
rect -3847 20602 -3834 20648
rect -3780 20602 -3767 20648
rect -3847 20569 -3767 20602
rect -3663 20648 -3583 20661
rect -3663 20602 -3650 20648
rect -3596 20602 -3583 20648
rect -3663 20569 -3583 20602
rect -3479 20648 -3399 20661
rect -3479 20602 -3466 20648
rect -3412 20602 -3399 20648
rect -3479 20569 -3399 20602
rect -3847 20036 -3767 20069
rect -3847 19990 -3834 20036
rect -3780 19990 -3767 20036
rect -3847 19977 -3767 19990
rect -3663 20036 -3583 20069
rect -3663 19990 -3650 20036
rect -3596 19990 -3583 20036
rect -3663 19977 -3583 19990
rect -3479 20036 -3399 20069
rect -3479 19990 -3466 20036
rect -3412 19990 -3399 20036
rect -3479 19977 -3399 19990
rect -2361 20649 -2281 20662
rect -2361 20603 -2348 20649
rect -2294 20603 -2281 20649
rect -2361 20570 -2281 20603
rect -2177 20649 -2097 20662
rect -2177 20603 -2164 20649
rect -2110 20603 -2097 20649
rect -2177 20570 -2097 20603
rect -1993 20649 -1913 20662
rect -1993 20603 -1980 20649
rect -1926 20603 -1913 20649
rect -1993 20570 -1913 20603
rect -2361 20037 -2281 20070
rect -2361 19991 -2348 20037
rect -2294 19991 -2281 20037
rect -2361 19978 -2281 19991
rect -2177 20037 -2097 20070
rect -2177 19991 -2164 20037
rect -2110 19991 -2097 20037
rect -2177 19978 -2097 19991
rect -1993 20037 -1913 20070
rect -1993 19991 -1980 20037
rect -1926 19991 -1913 20037
rect -1993 19978 -1913 19991
rect 195 20648 275 20661
rect 195 20602 208 20648
rect 262 20602 275 20648
rect 195 20569 275 20602
rect 379 20648 459 20661
rect 379 20602 392 20648
rect 446 20602 459 20648
rect 379 20569 459 20602
rect 563 20648 643 20661
rect 563 20602 576 20648
rect 630 20602 643 20648
rect 563 20569 643 20602
rect 195 20036 275 20069
rect 195 19990 208 20036
rect 262 19990 275 20036
rect 195 19977 275 19990
rect 379 20036 459 20069
rect 379 19990 392 20036
rect 446 19990 459 20036
rect 379 19977 459 19990
rect 563 20036 643 20069
rect 563 19990 576 20036
rect 630 19990 643 20036
rect 563 19977 643 19990
rect 1681 20649 1761 20662
rect 1681 20603 1694 20649
rect 1748 20603 1761 20649
rect 1681 20570 1761 20603
rect 1865 20649 1945 20662
rect 1865 20603 1878 20649
rect 1932 20603 1945 20649
rect 1865 20570 1945 20603
rect 2049 20649 2129 20662
rect 2049 20603 2062 20649
rect 2116 20603 2129 20649
rect 2049 20570 2129 20603
rect 1681 20037 1761 20070
rect 1681 19991 1694 20037
rect 1748 19991 1761 20037
rect 1681 19978 1761 19991
rect 1865 20037 1945 20070
rect 1865 19991 1878 20037
rect 1932 19991 1945 20037
rect 1865 19978 1945 19991
rect 2049 20037 2129 20070
rect 2049 19991 2062 20037
rect 2116 19991 2129 20037
rect 2049 19978 2129 19991
rect 4237 20648 4317 20661
rect 4237 20602 4250 20648
rect 4304 20602 4317 20648
rect 4237 20569 4317 20602
rect 4421 20648 4501 20661
rect 4421 20602 4434 20648
rect 4488 20602 4501 20648
rect 4421 20569 4501 20602
rect 4605 20648 4685 20661
rect 4605 20602 4618 20648
rect 4672 20602 4685 20648
rect 4605 20569 4685 20602
rect 4237 20036 4317 20069
rect 4237 19990 4250 20036
rect 4304 19990 4317 20036
rect 4237 19977 4317 19990
rect 4421 20036 4501 20069
rect 4421 19990 4434 20036
rect 4488 19990 4501 20036
rect 4421 19977 4501 19990
rect 4605 20036 4685 20069
rect 4605 19990 4618 20036
rect 4672 19990 4685 20036
rect 4605 19977 4685 19990
rect 5723 20649 5803 20662
rect 5723 20603 5736 20649
rect 5790 20603 5803 20649
rect 5723 20570 5803 20603
rect 5907 20649 5987 20662
rect 5907 20603 5920 20649
rect 5974 20603 5987 20649
rect 5907 20570 5987 20603
rect 6091 20649 6171 20662
rect 6091 20603 6104 20649
rect 6158 20603 6171 20649
rect 6091 20570 6171 20603
rect 5723 20037 5803 20070
rect 5723 19991 5736 20037
rect 5790 19991 5803 20037
rect 5723 19978 5803 19991
rect 5907 20037 5987 20070
rect 5907 19991 5920 20037
rect 5974 19991 5987 20037
rect 5907 19978 5987 19991
rect 6091 20037 6171 20070
rect 6091 19991 6104 20037
rect 6158 19991 6171 20037
rect 6091 19978 6171 19991
rect 8279 20648 8359 20661
rect 8279 20602 8292 20648
rect 8346 20602 8359 20648
rect 8279 20569 8359 20602
rect 8463 20648 8543 20661
rect 8463 20602 8476 20648
rect 8530 20602 8543 20648
rect 8463 20569 8543 20602
rect 8647 20648 8727 20661
rect 8647 20602 8660 20648
rect 8714 20602 8727 20648
rect 8647 20569 8727 20602
rect 8279 20036 8359 20069
rect 8279 19990 8292 20036
rect 8346 19990 8359 20036
rect 8279 19977 8359 19990
rect 8463 20036 8543 20069
rect 8463 19990 8476 20036
rect 8530 19990 8543 20036
rect 8463 19977 8543 19990
rect 8647 20036 8727 20069
rect 8647 19990 8660 20036
rect 8714 19990 8727 20036
rect 8647 19977 8727 19990
rect 9765 20649 9845 20662
rect 9765 20603 9778 20649
rect 9832 20603 9845 20649
rect 9765 20570 9845 20603
rect 9949 20649 10029 20662
rect 9949 20603 9962 20649
rect 10016 20603 10029 20649
rect 9949 20570 10029 20603
rect 10133 20649 10213 20662
rect 10133 20603 10146 20649
rect 10200 20603 10213 20649
rect 10133 20570 10213 20603
rect 9765 20037 9845 20070
rect 9765 19991 9778 20037
rect 9832 19991 9845 20037
rect 9765 19978 9845 19991
rect 9949 20037 10029 20070
rect 9949 19991 9962 20037
rect 10016 19991 10029 20037
rect 9949 19978 10029 19991
rect 10133 20037 10213 20070
rect 10133 19991 10146 20037
rect 10200 19991 10213 20037
rect 10133 19978 10213 19991
rect 12321 20648 12401 20661
rect 12321 20602 12334 20648
rect 12388 20602 12401 20648
rect 12321 20569 12401 20602
rect 12505 20648 12585 20661
rect 12505 20602 12518 20648
rect 12572 20602 12585 20648
rect 12505 20569 12585 20602
rect 12689 20648 12769 20661
rect 12689 20602 12702 20648
rect 12756 20602 12769 20648
rect 12689 20569 12769 20602
rect 12321 20036 12401 20069
rect 12321 19990 12334 20036
rect 12388 19990 12401 20036
rect 12321 19977 12401 19990
rect 12505 20036 12585 20069
rect 12505 19990 12518 20036
rect 12572 19990 12585 20036
rect 12505 19977 12585 19990
rect 12689 20036 12769 20069
rect 12689 19990 12702 20036
rect 12756 19990 12769 20036
rect 12689 19977 12769 19990
rect 13807 20649 13887 20662
rect 13807 20603 13820 20649
rect 13874 20603 13887 20649
rect 13807 20570 13887 20603
rect 13991 20649 14071 20662
rect 13991 20603 14004 20649
rect 14058 20603 14071 20649
rect 13991 20570 14071 20603
rect 14175 20649 14255 20662
rect 14175 20603 14188 20649
rect 14242 20603 14255 20649
rect 14175 20570 14255 20603
rect 13807 20037 13887 20070
rect 13807 19991 13820 20037
rect 13874 19991 13887 20037
rect 13807 19978 13887 19991
rect 13991 20037 14071 20070
rect 13991 19991 14004 20037
rect 14058 19991 14071 20037
rect 13991 19978 14071 19991
rect 14175 20037 14255 20070
rect 14175 19991 14188 20037
rect 14242 19991 14255 20037
rect 14175 19978 14255 19991
rect 16363 20648 16443 20661
rect 16363 20602 16376 20648
rect 16430 20602 16443 20648
rect 16363 20569 16443 20602
rect 16547 20648 16627 20661
rect 16547 20602 16560 20648
rect 16614 20602 16627 20648
rect 16547 20569 16627 20602
rect 16731 20648 16811 20661
rect 16731 20602 16744 20648
rect 16798 20602 16811 20648
rect 16731 20569 16811 20602
rect 16363 20036 16443 20069
rect 16363 19990 16376 20036
rect 16430 19990 16443 20036
rect 16363 19977 16443 19990
rect 16547 20036 16627 20069
rect 16547 19990 16560 20036
rect 16614 19990 16627 20036
rect 16547 19977 16627 19990
rect 16731 20036 16811 20069
rect 16731 19990 16744 20036
rect 16798 19990 16811 20036
rect 16731 19977 16811 19990
rect 17849 20649 17929 20662
rect 17849 20603 17862 20649
rect 17916 20603 17929 20649
rect 17849 20570 17929 20603
rect 18033 20649 18113 20662
rect 18033 20603 18046 20649
rect 18100 20603 18113 20649
rect 18033 20570 18113 20603
rect 18217 20649 18297 20662
rect 18217 20603 18230 20649
rect 18284 20603 18297 20649
rect 18217 20570 18297 20603
rect 17849 20037 17929 20070
rect 17849 19991 17862 20037
rect 17916 19991 17929 20037
rect 17849 19978 17929 19991
rect 18033 20037 18113 20070
rect 18033 19991 18046 20037
rect 18100 19991 18113 20037
rect 18033 19978 18113 19991
rect 18217 20037 18297 20070
rect 18217 19991 18230 20037
rect 18284 19991 18297 20037
rect 18217 19978 18297 19991
rect -7889 19491 -7809 19504
rect -7889 19445 -7876 19491
rect -7822 19445 -7809 19491
rect -7889 19412 -7809 19445
rect -7705 19491 -7625 19504
rect -7705 19445 -7692 19491
rect -7638 19445 -7625 19491
rect -7705 19412 -7625 19445
rect -7521 19491 -7441 19504
rect -7521 19445 -7508 19491
rect -7454 19445 -7441 19491
rect -7521 19412 -7441 19445
rect -7889 19179 -7809 19212
rect -7889 19133 -7876 19179
rect -7822 19133 -7809 19179
rect -7889 19120 -7809 19133
rect -7705 19179 -7625 19212
rect -7705 19133 -7692 19179
rect -7638 19133 -7625 19179
rect -7705 19120 -7625 19133
rect -7521 19179 -7441 19212
rect -7521 19133 -7508 19179
rect -7454 19133 -7441 19179
rect -7521 19120 -7441 19133
rect -6403 19492 -6323 19505
rect -6403 19446 -6390 19492
rect -6336 19446 -6323 19492
rect -6403 19413 -6323 19446
rect -6219 19492 -6139 19505
rect -6219 19446 -6206 19492
rect -6152 19446 -6139 19492
rect -6219 19413 -6139 19446
rect -6035 19492 -5955 19505
rect -6035 19446 -6022 19492
rect -5968 19446 -5955 19492
rect -6035 19413 -5955 19446
rect -6403 19180 -6323 19213
rect -6403 19134 -6390 19180
rect -6336 19134 -6323 19180
rect -6403 19121 -6323 19134
rect -6219 19180 -6139 19213
rect -6219 19134 -6206 19180
rect -6152 19134 -6139 19180
rect -6219 19121 -6139 19134
rect -6035 19180 -5955 19213
rect -6035 19134 -6022 19180
rect -5968 19134 -5955 19180
rect -6035 19121 -5955 19134
rect -3847 19488 -3767 19501
rect -3847 19442 -3834 19488
rect -3780 19442 -3767 19488
rect -3847 19409 -3767 19442
rect -3663 19488 -3583 19501
rect -3663 19442 -3650 19488
rect -3596 19442 -3583 19488
rect -3663 19409 -3583 19442
rect -3479 19488 -3399 19501
rect -3479 19442 -3466 19488
rect -3412 19442 -3399 19488
rect -3479 19409 -3399 19442
rect -3847 19176 -3767 19209
rect -3847 19130 -3834 19176
rect -3780 19130 -3767 19176
rect -3847 19117 -3767 19130
rect -3663 19176 -3583 19209
rect -3663 19130 -3650 19176
rect -3596 19130 -3583 19176
rect -3663 19117 -3583 19130
rect -3479 19176 -3399 19209
rect -3479 19130 -3466 19176
rect -3412 19130 -3399 19176
rect -3479 19117 -3399 19130
rect -2361 19489 -2281 19502
rect -2361 19443 -2348 19489
rect -2294 19443 -2281 19489
rect -2361 19410 -2281 19443
rect -2177 19489 -2097 19502
rect -2177 19443 -2164 19489
rect -2110 19443 -2097 19489
rect -2177 19410 -2097 19443
rect -1993 19489 -1913 19502
rect -1993 19443 -1980 19489
rect -1926 19443 -1913 19489
rect -1993 19410 -1913 19443
rect -2361 19177 -2281 19210
rect -2361 19131 -2348 19177
rect -2294 19131 -2281 19177
rect -2361 19118 -2281 19131
rect -2177 19177 -2097 19210
rect -2177 19131 -2164 19177
rect -2110 19131 -2097 19177
rect -2177 19118 -2097 19131
rect -1993 19177 -1913 19210
rect -1993 19131 -1980 19177
rect -1926 19131 -1913 19177
rect -1993 19118 -1913 19131
rect 195 19488 275 19501
rect 195 19442 208 19488
rect 262 19442 275 19488
rect 195 19409 275 19442
rect 379 19488 459 19501
rect 379 19442 392 19488
rect 446 19442 459 19488
rect 379 19409 459 19442
rect 563 19488 643 19501
rect 563 19442 576 19488
rect 630 19442 643 19488
rect 563 19409 643 19442
rect 195 19176 275 19209
rect 195 19130 208 19176
rect 262 19130 275 19176
rect 195 19117 275 19130
rect 379 19176 459 19209
rect 379 19130 392 19176
rect 446 19130 459 19176
rect 379 19117 459 19130
rect 563 19176 643 19209
rect 563 19130 576 19176
rect 630 19130 643 19176
rect 563 19117 643 19130
rect 1681 19489 1761 19502
rect 1681 19443 1694 19489
rect 1748 19443 1761 19489
rect 1681 19410 1761 19443
rect 1865 19489 1945 19502
rect 1865 19443 1878 19489
rect 1932 19443 1945 19489
rect 1865 19410 1945 19443
rect 2049 19489 2129 19502
rect 2049 19443 2062 19489
rect 2116 19443 2129 19489
rect 2049 19410 2129 19443
rect 1681 19177 1761 19210
rect 1681 19131 1694 19177
rect 1748 19131 1761 19177
rect 1681 19118 1761 19131
rect 1865 19177 1945 19210
rect 1865 19131 1878 19177
rect 1932 19131 1945 19177
rect 1865 19118 1945 19131
rect 2049 19177 2129 19210
rect 2049 19131 2062 19177
rect 2116 19131 2129 19177
rect 2049 19118 2129 19131
rect 4237 19488 4317 19501
rect 4237 19442 4250 19488
rect 4304 19442 4317 19488
rect 4237 19409 4317 19442
rect 4421 19488 4501 19501
rect 4421 19442 4434 19488
rect 4488 19442 4501 19488
rect 4421 19409 4501 19442
rect 4605 19488 4685 19501
rect 4605 19442 4618 19488
rect 4672 19442 4685 19488
rect 4605 19409 4685 19442
rect 4237 19176 4317 19209
rect 4237 19130 4250 19176
rect 4304 19130 4317 19176
rect 4237 19117 4317 19130
rect 4421 19176 4501 19209
rect 4421 19130 4434 19176
rect 4488 19130 4501 19176
rect 4421 19117 4501 19130
rect 4605 19176 4685 19209
rect 4605 19130 4618 19176
rect 4672 19130 4685 19176
rect 4605 19117 4685 19130
rect 5723 19489 5803 19502
rect 5723 19443 5736 19489
rect 5790 19443 5803 19489
rect 5723 19410 5803 19443
rect 5907 19489 5987 19502
rect 5907 19443 5920 19489
rect 5974 19443 5987 19489
rect 5907 19410 5987 19443
rect 6091 19489 6171 19502
rect 6091 19443 6104 19489
rect 6158 19443 6171 19489
rect 6091 19410 6171 19443
rect 5723 19177 5803 19210
rect 5723 19131 5736 19177
rect 5790 19131 5803 19177
rect 5723 19118 5803 19131
rect 5907 19177 5987 19210
rect 5907 19131 5920 19177
rect 5974 19131 5987 19177
rect 5907 19118 5987 19131
rect 6091 19177 6171 19210
rect 6091 19131 6104 19177
rect 6158 19131 6171 19177
rect 6091 19118 6171 19131
rect 8279 19488 8359 19501
rect 8279 19442 8292 19488
rect 8346 19442 8359 19488
rect 8279 19409 8359 19442
rect 8463 19488 8543 19501
rect 8463 19442 8476 19488
rect 8530 19442 8543 19488
rect 8463 19409 8543 19442
rect 8647 19488 8727 19501
rect 8647 19442 8660 19488
rect 8714 19442 8727 19488
rect 8647 19409 8727 19442
rect 8279 19176 8359 19209
rect 8279 19130 8292 19176
rect 8346 19130 8359 19176
rect 8279 19117 8359 19130
rect 8463 19176 8543 19209
rect 8463 19130 8476 19176
rect 8530 19130 8543 19176
rect 8463 19117 8543 19130
rect 8647 19176 8727 19209
rect 8647 19130 8660 19176
rect 8714 19130 8727 19176
rect 8647 19117 8727 19130
rect 9765 19489 9845 19502
rect 9765 19443 9778 19489
rect 9832 19443 9845 19489
rect 9765 19410 9845 19443
rect 9949 19489 10029 19502
rect 9949 19443 9962 19489
rect 10016 19443 10029 19489
rect 9949 19410 10029 19443
rect 10133 19489 10213 19502
rect 10133 19443 10146 19489
rect 10200 19443 10213 19489
rect 10133 19410 10213 19443
rect 9765 19177 9845 19210
rect 9765 19131 9778 19177
rect 9832 19131 9845 19177
rect 9765 19118 9845 19131
rect 9949 19177 10029 19210
rect 9949 19131 9962 19177
rect 10016 19131 10029 19177
rect 9949 19118 10029 19131
rect 10133 19177 10213 19210
rect 10133 19131 10146 19177
rect 10200 19131 10213 19177
rect 10133 19118 10213 19131
rect 12321 19488 12401 19501
rect 12321 19442 12334 19488
rect 12388 19442 12401 19488
rect 12321 19409 12401 19442
rect 12505 19488 12585 19501
rect 12505 19442 12518 19488
rect 12572 19442 12585 19488
rect 12505 19409 12585 19442
rect 12689 19488 12769 19501
rect 12689 19442 12702 19488
rect 12756 19442 12769 19488
rect 12689 19409 12769 19442
rect 12321 19176 12401 19209
rect 12321 19130 12334 19176
rect 12388 19130 12401 19176
rect 12321 19117 12401 19130
rect 12505 19176 12585 19209
rect 12505 19130 12518 19176
rect 12572 19130 12585 19176
rect 12505 19117 12585 19130
rect 12689 19176 12769 19209
rect 12689 19130 12702 19176
rect 12756 19130 12769 19176
rect 12689 19117 12769 19130
rect 13807 19489 13887 19502
rect 13807 19443 13820 19489
rect 13874 19443 13887 19489
rect 13807 19410 13887 19443
rect 13991 19489 14071 19502
rect 13991 19443 14004 19489
rect 14058 19443 14071 19489
rect 13991 19410 14071 19443
rect 14175 19489 14255 19502
rect 14175 19443 14188 19489
rect 14242 19443 14255 19489
rect 14175 19410 14255 19443
rect 13807 19177 13887 19210
rect 13807 19131 13820 19177
rect 13874 19131 13887 19177
rect 13807 19118 13887 19131
rect 13991 19177 14071 19210
rect 13991 19131 14004 19177
rect 14058 19131 14071 19177
rect 13991 19118 14071 19131
rect 14175 19177 14255 19210
rect 14175 19131 14188 19177
rect 14242 19131 14255 19177
rect 14175 19118 14255 19131
rect 16363 19488 16443 19501
rect 16363 19442 16376 19488
rect 16430 19442 16443 19488
rect 16363 19409 16443 19442
rect 16547 19488 16627 19501
rect 16547 19442 16560 19488
rect 16614 19442 16627 19488
rect 16547 19409 16627 19442
rect 16731 19488 16811 19501
rect 16731 19442 16744 19488
rect 16798 19442 16811 19488
rect 16731 19409 16811 19442
rect 16363 19176 16443 19209
rect 16363 19130 16376 19176
rect 16430 19130 16443 19176
rect 16363 19117 16443 19130
rect 16547 19176 16627 19209
rect 16547 19130 16560 19176
rect 16614 19130 16627 19176
rect 16547 19117 16627 19130
rect 16731 19176 16811 19209
rect 16731 19130 16744 19176
rect 16798 19130 16811 19176
rect 16731 19117 16811 19130
rect 17849 19489 17929 19502
rect 17849 19443 17862 19489
rect 17916 19443 17929 19489
rect 17849 19410 17929 19443
rect 18033 19489 18113 19502
rect 18033 19443 18046 19489
rect 18100 19443 18113 19489
rect 18033 19410 18113 19443
rect 18217 19489 18297 19502
rect 18217 19443 18230 19489
rect 18284 19443 18297 19489
rect 18217 19410 18297 19443
rect 17849 19177 17929 19210
rect 17849 19131 17862 19177
rect 17916 19131 17929 19177
rect 17849 19118 17929 19131
rect 18033 19177 18113 19210
rect 18033 19131 18046 19177
rect 18100 19131 18113 19177
rect 18033 19118 18113 19131
rect 18217 19177 18297 19210
rect 18217 19131 18230 19177
rect 18284 19131 18297 19177
rect 18217 19118 18297 19131
rect -7889 18446 -7809 18459
rect -7889 18400 -7876 18446
rect -7822 18400 -7809 18446
rect -7889 18367 -7809 18400
rect -7705 18446 -7625 18459
rect -7705 18400 -7692 18446
rect -7638 18400 -7625 18446
rect -7705 18367 -7625 18400
rect -7521 18446 -7441 18459
rect -7521 18400 -7508 18446
rect -7454 18400 -7441 18446
rect -7521 18367 -7441 18400
rect -7889 17834 -7809 17867
rect -7889 17788 -7876 17834
rect -7822 17788 -7809 17834
rect -7889 17775 -7809 17788
rect -7705 17834 -7625 17867
rect -7705 17788 -7692 17834
rect -7638 17788 -7625 17834
rect -7705 17775 -7625 17788
rect -7521 17834 -7441 17867
rect -7521 17788 -7508 17834
rect -7454 17788 -7441 17834
rect -7521 17775 -7441 17788
rect -3847 18443 -3767 18456
rect -3847 18397 -3834 18443
rect -3780 18397 -3767 18443
rect -3847 18364 -3767 18397
rect -3663 18443 -3583 18456
rect -3663 18397 -3650 18443
rect -3596 18397 -3583 18443
rect -3663 18364 -3583 18397
rect -3479 18443 -3399 18456
rect -3479 18397 -3466 18443
rect -3412 18397 -3399 18443
rect -3479 18364 -3399 18397
rect -3847 17831 -3767 17864
rect -3847 17785 -3834 17831
rect -3780 17785 -3767 17831
rect -3847 17772 -3767 17785
rect -3663 17831 -3583 17864
rect -3663 17785 -3650 17831
rect -3596 17785 -3583 17831
rect -3663 17772 -3583 17785
rect -3479 17831 -3399 17864
rect -3479 17785 -3466 17831
rect -3412 17785 -3399 17831
rect -3479 17772 -3399 17785
rect 195 18443 275 18456
rect 195 18397 208 18443
rect 262 18397 275 18443
rect 195 18364 275 18397
rect 379 18443 459 18456
rect 379 18397 392 18443
rect 446 18397 459 18443
rect 379 18364 459 18397
rect 563 18443 643 18456
rect 563 18397 576 18443
rect 630 18397 643 18443
rect 563 18364 643 18397
rect 195 17831 275 17864
rect 195 17785 208 17831
rect 262 17785 275 17831
rect 195 17772 275 17785
rect 379 17831 459 17864
rect 379 17785 392 17831
rect 446 17785 459 17831
rect 379 17772 459 17785
rect 563 17831 643 17864
rect 563 17785 576 17831
rect 630 17785 643 17831
rect 563 17772 643 17785
rect 4237 18443 4317 18456
rect 4237 18397 4250 18443
rect 4304 18397 4317 18443
rect 4237 18364 4317 18397
rect 4421 18443 4501 18456
rect 4421 18397 4434 18443
rect 4488 18397 4501 18443
rect 4421 18364 4501 18397
rect 4605 18443 4685 18456
rect 4605 18397 4618 18443
rect 4672 18397 4685 18443
rect 4605 18364 4685 18397
rect 4237 17831 4317 17864
rect 4237 17785 4250 17831
rect 4304 17785 4317 17831
rect 4237 17772 4317 17785
rect 4421 17831 4501 17864
rect 4421 17785 4434 17831
rect 4488 17785 4501 17831
rect 4421 17772 4501 17785
rect 4605 17831 4685 17864
rect 4605 17785 4618 17831
rect 4672 17785 4685 17831
rect 4605 17772 4685 17785
rect 8279 18443 8359 18456
rect 8279 18397 8292 18443
rect 8346 18397 8359 18443
rect 8279 18364 8359 18397
rect 8463 18443 8543 18456
rect 8463 18397 8476 18443
rect 8530 18397 8543 18443
rect 8463 18364 8543 18397
rect 8647 18443 8727 18456
rect 8647 18397 8660 18443
rect 8714 18397 8727 18443
rect 8647 18364 8727 18397
rect 8279 17831 8359 17864
rect 8279 17785 8292 17831
rect 8346 17785 8359 17831
rect 8279 17772 8359 17785
rect 8463 17831 8543 17864
rect 8463 17785 8476 17831
rect 8530 17785 8543 17831
rect 8463 17772 8543 17785
rect 8647 17831 8727 17864
rect 8647 17785 8660 17831
rect 8714 17785 8727 17831
rect 8647 17772 8727 17785
rect 12321 18443 12401 18456
rect 12321 18397 12334 18443
rect 12388 18397 12401 18443
rect 12321 18364 12401 18397
rect 12505 18443 12585 18456
rect 12505 18397 12518 18443
rect 12572 18397 12585 18443
rect 12505 18364 12585 18397
rect 12689 18443 12769 18456
rect 12689 18397 12702 18443
rect 12756 18397 12769 18443
rect 12689 18364 12769 18397
rect 12321 17831 12401 17864
rect 12321 17785 12334 17831
rect 12388 17785 12401 17831
rect 12321 17772 12401 17785
rect 12505 17831 12585 17864
rect 12505 17785 12518 17831
rect 12572 17785 12585 17831
rect 12505 17772 12585 17785
rect 12689 17831 12769 17864
rect 12689 17785 12702 17831
rect 12756 17785 12769 17831
rect 12689 17772 12769 17785
rect 16363 18443 16443 18456
rect 16363 18397 16376 18443
rect 16430 18397 16443 18443
rect 16363 18364 16443 18397
rect 16547 18443 16627 18456
rect 16547 18397 16560 18443
rect 16614 18397 16627 18443
rect 16547 18364 16627 18397
rect 16731 18443 16811 18456
rect 16731 18397 16744 18443
rect 16798 18397 16811 18443
rect 16731 18364 16811 18397
rect 16363 17831 16443 17864
rect 16363 17785 16376 17831
rect 16430 17785 16443 17831
rect 16363 17772 16443 17785
rect 16547 17831 16627 17864
rect 16547 17785 16560 17831
rect 16614 17785 16627 17831
rect 16547 17772 16627 17785
rect 16731 17831 16811 17864
rect 16731 17785 16744 17831
rect 16798 17785 16811 17831
rect 16731 17772 16811 17785
rect -7889 17286 -7809 17299
rect -7889 17240 -7876 17286
rect -7822 17240 -7809 17286
rect -7889 17207 -7809 17240
rect -7705 17286 -7625 17299
rect -7705 17240 -7692 17286
rect -7638 17240 -7625 17286
rect -7705 17207 -7625 17240
rect -7521 17286 -7441 17299
rect -7521 17240 -7508 17286
rect -7454 17240 -7441 17286
rect -7521 17207 -7441 17240
rect -7889 16974 -7809 17007
rect -7889 16928 -7876 16974
rect -7822 16928 -7809 16974
rect -7889 16915 -7809 16928
rect -7705 16974 -7625 17007
rect -7705 16928 -7692 16974
rect -7638 16928 -7625 16974
rect -7705 16915 -7625 16928
rect -7521 16974 -7441 17007
rect -7521 16928 -7508 16974
rect -7454 16928 -7441 16974
rect -7521 16915 -7441 16928
rect -3847 17283 -3767 17296
rect -3847 17237 -3834 17283
rect -3780 17237 -3767 17283
rect -3847 17204 -3767 17237
rect -3663 17283 -3583 17296
rect -3663 17237 -3650 17283
rect -3596 17237 -3583 17283
rect -3663 17204 -3583 17237
rect -3479 17283 -3399 17296
rect -3479 17237 -3466 17283
rect -3412 17237 -3399 17283
rect -3479 17204 -3399 17237
rect -3847 16971 -3767 17004
rect -3847 16925 -3834 16971
rect -3780 16925 -3767 16971
rect -3847 16912 -3767 16925
rect -3663 16971 -3583 17004
rect -3663 16925 -3650 16971
rect -3596 16925 -3583 16971
rect -3663 16912 -3583 16925
rect -3479 16971 -3399 17004
rect -3479 16925 -3466 16971
rect -3412 16925 -3399 16971
rect -3479 16912 -3399 16925
rect 195 17283 275 17296
rect 195 17237 208 17283
rect 262 17237 275 17283
rect 195 17204 275 17237
rect 379 17283 459 17296
rect 379 17237 392 17283
rect 446 17237 459 17283
rect 379 17204 459 17237
rect 563 17283 643 17296
rect 563 17237 576 17283
rect 630 17237 643 17283
rect 563 17204 643 17237
rect 195 16971 275 17004
rect 195 16925 208 16971
rect 262 16925 275 16971
rect 195 16912 275 16925
rect 379 16971 459 17004
rect 379 16925 392 16971
rect 446 16925 459 16971
rect 379 16912 459 16925
rect 563 16971 643 17004
rect 563 16925 576 16971
rect 630 16925 643 16971
rect 563 16912 643 16925
rect 4237 17283 4317 17296
rect 4237 17237 4250 17283
rect 4304 17237 4317 17283
rect 4237 17204 4317 17237
rect 4421 17283 4501 17296
rect 4421 17237 4434 17283
rect 4488 17237 4501 17283
rect 4421 17204 4501 17237
rect 4605 17283 4685 17296
rect 4605 17237 4618 17283
rect 4672 17237 4685 17283
rect 4605 17204 4685 17237
rect 4237 16971 4317 17004
rect 4237 16925 4250 16971
rect 4304 16925 4317 16971
rect 4237 16912 4317 16925
rect 4421 16971 4501 17004
rect 4421 16925 4434 16971
rect 4488 16925 4501 16971
rect 4421 16912 4501 16925
rect 4605 16971 4685 17004
rect 4605 16925 4618 16971
rect 4672 16925 4685 16971
rect 4605 16912 4685 16925
rect 8279 17283 8359 17296
rect 8279 17237 8292 17283
rect 8346 17237 8359 17283
rect 8279 17204 8359 17237
rect 8463 17283 8543 17296
rect 8463 17237 8476 17283
rect 8530 17237 8543 17283
rect 8463 17204 8543 17237
rect 8647 17283 8727 17296
rect 8647 17237 8660 17283
rect 8714 17237 8727 17283
rect 8647 17204 8727 17237
rect 8279 16971 8359 17004
rect 8279 16925 8292 16971
rect 8346 16925 8359 16971
rect 8279 16912 8359 16925
rect 8463 16971 8543 17004
rect 8463 16925 8476 16971
rect 8530 16925 8543 16971
rect 8463 16912 8543 16925
rect 8647 16971 8727 17004
rect 8647 16925 8660 16971
rect 8714 16925 8727 16971
rect 8647 16912 8727 16925
rect 12321 17283 12401 17296
rect 12321 17237 12334 17283
rect 12388 17237 12401 17283
rect 12321 17204 12401 17237
rect 12505 17283 12585 17296
rect 12505 17237 12518 17283
rect 12572 17237 12585 17283
rect 12505 17204 12585 17237
rect 12689 17283 12769 17296
rect 12689 17237 12702 17283
rect 12756 17237 12769 17283
rect 12689 17204 12769 17237
rect 12321 16971 12401 17004
rect 12321 16925 12334 16971
rect 12388 16925 12401 16971
rect 12321 16912 12401 16925
rect 12505 16971 12585 17004
rect 12505 16925 12518 16971
rect 12572 16925 12585 16971
rect 12505 16912 12585 16925
rect 12689 16971 12769 17004
rect 12689 16925 12702 16971
rect 12756 16925 12769 16971
rect 12689 16912 12769 16925
rect 16363 17283 16443 17296
rect 16363 17237 16376 17283
rect 16430 17237 16443 17283
rect 16363 17204 16443 17237
rect 16547 17283 16627 17296
rect 16547 17237 16560 17283
rect 16614 17237 16627 17283
rect 16547 17204 16627 17237
rect 16731 17283 16811 17296
rect 16731 17237 16744 17283
rect 16798 17237 16811 17283
rect 16731 17204 16811 17237
rect 16363 16971 16443 17004
rect 16363 16925 16376 16971
rect 16430 16925 16443 16971
rect 16363 16912 16443 16925
rect 16547 16971 16627 17004
rect 16547 16925 16560 16971
rect 16614 16925 16627 16971
rect 16547 16912 16627 16925
rect 16731 16971 16811 17004
rect 16731 16925 16744 16971
rect 16798 16925 16811 16971
rect 16731 16912 16811 16925
rect -11901 15482 -11821 15495
rect -11901 15436 -11888 15482
rect -11834 15436 -11821 15482
rect -11901 15403 -11821 15436
rect -11717 15482 -11637 15495
rect -11717 15436 -11704 15482
rect -11650 15436 -11637 15482
rect -11717 15403 -11637 15436
rect -11533 15482 -11453 15495
rect -11533 15436 -11520 15482
rect -11466 15436 -11453 15482
rect -11533 15403 -11453 15436
rect -11901 14870 -11821 14903
rect -11901 14824 -11888 14870
rect -11834 14824 -11821 14870
rect -11901 14811 -11821 14824
rect -11717 14870 -11637 14903
rect -11717 14824 -11704 14870
rect -11650 14824 -11637 14870
rect -11717 14811 -11637 14824
rect -11533 14870 -11453 14903
rect -11533 14824 -11520 14870
rect -11466 14824 -11453 14870
rect -11533 14811 -11453 14824
rect -7889 15482 -7809 15495
rect -7889 15436 -7876 15482
rect -7822 15436 -7809 15482
rect -7889 15403 -7809 15436
rect -7705 15482 -7625 15495
rect -7705 15436 -7692 15482
rect -7638 15436 -7625 15482
rect -7705 15403 -7625 15436
rect -7521 15482 -7441 15495
rect -7521 15436 -7508 15482
rect -7454 15436 -7441 15482
rect -7521 15403 -7441 15436
rect -7889 14870 -7809 14903
rect -7889 14824 -7876 14870
rect -7822 14824 -7809 14870
rect -7889 14811 -7809 14824
rect -7705 14870 -7625 14903
rect -7705 14824 -7692 14870
rect -7638 14824 -7625 14870
rect -7705 14811 -7625 14824
rect -7521 14870 -7441 14903
rect -7521 14824 -7508 14870
rect -7454 14824 -7441 14870
rect -7521 14811 -7441 14824
rect -3847 15482 -3767 15495
rect -3847 15436 -3834 15482
rect -3780 15436 -3767 15482
rect -3847 15403 -3767 15436
rect -3663 15482 -3583 15495
rect -3663 15436 -3650 15482
rect -3596 15436 -3583 15482
rect -3663 15403 -3583 15436
rect -3479 15482 -3399 15495
rect -3479 15436 -3466 15482
rect -3412 15436 -3399 15482
rect -3479 15403 -3399 15436
rect -3847 14870 -3767 14903
rect -3847 14824 -3834 14870
rect -3780 14824 -3767 14870
rect -3847 14811 -3767 14824
rect -3663 14870 -3583 14903
rect -3663 14824 -3650 14870
rect -3596 14824 -3583 14870
rect -3663 14811 -3583 14824
rect -3479 14870 -3399 14903
rect -3479 14824 -3466 14870
rect -3412 14824 -3399 14870
rect -3479 14811 -3399 14824
rect 195 15482 275 15495
rect 195 15436 208 15482
rect 262 15436 275 15482
rect 195 15403 275 15436
rect 379 15482 459 15495
rect 379 15436 392 15482
rect 446 15436 459 15482
rect 379 15403 459 15436
rect 563 15482 643 15495
rect 563 15436 576 15482
rect 630 15436 643 15482
rect 563 15403 643 15436
rect 195 14870 275 14903
rect 195 14824 208 14870
rect 262 14824 275 14870
rect 195 14811 275 14824
rect 379 14870 459 14903
rect 379 14824 392 14870
rect 446 14824 459 14870
rect 379 14811 459 14824
rect 563 14870 643 14903
rect 563 14824 576 14870
rect 630 14824 643 14870
rect 563 14811 643 14824
rect 4237 15482 4317 15495
rect 4237 15436 4250 15482
rect 4304 15436 4317 15482
rect 4237 15403 4317 15436
rect 4421 15482 4501 15495
rect 4421 15436 4434 15482
rect 4488 15436 4501 15482
rect 4421 15403 4501 15436
rect 4605 15482 4685 15495
rect 4605 15436 4618 15482
rect 4672 15436 4685 15482
rect 4605 15403 4685 15436
rect 4237 14870 4317 14903
rect 4237 14824 4250 14870
rect 4304 14824 4317 14870
rect 4237 14811 4317 14824
rect 4421 14870 4501 14903
rect 4421 14824 4434 14870
rect 4488 14824 4501 14870
rect 4421 14811 4501 14824
rect 4605 14870 4685 14903
rect 4605 14824 4618 14870
rect 4672 14824 4685 14870
rect 4605 14811 4685 14824
rect 8279 15482 8359 15495
rect 8279 15436 8292 15482
rect 8346 15436 8359 15482
rect 8279 15403 8359 15436
rect 8463 15482 8543 15495
rect 8463 15436 8476 15482
rect 8530 15436 8543 15482
rect 8463 15403 8543 15436
rect 8647 15482 8727 15495
rect 8647 15436 8660 15482
rect 8714 15436 8727 15482
rect 8647 15403 8727 15436
rect 8279 14870 8359 14903
rect 8279 14824 8292 14870
rect 8346 14824 8359 14870
rect 8279 14811 8359 14824
rect 8463 14870 8543 14903
rect 8463 14824 8476 14870
rect 8530 14824 8543 14870
rect 8463 14811 8543 14824
rect 8647 14870 8727 14903
rect 8647 14824 8660 14870
rect 8714 14824 8727 14870
rect 8647 14811 8727 14824
rect 12321 15482 12401 15495
rect 12321 15436 12334 15482
rect 12388 15436 12401 15482
rect 12321 15403 12401 15436
rect 12505 15482 12585 15495
rect 12505 15436 12518 15482
rect 12572 15436 12585 15482
rect 12505 15403 12585 15436
rect 12689 15482 12769 15495
rect 12689 15436 12702 15482
rect 12756 15436 12769 15482
rect 12689 15403 12769 15436
rect 12321 14870 12401 14903
rect 12321 14824 12334 14870
rect 12388 14824 12401 14870
rect 12321 14811 12401 14824
rect 12505 14870 12585 14903
rect 12505 14824 12518 14870
rect 12572 14824 12585 14870
rect 12505 14811 12585 14824
rect 12689 14870 12769 14903
rect 12689 14824 12702 14870
rect 12756 14824 12769 14870
rect 12689 14811 12769 14824
rect -11901 14322 -11821 14335
rect -11901 14276 -11888 14322
rect -11834 14276 -11821 14322
rect -11901 14243 -11821 14276
rect -11717 14322 -11637 14335
rect -11717 14276 -11704 14322
rect -11650 14276 -11637 14322
rect -11717 14243 -11637 14276
rect -11533 14322 -11453 14335
rect -11533 14276 -11520 14322
rect -11466 14276 -11453 14322
rect -11533 14243 -11453 14276
rect -11901 14010 -11821 14043
rect -11901 13964 -11888 14010
rect -11834 13964 -11821 14010
rect -11901 13951 -11821 13964
rect -11717 14010 -11637 14043
rect -11717 13964 -11704 14010
rect -11650 13964 -11637 14010
rect -11717 13951 -11637 13964
rect -11533 14010 -11453 14043
rect -11533 13964 -11520 14010
rect -11466 13964 -11453 14010
rect -11533 13951 -11453 13964
rect -7889 14322 -7809 14335
rect -7889 14276 -7876 14322
rect -7822 14276 -7809 14322
rect -7889 14243 -7809 14276
rect -7705 14322 -7625 14335
rect -7705 14276 -7692 14322
rect -7638 14276 -7625 14322
rect -7705 14243 -7625 14276
rect -7521 14322 -7441 14335
rect -7521 14276 -7508 14322
rect -7454 14276 -7441 14322
rect -7521 14243 -7441 14276
rect -7889 14010 -7809 14043
rect -7889 13964 -7876 14010
rect -7822 13964 -7809 14010
rect -7889 13951 -7809 13964
rect -7705 14010 -7625 14043
rect -7705 13964 -7692 14010
rect -7638 13964 -7625 14010
rect -7705 13951 -7625 13964
rect -7521 14010 -7441 14043
rect -7521 13964 -7508 14010
rect -7454 13964 -7441 14010
rect -7521 13951 -7441 13964
rect -3847 14322 -3767 14335
rect -3847 14276 -3834 14322
rect -3780 14276 -3767 14322
rect -3847 14243 -3767 14276
rect -3663 14322 -3583 14335
rect -3663 14276 -3650 14322
rect -3596 14276 -3583 14322
rect -3663 14243 -3583 14276
rect -3479 14322 -3399 14335
rect -3479 14276 -3466 14322
rect -3412 14276 -3399 14322
rect -3479 14243 -3399 14276
rect -3847 14010 -3767 14043
rect -3847 13964 -3834 14010
rect -3780 13964 -3767 14010
rect -3847 13951 -3767 13964
rect -3663 14010 -3583 14043
rect -3663 13964 -3650 14010
rect -3596 13964 -3583 14010
rect -3663 13951 -3583 13964
rect -3479 14010 -3399 14043
rect -3479 13964 -3466 14010
rect -3412 13964 -3399 14010
rect -3479 13951 -3399 13964
rect 195 14322 275 14335
rect 195 14276 208 14322
rect 262 14276 275 14322
rect 195 14243 275 14276
rect 379 14322 459 14335
rect 379 14276 392 14322
rect 446 14276 459 14322
rect 379 14243 459 14276
rect 563 14322 643 14335
rect 563 14276 576 14322
rect 630 14276 643 14322
rect 563 14243 643 14276
rect 195 14010 275 14043
rect 195 13964 208 14010
rect 262 13964 275 14010
rect 195 13951 275 13964
rect 379 14010 459 14043
rect 379 13964 392 14010
rect 446 13964 459 14010
rect 379 13951 459 13964
rect 563 14010 643 14043
rect 563 13964 576 14010
rect 630 13964 643 14010
rect 563 13951 643 13964
rect 4237 14322 4317 14335
rect 4237 14276 4250 14322
rect 4304 14276 4317 14322
rect 4237 14243 4317 14276
rect 4421 14322 4501 14335
rect 4421 14276 4434 14322
rect 4488 14276 4501 14322
rect 4421 14243 4501 14276
rect 4605 14322 4685 14335
rect 4605 14276 4618 14322
rect 4672 14276 4685 14322
rect 4605 14243 4685 14276
rect 4237 14010 4317 14043
rect 4237 13964 4250 14010
rect 4304 13964 4317 14010
rect 4237 13951 4317 13964
rect 4421 14010 4501 14043
rect 4421 13964 4434 14010
rect 4488 13964 4501 14010
rect 4421 13951 4501 13964
rect 4605 14010 4685 14043
rect 4605 13964 4618 14010
rect 4672 13964 4685 14010
rect 4605 13951 4685 13964
rect 8279 14322 8359 14335
rect 8279 14276 8292 14322
rect 8346 14276 8359 14322
rect 8279 14243 8359 14276
rect 8463 14322 8543 14335
rect 8463 14276 8476 14322
rect 8530 14276 8543 14322
rect 8463 14243 8543 14276
rect 8647 14322 8727 14335
rect 8647 14276 8660 14322
rect 8714 14276 8727 14322
rect 8647 14243 8727 14276
rect 8279 14010 8359 14043
rect 8279 13964 8292 14010
rect 8346 13964 8359 14010
rect 8279 13951 8359 13964
rect 8463 14010 8543 14043
rect 8463 13964 8476 14010
rect 8530 13964 8543 14010
rect 8463 13951 8543 13964
rect 8647 14010 8727 14043
rect 8647 13964 8660 14010
rect 8714 13964 8727 14010
rect 8647 13951 8727 13964
rect 12321 14322 12401 14335
rect 12321 14276 12334 14322
rect 12388 14276 12401 14322
rect 12321 14243 12401 14276
rect 12505 14322 12585 14335
rect 12505 14276 12518 14322
rect 12572 14276 12585 14322
rect 12505 14243 12585 14276
rect 12689 14322 12769 14335
rect 12689 14276 12702 14322
rect 12756 14276 12769 14322
rect 12689 14243 12769 14276
rect 12321 14010 12401 14043
rect 12321 13964 12334 14010
rect 12388 13964 12401 14010
rect 12321 13951 12401 13964
rect 12505 14010 12585 14043
rect 12505 13964 12518 14010
rect 12572 13964 12585 14010
rect 12505 13951 12585 13964
rect 12689 14010 12769 14043
rect 12689 13964 12702 14010
rect 12756 13964 12769 14010
rect 12689 13951 12769 13964
rect -11901 13277 -11821 13290
rect -11901 13231 -11888 13277
rect -11834 13231 -11821 13277
rect -11901 13198 -11821 13231
rect -11717 13277 -11637 13290
rect -11717 13231 -11704 13277
rect -11650 13231 -11637 13277
rect -11717 13198 -11637 13231
rect -11533 13277 -11453 13290
rect -11533 13231 -11520 13277
rect -11466 13231 -11453 13277
rect -11533 13198 -11453 13231
rect -11901 12665 -11821 12698
rect -11901 12619 -11888 12665
rect -11834 12619 -11821 12665
rect -11901 12606 -11821 12619
rect -11717 12665 -11637 12698
rect -11717 12619 -11704 12665
rect -11650 12619 -11637 12665
rect -11717 12606 -11637 12619
rect -11533 12665 -11453 12698
rect -11533 12619 -11520 12665
rect -11466 12619 -11453 12665
rect -11533 12606 -11453 12619
rect -10415 13277 -10335 13290
rect -10415 13231 -10402 13277
rect -10348 13231 -10335 13277
rect -10415 13198 -10335 13231
rect -10231 13277 -10151 13290
rect -10231 13231 -10218 13277
rect -10164 13231 -10151 13277
rect -10231 13198 -10151 13231
rect -10047 13277 -9967 13290
rect -10047 13231 -10034 13277
rect -9980 13231 -9967 13277
rect -10047 13198 -9967 13231
rect -10415 12665 -10335 12698
rect -10415 12619 -10402 12665
rect -10348 12619 -10335 12665
rect -10415 12606 -10335 12619
rect -10231 12665 -10151 12698
rect -10231 12619 -10218 12665
rect -10164 12619 -10151 12665
rect -10231 12606 -10151 12619
rect -10047 12665 -9967 12698
rect -10047 12619 -10034 12665
rect -9980 12619 -9967 12665
rect -10047 12606 -9967 12619
rect -7889 13277 -7809 13290
rect -7889 13231 -7876 13277
rect -7822 13231 -7809 13277
rect -7889 13198 -7809 13231
rect -7705 13277 -7625 13290
rect -7705 13231 -7692 13277
rect -7638 13231 -7625 13277
rect -7705 13198 -7625 13231
rect -7521 13277 -7441 13290
rect -7521 13231 -7508 13277
rect -7454 13231 -7441 13277
rect -7521 13198 -7441 13231
rect -7889 12665 -7809 12698
rect -7889 12619 -7876 12665
rect -7822 12619 -7809 12665
rect -7889 12606 -7809 12619
rect -7705 12665 -7625 12698
rect -7705 12619 -7692 12665
rect -7638 12619 -7625 12665
rect -7705 12606 -7625 12619
rect -7521 12665 -7441 12698
rect -7521 12619 -7508 12665
rect -7454 12619 -7441 12665
rect -7521 12606 -7441 12619
rect -6403 13277 -6323 13290
rect -6403 13231 -6390 13277
rect -6336 13231 -6323 13277
rect -6403 13198 -6323 13231
rect -6219 13277 -6139 13290
rect -6219 13231 -6206 13277
rect -6152 13231 -6139 13277
rect -6219 13198 -6139 13231
rect -6035 13277 -5955 13290
rect -6035 13231 -6022 13277
rect -5968 13231 -5955 13277
rect -6035 13198 -5955 13231
rect -6403 12665 -6323 12698
rect -6403 12619 -6390 12665
rect -6336 12619 -6323 12665
rect -6403 12606 -6323 12619
rect -6219 12665 -6139 12698
rect -6219 12619 -6206 12665
rect -6152 12619 -6139 12665
rect -6219 12606 -6139 12619
rect -6035 12665 -5955 12698
rect -6035 12619 -6022 12665
rect -5968 12619 -5955 12665
rect -6035 12606 -5955 12619
rect -3847 13277 -3767 13290
rect -3847 13231 -3834 13277
rect -3780 13231 -3767 13277
rect -3847 13198 -3767 13231
rect -3663 13277 -3583 13290
rect -3663 13231 -3650 13277
rect -3596 13231 -3583 13277
rect -3663 13198 -3583 13231
rect -3479 13277 -3399 13290
rect -3479 13231 -3466 13277
rect -3412 13231 -3399 13277
rect -3479 13198 -3399 13231
rect -3847 12665 -3767 12698
rect -3847 12619 -3834 12665
rect -3780 12619 -3767 12665
rect -3847 12606 -3767 12619
rect -3663 12665 -3583 12698
rect -3663 12619 -3650 12665
rect -3596 12619 -3583 12665
rect -3663 12606 -3583 12619
rect -3479 12665 -3399 12698
rect -3479 12619 -3466 12665
rect -3412 12619 -3399 12665
rect -3479 12606 -3399 12619
rect -2361 13277 -2281 13290
rect -2361 13231 -2348 13277
rect -2294 13231 -2281 13277
rect -2361 13198 -2281 13231
rect -2177 13277 -2097 13290
rect -2177 13231 -2164 13277
rect -2110 13231 -2097 13277
rect -2177 13198 -2097 13231
rect -1993 13277 -1913 13290
rect -1993 13231 -1980 13277
rect -1926 13231 -1913 13277
rect -1993 13198 -1913 13231
rect -2361 12665 -2281 12698
rect -2361 12619 -2348 12665
rect -2294 12619 -2281 12665
rect -2361 12606 -2281 12619
rect -2177 12665 -2097 12698
rect -2177 12619 -2164 12665
rect -2110 12619 -2097 12665
rect -2177 12606 -2097 12619
rect -1993 12665 -1913 12698
rect -1993 12619 -1980 12665
rect -1926 12619 -1913 12665
rect -1993 12606 -1913 12619
rect 195 13277 275 13290
rect 195 13231 208 13277
rect 262 13231 275 13277
rect 195 13198 275 13231
rect 379 13277 459 13290
rect 379 13231 392 13277
rect 446 13231 459 13277
rect 379 13198 459 13231
rect 563 13277 643 13290
rect 563 13231 576 13277
rect 630 13231 643 13277
rect 563 13198 643 13231
rect 195 12665 275 12698
rect 195 12619 208 12665
rect 262 12619 275 12665
rect 195 12606 275 12619
rect 379 12665 459 12698
rect 379 12619 392 12665
rect 446 12619 459 12665
rect 379 12606 459 12619
rect 563 12665 643 12698
rect 563 12619 576 12665
rect 630 12619 643 12665
rect 563 12606 643 12619
rect 1681 13277 1761 13290
rect 1681 13231 1694 13277
rect 1748 13231 1761 13277
rect 1681 13198 1761 13231
rect 1865 13277 1945 13290
rect 1865 13231 1878 13277
rect 1932 13231 1945 13277
rect 1865 13198 1945 13231
rect 2049 13277 2129 13290
rect 2049 13231 2062 13277
rect 2116 13231 2129 13277
rect 2049 13198 2129 13231
rect 1681 12665 1761 12698
rect 1681 12619 1694 12665
rect 1748 12619 1761 12665
rect 1681 12606 1761 12619
rect 1865 12665 1945 12698
rect 1865 12619 1878 12665
rect 1932 12619 1945 12665
rect 1865 12606 1945 12619
rect 2049 12665 2129 12698
rect 2049 12619 2062 12665
rect 2116 12619 2129 12665
rect 2049 12606 2129 12619
rect 4237 13277 4317 13290
rect 4237 13231 4250 13277
rect 4304 13231 4317 13277
rect 4237 13198 4317 13231
rect 4421 13277 4501 13290
rect 4421 13231 4434 13277
rect 4488 13231 4501 13277
rect 4421 13198 4501 13231
rect 4605 13277 4685 13290
rect 4605 13231 4618 13277
rect 4672 13231 4685 13277
rect 4605 13198 4685 13231
rect 4237 12665 4317 12698
rect 4237 12619 4250 12665
rect 4304 12619 4317 12665
rect 4237 12606 4317 12619
rect 4421 12665 4501 12698
rect 4421 12619 4434 12665
rect 4488 12619 4501 12665
rect 4421 12606 4501 12619
rect 4605 12665 4685 12698
rect 4605 12619 4618 12665
rect 4672 12619 4685 12665
rect 4605 12606 4685 12619
rect 5723 13277 5803 13290
rect 5723 13231 5736 13277
rect 5790 13231 5803 13277
rect 5723 13198 5803 13231
rect 5907 13277 5987 13290
rect 5907 13231 5920 13277
rect 5974 13231 5987 13277
rect 5907 13198 5987 13231
rect 6091 13277 6171 13290
rect 6091 13231 6104 13277
rect 6158 13231 6171 13277
rect 6091 13198 6171 13231
rect 5723 12665 5803 12698
rect 5723 12619 5736 12665
rect 5790 12619 5803 12665
rect 5723 12606 5803 12619
rect 5907 12665 5987 12698
rect 5907 12619 5920 12665
rect 5974 12619 5987 12665
rect 5907 12606 5987 12619
rect 6091 12665 6171 12698
rect 6091 12619 6104 12665
rect 6158 12619 6171 12665
rect 6091 12606 6171 12619
rect 8279 13277 8359 13290
rect 8279 13231 8292 13277
rect 8346 13231 8359 13277
rect 8279 13198 8359 13231
rect 8463 13277 8543 13290
rect 8463 13231 8476 13277
rect 8530 13231 8543 13277
rect 8463 13198 8543 13231
rect 8647 13277 8727 13290
rect 8647 13231 8660 13277
rect 8714 13231 8727 13277
rect 8647 13198 8727 13231
rect 8279 12665 8359 12698
rect 8279 12619 8292 12665
rect 8346 12619 8359 12665
rect 8279 12606 8359 12619
rect 8463 12665 8543 12698
rect 8463 12619 8476 12665
rect 8530 12619 8543 12665
rect 8463 12606 8543 12619
rect 8647 12665 8727 12698
rect 8647 12619 8660 12665
rect 8714 12619 8727 12665
rect 8647 12606 8727 12619
rect 9765 13277 9845 13290
rect 9765 13231 9778 13277
rect 9832 13231 9845 13277
rect 9765 13198 9845 13231
rect 9949 13277 10029 13290
rect 9949 13231 9962 13277
rect 10016 13231 10029 13277
rect 9949 13198 10029 13231
rect 10133 13277 10213 13290
rect 10133 13231 10146 13277
rect 10200 13231 10213 13277
rect 10133 13198 10213 13231
rect 9765 12665 9845 12698
rect 9765 12619 9778 12665
rect 9832 12619 9845 12665
rect 9765 12606 9845 12619
rect 9949 12665 10029 12698
rect 9949 12619 9962 12665
rect 10016 12619 10029 12665
rect 9949 12606 10029 12619
rect 10133 12665 10213 12698
rect 10133 12619 10146 12665
rect 10200 12619 10213 12665
rect 10133 12606 10213 12619
rect 12321 13277 12401 13290
rect 12321 13231 12334 13277
rect 12388 13231 12401 13277
rect 12321 13198 12401 13231
rect 12505 13277 12585 13290
rect 12505 13231 12518 13277
rect 12572 13231 12585 13277
rect 12505 13198 12585 13231
rect 12689 13277 12769 13290
rect 12689 13231 12702 13277
rect 12756 13231 12769 13277
rect 12689 13198 12769 13231
rect 12321 12665 12401 12698
rect 12321 12619 12334 12665
rect 12388 12619 12401 12665
rect 12321 12606 12401 12619
rect 12505 12665 12585 12698
rect 12505 12619 12518 12665
rect 12572 12619 12585 12665
rect 12505 12606 12585 12619
rect 12689 12665 12769 12698
rect 12689 12619 12702 12665
rect 12756 12619 12769 12665
rect 12689 12606 12769 12619
rect 13807 13277 13887 13290
rect 13807 13231 13820 13277
rect 13874 13231 13887 13277
rect 13807 13198 13887 13231
rect 13991 13277 14071 13290
rect 13991 13231 14004 13277
rect 14058 13231 14071 13277
rect 13991 13198 14071 13231
rect 14175 13277 14255 13290
rect 14175 13231 14188 13277
rect 14242 13231 14255 13277
rect 14175 13198 14255 13231
rect 13807 12665 13887 12698
rect 13807 12619 13820 12665
rect 13874 12619 13887 12665
rect 13807 12606 13887 12619
rect 13991 12665 14071 12698
rect 13991 12619 14004 12665
rect 14058 12619 14071 12665
rect 13991 12606 14071 12619
rect 14175 12665 14255 12698
rect 14175 12619 14188 12665
rect 14242 12619 14255 12665
rect 14175 12606 14255 12619
rect -11901 12117 -11821 12130
rect -11901 12071 -11888 12117
rect -11834 12071 -11821 12117
rect -11901 12038 -11821 12071
rect -11717 12117 -11637 12130
rect -11717 12071 -11704 12117
rect -11650 12071 -11637 12117
rect -11717 12038 -11637 12071
rect -11533 12117 -11453 12130
rect -11533 12071 -11520 12117
rect -11466 12071 -11453 12117
rect -11533 12038 -11453 12071
rect -11901 11805 -11821 11838
rect -11901 11759 -11888 11805
rect -11834 11759 -11821 11805
rect -11901 11746 -11821 11759
rect -11717 11805 -11637 11838
rect -11717 11759 -11704 11805
rect -11650 11759 -11637 11805
rect -11717 11746 -11637 11759
rect -11533 11805 -11453 11838
rect -11533 11759 -11520 11805
rect -11466 11759 -11453 11805
rect -11533 11746 -11453 11759
rect -10415 12117 -10335 12130
rect -10415 12071 -10402 12117
rect -10348 12071 -10335 12117
rect -10415 12038 -10335 12071
rect -10231 12117 -10151 12130
rect -10231 12071 -10218 12117
rect -10164 12071 -10151 12117
rect -10231 12038 -10151 12071
rect -10047 12117 -9967 12130
rect -10047 12071 -10034 12117
rect -9980 12071 -9967 12117
rect -10047 12038 -9967 12071
rect -10415 11805 -10335 11838
rect -10415 11759 -10402 11805
rect -10348 11759 -10335 11805
rect -10415 11746 -10335 11759
rect -10231 11805 -10151 11838
rect -10231 11759 -10218 11805
rect -10164 11759 -10151 11805
rect -10231 11746 -10151 11759
rect -10047 11805 -9967 11838
rect -10047 11759 -10034 11805
rect -9980 11759 -9967 11805
rect -10047 11746 -9967 11759
rect -7889 12117 -7809 12130
rect -7889 12071 -7876 12117
rect -7822 12071 -7809 12117
rect -7889 12038 -7809 12071
rect -7705 12117 -7625 12130
rect -7705 12071 -7692 12117
rect -7638 12071 -7625 12117
rect -7705 12038 -7625 12071
rect -7521 12117 -7441 12130
rect -7521 12071 -7508 12117
rect -7454 12071 -7441 12117
rect -7521 12038 -7441 12071
rect -7889 11805 -7809 11838
rect -7889 11759 -7876 11805
rect -7822 11759 -7809 11805
rect -7889 11746 -7809 11759
rect -7705 11805 -7625 11838
rect -7705 11759 -7692 11805
rect -7638 11759 -7625 11805
rect -7705 11746 -7625 11759
rect -7521 11805 -7441 11838
rect -7521 11759 -7508 11805
rect -7454 11759 -7441 11805
rect -7521 11746 -7441 11759
rect -6403 12117 -6323 12130
rect -6403 12071 -6390 12117
rect -6336 12071 -6323 12117
rect -6403 12038 -6323 12071
rect -6219 12117 -6139 12130
rect -6219 12071 -6206 12117
rect -6152 12071 -6139 12117
rect -6219 12038 -6139 12071
rect -6035 12117 -5955 12130
rect -6035 12071 -6022 12117
rect -5968 12071 -5955 12117
rect -6035 12038 -5955 12071
rect -6403 11805 -6323 11838
rect -6403 11759 -6390 11805
rect -6336 11759 -6323 11805
rect -6403 11746 -6323 11759
rect -6219 11805 -6139 11838
rect -6219 11759 -6206 11805
rect -6152 11759 -6139 11805
rect -6219 11746 -6139 11759
rect -6035 11805 -5955 11838
rect -6035 11759 -6022 11805
rect -5968 11759 -5955 11805
rect -6035 11746 -5955 11759
rect -3847 12117 -3767 12130
rect -3847 12071 -3834 12117
rect -3780 12071 -3767 12117
rect -3847 12038 -3767 12071
rect -3663 12117 -3583 12130
rect -3663 12071 -3650 12117
rect -3596 12071 -3583 12117
rect -3663 12038 -3583 12071
rect -3479 12117 -3399 12130
rect -3479 12071 -3466 12117
rect -3412 12071 -3399 12117
rect -3479 12038 -3399 12071
rect -3847 11805 -3767 11838
rect -3847 11759 -3834 11805
rect -3780 11759 -3767 11805
rect -3847 11746 -3767 11759
rect -3663 11805 -3583 11838
rect -3663 11759 -3650 11805
rect -3596 11759 -3583 11805
rect -3663 11746 -3583 11759
rect -3479 11805 -3399 11838
rect -3479 11759 -3466 11805
rect -3412 11759 -3399 11805
rect -3479 11746 -3399 11759
rect -2361 12117 -2281 12130
rect -2361 12071 -2348 12117
rect -2294 12071 -2281 12117
rect -2361 12038 -2281 12071
rect -2177 12117 -2097 12130
rect -2177 12071 -2164 12117
rect -2110 12071 -2097 12117
rect -2177 12038 -2097 12071
rect -1993 12117 -1913 12130
rect -1993 12071 -1980 12117
rect -1926 12071 -1913 12117
rect -1993 12038 -1913 12071
rect -2361 11805 -2281 11838
rect -2361 11759 -2348 11805
rect -2294 11759 -2281 11805
rect -2361 11746 -2281 11759
rect -2177 11805 -2097 11838
rect -2177 11759 -2164 11805
rect -2110 11759 -2097 11805
rect -2177 11746 -2097 11759
rect -1993 11805 -1913 11838
rect -1993 11759 -1980 11805
rect -1926 11759 -1913 11805
rect -1993 11746 -1913 11759
rect 195 12117 275 12130
rect 195 12071 208 12117
rect 262 12071 275 12117
rect 195 12038 275 12071
rect 379 12117 459 12130
rect 379 12071 392 12117
rect 446 12071 459 12117
rect 379 12038 459 12071
rect 563 12117 643 12130
rect 563 12071 576 12117
rect 630 12071 643 12117
rect 563 12038 643 12071
rect 195 11805 275 11838
rect 195 11759 208 11805
rect 262 11759 275 11805
rect 195 11746 275 11759
rect 379 11805 459 11838
rect 379 11759 392 11805
rect 446 11759 459 11805
rect 379 11746 459 11759
rect 563 11805 643 11838
rect 563 11759 576 11805
rect 630 11759 643 11805
rect 563 11746 643 11759
rect 1681 12117 1761 12130
rect 1681 12071 1694 12117
rect 1748 12071 1761 12117
rect 1681 12038 1761 12071
rect 1865 12117 1945 12130
rect 1865 12071 1878 12117
rect 1932 12071 1945 12117
rect 1865 12038 1945 12071
rect 2049 12117 2129 12130
rect 2049 12071 2062 12117
rect 2116 12071 2129 12117
rect 2049 12038 2129 12071
rect 1681 11805 1761 11838
rect 1681 11759 1694 11805
rect 1748 11759 1761 11805
rect 1681 11746 1761 11759
rect 1865 11805 1945 11838
rect 1865 11759 1878 11805
rect 1932 11759 1945 11805
rect 1865 11746 1945 11759
rect 2049 11805 2129 11838
rect 2049 11759 2062 11805
rect 2116 11759 2129 11805
rect 2049 11746 2129 11759
rect 4237 12117 4317 12130
rect 4237 12071 4250 12117
rect 4304 12071 4317 12117
rect 4237 12038 4317 12071
rect 4421 12117 4501 12130
rect 4421 12071 4434 12117
rect 4488 12071 4501 12117
rect 4421 12038 4501 12071
rect 4605 12117 4685 12130
rect 4605 12071 4618 12117
rect 4672 12071 4685 12117
rect 4605 12038 4685 12071
rect 4237 11805 4317 11838
rect 4237 11759 4250 11805
rect 4304 11759 4317 11805
rect 4237 11746 4317 11759
rect 4421 11805 4501 11838
rect 4421 11759 4434 11805
rect 4488 11759 4501 11805
rect 4421 11746 4501 11759
rect 4605 11805 4685 11838
rect 4605 11759 4618 11805
rect 4672 11759 4685 11805
rect 4605 11746 4685 11759
rect 5723 12117 5803 12130
rect 5723 12071 5736 12117
rect 5790 12071 5803 12117
rect 5723 12038 5803 12071
rect 5907 12117 5987 12130
rect 5907 12071 5920 12117
rect 5974 12071 5987 12117
rect 5907 12038 5987 12071
rect 6091 12117 6171 12130
rect 6091 12071 6104 12117
rect 6158 12071 6171 12117
rect 6091 12038 6171 12071
rect 5723 11805 5803 11838
rect 5723 11759 5736 11805
rect 5790 11759 5803 11805
rect 5723 11746 5803 11759
rect 5907 11805 5987 11838
rect 5907 11759 5920 11805
rect 5974 11759 5987 11805
rect 5907 11746 5987 11759
rect 6091 11805 6171 11838
rect 6091 11759 6104 11805
rect 6158 11759 6171 11805
rect 6091 11746 6171 11759
rect 8279 12117 8359 12130
rect 8279 12071 8292 12117
rect 8346 12071 8359 12117
rect 8279 12038 8359 12071
rect 8463 12117 8543 12130
rect 8463 12071 8476 12117
rect 8530 12071 8543 12117
rect 8463 12038 8543 12071
rect 8647 12117 8727 12130
rect 8647 12071 8660 12117
rect 8714 12071 8727 12117
rect 8647 12038 8727 12071
rect 8279 11805 8359 11838
rect 8279 11759 8292 11805
rect 8346 11759 8359 11805
rect 8279 11746 8359 11759
rect 8463 11805 8543 11838
rect 8463 11759 8476 11805
rect 8530 11759 8543 11805
rect 8463 11746 8543 11759
rect 8647 11805 8727 11838
rect 8647 11759 8660 11805
rect 8714 11759 8727 11805
rect 8647 11746 8727 11759
rect 9765 12117 9845 12130
rect 9765 12071 9778 12117
rect 9832 12071 9845 12117
rect 9765 12038 9845 12071
rect 9949 12117 10029 12130
rect 9949 12071 9962 12117
rect 10016 12071 10029 12117
rect 9949 12038 10029 12071
rect 10133 12117 10213 12130
rect 10133 12071 10146 12117
rect 10200 12071 10213 12117
rect 10133 12038 10213 12071
rect 9765 11805 9845 11838
rect 9765 11759 9778 11805
rect 9832 11759 9845 11805
rect 9765 11746 9845 11759
rect 9949 11805 10029 11838
rect 9949 11759 9962 11805
rect 10016 11759 10029 11805
rect 9949 11746 10029 11759
rect 10133 11805 10213 11838
rect 10133 11759 10146 11805
rect 10200 11759 10213 11805
rect 10133 11746 10213 11759
rect 12321 12117 12401 12130
rect 12321 12071 12334 12117
rect 12388 12071 12401 12117
rect 12321 12038 12401 12071
rect 12505 12117 12585 12130
rect 12505 12071 12518 12117
rect 12572 12071 12585 12117
rect 12505 12038 12585 12071
rect 12689 12117 12769 12130
rect 12689 12071 12702 12117
rect 12756 12071 12769 12117
rect 12689 12038 12769 12071
rect 12321 11805 12401 11838
rect 12321 11759 12334 11805
rect 12388 11759 12401 11805
rect 12321 11746 12401 11759
rect 12505 11805 12585 11838
rect 12505 11759 12518 11805
rect 12572 11759 12585 11805
rect 12505 11746 12585 11759
rect 12689 11805 12769 11838
rect 12689 11759 12702 11805
rect 12756 11759 12769 11805
rect 12689 11746 12769 11759
rect 13807 12117 13887 12130
rect 13807 12071 13820 12117
rect 13874 12071 13887 12117
rect 13807 12038 13887 12071
rect 13991 12117 14071 12130
rect 13991 12071 14004 12117
rect 14058 12071 14071 12117
rect 13991 12038 14071 12071
rect 14175 12117 14255 12130
rect 14175 12071 14188 12117
rect 14242 12071 14255 12117
rect 14175 12038 14255 12071
rect 13807 11805 13887 11838
rect 13807 11759 13820 11805
rect 13874 11759 13887 11805
rect 13807 11746 13887 11759
rect 13991 11805 14071 11838
rect 13991 11759 14004 11805
rect 14058 11759 14071 11805
rect 13991 11746 14071 11759
rect 14175 11805 14255 11838
rect 14175 11759 14188 11805
rect 14242 11759 14255 11805
rect 14175 11746 14255 11759
rect -11901 11072 -11821 11085
rect -11901 11026 -11888 11072
rect -11834 11026 -11821 11072
rect -11901 10993 -11821 11026
rect -11717 11072 -11637 11085
rect -11717 11026 -11704 11072
rect -11650 11026 -11637 11072
rect -11717 10993 -11637 11026
rect -11533 11072 -11453 11085
rect -11533 11026 -11520 11072
rect -11466 11026 -11453 11072
rect -11533 10993 -11453 11026
rect -11901 10460 -11821 10493
rect -11901 10414 -11888 10460
rect -11834 10414 -11821 10460
rect -11901 10401 -11821 10414
rect -11717 10460 -11637 10493
rect -11717 10414 -11704 10460
rect -11650 10414 -11637 10460
rect -11717 10401 -11637 10414
rect -11533 10460 -11453 10493
rect -11533 10414 -11520 10460
rect -11466 10414 -11453 10460
rect -11533 10401 -11453 10414
rect -10415 11073 -10335 11086
rect -10415 11027 -10402 11073
rect -10348 11027 -10335 11073
rect -10415 10994 -10335 11027
rect -10231 11073 -10151 11086
rect -10231 11027 -10218 11073
rect -10164 11027 -10151 11073
rect -10231 10994 -10151 11027
rect -10047 11073 -9967 11086
rect -10047 11027 -10034 11073
rect -9980 11027 -9967 11073
rect -10047 10994 -9967 11027
rect -10415 10461 -10335 10494
rect -10415 10415 -10402 10461
rect -10348 10415 -10335 10461
rect -10415 10402 -10335 10415
rect -10231 10461 -10151 10494
rect -10231 10415 -10218 10461
rect -10164 10415 -10151 10461
rect -10231 10402 -10151 10415
rect -10047 10461 -9967 10494
rect -10047 10415 -10034 10461
rect -9980 10415 -9967 10461
rect -10047 10402 -9967 10415
rect -7889 11072 -7809 11085
rect -7889 11026 -7876 11072
rect -7822 11026 -7809 11072
rect -7889 10993 -7809 11026
rect -7705 11072 -7625 11085
rect -7705 11026 -7692 11072
rect -7638 11026 -7625 11072
rect -7705 10993 -7625 11026
rect -7521 11072 -7441 11085
rect -7521 11026 -7508 11072
rect -7454 11026 -7441 11072
rect -7521 10993 -7441 11026
rect -7889 10460 -7809 10493
rect -7889 10414 -7876 10460
rect -7822 10414 -7809 10460
rect -7889 10401 -7809 10414
rect -7705 10460 -7625 10493
rect -7705 10414 -7692 10460
rect -7638 10414 -7625 10460
rect -7705 10401 -7625 10414
rect -7521 10460 -7441 10493
rect -7521 10414 -7508 10460
rect -7454 10414 -7441 10460
rect -7521 10401 -7441 10414
rect -6403 11073 -6323 11086
rect -6403 11027 -6390 11073
rect -6336 11027 -6323 11073
rect -6403 10994 -6323 11027
rect -6219 11073 -6139 11086
rect -6219 11027 -6206 11073
rect -6152 11027 -6139 11073
rect -6219 10994 -6139 11027
rect -6035 11073 -5955 11086
rect -6035 11027 -6022 11073
rect -5968 11027 -5955 11073
rect -6035 10994 -5955 11027
rect -6403 10461 -6323 10494
rect -6403 10415 -6390 10461
rect -6336 10415 -6323 10461
rect -6403 10402 -6323 10415
rect -6219 10461 -6139 10494
rect -6219 10415 -6206 10461
rect -6152 10415 -6139 10461
rect -6219 10402 -6139 10415
rect -6035 10461 -5955 10494
rect -6035 10415 -6022 10461
rect -5968 10415 -5955 10461
rect -6035 10402 -5955 10415
rect -3847 11072 -3767 11085
rect -3847 11026 -3834 11072
rect -3780 11026 -3767 11072
rect -3847 10993 -3767 11026
rect -3663 11072 -3583 11085
rect -3663 11026 -3650 11072
rect -3596 11026 -3583 11072
rect -3663 10993 -3583 11026
rect -3479 11072 -3399 11085
rect -3479 11026 -3466 11072
rect -3412 11026 -3399 11072
rect -3479 10993 -3399 11026
rect -3847 10460 -3767 10493
rect -3847 10414 -3834 10460
rect -3780 10414 -3767 10460
rect -3847 10401 -3767 10414
rect -3663 10460 -3583 10493
rect -3663 10414 -3650 10460
rect -3596 10414 -3583 10460
rect -3663 10401 -3583 10414
rect -3479 10460 -3399 10493
rect -3479 10414 -3466 10460
rect -3412 10414 -3399 10460
rect -3479 10401 -3399 10414
rect -2361 11073 -2281 11086
rect -2361 11027 -2348 11073
rect -2294 11027 -2281 11073
rect -2361 10994 -2281 11027
rect -2177 11073 -2097 11086
rect -2177 11027 -2164 11073
rect -2110 11027 -2097 11073
rect -2177 10994 -2097 11027
rect -1993 11073 -1913 11086
rect -1993 11027 -1980 11073
rect -1926 11027 -1913 11073
rect -1993 10994 -1913 11027
rect -2361 10461 -2281 10494
rect -2361 10415 -2348 10461
rect -2294 10415 -2281 10461
rect -2361 10402 -2281 10415
rect -2177 10461 -2097 10494
rect -2177 10415 -2164 10461
rect -2110 10415 -2097 10461
rect -2177 10402 -2097 10415
rect -1993 10461 -1913 10494
rect -1993 10415 -1980 10461
rect -1926 10415 -1913 10461
rect -1993 10402 -1913 10415
rect 195 11072 275 11085
rect 195 11026 208 11072
rect 262 11026 275 11072
rect 195 10993 275 11026
rect 379 11072 459 11085
rect 379 11026 392 11072
rect 446 11026 459 11072
rect 379 10993 459 11026
rect 563 11072 643 11085
rect 563 11026 576 11072
rect 630 11026 643 11072
rect 563 10993 643 11026
rect 195 10460 275 10493
rect 195 10414 208 10460
rect 262 10414 275 10460
rect 195 10401 275 10414
rect 379 10460 459 10493
rect 379 10414 392 10460
rect 446 10414 459 10460
rect 379 10401 459 10414
rect 563 10460 643 10493
rect 563 10414 576 10460
rect 630 10414 643 10460
rect 563 10401 643 10414
rect 1681 11073 1761 11086
rect 1681 11027 1694 11073
rect 1748 11027 1761 11073
rect 1681 10994 1761 11027
rect 1865 11073 1945 11086
rect 1865 11027 1878 11073
rect 1932 11027 1945 11073
rect 1865 10994 1945 11027
rect 2049 11073 2129 11086
rect 2049 11027 2062 11073
rect 2116 11027 2129 11073
rect 2049 10994 2129 11027
rect 1681 10461 1761 10494
rect 1681 10415 1694 10461
rect 1748 10415 1761 10461
rect 1681 10402 1761 10415
rect 1865 10461 1945 10494
rect 1865 10415 1878 10461
rect 1932 10415 1945 10461
rect 1865 10402 1945 10415
rect 2049 10461 2129 10494
rect 2049 10415 2062 10461
rect 2116 10415 2129 10461
rect 2049 10402 2129 10415
rect 4237 11072 4317 11085
rect 4237 11026 4250 11072
rect 4304 11026 4317 11072
rect 4237 10993 4317 11026
rect 4421 11072 4501 11085
rect 4421 11026 4434 11072
rect 4488 11026 4501 11072
rect 4421 10993 4501 11026
rect 4605 11072 4685 11085
rect 4605 11026 4618 11072
rect 4672 11026 4685 11072
rect 4605 10993 4685 11026
rect 4237 10460 4317 10493
rect 4237 10414 4250 10460
rect 4304 10414 4317 10460
rect 4237 10401 4317 10414
rect 4421 10460 4501 10493
rect 4421 10414 4434 10460
rect 4488 10414 4501 10460
rect 4421 10401 4501 10414
rect 4605 10460 4685 10493
rect 4605 10414 4618 10460
rect 4672 10414 4685 10460
rect 4605 10401 4685 10414
rect 5723 11073 5803 11086
rect 5723 11027 5736 11073
rect 5790 11027 5803 11073
rect 5723 10994 5803 11027
rect 5907 11073 5987 11086
rect 5907 11027 5920 11073
rect 5974 11027 5987 11073
rect 5907 10994 5987 11027
rect 6091 11073 6171 11086
rect 6091 11027 6104 11073
rect 6158 11027 6171 11073
rect 6091 10994 6171 11027
rect 5723 10461 5803 10494
rect 5723 10415 5736 10461
rect 5790 10415 5803 10461
rect 5723 10402 5803 10415
rect 5907 10461 5987 10494
rect 5907 10415 5920 10461
rect 5974 10415 5987 10461
rect 5907 10402 5987 10415
rect 6091 10461 6171 10494
rect 6091 10415 6104 10461
rect 6158 10415 6171 10461
rect 6091 10402 6171 10415
rect 8279 11072 8359 11085
rect 8279 11026 8292 11072
rect 8346 11026 8359 11072
rect 8279 10993 8359 11026
rect 8463 11072 8543 11085
rect 8463 11026 8476 11072
rect 8530 11026 8543 11072
rect 8463 10993 8543 11026
rect 8647 11072 8727 11085
rect 8647 11026 8660 11072
rect 8714 11026 8727 11072
rect 8647 10993 8727 11026
rect 8279 10460 8359 10493
rect 8279 10414 8292 10460
rect 8346 10414 8359 10460
rect 8279 10401 8359 10414
rect 8463 10460 8543 10493
rect 8463 10414 8476 10460
rect 8530 10414 8543 10460
rect 8463 10401 8543 10414
rect 8647 10460 8727 10493
rect 8647 10414 8660 10460
rect 8714 10414 8727 10460
rect 8647 10401 8727 10414
rect 9765 11073 9845 11086
rect 9765 11027 9778 11073
rect 9832 11027 9845 11073
rect 9765 10994 9845 11027
rect 9949 11073 10029 11086
rect 9949 11027 9962 11073
rect 10016 11027 10029 11073
rect 9949 10994 10029 11027
rect 10133 11073 10213 11086
rect 10133 11027 10146 11073
rect 10200 11027 10213 11073
rect 10133 10994 10213 11027
rect 9765 10461 9845 10494
rect 9765 10415 9778 10461
rect 9832 10415 9845 10461
rect 9765 10402 9845 10415
rect 9949 10461 10029 10494
rect 9949 10415 9962 10461
rect 10016 10415 10029 10461
rect 9949 10402 10029 10415
rect 10133 10461 10213 10494
rect 10133 10415 10146 10461
rect 10200 10415 10213 10461
rect 10133 10402 10213 10415
rect 12321 11072 12401 11085
rect 12321 11026 12334 11072
rect 12388 11026 12401 11072
rect 12321 10993 12401 11026
rect 12505 11072 12585 11085
rect 12505 11026 12518 11072
rect 12572 11026 12585 11072
rect 12505 10993 12585 11026
rect 12689 11072 12769 11085
rect 12689 11026 12702 11072
rect 12756 11026 12769 11072
rect 12689 10993 12769 11026
rect 12321 10460 12401 10493
rect 12321 10414 12334 10460
rect 12388 10414 12401 10460
rect 12321 10401 12401 10414
rect 12505 10460 12585 10493
rect 12505 10414 12518 10460
rect 12572 10414 12585 10460
rect 12505 10401 12585 10414
rect 12689 10460 12769 10493
rect 12689 10414 12702 10460
rect 12756 10414 12769 10460
rect 12689 10401 12769 10414
rect 13807 11073 13887 11086
rect 13807 11027 13820 11073
rect 13874 11027 13887 11073
rect 13807 10994 13887 11027
rect 13991 11073 14071 11086
rect 13991 11027 14004 11073
rect 14058 11027 14071 11073
rect 13991 10994 14071 11027
rect 14175 11073 14255 11086
rect 14175 11027 14188 11073
rect 14242 11027 14255 11073
rect 14175 10994 14255 11027
rect 13807 10461 13887 10494
rect 13807 10415 13820 10461
rect 13874 10415 13887 10461
rect 13807 10402 13887 10415
rect 13991 10461 14071 10494
rect 13991 10415 14004 10461
rect 14058 10415 14071 10461
rect 13991 10402 14071 10415
rect 14175 10461 14255 10494
rect 14175 10415 14188 10461
rect 14242 10415 14255 10461
rect 14175 10402 14255 10415
rect -11901 9912 -11821 9925
rect -11901 9866 -11888 9912
rect -11834 9866 -11821 9912
rect -11901 9833 -11821 9866
rect -11717 9912 -11637 9925
rect -11717 9866 -11704 9912
rect -11650 9866 -11637 9912
rect -11717 9833 -11637 9866
rect -11533 9912 -11453 9925
rect -11533 9866 -11520 9912
rect -11466 9866 -11453 9912
rect -11533 9833 -11453 9866
rect -11901 9600 -11821 9633
rect -11901 9554 -11888 9600
rect -11834 9554 -11821 9600
rect -11901 9541 -11821 9554
rect -11717 9600 -11637 9633
rect -11717 9554 -11704 9600
rect -11650 9554 -11637 9600
rect -11717 9541 -11637 9554
rect -11533 9600 -11453 9633
rect -11533 9554 -11520 9600
rect -11466 9554 -11453 9600
rect -11533 9541 -11453 9554
rect -10415 9913 -10335 9926
rect -10415 9867 -10402 9913
rect -10348 9867 -10335 9913
rect -10415 9834 -10335 9867
rect -10231 9913 -10151 9926
rect -10231 9867 -10218 9913
rect -10164 9867 -10151 9913
rect -10231 9834 -10151 9867
rect -10047 9913 -9967 9926
rect -10047 9867 -10034 9913
rect -9980 9867 -9967 9913
rect -10047 9834 -9967 9867
rect -10415 9601 -10335 9634
rect -10415 9555 -10402 9601
rect -10348 9555 -10335 9601
rect -10415 9542 -10335 9555
rect -10231 9601 -10151 9634
rect -10231 9555 -10218 9601
rect -10164 9555 -10151 9601
rect -10231 9542 -10151 9555
rect -10047 9601 -9967 9634
rect -10047 9555 -10034 9601
rect -9980 9555 -9967 9601
rect -10047 9542 -9967 9555
rect -7889 9912 -7809 9925
rect -7889 9866 -7876 9912
rect -7822 9866 -7809 9912
rect -7889 9833 -7809 9866
rect -7705 9912 -7625 9925
rect -7705 9866 -7692 9912
rect -7638 9866 -7625 9912
rect -7705 9833 -7625 9866
rect -7521 9912 -7441 9925
rect -7521 9866 -7508 9912
rect -7454 9866 -7441 9912
rect -7521 9833 -7441 9866
rect -7889 9600 -7809 9633
rect -7889 9554 -7876 9600
rect -7822 9554 -7809 9600
rect -7889 9541 -7809 9554
rect -7705 9600 -7625 9633
rect -7705 9554 -7692 9600
rect -7638 9554 -7625 9600
rect -7705 9541 -7625 9554
rect -7521 9600 -7441 9633
rect -7521 9554 -7508 9600
rect -7454 9554 -7441 9600
rect -7521 9541 -7441 9554
rect -6403 9913 -6323 9926
rect -6403 9867 -6390 9913
rect -6336 9867 -6323 9913
rect -6403 9834 -6323 9867
rect -6219 9913 -6139 9926
rect -6219 9867 -6206 9913
rect -6152 9867 -6139 9913
rect -6219 9834 -6139 9867
rect -6035 9913 -5955 9926
rect -6035 9867 -6022 9913
rect -5968 9867 -5955 9913
rect -6035 9834 -5955 9867
rect -6403 9601 -6323 9634
rect -6403 9555 -6390 9601
rect -6336 9555 -6323 9601
rect -6403 9542 -6323 9555
rect -6219 9601 -6139 9634
rect -6219 9555 -6206 9601
rect -6152 9555 -6139 9601
rect -6219 9542 -6139 9555
rect -6035 9601 -5955 9634
rect -6035 9555 -6022 9601
rect -5968 9555 -5955 9601
rect -6035 9542 -5955 9555
rect -3847 9912 -3767 9925
rect -3847 9866 -3834 9912
rect -3780 9866 -3767 9912
rect -3847 9833 -3767 9866
rect -3663 9912 -3583 9925
rect -3663 9866 -3650 9912
rect -3596 9866 -3583 9912
rect -3663 9833 -3583 9866
rect -3479 9912 -3399 9925
rect -3479 9866 -3466 9912
rect -3412 9866 -3399 9912
rect -3479 9833 -3399 9866
rect -3847 9600 -3767 9633
rect -3847 9554 -3834 9600
rect -3780 9554 -3767 9600
rect -3847 9541 -3767 9554
rect -3663 9600 -3583 9633
rect -3663 9554 -3650 9600
rect -3596 9554 -3583 9600
rect -3663 9541 -3583 9554
rect -3479 9600 -3399 9633
rect -3479 9554 -3466 9600
rect -3412 9554 -3399 9600
rect -3479 9541 -3399 9554
rect -2361 9913 -2281 9926
rect -2361 9867 -2348 9913
rect -2294 9867 -2281 9913
rect -2361 9834 -2281 9867
rect -2177 9913 -2097 9926
rect -2177 9867 -2164 9913
rect -2110 9867 -2097 9913
rect -2177 9834 -2097 9867
rect -1993 9913 -1913 9926
rect -1993 9867 -1980 9913
rect -1926 9867 -1913 9913
rect -1993 9834 -1913 9867
rect -2361 9601 -2281 9634
rect -2361 9555 -2348 9601
rect -2294 9555 -2281 9601
rect -2361 9542 -2281 9555
rect -2177 9601 -2097 9634
rect -2177 9555 -2164 9601
rect -2110 9555 -2097 9601
rect -2177 9542 -2097 9555
rect -1993 9601 -1913 9634
rect -1993 9555 -1980 9601
rect -1926 9555 -1913 9601
rect -1993 9542 -1913 9555
rect 195 9912 275 9925
rect 195 9866 208 9912
rect 262 9866 275 9912
rect 195 9833 275 9866
rect 379 9912 459 9925
rect 379 9866 392 9912
rect 446 9866 459 9912
rect 379 9833 459 9866
rect 563 9912 643 9925
rect 563 9866 576 9912
rect 630 9866 643 9912
rect 563 9833 643 9866
rect 195 9600 275 9633
rect 195 9554 208 9600
rect 262 9554 275 9600
rect 195 9541 275 9554
rect 379 9600 459 9633
rect 379 9554 392 9600
rect 446 9554 459 9600
rect 379 9541 459 9554
rect 563 9600 643 9633
rect 563 9554 576 9600
rect 630 9554 643 9600
rect 563 9541 643 9554
rect 1681 9913 1761 9926
rect 1681 9867 1694 9913
rect 1748 9867 1761 9913
rect 1681 9834 1761 9867
rect 1865 9913 1945 9926
rect 1865 9867 1878 9913
rect 1932 9867 1945 9913
rect 1865 9834 1945 9867
rect 2049 9913 2129 9926
rect 2049 9867 2062 9913
rect 2116 9867 2129 9913
rect 2049 9834 2129 9867
rect 1681 9601 1761 9634
rect 1681 9555 1694 9601
rect 1748 9555 1761 9601
rect 1681 9542 1761 9555
rect 1865 9601 1945 9634
rect 1865 9555 1878 9601
rect 1932 9555 1945 9601
rect 1865 9542 1945 9555
rect 2049 9601 2129 9634
rect 2049 9555 2062 9601
rect 2116 9555 2129 9601
rect 2049 9542 2129 9555
rect 4237 9912 4317 9925
rect 4237 9866 4250 9912
rect 4304 9866 4317 9912
rect 4237 9833 4317 9866
rect 4421 9912 4501 9925
rect 4421 9866 4434 9912
rect 4488 9866 4501 9912
rect 4421 9833 4501 9866
rect 4605 9912 4685 9925
rect 4605 9866 4618 9912
rect 4672 9866 4685 9912
rect 4605 9833 4685 9866
rect 4237 9600 4317 9633
rect 4237 9554 4250 9600
rect 4304 9554 4317 9600
rect 4237 9541 4317 9554
rect 4421 9600 4501 9633
rect 4421 9554 4434 9600
rect 4488 9554 4501 9600
rect 4421 9541 4501 9554
rect 4605 9600 4685 9633
rect 4605 9554 4618 9600
rect 4672 9554 4685 9600
rect 4605 9541 4685 9554
rect 5723 9913 5803 9926
rect 5723 9867 5736 9913
rect 5790 9867 5803 9913
rect 5723 9834 5803 9867
rect 5907 9913 5987 9926
rect 5907 9867 5920 9913
rect 5974 9867 5987 9913
rect 5907 9834 5987 9867
rect 6091 9913 6171 9926
rect 6091 9867 6104 9913
rect 6158 9867 6171 9913
rect 6091 9834 6171 9867
rect 5723 9601 5803 9634
rect 5723 9555 5736 9601
rect 5790 9555 5803 9601
rect 5723 9542 5803 9555
rect 5907 9601 5987 9634
rect 5907 9555 5920 9601
rect 5974 9555 5987 9601
rect 5907 9542 5987 9555
rect 6091 9601 6171 9634
rect 6091 9555 6104 9601
rect 6158 9555 6171 9601
rect 6091 9542 6171 9555
rect 8279 9912 8359 9925
rect 8279 9866 8292 9912
rect 8346 9866 8359 9912
rect 8279 9833 8359 9866
rect 8463 9912 8543 9925
rect 8463 9866 8476 9912
rect 8530 9866 8543 9912
rect 8463 9833 8543 9866
rect 8647 9912 8727 9925
rect 8647 9866 8660 9912
rect 8714 9866 8727 9912
rect 8647 9833 8727 9866
rect 8279 9600 8359 9633
rect 8279 9554 8292 9600
rect 8346 9554 8359 9600
rect 8279 9541 8359 9554
rect 8463 9600 8543 9633
rect 8463 9554 8476 9600
rect 8530 9554 8543 9600
rect 8463 9541 8543 9554
rect 8647 9600 8727 9633
rect 8647 9554 8660 9600
rect 8714 9554 8727 9600
rect 8647 9541 8727 9554
rect 9765 9913 9845 9926
rect 9765 9867 9778 9913
rect 9832 9867 9845 9913
rect 9765 9834 9845 9867
rect 9949 9913 10029 9926
rect 9949 9867 9962 9913
rect 10016 9867 10029 9913
rect 9949 9834 10029 9867
rect 10133 9913 10213 9926
rect 10133 9867 10146 9913
rect 10200 9867 10213 9913
rect 10133 9834 10213 9867
rect 9765 9601 9845 9634
rect 9765 9555 9778 9601
rect 9832 9555 9845 9601
rect 9765 9542 9845 9555
rect 9949 9601 10029 9634
rect 9949 9555 9962 9601
rect 10016 9555 10029 9601
rect 9949 9542 10029 9555
rect 10133 9601 10213 9634
rect 10133 9555 10146 9601
rect 10200 9555 10213 9601
rect 10133 9542 10213 9555
rect 12321 9912 12401 9925
rect 12321 9866 12334 9912
rect 12388 9866 12401 9912
rect 12321 9833 12401 9866
rect 12505 9912 12585 9925
rect 12505 9866 12518 9912
rect 12572 9866 12585 9912
rect 12505 9833 12585 9866
rect 12689 9912 12769 9925
rect 12689 9866 12702 9912
rect 12756 9866 12769 9912
rect 12689 9833 12769 9866
rect 12321 9600 12401 9633
rect 12321 9554 12334 9600
rect 12388 9554 12401 9600
rect 12321 9541 12401 9554
rect 12505 9600 12585 9633
rect 12505 9554 12518 9600
rect 12572 9554 12585 9600
rect 12505 9541 12585 9554
rect 12689 9600 12769 9633
rect 12689 9554 12702 9600
rect 12756 9554 12769 9600
rect 12689 9541 12769 9554
rect 13807 9913 13887 9926
rect 13807 9867 13820 9913
rect 13874 9867 13887 9913
rect 13807 9834 13887 9867
rect 13991 9913 14071 9926
rect 13991 9867 14004 9913
rect 14058 9867 14071 9913
rect 13991 9834 14071 9867
rect 14175 9913 14255 9926
rect 14175 9867 14188 9913
rect 14242 9867 14255 9913
rect 14175 9834 14255 9867
rect 13807 9601 13887 9634
rect 13807 9555 13820 9601
rect 13874 9555 13887 9601
rect 13807 9542 13887 9555
rect 13991 9601 14071 9634
rect 13991 9555 14004 9601
rect 14058 9555 14071 9601
rect 13991 9542 14071 9555
rect 14175 9601 14255 9634
rect 14175 9555 14188 9601
rect 14242 9555 14255 9601
rect 14175 9542 14255 9555
rect -11901 8867 -11821 8880
rect -11901 8821 -11888 8867
rect -11834 8821 -11821 8867
rect -11901 8788 -11821 8821
rect -11717 8867 -11637 8880
rect -11717 8821 -11704 8867
rect -11650 8821 -11637 8867
rect -11717 8788 -11637 8821
rect -11533 8867 -11453 8880
rect -11533 8821 -11520 8867
rect -11466 8821 -11453 8867
rect -11533 8788 -11453 8821
rect -11901 8255 -11821 8288
rect -11901 8209 -11888 8255
rect -11834 8209 -11821 8255
rect -11901 8196 -11821 8209
rect -11717 8255 -11637 8288
rect -11717 8209 -11704 8255
rect -11650 8209 -11637 8255
rect -11717 8196 -11637 8209
rect -11533 8255 -11453 8288
rect -11533 8209 -11520 8255
rect -11466 8209 -11453 8255
rect -11533 8196 -11453 8209
rect -7889 8867 -7809 8880
rect -7889 8821 -7876 8867
rect -7822 8821 -7809 8867
rect -7889 8788 -7809 8821
rect -7705 8867 -7625 8880
rect -7705 8821 -7692 8867
rect -7638 8821 -7625 8867
rect -7705 8788 -7625 8821
rect -7521 8867 -7441 8880
rect -7521 8821 -7508 8867
rect -7454 8821 -7441 8867
rect -7521 8788 -7441 8821
rect -7889 8255 -7809 8288
rect -7889 8209 -7876 8255
rect -7822 8209 -7809 8255
rect -7889 8196 -7809 8209
rect -7705 8255 -7625 8288
rect -7705 8209 -7692 8255
rect -7638 8209 -7625 8255
rect -7705 8196 -7625 8209
rect -7521 8255 -7441 8288
rect -7521 8209 -7508 8255
rect -7454 8209 -7441 8255
rect -7521 8196 -7441 8209
rect -3847 8867 -3767 8880
rect -3847 8821 -3834 8867
rect -3780 8821 -3767 8867
rect -3847 8788 -3767 8821
rect -3663 8867 -3583 8880
rect -3663 8821 -3650 8867
rect -3596 8821 -3583 8867
rect -3663 8788 -3583 8821
rect -3479 8867 -3399 8880
rect -3479 8821 -3466 8867
rect -3412 8821 -3399 8867
rect -3479 8788 -3399 8821
rect -3847 8255 -3767 8288
rect -3847 8209 -3834 8255
rect -3780 8209 -3767 8255
rect -3847 8196 -3767 8209
rect -3663 8255 -3583 8288
rect -3663 8209 -3650 8255
rect -3596 8209 -3583 8255
rect -3663 8196 -3583 8209
rect -3479 8255 -3399 8288
rect -3479 8209 -3466 8255
rect -3412 8209 -3399 8255
rect -3479 8196 -3399 8209
rect 195 8867 275 8880
rect 195 8821 208 8867
rect 262 8821 275 8867
rect 195 8788 275 8821
rect 379 8867 459 8880
rect 379 8821 392 8867
rect 446 8821 459 8867
rect 379 8788 459 8821
rect 563 8867 643 8880
rect 563 8821 576 8867
rect 630 8821 643 8867
rect 563 8788 643 8821
rect 195 8255 275 8288
rect 195 8209 208 8255
rect 262 8209 275 8255
rect 195 8196 275 8209
rect 379 8255 459 8288
rect 379 8209 392 8255
rect 446 8209 459 8255
rect 379 8196 459 8209
rect 563 8255 643 8288
rect 563 8209 576 8255
rect 630 8209 643 8255
rect 563 8196 643 8209
rect 4237 8867 4317 8880
rect 4237 8821 4250 8867
rect 4304 8821 4317 8867
rect 4237 8788 4317 8821
rect 4421 8867 4501 8880
rect 4421 8821 4434 8867
rect 4488 8821 4501 8867
rect 4421 8788 4501 8821
rect 4605 8867 4685 8880
rect 4605 8821 4618 8867
rect 4672 8821 4685 8867
rect 4605 8788 4685 8821
rect 4237 8255 4317 8288
rect 4237 8209 4250 8255
rect 4304 8209 4317 8255
rect 4237 8196 4317 8209
rect 4421 8255 4501 8288
rect 4421 8209 4434 8255
rect 4488 8209 4501 8255
rect 4421 8196 4501 8209
rect 4605 8255 4685 8288
rect 4605 8209 4618 8255
rect 4672 8209 4685 8255
rect 4605 8196 4685 8209
rect 8279 8867 8359 8880
rect 8279 8821 8292 8867
rect 8346 8821 8359 8867
rect 8279 8788 8359 8821
rect 8463 8867 8543 8880
rect 8463 8821 8476 8867
rect 8530 8821 8543 8867
rect 8463 8788 8543 8821
rect 8647 8867 8727 8880
rect 8647 8821 8660 8867
rect 8714 8821 8727 8867
rect 8647 8788 8727 8821
rect 8279 8255 8359 8288
rect 8279 8209 8292 8255
rect 8346 8209 8359 8255
rect 8279 8196 8359 8209
rect 8463 8255 8543 8288
rect 8463 8209 8476 8255
rect 8530 8209 8543 8255
rect 8463 8196 8543 8209
rect 8647 8255 8727 8288
rect 8647 8209 8660 8255
rect 8714 8209 8727 8255
rect 8647 8196 8727 8209
rect 12321 8867 12401 8880
rect 12321 8821 12334 8867
rect 12388 8821 12401 8867
rect 12321 8788 12401 8821
rect 12505 8867 12585 8880
rect 12505 8821 12518 8867
rect 12572 8821 12585 8867
rect 12505 8788 12585 8821
rect 12689 8867 12769 8880
rect 12689 8821 12702 8867
rect 12756 8821 12769 8867
rect 12689 8788 12769 8821
rect 12321 8255 12401 8288
rect 12321 8209 12334 8255
rect 12388 8209 12401 8255
rect 12321 8196 12401 8209
rect 12505 8255 12585 8288
rect 12505 8209 12518 8255
rect 12572 8209 12585 8255
rect 12505 8196 12585 8209
rect 12689 8255 12769 8288
rect 12689 8209 12702 8255
rect 12756 8209 12769 8255
rect 12689 8196 12769 8209
rect -11901 7707 -11821 7720
rect -11901 7661 -11888 7707
rect -11834 7661 -11821 7707
rect -11901 7628 -11821 7661
rect -11717 7707 -11637 7720
rect -11717 7661 -11704 7707
rect -11650 7661 -11637 7707
rect -11717 7628 -11637 7661
rect -11533 7707 -11453 7720
rect -11533 7661 -11520 7707
rect -11466 7661 -11453 7707
rect -11533 7628 -11453 7661
rect -11901 7395 -11821 7428
rect -11901 7349 -11888 7395
rect -11834 7349 -11821 7395
rect -11901 7336 -11821 7349
rect -11717 7395 -11637 7428
rect -11717 7349 -11704 7395
rect -11650 7349 -11637 7395
rect -11717 7336 -11637 7349
rect -11533 7395 -11453 7428
rect -11533 7349 -11520 7395
rect -11466 7349 -11453 7395
rect -11533 7336 -11453 7349
rect -7889 7707 -7809 7720
rect -7889 7661 -7876 7707
rect -7822 7661 -7809 7707
rect -7889 7628 -7809 7661
rect -7705 7707 -7625 7720
rect -7705 7661 -7692 7707
rect -7638 7661 -7625 7707
rect -7705 7628 -7625 7661
rect -7521 7707 -7441 7720
rect -7521 7661 -7508 7707
rect -7454 7661 -7441 7707
rect -7521 7628 -7441 7661
rect -7889 7395 -7809 7428
rect -7889 7349 -7876 7395
rect -7822 7349 -7809 7395
rect -7889 7336 -7809 7349
rect -7705 7395 -7625 7428
rect -7705 7349 -7692 7395
rect -7638 7349 -7625 7395
rect -7705 7336 -7625 7349
rect -7521 7395 -7441 7428
rect -7521 7349 -7508 7395
rect -7454 7349 -7441 7395
rect -7521 7336 -7441 7349
rect -3847 7707 -3767 7720
rect -3847 7661 -3834 7707
rect -3780 7661 -3767 7707
rect -3847 7628 -3767 7661
rect -3663 7707 -3583 7720
rect -3663 7661 -3650 7707
rect -3596 7661 -3583 7707
rect -3663 7628 -3583 7661
rect -3479 7707 -3399 7720
rect -3479 7661 -3466 7707
rect -3412 7661 -3399 7707
rect -3479 7628 -3399 7661
rect -3847 7395 -3767 7428
rect -3847 7349 -3834 7395
rect -3780 7349 -3767 7395
rect -3847 7336 -3767 7349
rect -3663 7395 -3583 7428
rect -3663 7349 -3650 7395
rect -3596 7349 -3583 7395
rect -3663 7336 -3583 7349
rect -3479 7395 -3399 7428
rect -3479 7349 -3466 7395
rect -3412 7349 -3399 7395
rect -3479 7336 -3399 7349
rect 195 7707 275 7720
rect 195 7661 208 7707
rect 262 7661 275 7707
rect 195 7628 275 7661
rect 379 7707 459 7720
rect 379 7661 392 7707
rect 446 7661 459 7707
rect 379 7628 459 7661
rect 563 7707 643 7720
rect 563 7661 576 7707
rect 630 7661 643 7707
rect 563 7628 643 7661
rect 195 7395 275 7428
rect 195 7349 208 7395
rect 262 7349 275 7395
rect 195 7336 275 7349
rect 379 7395 459 7428
rect 379 7349 392 7395
rect 446 7349 459 7395
rect 379 7336 459 7349
rect 563 7395 643 7428
rect 563 7349 576 7395
rect 630 7349 643 7395
rect 563 7336 643 7349
rect 4237 7707 4317 7720
rect 4237 7661 4250 7707
rect 4304 7661 4317 7707
rect 4237 7628 4317 7661
rect 4421 7707 4501 7720
rect 4421 7661 4434 7707
rect 4488 7661 4501 7707
rect 4421 7628 4501 7661
rect 4605 7707 4685 7720
rect 4605 7661 4618 7707
rect 4672 7661 4685 7707
rect 4605 7628 4685 7661
rect 4237 7395 4317 7428
rect 4237 7349 4250 7395
rect 4304 7349 4317 7395
rect 4237 7336 4317 7349
rect 4421 7395 4501 7428
rect 4421 7349 4434 7395
rect 4488 7349 4501 7395
rect 4421 7336 4501 7349
rect 4605 7395 4685 7428
rect 4605 7349 4618 7395
rect 4672 7349 4685 7395
rect 4605 7336 4685 7349
rect 8279 7707 8359 7720
rect 8279 7661 8292 7707
rect 8346 7661 8359 7707
rect 8279 7628 8359 7661
rect 8463 7707 8543 7720
rect 8463 7661 8476 7707
rect 8530 7661 8543 7707
rect 8463 7628 8543 7661
rect 8647 7707 8727 7720
rect 8647 7661 8660 7707
rect 8714 7661 8727 7707
rect 8647 7628 8727 7661
rect 8279 7395 8359 7428
rect 8279 7349 8292 7395
rect 8346 7349 8359 7395
rect 8279 7336 8359 7349
rect 8463 7395 8543 7428
rect 8463 7349 8476 7395
rect 8530 7349 8543 7395
rect 8463 7336 8543 7349
rect 8647 7395 8727 7428
rect 8647 7349 8660 7395
rect 8714 7349 8727 7395
rect 8647 7336 8727 7349
rect 12321 7707 12401 7720
rect 12321 7661 12334 7707
rect 12388 7661 12401 7707
rect 12321 7628 12401 7661
rect 12505 7707 12585 7720
rect 12505 7661 12518 7707
rect 12572 7661 12585 7707
rect 12505 7628 12585 7661
rect 12689 7707 12769 7720
rect 12689 7661 12702 7707
rect 12756 7661 12769 7707
rect 12689 7628 12769 7661
rect 12321 7395 12401 7428
rect 12321 7349 12334 7395
rect 12388 7349 12401 7395
rect 12321 7336 12401 7349
rect 12505 7395 12585 7428
rect 12505 7349 12518 7395
rect 12572 7349 12585 7395
rect 12505 7336 12585 7349
rect 12689 7395 12769 7428
rect 12689 7349 12702 7395
rect 12756 7349 12769 7395
rect 12689 7336 12769 7349
rect -10831 5220 -10771 5270
rect -10661 5220 -10601 5270
rect -10491 5220 -10431 5270
rect -10321 5220 -10261 5270
rect -10151 5220 -10091 5270
rect -10831 4860 -10771 4880
rect -10661 4860 -10601 4880
rect -10491 4860 -10431 4880
rect -10321 4860 -10261 4880
rect -10831 4850 -10261 4860
rect -10831 4823 -10201 4850
rect -10831 4800 -10274 4823
rect -10661 4620 -10601 4800
rect -10321 4777 -10274 4800
rect -10228 4777 -10201 4823
rect -10321 4750 -10201 4777
rect -10321 4620 -10261 4750
rect -10151 4700 -10091 4880
rect -10831 4560 -10261 4620
rect -10211 4673 -10091 4700
rect -10211 4627 -10184 4673
rect -10138 4627 -10091 4673
rect -10211 4600 -10091 4627
rect -10831 4540 -10771 4560
rect -10661 4540 -10601 4560
rect -10491 4540 -10431 4560
rect -10321 4540 -10261 4560
rect -10151 4540 -10091 4600
rect -8431 4946 -8351 4959
rect -8431 4900 -8418 4946
rect -8364 4900 -8351 4946
rect -8431 4867 -8351 4900
rect -8431 4634 -8351 4667
rect -8431 4588 -8418 4634
rect -8364 4588 -8351 4634
rect -8431 4575 -8351 4588
rect -7971 4946 -7891 4959
rect -7971 4900 -7958 4946
rect -7904 4900 -7891 4946
rect -7971 4867 -7891 4900
rect -7971 4634 -7891 4667
rect -7971 4588 -7958 4634
rect -7904 4588 -7891 4634
rect -7971 4575 -7891 4588
rect -10831 4320 -10771 4370
rect -10661 4320 -10601 4370
rect -10491 4320 -10431 4370
rect -10321 4320 -10261 4370
rect -10151 4320 -10091 4370
rect -9401 4362 -9321 4406
rect -9401 3529 -9321 3562
rect -9401 3483 -9388 3529
rect -9334 3483 -9321 3529
rect -9401 3470 -9321 3483
rect -8431 4126 -8351 4139
rect -8431 4080 -8418 4126
rect -8364 4080 -8351 4126
rect -8431 4047 -8351 4080
rect -8431 3814 -8351 3847
rect -8431 3768 -8418 3814
rect -8364 3768 -8351 3814
rect -8431 3755 -8351 3768
rect -7971 4126 -7891 4139
rect -7971 4080 -7958 4126
rect -7904 4080 -7891 4126
rect -7971 4047 -7891 4080
rect -7971 3814 -7891 3847
rect -7971 3768 -7958 3814
rect -7904 3768 -7891 3814
rect -7971 3755 -7891 3768
rect -7001 4362 -6921 4406
rect -7001 3529 -6921 3562
rect -7001 3483 -6988 3529
rect -6934 3483 -6921 3529
rect -7001 3470 -6921 3483
rect -9401 3193 -9321 3206
rect -9401 3147 -9388 3193
rect -9334 3147 -9321 3193
rect -9401 3114 -9321 3147
rect -9401 2670 -9321 2714
rect -7001 3193 -6921 3206
rect -7001 3147 -6988 3193
rect -6934 3147 -6921 3193
rect -7001 3114 -6921 3147
rect -7001 2670 -6921 2714
rect -10949 1756 -10869 1769
rect -10949 1710 -10936 1756
rect -10882 1710 -10869 1756
rect -10949 1677 -10869 1710
rect -10949 1484 -10869 1517
rect -10949 1438 -10936 1484
rect -10882 1438 -10869 1484
rect -10949 1425 -10869 1438
rect -10089 1756 -10009 1769
rect -10089 1710 -10076 1756
rect -10022 1710 -10009 1756
rect -10089 1677 -10009 1710
rect -10089 1484 -10009 1517
rect -10089 1438 -10076 1484
rect -10022 1438 -10009 1484
rect -10089 1425 -10009 1438
rect -9629 1776 -9429 1789
rect -9629 1730 -9616 1776
rect -9442 1730 -9429 1776
rect -9629 1697 -9429 1730
rect -9325 1776 -9125 1789
rect -9325 1730 -9312 1776
rect -9138 1730 -9125 1776
rect -9325 1697 -9125 1730
rect -9021 1776 -8821 1789
rect -9021 1730 -9008 1776
rect -8834 1730 -8821 1776
rect -9021 1697 -8821 1730
rect -8717 1776 -8517 1789
rect -8717 1730 -8704 1776
rect -8530 1730 -8517 1776
rect -8717 1697 -8517 1730
rect -8413 1776 -8213 1789
rect -8413 1730 -8400 1776
rect -8226 1730 -8213 1776
rect -8413 1697 -8213 1730
rect -8109 1776 -7909 1789
rect -8109 1730 -8096 1776
rect -7922 1730 -7909 1776
rect -8109 1697 -7909 1730
rect -7805 1776 -7605 1789
rect -7805 1730 -7792 1776
rect -7618 1730 -7605 1776
rect -7805 1697 -7605 1730
rect -7501 1776 -7301 1789
rect -7501 1730 -7488 1776
rect -7314 1730 -7301 1776
rect -7501 1697 -7301 1730
rect -7197 1776 -6997 1789
rect -7197 1730 -7184 1776
rect -7010 1730 -6997 1776
rect -7197 1697 -6997 1730
rect -6893 1776 -6693 1789
rect -6893 1730 -6880 1776
rect -6706 1730 -6693 1776
rect -6893 1697 -6693 1730
rect -9629 1464 -9429 1497
rect -9629 1418 -9616 1464
rect -9442 1418 -9429 1464
rect -9629 1405 -9429 1418
rect -9325 1464 -9125 1497
rect -9325 1418 -9312 1464
rect -9138 1418 -9125 1464
rect -9325 1405 -9125 1418
rect -9021 1464 -8821 1497
rect -9021 1418 -9008 1464
rect -8834 1418 -8821 1464
rect -9021 1405 -8821 1418
rect -8717 1464 -8517 1497
rect -8717 1418 -8704 1464
rect -8530 1418 -8517 1464
rect -8717 1405 -8517 1418
rect -8413 1464 -8213 1497
rect -8413 1418 -8400 1464
rect -8226 1418 -8213 1464
rect -8413 1405 -8213 1418
rect -8109 1464 -7909 1497
rect -8109 1418 -8096 1464
rect -7922 1418 -7909 1464
rect -8109 1405 -7909 1418
rect -7805 1464 -7605 1497
rect -7805 1418 -7792 1464
rect -7618 1418 -7605 1464
rect -7805 1405 -7605 1418
rect -7501 1464 -7301 1497
rect -7501 1418 -7488 1464
rect -7314 1418 -7301 1464
rect -7501 1405 -7301 1418
rect -7197 1464 -6997 1497
rect -7197 1418 -7184 1464
rect -7010 1418 -6997 1464
rect -7197 1405 -6997 1418
rect -6893 1464 -6693 1497
rect -6893 1418 -6880 1464
rect -6706 1418 -6693 1464
rect -6893 1405 -6693 1418
rect -6313 1756 -6233 1769
rect -6313 1710 -6300 1756
rect -6246 1710 -6233 1756
rect -6313 1677 -6233 1710
rect -6313 1484 -6233 1517
rect -6313 1438 -6300 1484
rect -6246 1438 -6233 1484
rect -6313 1425 -6233 1438
rect -5453 1756 -5373 1769
rect -5453 1710 -5440 1756
rect -5386 1710 -5373 1756
rect -5453 1677 -5373 1710
rect -5453 1484 -5373 1517
rect -5453 1438 -5440 1484
rect -5386 1438 -5373 1484
rect -5453 1425 -5373 1438
rect -9767 820 -9567 833
rect -9767 774 -9754 820
rect -9580 774 -9567 820
rect -9767 741 -9567 774
rect -9463 820 -9263 833
rect -9463 774 -9450 820
rect -9276 774 -9263 820
rect -9463 741 -9263 774
rect -9159 820 -8959 833
rect -9159 774 -9146 820
rect -8972 774 -8959 820
rect -9159 741 -8959 774
rect -8855 820 -8655 833
rect -8855 774 -8842 820
rect -8668 774 -8655 820
rect -8855 741 -8655 774
rect -8551 820 -8351 833
rect -8551 774 -8538 820
rect -8364 774 -8351 820
rect -8551 741 -8351 774
rect -9767 308 -9567 341
rect -9767 262 -9754 308
rect -9580 262 -9567 308
rect -9767 249 -9567 262
rect -9463 308 -9263 341
rect -9463 262 -9450 308
rect -9276 262 -9263 308
rect -9463 249 -9263 262
rect -9159 308 -8959 341
rect -9159 262 -9146 308
rect -8972 262 -8959 308
rect -9159 249 -8959 262
rect -8855 308 -8655 341
rect -8855 262 -8842 308
rect -8668 262 -8655 308
rect -8855 249 -8655 262
rect -8551 308 -8351 341
rect -8551 262 -8538 308
rect -8364 262 -8351 308
rect -8551 249 -8351 262
rect -7971 820 -7771 833
rect -7971 774 -7958 820
rect -7784 774 -7771 820
rect -7971 741 -7771 774
rect -7667 820 -7467 833
rect -7667 774 -7654 820
rect -7480 774 -7467 820
rect -7667 741 -7467 774
rect -7363 820 -7163 833
rect -7363 774 -7350 820
rect -7176 774 -7163 820
rect -7363 741 -7163 774
rect -7059 820 -6859 833
rect -7059 774 -7046 820
rect -6872 774 -6859 820
rect -7059 741 -6859 774
rect -6755 820 -6555 833
rect -6755 774 -6742 820
rect -6568 774 -6555 820
rect -6755 741 -6555 774
rect -7971 308 -7771 341
rect -7971 262 -7958 308
rect -7784 262 -7771 308
rect -7971 249 -7771 262
rect -7667 308 -7467 341
rect -7667 262 -7654 308
rect -7480 262 -7467 308
rect -7667 249 -7467 262
rect -7363 308 -7163 341
rect -7363 262 -7350 308
rect -7176 262 -7163 308
rect -7363 249 -7163 262
rect -7059 308 -6859 341
rect -7059 262 -7046 308
rect -6872 262 -6859 308
rect -7059 249 -6859 262
rect -6755 308 -6555 341
rect -6755 262 -6742 308
rect -6568 262 -6555 308
rect -6755 249 -6555 262
rect -9933 -665 -9733 -652
rect -9933 -711 -9920 -665
rect -9746 -711 -9733 -665
rect -9933 -744 -9733 -711
rect -9629 -665 -9429 -652
rect -9629 -711 -9616 -665
rect -9442 -711 -9429 -665
rect -9629 -744 -9429 -711
rect -9325 -665 -9125 -652
rect -9325 -711 -9312 -665
rect -9138 -711 -9125 -665
rect -9325 -744 -9125 -711
rect -9021 -665 -8821 -652
rect -9021 -711 -9008 -665
rect -8834 -711 -8821 -665
rect -9021 -744 -8821 -711
rect -8717 -665 -8517 -652
rect -8717 -711 -8704 -665
rect -8530 -711 -8517 -665
rect -8717 -744 -8517 -711
rect -8413 -665 -8213 -652
rect -8413 -711 -8400 -665
rect -8226 -711 -8213 -665
rect -8413 -744 -8213 -711
rect -8109 -665 -7909 -652
rect -8109 -711 -8096 -665
rect -7922 -711 -7909 -665
rect -8109 -744 -7909 -711
rect -7805 -665 -7605 -652
rect -7805 -711 -7792 -665
rect -7618 -711 -7605 -665
rect -7805 -744 -7605 -711
rect -7501 -665 -7301 -652
rect -7501 -711 -7488 -665
rect -7314 -711 -7301 -665
rect -7501 -744 -7301 -711
rect -7197 -665 -6997 -652
rect -7197 -711 -7184 -665
rect -7010 -711 -6997 -665
rect -7197 -744 -6997 -711
rect -6893 -665 -6693 -652
rect -6893 -711 -6880 -665
rect -6706 -711 -6693 -665
rect -6893 -744 -6693 -711
rect -6589 -665 -6389 -652
rect -6589 -711 -6576 -665
rect -6402 -711 -6389 -665
rect -6589 -744 -6389 -711
rect -9933 -1077 -9733 -1044
rect -9933 -1123 -9920 -1077
rect -9746 -1123 -9733 -1077
rect -9933 -1136 -9733 -1123
rect -9629 -1077 -9429 -1044
rect -9629 -1123 -9616 -1077
rect -9442 -1123 -9429 -1077
rect -9629 -1136 -9429 -1123
rect -9325 -1077 -9125 -1044
rect -9325 -1123 -9312 -1077
rect -9138 -1123 -9125 -1077
rect -9325 -1136 -9125 -1123
rect -9021 -1077 -8821 -1044
rect -9021 -1123 -9008 -1077
rect -8834 -1123 -8821 -1077
rect -9021 -1136 -8821 -1123
rect -8717 -1077 -8517 -1044
rect -8717 -1123 -8704 -1077
rect -8530 -1123 -8517 -1077
rect -8717 -1136 -8517 -1123
rect -8413 -1077 -8213 -1044
rect -8413 -1123 -8400 -1077
rect -8226 -1123 -8213 -1077
rect -8413 -1136 -8213 -1123
rect -8109 -1077 -7909 -1044
rect -8109 -1123 -8096 -1077
rect -7922 -1123 -7909 -1077
rect -8109 -1136 -7909 -1123
rect -7805 -1077 -7605 -1044
rect -7805 -1123 -7792 -1077
rect -7618 -1123 -7605 -1077
rect -7805 -1136 -7605 -1123
rect -7501 -1077 -7301 -1044
rect -7501 -1123 -7488 -1077
rect -7314 -1123 -7301 -1077
rect -7501 -1136 -7301 -1123
rect -7197 -1077 -6997 -1044
rect -7197 -1123 -7184 -1077
rect -7010 -1123 -6997 -1077
rect -7197 -1136 -6997 -1123
rect -6893 -1077 -6693 -1044
rect -6893 -1123 -6880 -1077
rect -6706 -1123 -6693 -1077
rect -6893 -1136 -6693 -1123
rect -6589 -1077 -6389 -1044
rect -6589 -1123 -6576 -1077
rect -6402 -1123 -6389 -1077
rect -6589 -1136 -6389 -1123
rect -9271 -1138 -9181 -1136
rect -9933 -1628 -9733 -1615
rect -9933 -1674 -9920 -1628
rect -9746 -1674 -9733 -1628
rect -9933 -1707 -9733 -1674
rect -9629 -1628 -9429 -1615
rect -9629 -1674 -9616 -1628
rect -9442 -1674 -9429 -1628
rect -9629 -1707 -9429 -1674
rect -9325 -1628 -9125 -1615
rect -9325 -1674 -9312 -1628
rect -9138 -1674 -9125 -1628
rect -9325 -1707 -9125 -1674
rect -9021 -1628 -8821 -1615
rect -9021 -1674 -9008 -1628
rect -8834 -1674 -8821 -1628
rect -9021 -1707 -8821 -1674
rect -8717 -1628 -8517 -1615
rect -8717 -1674 -8704 -1628
rect -8530 -1674 -8517 -1628
rect -8717 -1707 -8517 -1674
rect -8413 -1628 -8213 -1615
rect -8413 -1674 -8400 -1628
rect -8226 -1674 -8213 -1628
rect -8413 -1707 -8213 -1674
rect -8109 -1628 -7909 -1615
rect -8109 -1674 -8096 -1628
rect -7922 -1674 -7909 -1628
rect -8109 -1707 -7909 -1674
rect -7805 -1628 -7605 -1615
rect -7805 -1674 -7792 -1628
rect -7618 -1674 -7605 -1628
rect -7805 -1707 -7605 -1674
rect -7501 -1628 -7301 -1615
rect -7501 -1674 -7488 -1628
rect -7314 -1674 -7301 -1628
rect -7501 -1707 -7301 -1674
rect -7197 -1628 -6997 -1615
rect -7197 -1674 -7184 -1628
rect -7010 -1674 -6997 -1628
rect -7197 -1707 -6997 -1674
rect -6893 -1628 -6693 -1615
rect -6893 -1674 -6880 -1628
rect -6706 -1674 -6693 -1628
rect -6893 -1707 -6693 -1674
rect -6589 -1628 -6389 -1615
rect -6589 -1674 -6576 -1628
rect -6402 -1674 -6389 -1628
rect -6589 -1707 -6389 -1674
rect -9933 -2040 -9733 -2007
rect -9933 -2086 -9920 -2040
rect -9746 -2086 -9733 -2040
rect -9933 -2099 -9733 -2086
rect -9629 -2040 -9429 -2007
rect -9629 -2086 -9616 -2040
rect -9442 -2086 -9429 -2040
rect -9629 -2099 -9429 -2086
rect -9325 -2040 -9125 -2007
rect -9325 -2086 -9312 -2040
rect -9138 -2086 -9125 -2040
rect -9325 -2099 -9125 -2086
rect -9021 -2040 -8821 -2007
rect -9021 -2086 -9008 -2040
rect -8834 -2086 -8821 -2040
rect -9021 -2099 -8821 -2086
rect -8717 -2040 -8517 -2007
rect -8717 -2086 -8704 -2040
rect -8530 -2086 -8517 -2040
rect -8717 -2099 -8517 -2086
rect -8413 -2040 -8213 -2007
rect -8413 -2086 -8400 -2040
rect -8226 -2086 -8213 -2040
rect -8413 -2099 -8213 -2086
rect -8109 -2040 -7909 -2007
rect -8109 -2086 -8096 -2040
rect -7922 -2086 -7909 -2040
rect -8109 -2099 -7909 -2086
rect -7805 -2040 -7605 -2007
rect -7805 -2086 -7792 -2040
rect -7618 -2086 -7605 -2040
rect -7805 -2099 -7605 -2086
rect -7501 -2040 -7301 -2007
rect -7501 -2086 -7488 -2040
rect -7314 -2086 -7301 -2040
rect -7501 -2099 -7301 -2086
rect -7197 -2040 -6997 -2007
rect -7197 -2086 -7184 -2040
rect -7010 -2086 -6997 -2040
rect -7197 -2099 -6997 -2086
rect -6893 -2040 -6693 -2007
rect -6893 -2086 -6880 -2040
rect -6706 -2086 -6693 -2040
rect -6893 -2099 -6693 -2086
rect -6589 -2040 -6389 -2007
rect -6589 -2086 -6576 -2040
rect -6402 -2086 -6389 -2040
rect -6589 -2099 -6389 -2086
rect -8385 -2554 -8305 -2541
rect -8385 -2600 -8372 -2554
rect -8318 -2600 -8305 -2554
rect -8385 -2633 -8305 -2600
rect -8201 -2554 -8121 -2541
rect -8201 -2600 -8188 -2554
rect -8134 -2600 -8121 -2554
rect -8201 -2633 -8121 -2600
rect -8017 -2554 -7937 -2541
rect -8017 -2600 -8004 -2554
rect -7950 -2600 -7937 -2554
rect -8017 -2633 -7937 -2600
rect -8385 -2826 -8305 -2793
rect -8385 -2872 -8372 -2826
rect -8318 -2872 -8305 -2826
rect -8385 -2885 -8305 -2872
rect -8201 -2826 -8121 -2793
rect -8201 -2872 -8188 -2826
rect -8134 -2872 -8121 -2826
rect -8201 -2885 -8121 -2872
rect -8017 -2826 -7937 -2793
rect -8017 -2872 -8004 -2826
rect -7950 -2872 -7937 -2826
rect -8017 -2885 -7937 -2872
<< polycontact >>
rect 40608 38440 40654 38486
rect 40698 38290 40744 38336
rect -4618 37317 -4564 37363
rect -4434 37317 -4380 37363
rect -4250 37317 -4196 37363
rect -4618 36705 -4564 36751
rect -4434 36705 -4380 36751
rect -4250 36705 -4196 36751
rect 4854 37317 4908 37363
rect 5038 37317 5092 37363
rect 5222 37317 5276 37363
rect 4854 36705 4908 36751
rect 5038 36705 5092 36751
rect 5222 36705 5276 36751
rect 14326 37318 14380 37364
rect 14510 37318 14564 37364
rect 14694 37318 14748 37364
rect 14326 36706 14380 36752
rect 14510 36706 14564 36752
rect 14694 36706 14748 36752
rect 23798 37318 23852 37364
rect 23982 37318 24036 37364
rect 24166 37318 24220 37364
rect 23798 36706 23852 36752
rect 23982 36706 24036 36752
rect 24166 36706 24220 36752
rect 33270 37318 33324 37364
rect 33454 37318 33508 37364
rect 33638 37318 33692 37364
rect 33270 36706 33324 36752
rect 33454 36706 33508 36752
rect 33638 36706 33692 36752
rect 42742 37318 42796 37364
rect 42926 37318 42980 37364
rect 43110 37318 43164 37364
rect 42742 36706 42796 36752
rect 42926 36706 42980 36752
rect 43110 36706 43164 36752
rect -4618 36157 -4564 36203
rect -4434 36157 -4380 36203
rect -4250 36157 -4196 36203
rect -4618 35845 -4564 35891
rect -4434 35845 -4380 35891
rect -4250 35845 -4196 35891
rect 4854 36157 4908 36203
rect 5038 36157 5092 36203
rect 5222 36157 5276 36203
rect 4854 35845 4908 35891
rect 5038 35845 5092 35891
rect 5222 35845 5276 35891
rect 14326 36158 14380 36204
rect 14510 36158 14564 36204
rect 14694 36158 14748 36204
rect 14326 35846 14380 35892
rect 14510 35846 14564 35892
rect 14694 35846 14748 35892
rect 23798 36158 23852 36204
rect 23982 36158 24036 36204
rect 24166 36158 24220 36204
rect 23798 35846 23852 35892
rect 23982 35846 24036 35892
rect 24166 35846 24220 35892
rect 33270 36158 33324 36204
rect 33454 36158 33508 36204
rect 33638 36158 33692 36204
rect 33270 35846 33324 35892
rect 33454 35846 33508 35892
rect 33638 35846 33692 35892
rect 42742 36158 42796 36204
rect 42926 36158 42980 36204
rect 43110 36158 43164 36204
rect 42742 35846 42796 35892
rect 42926 35846 42980 35892
rect 43110 35846 43164 35892
rect -4618 35112 -4564 35158
rect -4434 35112 -4380 35158
rect -4250 35112 -4196 35158
rect -4618 34500 -4564 34546
rect -4434 34500 -4380 34546
rect -4250 34500 -4196 34546
rect -3132 35112 -3078 35158
rect -2948 35112 -2894 35158
rect -2764 35112 -2710 35158
rect -3132 34500 -3078 34546
rect -2948 34500 -2894 34546
rect -2764 34500 -2710 34546
rect 4854 35112 4908 35158
rect 5038 35112 5092 35158
rect 5222 35112 5276 35158
rect 4854 34500 4908 34546
rect 5038 34500 5092 34546
rect 5222 34500 5276 34546
rect 6340 35112 6394 35158
rect 6524 35112 6578 35158
rect 6708 35112 6762 35158
rect 6340 34500 6394 34546
rect 6524 34500 6578 34546
rect 6708 34500 6762 34546
rect 14326 35113 14380 35159
rect 14510 35113 14564 35159
rect 14694 35113 14748 35159
rect 14326 34501 14380 34547
rect 14510 34501 14564 34547
rect 14694 34501 14748 34547
rect 15812 35113 15866 35159
rect 15996 35113 16050 35159
rect 16180 35113 16234 35159
rect 15812 34501 15866 34547
rect 15996 34501 16050 34547
rect 16180 34501 16234 34547
rect 23798 35113 23852 35159
rect 23982 35113 24036 35159
rect 24166 35113 24220 35159
rect 23798 34501 23852 34547
rect 23982 34501 24036 34547
rect 24166 34501 24220 34547
rect 25284 35113 25338 35159
rect 25468 35113 25522 35159
rect 25652 35113 25706 35159
rect 25284 34501 25338 34547
rect 25468 34501 25522 34547
rect 25652 34501 25706 34547
rect 33270 35113 33324 35159
rect 33454 35113 33508 35159
rect 33638 35113 33692 35159
rect 33270 34501 33324 34547
rect 33454 34501 33508 34547
rect 33638 34501 33692 34547
rect 34756 35113 34810 35159
rect 34940 35113 34994 35159
rect 35124 35113 35178 35159
rect 34756 34501 34810 34547
rect 34940 34501 34994 34547
rect 35124 34501 35178 34547
rect 42742 35113 42796 35159
rect 42926 35113 42980 35159
rect 43110 35113 43164 35159
rect 42742 34501 42796 34547
rect 42926 34501 42980 34547
rect 43110 34501 43164 34547
rect 44228 35113 44282 35159
rect 44412 35113 44466 35159
rect 44596 35113 44650 35159
rect 44228 34501 44282 34547
rect 44412 34501 44466 34547
rect 44596 34501 44650 34547
rect -4618 33952 -4564 33998
rect -4434 33952 -4380 33998
rect -4250 33952 -4196 33998
rect -4618 33640 -4564 33686
rect -4434 33640 -4380 33686
rect -4250 33640 -4196 33686
rect -3132 33952 -3078 33998
rect -2948 33952 -2894 33998
rect -2764 33952 -2710 33998
rect -3132 33640 -3078 33686
rect -2948 33640 -2894 33686
rect -2764 33640 -2710 33686
rect 4854 33952 4908 33998
rect 5038 33952 5092 33998
rect 5222 33952 5276 33998
rect 4854 33640 4908 33686
rect 5038 33640 5092 33686
rect 5222 33640 5276 33686
rect 6340 33952 6394 33998
rect 6524 33952 6578 33998
rect 6708 33952 6762 33998
rect 6340 33640 6394 33686
rect 6524 33640 6578 33686
rect 6708 33640 6762 33686
rect 14326 33953 14380 33999
rect 14510 33953 14564 33999
rect 14694 33953 14748 33999
rect 14326 33641 14380 33687
rect 14510 33641 14564 33687
rect 14694 33641 14748 33687
rect 15812 33953 15866 33999
rect 15996 33953 16050 33999
rect 16180 33953 16234 33999
rect 15812 33641 15866 33687
rect 15996 33641 16050 33687
rect 16180 33641 16234 33687
rect 23798 33953 23852 33999
rect 23982 33953 24036 33999
rect 24166 33953 24220 33999
rect 23798 33641 23852 33687
rect 23982 33641 24036 33687
rect 24166 33641 24220 33687
rect 25284 33953 25338 33999
rect 25468 33953 25522 33999
rect 25652 33953 25706 33999
rect 25284 33641 25338 33687
rect 25468 33641 25522 33687
rect 25652 33641 25706 33687
rect 33270 33953 33324 33999
rect 33454 33953 33508 33999
rect 33638 33953 33692 33999
rect 33270 33641 33324 33687
rect 33454 33641 33508 33687
rect 33638 33641 33692 33687
rect 34756 33953 34810 33999
rect 34940 33953 34994 33999
rect 35124 33953 35178 33999
rect 34756 33641 34810 33687
rect 34940 33641 34994 33687
rect 35124 33641 35178 33687
rect 42742 33953 42796 33999
rect 42926 33953 42980 33999
rect 43110 33953 43164 33999
rect 42742 33641 42796 33687
rect 42926 33641 42980 33687
rect 43110 33641 43164 33687
rect 44228 33953 44282 33999
rect 44412 33953 44466 33999
rect 44596 33953 44650 33999
rect 44228 33641 44282 33687
rect 44412 33641 44466 33687
rect 44596 33641 44650 33687
rect -4618 32907 -4564 32953
rect -4434 32907 -4380 32953
rect -4250 32907 -4196 32953
rect -4618 32295 -4564 32341
rect -4434 32295 -4380 32341
rect -4250 32295 -4196 32341
rect -3132 32908 -3078 32954
rect -2948 32908 -2894 32954
rect -2764 32908 -2710 32954
rect -3132 32296 -3078 32342
rect -2948 32296 -2894 32342
rect -2764 32296 -2710 32342
rect 4854 32907 4908 32953
rect 5038 32907 5092 32953
rect 5222 32907 5276 32953
rect 4854 32295 4908 32341
rect 5038 32295 5092 32341
rect 5222 32295 5276 32341
rect 6340 32908 6394 32954
rect 6524 32908 6578 32954
rect 6708 32908 6762 32954
rect 6340 32296 6394 32342
rect 6524 32296 6578 32342
rect 6708 32296 6762 32342
rect 14326 32908 14380 32954
rect 14510 32908 14564 32954
rect 14694 32908 14748 32954
rect 14326 32296 14380 32342
rect 14510 32296 14564 32342
rect 14694 32296 14748 32342
rect 15812 32909 15866 32955
rect 15996 32909 16050 32955
rect 16180 32909 16234 32955
rect 15812 32297 15866 32343
rect 15996 32297 16050 32343
rect 16180 32297 16234 32343
rect 23798 32908 23852 32954
rect 23982 32908 24036 32954
rect 24166 32908 24220 32954
rect 23798 32296 23852 32342
rect 23982 32296 24036 32342
rect 24166 32296 24220 32342
rect 25284 32909 25338 32955
rect 25468 32909 25522 32955
rect 25652 32909 25706 32955
rect 25284 32297 25338 32343
rect 25468 32297 25522 32343
rect 25652 32297 25706 32343
rect 33270 32908 33324 32954
rect 33454 32908 33508 32954
rect 33638 32908 33692 32954
rect 33270 32296 33324 32342
rect 33454 32296 33508 32342
rect 33638 32296 33692 32342
rect 34756 32909 34810 32955
rect 34940 32909 34994 32955
rect 35124 32909 35178 32955
rect 34756 32297 34810 32343
rect 34940 32297 34994 32343
rect 35124 32297 35178 32343
rect 42742 32908 42796 32954
rect 42926 32908 42980 32954
rect 43110 32908 43164 32954
rect 42742 32296 42796 32342
rect 42926 32296 42980 32342
rect 43110 32296 43164 32342
rect 44228 32909 44282 32955
rect 44412 32909 44466 32955
rect 44596 32909 44650 32955
rect 44228 32297 44282 32343
rect 44412 32297 44466 32343
rect 44596 32297 44650 32343
rect -9760 31792 -9686 31838
rect -9760 31080 -9686 31126
rect -8872 31792 -8798 31838
rect -8872 31080 -8798 31126
rect -8392 31792 -8318 31838
rect -8392 31080 -8318 31126
rect -4618 31747 -4564 31793
rect -4434 31747 -4380 31793
rect -4250 31747 -4196 31793
rect -4618 31435 -4564 31481
rect -4434 31435 -4380 31481
rect -4250 31435 -4196 31481
rect -3132 31748 -3078 31794
rect -2948 31748 -2894 31794
rect -2764 31748 -2710 31794
rect -3132 31436 -3078 31482
rect -2948 31436 -2894 31482
rect -2764 31436 -2710 31482
rect -288 31792 -214 31838
rect -288 31080 -214 31126
rect 600 31792 674 31838
rect 600 31080 674 31126
rect 1080 31792 1154 31838
rect 1080 31080 1154 31126
rect 4854 31747 4908 31793
rect 5038 31747 5092 31793
rect 5222 31747 5276 31793
rect 4854 31435 4908 31481
rect 5038 31435 5092 31481
rect 5222 31435 5276 31481
rect 6340 31748 6394 31794
rect 6524 31748 6578 31794
rect 6708 31748 6762 31794
rect 6340 31436 6394 31482
rect 6524 31436 6578 31482
rect 6708 31436 6762 31482
rect 9184 31793 9258 31839
rect 9184 31081 9258 31127
rect 10072 31793 10146 31839
rect 10072 31081 10146 31127
rect 10552 31793 10626 31839
rect 10552 31081 10626 31127
rect 14326 31748 14380 31794
rect 14510 31748 14564 31794
rect 14694 31748 14748 31794
rect 14326 31436 14380 31482
rect 14510 31436 14564 31482
rect 14694 31436 14748 31482
rect 15812 31749 15866 31795
rect 15996 31749 16050 31795
rect 16180 31749 16234 31795
rect 15812 31437 15866 31483
rect 15996 31437 16050 31483
rect 16180 31437 16234 31483
rect 18656 31793 18730 31839
rect 18656 31081 18730 31127
rect 19544 31793 19618 31839
rect 19544 31081 19618 31127
rect 20024 31793 20098 31839
rect 20024 31081 20098 31127
rect 23798 31748 23852 31794
rect 23982 31748 24036 31794
rect 24166 31748 24220 31794
rect 23798 31436 23852 31482
rect 23982 31436 24036 31482
rect 24166 31436 24220 31482
rect 25284 31749 25338 31795
rect 25468 31749 25522 31795
rect 25652 31749 25706 31795
rect 25284 31437 25338 31483
rect 25468 31437 25522 31483
rect 25652 31437 25706 31483
rect 28128 31793 28202 31839
rect 28128 31081 28202 31127
rect 29016 31793 29090 31839
rect 29016 31081 29090 31127
rect 29496 31793 29570 31839
rect 29496 31081 29570 31127
rect 33270 31748 33324 31794
rect 33454 31748 33508 31794
rect 33638 31748 33692 31794
rect 33270 31436 33324 31482
rect 33454 31436 33508 31482
rect 33638 31436 33692 31482
rect 34756 31749 34810 31795
rect 34940 31749 34994 31795
rect 35124 31749 35178 31795
rect 34756 31437 34810 31483
rect 34940 31437 34994 31483
rect 35124 31437 35178 31483
rect 37600 31793 37674 31839
rect 37600 31081 37674 31127
rect 38488 31793 38562 31839
rect 38488 31081 38562 31127
rect 38968 31793 39042 31839
rect 38968 31081 39042 31127
rect 42742 31748 42796 31794
rect 42926 31748 42980 31794
rect 43110 31748 43164 31794
rect 42742 31436 42796 31482
rect 42926 31436 42980 31482
rect 43110 31436 43164 31482
rect 44228 31749 44282 31795
rect 44412 31749 44466 31795
rect 44596 31749 44650 31795
rect 44228 31437 44282 31483
rect 44412 31437 44466 31483
rect 44596 31437 44650 31483
rect -10654 30372 -10580 30418
rect -10654 29660 -10580 29706
rect -9760 30672 -9686 30718
rect -9556 30672 -9482 30718
rect -9760 30360 -9686 30406
rect -9556 30360 -9482 30406
rect -9076 30672 -9002 30718
rect -8872 30672 -8798 30718
rect -9076 30360 -9002 30406
rect -8872 30360 -8798 30406
rect -8392 30672 -8318 30718
rect -8392 30360 -8318 30406
rect -7532 30616 -7458 30662
rect -7328 30616 -7254 30662
rect -7532 29904 -7458 29950
rect -7328 29904 -7254 29950
rect -6848 30616 -6774 30662
rect -6644 30616 -6570 30662
rect -6848 29904 -6774 29950
rect -6644 29904 -6570 29950
rect -6164 30616 -6090 30662
rect -6164 29904 -6090 29950
rect -4618 30702 -4564 30748
rect -4434 30702 -4380 30748
rect -4250 30702 -4196 30748
rect -4618 30090 -4564 30136
rect -4434 30090 -4380 30136
rect -4250 30090 -4196 30136
rect -10654 29252 -10580 29298
rect -10654 28940 -10580 28986
rect -9760 29452 -9686 29498
rect -9760 28740 -9686 28786
rect -8872 29452 -8798 29498
rect -8872 28740 -8798 28786
rect -8392 29452 -8318 29498
rect -8392 28740 -8318 28786
rect -7532 29496 -7458 29542
rect -7532 29184 -7458 29230
rect -6848 29496 -6774 29542
rect -6848 29184 -6774 29230
rect -6164 29496 -6090 29542
rect -6164 29184 -6090 29230
rect -4618 29542 -4564 29588
rect -4434 29542 -4380 29588
rect -4250 29542 -4196 29588
rect -4618 29230 -4564 29276
rect -4434 29230 -4380 29276
rect -4250 29230 -4196 29276
rect -1182 30372 -1108 30418
rect -1182 29660 -1108 29706
rect -288 30672 -214 30718
rect -84 30672 -10 30718
rect -288 30360 -214 30406
rect -84 30360 -10 30406
rect 396 30672 470 30718
rect 600 30672 674 30718
rect 396 30360 470 30406
rect 600 30360 674 30406
rect 1080 30672 1154 30718
rect 1080 30360 1154 30406
rect 1940 30616 2014 30662
rect 2144 30616 2218 30662
rect 1940 29904 2014 29950
rect 2144 29904 2218 29950
rect 2624 30616 2698 30662
rect 2828 30616 2902 30662
rect 2624 29904 2698 29950
rect 2828 29904 2902 29950
rect 3308 30616 3382 30662
rect 3308 29904 3382 29950
rect 4854 30702 4908 30748
rect 5038 30702 5092 30748
rect 5222 30702 5276 30748
rect 4854 30090 4908 30136
rect 5038 30090 5092 30136
rect 5222 30090 5276 30136
rect -1182 29252 -1108 29298
rect -1182 28940 -1108 28986
rect -288 29452 -214 29498
rect -288 28740 -214 28786
rect 600 29452 674 29498
rect 600 28740 674 28786
rect 1080 29452 1154 29498
rect 1080 28740 1154 28786
rect 1940 29496 2014 29542
rect 1940 29184 2014 29230
rect 2624 29496 2698 29542
rect 2624 29184 2698 29230
rect 3308 29496 3382 29542
rect 3308 29184 3382 29230
rect 4854 29542 4908 29588
rect 5038 29542 5092 29588
rect 5222 29542 5276 29588
rect 4854 29230 4908 29276
rect 5038 29230 5092 29276
rect 5222 29230 5276 29276
rect 8290 30373 8364 30419
rect 8290 29661 8364 29707
rect 9184 30673 9258 30719
rect 9388 30673 9462 30719
rect 9184 30361 9258 30407
rect 9388 30361 9462 30407
rect 9868 30673 9942 30719
rect 10072 30673 10146 30719
rect 9868 30361 9942 30407
rect 10072 30361 10146 30407
rect 10552 30673 10626 30719
rect 10552 30361 10626 30407
rect 11412 30617 11486 30663
rect 11616 30617 11690 30663
rect 11412 29905 11486 29951
rect 11616 29905 11690 29951
rect 12096 30617 12170 30663
rect 12300 30617 12374 30663
rect 12096 29905 12170 29951
rect 12300 29905 12374 29951
rect 12780 30617 12854 30663
rect 12780 29905 12854 29951
rect 14326 30703 14380 30749
rect 14510 30703 14564 30749
rect 14694 30703 14748 30749
rect 14326 30091 14380 30137
rect 14510 30091 14564 30137
rect 14694 30091 14748 30137
rect 8290 29253 8364 29299
rect 8290 28941 8364 28987
rect 9184 29453 9258 29499
rect 9184 28741 9258 28787
rect 10072 29453 10146 29499
rect 10072 28741 10146 28787
rect 10552 29453 10626 29499
rect 10552 28741 10626 28787
rect 11412 29497 11486 29543
rect 11412 29185 11486 29231
rect 12096 29497 12170 29543
rect 12096 29185 12170 29231
rect 12780 29497 12854 29543
rect 12780 29185 12854 29231
rect 14326 29543 14380 29589
rect 14510 29543 14564 29589
rect 14694 29543 14748 29589
rect 14326 29231 14380 29277
rect 14510 29231 14564 29277
rect 14694 29231 14748 29277
rect 17762 30373 17836 30419
rect 17762 29661 17836 29707
rect 18656 30673 18730 30719
rect 18860 30673 18934 30719
rect 18656 30361 18730 30407
rect 18860 30361 18934 30407
rect 19340 30673 19414 30719
rect 19544 30673 19618 30719
rect 19340 30361 19414 30407
rect 19544 30361 19618 30407
rect 20024 30673 20098 30719
rect 20024 30361 20098 30407
rect 20884 30617 20958 30663
rect 21088 30617 21162 30663
rect 20884 29905 20958 29951
rect 21088 29905 21162 29951
rect 21568 30617 21642 30663
rect 21772 30617 21846 30663
rect 21568 29905 21642 29951
rect 21772 29905 21846 29951
rect 22252 30617 22326 30663
rect 22252 29905 22326 29951
rect 23798 30703 23852 30749
rect 23982 30703 24036 30749
rect 24166 30703 24220 30749
rect 23798 30091 23852 30137
rect 23982 30091 24036 30137
rect 24166 30091 24220 30137
rect 17762 29253 17836 29299
rect 17762 28941 17836 28987
rect 18656 29453 18730 29499
rect 18656 28741 18730 28787
rect 19544 29453 19618 29499
rect 19544 28741 19618 28787
rect 20024 29453 20098 29499
rect 20024 28741 20098 28787
rect 20884 29497 20958 29543
rect 20884 29185 20958 29231
rect 21568 29497 21642 29543
rect 21568 29185 21642 29231
rect 22252 29497 22326 29543
rect 22252 29185 22326 29231
rect 23798 29543 23852 29589
rect 23982 29543 24036 29589
rect 24166 29543 24220 29589
rect 23798 29231 23852 29277
rect 23982 29231 24036 29277
rect 24166 29231 24220 29277
rect 27234 30373 27308 30419
rect 27234 29661 27308 29707
rect 28128 30673 28202 30719
rect 28332 30673 28406 30719
rect 28128 30361 28202 30407
rect 28332 30361 28406 30407
rect 28812 30673 28886 30719
rect 29016 30673 29090 30719
rect 28812 30361 28886 30407
rect 29016 30361 29090 30407
rect 29496 30673 29570 30719
rect 29496 30361 29570 30407
rect 30356 30617 30430 30663
rect 30560 30617 30634 30663
rect 30356 29905 30430 29951
rect 30560 29905 30634 29951
rect 31040 30617 31114 30663
rect 31244 30617 31318 30663
rect 31040 29905 31114 29951
rect 31244 29905 31318 29951
rect 31724 30617 31798 30663
rect 31724 29905 31798 29951
rect 33270 30703 33324 30749
rect 33454 30703 33508 30749
rect 33638 30703 33692 30749
rect 33270 30091 33324 30137
rect 33454 30091 33508 30137
rect 33638 30091 33692 30137
rect 27234 29253 27308 29299
rect 27234 28941 27308 28987
rect 28128 29453 28202 29499
rect 28128 28741 28202 28787
rect 29016 29453 29090 29499
rect 29016 28741 29090 28787
rect 29496 29453 29570 29499
rect 29496 28741 29570 28787
rect 30356 29497 30430 29543
rect 30356 29185 30430 29231
rect 31040 29497 31114 29543
rect 31040 29185 31114 29231
rect 31724 29497 31798 29543
rect 31724 29185 31798 29231
rect 33270 29543 33324 29589
rect 33454 29543 33508 29589
rect 33638 29543 33692 29589
rect 33270 29231 33324 29277
rect 33454 29231 33508 29277
rect 33638 29231 33692 29277
rect 36706 30373 36780 30419
rect 36706 29661 36780 29707
rect 37600 30673 37674 30719
rect 37804 30673 37878 30719
rect 37600 30361 37674 30407
rect 37804 30361 37878 30407
rect 38284 30673 38358 30719
rect 38488 30673 38562 30719
rect 38284 30361 38358 30407
rect 38488 30361 38562 30407
rect 38968 30673 39042 30719
rect 38968 30361 39042 30407
rect 39828 30617 39902 30663
rect 40032 30617 40106 30663
rect 39828 29905 39902 29951
rect 40032 29905 40106 29951
rect 40512 30617 40586 30663
rect 40716 30617 40790 30663
rect 40512 29905 40586 29951
rect 40716 29905 40790 29951
rect 41196 30617 41270 30663
rect 41196 29905 41270 29951
rect 42742 30703 42796 30749
rect 42926 30703 42980 30749
rect 43110 30703 43164 30749
rect 42742 30091 42796 30137
rect 42926 30091 42980 30137
rect 43110 30091 43164 30137
rect 36706 29253 36780 29299
rect 36706 28941 36780 28987
rect 37600 29453 37674 29499
rect 37600 28741 37674 28787
rect 38488 29453 38562 29499
rect 38488 28741 38562 28787
rect 38968 29453 39042 29499
rect 38968 28741 39042 28787
rect 39828 29497 39902 29543
rect 39828 29185 39902 29231
rect 40512 29497 40586 29543
rect 40512 29185 40586 29231
rect 41196 29497 41270 29543
rect 41196 29185 41270 29231
rect 42742 29543 42796 29589
rect 42926 29543 42980 29589
rect 43110 29543 43164 29589
rect 42742 29231 42796 29277
rect 42926 29231 42980 29277
rect 43110 29231 43164 29277
rect -12367 28442 -12293 28488
rect -12367 27730 -12293 27776
rect -9760 28332 -9686 28378
rect -9556 28332 -9482 28378
rect -9760 28020 -9686 28066
rect -9556 28020 -9482 28066
rect -9076 28332 -9002 28378
rect -8872 28332 -8798 28378
rect -9076 28020 -9002 28066
rect -8872 28020 -8798 28066
rect -8392 28332 -8318 28378
rect -8392 28020 -8318 28066
rect -288 28332 -214 28378
rect -84 28332 -10 28378
rect -288 28020 -214 28066
rect -84 28020 -10 28066
rect 396 28332 470 28378
rect 600 28332 674 28378
rect 396 28020 470 28066
rect 600 28020 674 28066
rect 1080 28332 1154 28378
rect 1080 28020 1154 28066
rect 9184 28333 9258 28379
rect 9388 28333 9462 28379
rect 9184 28021 9258 28067
rect 9388 28021 9462 28067
rect 9868 28333 9942 28379
rect 10072 28333 10146 28379
rect 9868 28021 9942 28067
rect 10072 28021 10146 28067
rect 10552 28333 10626 28379
rect 10552 28021 10626 28067
rect 18656 28333 18730 28379
rect 18860 28333 18934 28379
rect 18656 28021 18730 28067
rect 18860 28021 18934 28067
rect 19340 28333 19414 28379
rect 19544 28333 19618 28379
rect 19340 28021 19414 28067
rect 19544 28021 19618 28067
rect 20024 28333 20098 28379
rect 20024 28021 20098 28067
rect 28128 28333 28202 28379
rect 28332 28333 28406 28379
rect 28128 28021 28202 28067
rect 28332 28021 28406 28067
rect 28812 28333 28886 28379
rect 29016 28333 29090 28379
rect 28812 28021 28886 28067
rect 29016 28021 29090 28067
rect 29496 28333 29570 28379
rect 29496 28021 29570 28067
rect 37600 28333 37674 28379
rect 37804 28333 37878 28379
rect 37600 28021 37674 28067
rect 37804 28021 37878 28067
rect 38284 28333 38358 28379
rect 38488 28333 38562 28379
rect 38284 28021 38358 28067
rect 38488 28021 38562 28067
rect 38968 28333 39042 28379
rect 38968 28021 39042 28067
rect -12367 27322 -12293 27368
rect -12367 27010 -12293 27056
rect -7876 25015 -7822 25061
rect -7692 25015 -7638 25061
rect -7508 25015 -7454 25061
rect -7876 24403 -7822 24449
rect -7692 24403 -7638 24449
rect -7508 24403 -7454 24449
rect -3834 25012 -3780 25058
rect -3650 25012 -3596 25058
rect -3466 25012 -3412 25058
rect -3834 24400 -3780 24446
rect -3650 24400 -3596 24446
rect -3466 24400 -3412 24446
rect 208 25012 262 25058
rect 392 25012 446 25058
rect 576 25012 630 25058
rect 208 24400 262 24446
rect 392 24400 446 24446
rect 576 24400 630 24446
rect 4250 25012 4304 25058
rect 4434 25012 4488 25058
rect 4618 25012 4672 25058
rect 4250 24400 4304 24446
rect 4434 24400 4488 24446
rect 4618 24400 4672 24446
rect 8292 25012 8346 25058
rect 8476 25012 8530 25058
rect 8660 25012 8714 25058
rect 8292 24400 8346 24446
rect 8476 24400 8530 24446
rect 8660 24400 8714 24446
rect 12334 25012 12388 25058
rect 12518 25012 12572 25058
rect 12702 25012 12756 25058
rect 12334 24400 12388 24446
rect 12518 24400 12572 24446
rect 12702 24400 12756 24446
rect 16376 25012 16430 25058
rect 16560 25012 16614 25058
rect 16744 25012 16798 25058
rect 16376 24400 16430 24446
rect 16560 24400 16614 24446
rect 16744 24400 16798 24446
rect -7876 23855 -7822 23901
rect -7692 23855 -7638 23901
rect -7508 23855 -7454 23901
rect -7876 23543 -7822 23589
rect -7692 23543 -7638 23589
rect -7508 23543 -7454 23589
rect -3834 23852 -3780 23898
rect -3650 23852 -3596 23898
rect -3466 23852 -3412 23898
rect -3834 23540 -3780 23586
rect -3650 23540 -3596 23586
rect -3466 23540 -3412 23586
rect 208 23852 262 23898
rect 392 23852 446 23898
rect 576 23852 630 23898
rect 208 23540 262 23586
rect 392 23540 446 23586
rect 576 23540 630 23586
rect 4250 23852 4304 23898
rect 4434 23852 4488 23898
rect 4618 23852 4672 23898
rect 4250 23540 4304 23586
rect 4434 23540 4488 23586
rect 4618 23540 4672 23586
rect 8292 23852 8346 23898
rect 8476 23852 8530 23898
rect 8660 23852 8714 23898
rect 8292 23540 8346 23586
rect 8476 23540 8530 23586
rect 8660 23540 8714 23586
rect 12334 23852 12388 23898
rect 12518 23852 12572 23898
rect 12702 23852 12756 23898
rect 12334 23540 12388 23586
rect 12518 23540 12572 23586
rect 12702 23540 12756 23586
rect 16376 23852 16430 23898
rect 16560 23852 16614 23898
rect 16744 23852 16798 23898
rect 16376 23540 16430 23586
rect 16560 23540 16614 23586
rect 16744 23540 16798 23586
rect -7876 22810 -7822 22856
rect -7692 22810 -7638 22856
rect -7508 22810 -7454 22856
rect -7876 22198 -7822 22244
rect -7692 22198 -7638 22244
rect -7508 22198 -7454 22244
rect -6390 22810 -6336 22856
rect -6206 22810 -6152 22856
rect -6022 22810 -5968 22856
rect -6390 22198 -6336 22244
rect -6206 22198 -6152 22244
rect -6022 22198 -5968 22244
rect -3834 22807 -3780 22853
rect -3650 22807 -3596 22853
rect -3466 22807 -3412 22853
rect -3834 22195 -3780 22241
rect -3650 22195 -3596 22241
rect -3466 22195 -3412 22241
rect -2348 22807 -2294 22853
rect -2164 22807 -2110 22853
rect -1980 22807 -1926 22853
rect -2348 22195 -2294 22241
rect -2164 22195 -2110 22241
rect -1980 22195 -1926 22241
rect 208 22807 262 22853
rect 392 22807 446 22853
rect 576 22807 630 22853
rect 208 22195 262 22241
rect 392 22195 446 22241
rect 576 22195 630 22241
rect 1694 22807 1748 22853
rect 1878 22807 1932 22853
rect 2062 22807 2116 22853
rect 1694 22195 1748 22241
rect 1878 22195 1932 22241
rect 2062 22195 2116 22241
rect 4250 22807 4304 22853
rect 4434 22807 4488 22853
rect 4618 22807 4672 22853
rect 4250 22195 4304 22241
rect 4434 22195 4488 22241
rect 4618 22195 4672 22241
rect 5736 22807 5790 22853
rect 5920 22807 5974 22853
rect 6104 22807 6158 22853
rect 5736 22195 5790 22241
rect 5920 22195 5974 22241
rect 6104 22195 6158 22241
rect 8292 22807 8346 22853
rect 8476 22807 8530 22853
rect 8660 22807 8714 22853
rect 8292 22195 8346 22241
rect 8476 22195 8530 22241
rect 8660 22195 8714 22241
rect 9778 22807 9832 22853
rect 9962 22807 10016 22853
rect 10146 22807 10200 22853
rect 9778 22195 9832 22241
rect 9962 22195 10016 22241
rect 10146 22195 10200 22241
rect 12334 22807 12388 22853
rect 12518 22807 12572 22853
rect 12702 22807 12756 22853
rect 12334 22195 12388 22241
rect 12518 22195 12572 22241
rect 12702 22195 12756 22241
rect 13820 22807 13874 22853
rect 14004 22807 14058 22853
rect 14188 22807 14242 22853
rect 13820 22195 13874 22241
rect 14004 22195 14058 22241
rect 14188 22195 14242 22241
rect 16376 22807 16430 22853
rect 16560 22807 16614 22853
rect 16744 22807 16798 22853
rect 16376 22195 16430 22241
rect 16560 22195 16614 22241
rect 16744 22195 16798 22241
rect 17862 22807 17916 22853
rect 18046 22807 18100 22853
rect 18230 22807 18284 22853
rect 17862 22195 17916 22241
rect 18046 22195 18100 22241
rect 18230 22195 18284 22241
rect -7876 21650 -7822 21696
rect -7692 21650 -7638 21696
rect -7508 21650 -7454 21696
rect -7876 21338 -7822 21384
rect -7692 21338 -7638 21384
rect -7508 21338 -7454 21384
rect -6390 21650 -6336 21696
rect -6206 21650 -6152 21696
rect -6022 21650 -5968 21696
rect -6390 21338 -6336 21384
rect -6206 21338 -6152 21384
rect -6022 21338 -5968 21384
rect -3834 21647 -3780 21693
rect -3650 21647 -3596 21693
rect -3466 21647 -3412 21693
rect -3834 21335 -3780 21381
rect -3650 21335 -3596 21381
rect -3466 21335 -3412 21381
rect -2348 21647 -2294 21693
rect -2164 21647 -2110 21693
rect -1980 21647 -1926 21693
rect -2348 21335 -2294 21381
rect -2164 21335 -2110 21381
rect -1980 21335 -1926 21381
rect 208 21647 262 21693
rect 392 21647 446 21693
rect 576 21647 630 21693
rect 208 21335 262 21381
rect 392 21335 446 21381
rect 576 21335 630 21381
rect 1694 21647 1748 21693
rect 1878 21647 1932 21693
rect 2062 21647 2116 21693
rect 1694 21335 1748 21381
rect 1878 21335 1932 21381
rect 2062 21335 2116 21381
rect 4250 21647 4304 21693
rect 4434 21647 4488 21693
rect 4618 21647 4672 21693
rect 4250 21335 4304 21381
rect 4434 21335 4488 21381
rect 4618 21335 4672 21381
rect 5736 21647 5790 21693
rect 5920 21647 5974 21693
rect 6104 21647 6158 21693
rect 5736 21335 5790 21381
rect 5920 21335 5974 21381
rect 6104 21335 6158 21381
rect 8292 21647 8346 21693
rect 8476 21647 8530 21693
rect 8660 21647 8714 21693
rect 8292 21335 8346 21381
rect 8476 21335 8530 21381
rect 8660 21335 8714 21381
rect 9778 21647 9832 21693
rect 9962 21647 10016 21693
rect 10146 21647 10200 21693
rect 9778 21335 9832 21381
rect 9962 21335 10016 21381
rect 10146 21335 10200 21381
rect 12334 21647 12388 21693
rect 12518 21647 12572 21693
rect 12702 21647 12756 21693
rect 12334 21335 12388 21381
rect 12518 21335 12572 21381
rect 12702 21335 12756 21381
rect 13820 21647 13874 21693
rect 14004 21647 14058 21693
rect 14188 21647 14242 21693
rect 13820 21335 13874 21381
rect 14004 21335 14058 21381
rect 14188 21335 14242 21381
rect 16376 21647 16430 21693
rect 16560 21647 16614 21693
rect 16744 21647 16798 21693
rect 16376 21335 16430 21381
rect 16560 21335 16614 21381
rect 16744 21335 16798 21381
rect 17862 21647 17916 21693
rect 18046 21647 18100 21693
rect 18230 21647 18284 21693
rect 17862 21335 17916 21381
rect 18046 21335 18100 21381
rect 18230 21335 18284 21381
rect -7876 20605 -7822 20651
rect -7692 20605 -7638 20651
rect -7508 20605 -7454 20651
rect -7876 19993 -7822 20039
rect -7692 19993 -7638 20039
rect -7508 19993 -7454 20039
rect -6390 20606 -6336 20652
rect -6206 20606 -6152 20652
rect -6022 20606 -5968 20652
rect -6390 19994 -6336 20040
rect -6206 19994 -6152 20040
rect -6022 19994 -5968 20040
rect -3834 20602 -3780 20648
rect -3650 20602 -3596 20648
rect -3466 20602 -3412 20648
rect -3834 19990 -3780 20036
rect -3650 19990 -3596 20036
rect -3466 19990 -3412 20036
rect -2348 20603 -2294 20649
rect -2164 20603 -2110 20649
rect -1980 20603 -1926 20649
rect -2348 19991 -2294 20037
rect -2164 19991 -2110 20037
rect -1980 19991 -1926 20037
rect 208 20602 262 20648
rect 392 20602 446 20648
rect 576 20602 630 20648
rect 208 19990 262 20036
rect 392 19990 446 20036
rect 576 19990 630 20036
rect 1694 20603 1748 20649
rect 1878 20603 1932 20649
rect 2062 20603 2116 20649
rect 1694 19991 1748 20037
rect 1878 19991 1932 20037
rect 2062 19991 2116 20037
rect 4250 20602 4304 20648
rect 4434 20602 4488 20648
rect 4618 20602 4672 20648
rect 4250 19990 4304 20036
rect 4434 19990 4488 20036
rect 4618 19990 4672 20036
rect 5736 20603 5790 20649
rect 5920 20603 5974 20649
rect 6104 20603 6158 20649
rect 5736 19991 5790 20037
rect 5920 19991 5974 20037
rect 6104 19991 6158 20037
rect 8292 20602 8346 20648
rect 8476 20602 8530 20648
rect 8660 20602 8714 20648
rect 8292 19990 8346 20036
rect 8476 19990 8530 20036
rect 8660 19990 8714 20036
rect 9778 20603 9832 20649
rect 9962 20603 10016 20649
rect 10146 20603 10200 20649
rect 9778 19991 9832 20037
rect 9962 19991 10016 20037
rect 10146 19991 10200 20037
rect 12334 20602 12388 20648
rect 12518 20602 12572 20648
rect 12702 20602 12756 20648
rect 12334 19990 12388 20036
rect 12518 19990 12572 20036
rect 12702 19990 12756 20036
rect 13820 20603 13874 20649
rect 14004 20603 14058 20649
rect 14188 20603 14242 20649
rect 13820 19991 13874 20037
rect 14004 19991 14058 20037
rect 14188 19991 14242 20037
rect 16376 20602 16430 20648
rect 16560 20602 16614 20648
rect 16744 20602 16798 20648
rect 16376 19990 16430 20036
rect 16560 19990 16614 20036
rect 16744 19990 16798 20036
rect 17862 20603 17916 20649
rect 18046 20603 18100 20649
rect 18230 20603 18284 20649
rect 17862 19991 17916 20037
rect 18046 19991 18100 20037
rect 18230 19991 18284 20037
rect -7876 19445 -7822 19491
rect -7692 19445 -7638 19491
rect -7508 19445 -7454 19491
rect -7876 19133 -7822 19179
rect -7692 19133 -7638 19179
rect -7508 19133 -7454 19179
rect -6390 19446 -6336 19492
rect -6206 19446 -6152 19492
rect -6022 19446 -5968 19492
rect -6390 19134 -6336 19180
rect -6206 19134 -6152 19180
rect -6022 19134 -5968 19180
rect -3834 19442 -3780 19488
rect -3650 19442 -3596 19488
rect -3466 19442 -3412 19488
rect -3834 19130 -3780 19176
rect -3650 19130 -3596 19176
rect -3466 19130 -3412 19176
rect -2348 19443 -2294 19489
rect -2164 19443 -2110 19489
rect -1980 19443 -1926 19489
rect -2348 19131 -2294 19177
rect -2164 19131 -2110 19177
rect -1980 19131 -1926 19177
rect 208 19442 262 19488
rect 392 19442 446 19488
rect 576 19442 630 19488
rect 208 19130 262 19176
rect 392 19130 446 19176
rect 576 19130 630 19176
rect 1694 19443 1748 19489
rect 1878 19443 1932 19489
rect 2062 19443 2116 19489
rect 1694 19131 1748 19177
rect 1878 19131 1932 19177
rect 2062 19131 2116 19177
rect 4250 19442 4304 19488
rect 4434 19442 4488 19488
rect 4618 19442 4672 19488
rect 4250 19130 4304 19176
rect 4434 19130 4488 19176
rect 4618 19130 4672 19176
rect 5736 19443 5790 19489
rect 5920 19443 5974 19489
rect 6104 19443 6158 19489
rect 5736 19131 5790 19177
rect 5920 19131 5974 19177
rect 6104 19131 6158 19177
rect 8292 19442 8346 19488
rect 8476 19442 8530 19488
rect 8660 19442 8714 19488
rect 8292 19130 8346 19176
rect 8476 19130 8530 19176
rect 8660 19130 8714 19176
rect 9778 19443 9832 19489
rect 9962 19443 10016 19489
rect 10146 19443 10200 19489
rect 9778 19131 9832 19177
rect 9962 19131 10016 19177
rect 10146 19131 10200 19177
rect 12334 19442 12388 19488
rect 12518 19442 12572 19488
rect 12702 19442 12756 19488
rect 12334 19130 12388 19176
rect 12518 19130 12572 19176
rect 12702 19130 12756 19176
rect 13820 19443 13874 19489
rect 14004 19443 14058 19489
rect 14188 19443 14242 19489
rect 13820 19131 13874 19177
rect 14004 19131 14058 19177
rect 14188 19131 14242 19177
rect 16376 19442 16430 19488
rect 16560 19442 16614 19488
rect 16744 19442 16798 19488
rect 16376 19130 16430 19176
rect 16560 19130 16614 19176
rect 16744 19130 16798 19176
rect 17862 19443 17916 19489
rect 18046 19443 18100 19489
rect 18230 19443 18284 19489
rect 17862 19131 17916 19177
rect 18046 19131 18100 19177
rect 18230 19131 18284 19177
rect -7876 18400 -7822 18446
rect -7692 18400 -7638 18446
rect -7508 18400 -7454 18446
rect -7876 17788 -7822 17834
rect -7692 17788 -7638 17834
rect -7508 17788 -7454 17834
rect -3834 18397 -3780 18443
rect -3650 18397 -3596 18443
rect -3466 18397 -3412 18443
rect -3834 17785 -3780 17831
rect -3650 17785 -3596 17831
rect -3466 17785 -3412 17831
rect 208 18397 262 18443
rect 392 18397 446 18443
rect 576 18397 630 18443
rect 208 17785 262 17831
rect 392 17785 446 17831
rect 576 17785 630 17831
rect 4250 18397 4304 18443
rect 4434 18397 4488 18443
rect 4618 18397 4672 18443
rect 4250 17785 4304 17831
rect 4434 17785 4488 17831
rect 4618 17785 4672 17831
rect 8292 18397 8346 18443
rect 8476 18397 8530 18443
rect 8660 18397 8714 18443
rect 8292 17785 8346 17831
rect 8476 17785 8530 17831
rect 8660 17785 8714 17831
rect 12334 18397 12388 18443
rect 12518 18397 12572 18443
rect 12702 18397 12756 18443
rect 12334 17785 12388 17831
rect 12518 17785 12572 17831
rect 12702 17785 12756 17831
rect 16376 18397 16430 18443
rect 16560 18397 16614 18443
rect 16744 18397 16798 18443
rect 16376 17785 16430 17831
rect 16560 17785 16614 17831
rect 16744 17785 16798 17831
rect -7876 17240 -7822 17286
rect -7692 17240 -7638 17286
rect -7508 17240 -7454 17286
rect -7876 16928 -7822 16974
rect -7692 16928 -7638 16974
rect -7508 16928 -7454 16974
rect -3834 17237 -3780 17283
rect -3650 17237 -3596 17283
rect -3466 17237 -3412 17283
rect -3834 16925 -3780 16971
rect -3650 16925 -3596 16971
rect -3466 16925 -3412 16971
rect 208 17237 262 17283
rect 392 17237 446 17283
rect 576 17237 630 17283
rect 208 16925 262 16971
rect 392 16925 446 16971
rect 576 16925 630 16971
rect 4250 17237 4304 17283
rect 4434 17237 4488 17283
rect 4618 17237 4672 17283
rect 4250 16925 4304 16971
rect 4434 16925 4488 16971
rect 4618 16925 4672 16971
rect 8292 17237 8346 17283
rect 8476 17237 8530 17283
rect 8660 17237 8714 17283
rect 8292 16925 8346 16971
rect 8476 16925 8530 16971
rect 8660 16925 8714 16971
rect 12334 17237 12388 17283
rect 12518 17237 12572 17283
rect 12702 17237 12756 17283
rect 12334 16925 12388 16971
rect 12518 16925 12572 16971
rect 12702 16925 12756 16971
rect 16376 17237 16430 17283
rect 16560 17237 16614 17283
rect 16744 17237 16798 17283
rect 16376 16925 16430 16971
rect 16560 16925 16614 16971
rect 16744 16925 16798 16971
rect -11888 15436 -11834 15482
rect -11704 15436 -11650 15482
rect -11520 15436 -11466 15482
rect -11888 14824 -11834 14870
rect -11704 14824 -11650 14870
rect -11520 14824 -11466 14870
rect -7876 15436 -7822 15482
rect -7692 15436 -7638 15482
rect -7508 15436 -7454 15482
rect -7876 14824 -7822 14870
rect -7692 14824 -7638 14870
rect -7508 14824 -7454 14870
rect -3834 15436 -3780 15482
rect -3650 15436 -3596 15482
rect -3466 15436 -3412 15482
rect -3834 14824 -3780 14870
rect -3650 14824 -3596 14870
rect -3466 14824 -3412 14870
rect 208 15436 262 15482
rect 392 15436 446 15482
rect 576 15436 630 15482
rect 208 14824 262 14870
rect 392 14824 446 14870
rect 576 14824 630 14870
rect 4250 15436 4304 15482
rect 4434 15436 4488 15482
rect 4618 15436 4672 15482
rect 4250 14824 4304 14870
rect 4434 14824 4488 14870
rect 4618 14824 4672 14870
rect 8292 15436 8346 15482
rect 8476 15436 8530 15482
rect 8660 15436 8714 15482
rect 8292 14824 8346 14870
rect 8476 14824 8530 14870
rect 8660 14824 8714 14870
rect 12334 15436 12388 15482
rect 12518 15436 12572 15482
rect 12702 15436 12756 15482
rect 12334 14824 12388 14870
rect 12518 14824 12572 14870
rect 12702 14824 12756 14870
rect -11888 14276 -11834 14322
rect -11704 14276 -11650 14322
rect -11520 14276 -11466 14322
rect -11888 13964 -11834 14010
rect -11704 13964 -11650 14010
rect -11520 13964 -11466 14010
rect -7876 14276 -7822 14322
rect -7692 14276 -7638 14322
rect -7508 14276 -7454 14322
rect -7876 13964 -7822 14010
rect -7692 13964 -7638 14010
rect -7508 13964 -7454 14010
rect -3834 14276 -3780 14322
rect -3650 14276 -3596 14322
rect -3466 14276 -3412 14322
rect -3834 13964 -3780 14010
rect -3650 13964 -3596 14010
rect -3466 13964 -3412 14010
rect 208 14276 262 14322
rect 392 14276 446 14322
rect 576 14276 630 14322
rect 208 13964 262 14010
rect 392 13964 446 14010
rect 576 13964 630 14010
rect 4250 14276 4304 14322
rect 4434 14276 4488 14322
rect 4618 14276 4672 14322
rect 4250 13964 4304 14010
rect 4434 13964 4488 14010
rect 4618 13964 4672 14010
rect 8292 14276 8346 14322
rect 8476 14276 8530 14322
rect 8660 14276 8714 14322
rect 8292 13964 8346 14010
rect 8476 13964 8530 14010
rect 8660 13964 8714 14010
rect 12334 14276 12388 14322
rect 12518 14276 12572 14322
rect 12702 14276 12756 14322
rect 12334 13964 12388 14010
rect 12518 13964 12572 14010
rect 12702 13964 12756 14010
rect -11888 13231 -11834 13277
rect -11704 13231 -11650 13277
rect -11520 13231 -11466 13277
rect -11888 12619 -11834 12665
rect -11704 12619 -11650 12665
rect -11520 12619 -11466 12665
rect -10402 13231 -10348 13277
rect -10218 13231 -10164 13277
rect -10034 13231 -9980 13277
rect -10402 12619 -10348 12665
rect -10218 12619 -10164 12665
rect -10034 12619 -9980 12665
rect -7876 13231 -7822 13277
rect -7692 13231 -7638 13277
rect -7508 13231 -7454 13277
rect -7876 12619 -7822 12665
rect -7692 12619 -7638 12665
rect -7508 12619 -7454 12665
rect -6390 13231 -6336 13277
rect -6206 13231 -6152 13277
rect -6022 13231 -5968 13277
rect -6390 12619 -6336 12665
rect -6206 12619 -6152 12665
rect -6022 12619 -5968 12665
rect -3834 13231 -3780 13277
rect -3650 13231 -3596 13277
rect -3466 13231 -3412 13277
rect -3834 12619 -3780 12665
rect -3650 12619 -3596 12665
rect -3466 12619 -3412 12665
rect -2348 13231 -2294 13277
rect -2164 13231 -2110 13277
rect -1980 13231 -1926 13277
rect -2348 12619 -2294 12665
rect -2164 12619 -2110 12665
rect -1980 12619 -1926 12665
rect 208 13231 262 13277
rect 392 13231 446 13277
rect 576 13231 630 13277
rect 208 12619 262 12665
rect 392 12619 446 12665
rect 576 12619 630 12665
rect 1694 13231 1748 13277
rect 1878 13231 1932 13277
rect 2062 13231 2116 13277
rect 1694 12619 1748 12665
rect 1878 12619 1932 12665
rect 2062 12619 2116 12665
rect 4250 13231 4304 13277
rect 4434 13231 4488 13277
rect 4618 13231 4672 13277
rect 4250 12619 4304 12665
rect 4434 12619 4488 12665
rect 4618 12619 4672 12665
rect 5736 13231 5790 13277
rect 5920 13231 5974 13277
rect 6104 13231 6158 13277
rect 5736 12619 5790 12665
rect 5920 12619 5974 12665
rect 6104 12619 6158 12665
rect 8292 13231 8346 13277
rect 8476 13231 8530 13277
rect 8660 13231 8714 13277
rect 8292 12619 8346 12665
rect 8476 12619 8530 12665
rect 8660 12619 8714 12665
rect 9778 13231 9832 13277
rect 9962 13231 10016 13277
rect 10146 13231 10200 13277
rect 9778 12619 9832 12665
rect 9962 12619 10016 12665
rect 10146 12619 10200 12665
rect 12334 13231 12388 13277
rect 12518 13231 12572 13277
rect 12702 13231 12756 13277
rect 12334 12619 12388 12665
rect 12518 12619 12572 12665
rect 12702 12619 12756 12665
rect 13820 13231 13874 13277
rect 14004 13231 14058 13277
rect 14188 13231 14242 13277
rect 13820 12619 13874 12665
rect 14004 12619 14058 12665
rect 14188 12619 14242 12665
rect -11888 12071 -11834 12117
rect -11704 12071 -11650 12117
rect -11520 12071 -11466 12117
rect -11888 11759 -11834 11805
rect -11704 11759 -11650 11805
rect -11520 11759 -11466 11805
rect -10402 12071 -10348 12117
rect -10218 12071 -10164 12117
rect -10034 12071 -9980 12117
rect -10402 11759 -10348 11805
rect -10218 11759 -10164 11805
rect -10034 11759 -9980 11805
rect -7876 12071 -7822 12117
rect -7692 12071 -7638 12117
rect -7508 12071 -7454 12117
rect -7876 11759 -7822 11805
rect -7692 11759 -7638 11805
rect -7508 11759 -7454 11805
rect -6390 12071 -6336 12117
rect -6206 12071 -6152 12117
rect -6022 12071 -5968 12117
rect -6390 11759 -6336 11805
rect -6206 11759 -6152 11805
rect -6022 11759 -5968 11805
rect -3834 12071 -3780 12117
rect -3650 12071 -3596 12117
rect -3466 12071 -3412 12117
rect -3834 11759 -3780 11805
rect -3650 11759 -3596 11805
rect -3466 11759 -3412 11805
rect -2348 12071 -2294 12117
rect -2164 12071 -2110 12117
rect -1980 12071 -1926 12117
rect -2348 11759 -2294 11805
rect -2164 11759 -2110 11805
rect -1980 11759 -1926 11805
rect 208 12071 262 12117
rect 392 12071 446 12117
rect 576 12071 630 12117
rect 208 11759 262 11805
rect 392 11759 446 11805
rect 576 11759 630 11805
rect 1694 12071 1748 12117
rect 1878 12071 1932 12117
rect 2062 12071 2116 12117
rect 1694 11759 1748 11805
rect 1878 11759 1932 11805
rect 2062 11759 2116 11805
rect 4250 12071 4304 12117
rect 4434 12071 4488 12117
rect 4618 12071 4672 12117
rect 4250 11759 4304 11805
rect 4434 11759 4488 11805
rect 4618 11759 4672 11805
rect 5736 12071 5790 12117
rect 5920 12071 5974 12117
rect 6104 12071 6158 12117
rect 5736 11759 5790 11805
rect 5920 11759 5974 11805
rect 6104 11759 6158 11805
rect 8292 12071 8346 12117
rect 8476 12071 8530 12117
rect 8660 12071 8714 12117
rect 8292 11759 8346 11805
rect 8476 11759 8530 11805
rect 8660 11759 8714 11805
rect 9778 12071 9832 12117
rect 9962 12071 10016 12117
rect 10146 12071 10200 12117
rect 9778 11759 9832 11805
rect 9962 11759 10016 11805
rect 10146 11759 10200 11805
rect 12334 12071 12388 12117
rect 12518 12071 12572 12117
rect 12702 12071 12756 12117
rect 12334 11759 12388 11805
rect 12518 11759 12572 11805
rect 12702 11759 12756 11805
rect 13820 12071 13874 12117
rect 14004 12071 14058 12117
rect 14188 12071 14242 12117
rect 13820 11759 13874 11805
rect 14004 11759 14058 11805
rect 14188 11759 14242 11805
rect -11888 11026 -11834 11072
rect -11704 11026 -11650 11072
rect -11520 11026 -11466 11072
rect -11888 10414 -11834 10460
rect -11704 10414 -11650 10460
rect -11520 10414 -11466 10460
rect -10402 11027 -10348 11073
rect -10218 11027 -10164 11073
rect -10034 11027 -9980 11073
rect -10402 10415 -10348 10461
rect -10218 10415 -10164 10461
rect -10034 10415 -9980 10461
rect -7876 11026 -7822 11072
rect -7692 11026 -7638 11072
rect -7508 11026 -7454 11072
rect -7876 10414 -7822 10460
rect -7692 10414 -7638 10460
rect -7508 10414 -7454 10460
rect -6390 11027 -6336 11073
rect -6206 11027 -6152 11073
rect -6022 11027 -5968 11073
rect -6390 10415 -6336 10461
rect -6206 10415 -6152 10461
rect -6022 10415 -5968 10461
rect -3834 11026 -3780 11072
rect -3650 11026 -3596 11072
rect -3466 11026 -3412 11072
rect -3834 10414 -3780 10460
rect -3650 10414 -3596 10460
rect -3466 10414 -3412 10460
rect -2348 11027 -2294 11073
rect -2164 11027 -2110 11073
rect -1980 11027 -1926 11073
rect -2348 10415 -2294 10461
rect -2164 10415 -2110 10461
rect -1980 10415 -1926 10461
rect 208 11026 262 11072
rect 392 11026 446 11072
rect 576 11026 630 11072
rect 208 10414 262 10460
rect 392 10414 446 10460
rect 576 10414 630 10460
rect 1694 11027 1748 11073
rect 1878 11027 1932 11073
rect 2062 11027 2116 11073
rect 1694 10415 1748 10461
rect 1878 10415 1932 10461
rect 2062 10415 2116 10461
rect 4250 11026 4304 11072
rect 4434 11026 4488 11072
rect 4618 11026 4672 11072
rect 4250 10414 4304 10460
rect 4434 10414 4488 10460
rect 4618 10414 4672 10460
rect 5736 11027 5790 11073
rect 5920 11027 5974 11073
rect 6104 11027 6158 11073
rect 5736 10415 5790 10461
rect 5920 10415 5974 10461
rect 6104 10415 6158 10461
rect 8292 11026 8346 11072
rect 8476 11026 8530 11072
rect 8660 11026 8714 11072
rect 8292 10414 8346 10460
rect 8476 10414 8530 10460
rect 8660 10414 8714 10460
rect 9778 11027 9832 11073
rect 9962 11027 10016 11073
rect 10146 11027 10200 11073
rect 9778 10415 9832 10461
rect 9962 10415 10016 10461
rect 10146 10415 10200 10461
rect 12334 11026 12388 11072
rect 12518 11026 12572 11072
rect 12702 11026 12756 11072
rect 12334 10414 12388 10460
rect 12518 10414 12572 10460
rect 12702 10414 12756 10460
rect 13820 11027 13874 11073
rect 14004 11027 14058 11073
rect 14188 11027 14242 11073
rect 13820 10415 13874 10461
rect 14004 10415 14058 10461
rect 14188 10415 14242 10461
rect -11888 9866 -11834 9912
rect -11704 9866 -11650 9912
rect -11520 9866 -11466 9912
rect -11888 9554 -11834 9600
rect -11704 9554 -11650 9600
rect -11520 9554 -11466 9600
rect -10402 9867 -10348 9913
rect -10218 9867 -10164 9913
rect -10034 9867 -9980 9913
rect -10402 9555 -10348 9601
rect -10218 9555 -10164 9601
rect -10034 9555 -9980 9601
rect -7876 9866 -7822 9912
rect -7692 9866 -7638 9912
rect -7508 9866 -7454 9912
rect -7876 9554 -7822 9600
rect -7692 9554 -7638 9600
rect -7508 9554 -7454 9600
rect -6390 9867 -6336 9913
rect -6206 9867 -6152 9913
rect -6022 9867 -5968 9913
rect -6390 9555 -6336 9601
rect -6206 9555 -6152 9601
rect -6022 9555 -5968 9601
rect -3834 9866 -3780 9912
rect -3650 9866 -3596 9912
rect -3466 9866 -3412 9912
rect -3834 9554 -3780 9600
rect -3650 9554 -3596 9600
rect -3466 9554 -3412 9600
rect -2348 9867 -2294 9913
rect -2164 9867 -2110 9913
rect -1980 9867 -1926 9913
rect -2348 9555 -2294 9601
rect -2164 9555 -2110 9601
rect -1980 9555 -1926 9601
rect 208 9866 262 9912
rect 392 9866 446 9912
rect 576 9866 630 9912
rect 208 9554 262 9600
rect 392 9554 446 9600
rect 576 9554 630 9600
rect 1694 9867 1748 9913
rect 1878 9867 1932 9913
rect 2062 9867 2116 9913
rect 1694 9555 1748 9601
rect 1878 9555 1932 9601
rect 2062 9555 2116 9601
rect 4250 9866 4304 9912
rect 4434 9866 4488 9912
rect 4618 9866 4672 9912
rect 4250 9554 4304 9600
rect 4434 9554 4488 9600
rect 4618 9554 4672 9600
rect 5736 9867 5790 9913
rect 5920 9867 5974 9913
rect 6104 9867 6158 9913
rect 5736 9555 5790 9601
rect 5920 9555 5974 9601
rect 6104 9555 6158 9601
rect 8292 9866 8346 9912
rect 8476 9866 8530 9912
rect 8660 9866 8714 9912
rect 8292 9554 8346 9600
rect 8476 9554 8530 9600
rect 8660 9554 8714 9600
rect 9778 9867 9832 9913
rect 9962 9867 10016 9913
rect 10146 9867 10200 9913
rect 9778 9555 9832 9601
rect 9962 9555 10016 9601
rect 10146 9555 10200 9601
rect 12334 9866 12388 9912
rect 12518 9866 12572 9912
rect 12702 9866 12756 9912
rect 12334 9554 12388 9600
rect 12518 9554 12572 9600
rect 12702 9554 12756 9600
rect 13820 9867 13874 9913
rect 14004 9867 14058 9913
rect 14188 9867 14242 9913
rect 13820 9555 13874 9601
rect 14004 9555 14058 9601
rect 14188 9555 14242 9601
rect -11888 8821 -11834 8867
rect -11704 8821 -11650 8867
rect -11520 8821 -11466 8867
rect -11888 8209 -11834 8255
rect -11704 8209 -11650 8255
rect -11520 8209 -11466 8255
rect -7876 8821 -7822 8867
rect -7692 8821 -7638 8867
rect -7508 8821 -7454 8867
rect -7876 8209 -7822 8255
rect -7692 8209 -7638 8255
rect -7508 8209 -7454 8255
rect -3834 8821 -3780 8867
rect -3650 8821 -3596 8867
rect -3466 8821 -3412 8867
rect -3834 8209 -3780 8255
rect -3650 8209 -3596 8255
rect -3466 8209 -3412 8255
rect 208 8821 262 8867
rect 392 8821 446 8867
rect 576 8821 630 8867
rect 208 8209 262 8255
rect 392 8209 446 8255
rect 576 8209 630 8255
rect 4250 8821 4304 8867
rect 4434 8821 4488 8867
rect 4618 8821 4672 8867
rect 4250 8209 4304 8255
rect 4434 8209 4488 8255
rect 4618 8209 4672 8255
rect 8292 8821 8346 8867
rect 8476 8821 8530 8867
rect 8660 8821 8714 8867
rect 8292 8209 8346 8255
rect 8476 8209 8530 8255
rect 8660 8209 8714 8255
rect 12334 8821 12388 8867
rect 12518 8821 12572 8867
rect 12702 8821 12756 8867
rect 12334 8209 12388 8255
rect 12518 8209 12572 8255
rect 12702 8209 12756 8255
rect -11888 7661 -11834 7707
rect -11704 7661 -11650 7707
rect -11520 7661 -11466 7707
rect -11888 7349 -11834 7395
rect -11704 7349 -11650 7395
rect -11520 7349 -11466 7395
rect -7876 7661 -7822 7707
rect -7692 7661 -7638 7707
rect -7508 7661 -7454 7707
rect -7876 7349 -7822 7395
rect -7692 7349 -7638 7395
rect -7508 7349 -7454 7395
rect -3834 7661 -3780 7707
rect -3650 7661 -3596 7707
rect -3466 7661 -3412 7707
rect -3834 7349 -3780 7395
rect -3650 7349 -3596 7395
rect -3466 7349 -3412 7395
rect 208 7661 262 7707
rect 392 7661 446 7707
rect 576 7661 630 7707
rect 208 7349 262 7395
rect 392 7349 446 7395
rect 576 7349 630 7395
rect 4250 7661 4304 7707
rect 4434 7661 4488 7707
rect 4618 7661 4672 7707
rect 4250 7349 4304 7395
rect 4434 7349 4488 7395
rect 4618 7349 4672 7395
rect 8292 7661 8346 7707
rect 8476 7661 8530 7707
rect 8660 7661 8714 7707
rect 8292 7349 8346 7395
rect 8476 7349 8530 7395
rect 8660 7349 8714 7395
rect 12334 7661 12388 7707
rect 12518 7661 12572 7707
rect 12702 7661 12756 7707
rect 12334 7349 12388 7395
rect 12518 7349 12572 7395
rect 12702 7349 12756 7395
rect -10274 4777 -10228 4823
rect -10184 4627 -10138 4673
rect -8418 4900 -8364 4946
rect -8418 4588 -8364 4634
rect -7958 4900 -7904 4946
rect -7958 4588 -7904 4634
rect -9388 3483 -9334 3529
rect -8418 4080 -8364 4126
rect -8418 3768 -8364 3814
rect -7958 4080 -7904 4126
rect -7958 3768 -7904 3814
rect -6988 3483 -6934 3529
rect -9388 3147 -9334 3193
rect -6988 3147 -6934 3193
rect -10936 1710 -10882 1756
rect -10936 1438 -10882 1484
rect -10076 1710 -10022 1756
rect -10076 1438 -10022 1484
rect -9616 1730 -9442 1776
rect -9312 1730 -9138 1776
rect -9008 1730 -8834 1776
rect -8704 1730 -8530 1776
rect -8400 1730 -8226 1776
rect -8096 1730 -7922 1776
rect -7792 1730 -7618 1776
rect -7488 1730 -7314 1776
rect -7184 1730 -7010 1776
rect -6880 1730 -6706 1776
rect -9616 1418 -9442 1464
rect -9312 1418 -9138 1464
rect -9008 1418 -8834 1464
rect -8704 1418 -8530 1464
rect -8400 1418 -8226 1464
rect -8096 1418 -7922 1464
rect -7792 1418 -7618 1464
rect -7488 1418 -7314 1464
rect -7184 1418 -7010 1464
rect -6880 1418 -6706 1464
rect -6300 1710 -6246 1756
rect -6300 1438 -6246 1484
rect -5440 1710 -5386 1756
rect -5440 1438 -5386 1484
rect -9754 774 -9580 820
rect -9450 774 -9276 820
rect -9146 774 -8972 820
rect -8842 774 -8668 820
rect -8538 774 -8364 820
rect -9754 262 -9580 308
rect -9450 262 -9276 308
rect -9146 262 -8972 308
rect -8842 262 -8668 308
rect -8538 262 -8364 308
rect -7958 774 -7784 820
rect -7654 774 -7480 820
rect -7350 774 -7176 820
rect -7046 774 -6872 820
rect -6742 774 -6568 820
rect -7958 262 -7784 308
rect -7654 262 -7480 308
rect -7350 262 -7176 308
rect -7046 262 -6872 308
rect -6742 262 -6568 308
rect -9920 -711 -9746 -665
rect -9616 -711 -9442 -665
rect -9312 -711 -9138 -665
rect -9008 -711 -8834 -665
rect -8704 -711 -8530 -665
rect -8400 -711 -8226 -665
rect -8096 -711 -7922 -665
rect -7792 -711 -7618 -665
rect -7488 -711 -7314 -665
rect -7184 -711 -7010 -665
rect -6880 -711 -6706 -665
rect -6576 -711 -6402 -665
rect -9920 -1123 -9746 -1077
rect -9616 -1123 -9442 -1077
rect -9312 -1123 -9138 -1077
rect -9008 -1123 -8834 -1077
rect -8704 -1123 -8530 -1077
rect -8400 -1123 -8226 -1077
rect -8096 -1123 -7922 -1077
rect -7792 -1123 -7618 -1077
rect -7488 -1123 -7314 -1077
rect -7184 -1123 -7010 -1077
rect -6880 -1123 -6706 -1077
rect -6576 -1123 -6402 -1077
rect -9920 -1674 -9746 -1628
rect -9616 -1674 -9442 -1628
rect -9312 -1674 -9138 -1628
rect -9008 -1674 -8834 -1628
rect -8704 -1674 -8530 -1628
rect -8400 -1674 -8226 -1628
rect -8096 -1674 -7922 -1628
rect -7792 -1674 -7618 -1628
rect -7488 -1674 -7314 -1628
rect -7184 -1674 -7010 -1628
rect -6880 -1674 -6706 -1628
rect -6576 -1674 -6402 -1628
rect -9920 -2086 -9746 -2040
rect -9616 -2086 -9442 -2040
rect -9312 -2086 -9138 -2040
rect -9008 -2086 -8834 -2040
rect -8704 -2086 -8530 -2040
rect -8400 -2086 -8226 -2040
rect -8096 -2086 -7922 -2040
rect -7792 -2086 -7618 -2040
rect -7488 -2086 -7314 -2040
rect -7184 -2086 -7010 -2040
rect -6880 -2086 -6706 -2040
rect -6576 -2086 -6402 -2040
rect -8372 -2600 -8318 -2554
rect -8188 -2600 -8134 -2554
rect -8004 -2600 -7950 -2554
rect -8372 -2872 -8318 -2826
rect -8188 -2872 -8134 -2826
rect -8004 -2872 -7950 -2826
<< metal1 >>
rect 40726 39167 40972 39180
rect 40726 39093 40739 39167
rect 40957 39093 40972 39167
rect 39851 39021 40991 39093
rect 39851 38975 40103 39021
rect 40149 38975 40343 39021
rect 40389 38975 40583 39021
rect 40629 38975 40823 39021
rect 40869 38975 40991 39021
rect 39851 38953 40991 38975
rect 39971 38830 40021 38953
rect 39971 38596 39973 38830
rect 40019 38596 40021 38830
rect 40141 38855 40191 38883
rect 40141 38621 40143 38855
rect 40189 38621 40191 38855
rect 40141 38603 40191 38621
rect 40311 38830 40361 38953
rect 39971 38543 40021 38596
rect 40111 38599 40211 38603
rect 40111 38547 40135 38599
rect 40187 38547 40211 38599
rect 40111 38543 40211 38547
rect 40311 38596 40313 38830
rect 40359 38596 40361 38830
rect 40311 38543 40361 38596
rect 40481 38855 40531 38883
rect 40481 38621 40483 38855
rect 40529 38621 40531 38855
rect 40141 38493 40191 38543
rect 40481 38493 40531 38621
rect 40651 38830 40701 38953
rect 40651 38596 40653 38830
rect 40699 38596 40701 38830
rect 40651 38543 40701 38596
rect 40821 38830 40871 38883
rect 40821 38596 40823 38830
rect 40869 38596 40871 38830
rect 40821 38493 40871 38596
rect 40141 38433 40531 38493
rect 40581 38486 40871 38493
rect 40581 38440 40608 38486
rect 40654 38440 40871 38486
rect 40581 38433 40871 38440
rect 40141 38313 40191 38433
rect 40481 38313 40531 38433
rect 40141 38253 40531 38313
rect 40671 38339 40771 38343
rect 40671 38287 40695 38339
rect 40747 38287 40771 38339
rect 40671 38283 40771 38287
rect 39971 38141 40021 38203
rect 39971 38095 39973 38141
rect 40019 38095 40021 38141
rect 39971 37963 40021 38095
rect 40141 38141 40191 38253
rect 40141 38095 40143 38141
rect 40189 38095 40191 38141
rect 40141 38033 40191 38095
rect 40311 38141 40361 38203
rect 40311 38095 40313 38141
rect 40359 38095 40361 38141
rect 40311 37963 40361 38095
rect 40481 38141 40531 38253
rect 40481 38095 40483 38141
rect 40529 38095 40531 38141
rect 40481 38033 40531 38095
rect 40651 38141 40701 38203
rect 40651 38095 40653 38141
rect 40699 38095 40701 38141
rect 40651 37963 40701 38095
rect 40821 38141 40871 38433
rect 40821 38095 40823 38141
rect 40869 38095 40871 38141
rect 40821 38033 40871 38095
rect 39851 37941 40991 37963
rect 39851 37895 40103 37941
rect 40149 37895 40343 37941
rect 40389 37895 40583 37941
rect 40629 37895 40823 37941
rect 40869 37895 40991 37941
rect 39851 37823 40991 37895
rect 40723 37749 40737 37823
rect 40955 37749 40967 37823
rect 40723 37737 40967 37749
rect -5024 37619 -3477 37675
rect -5521 36598 -5433 36610
rect -5024 36598 -4968 37619
rect -4355 37567 -4269 37571
rect -4355 37511 -4343 37567
rect -4287 37511 -4269 37567
rect -4355 37499 -4269 37511
rect -4844 37354 -4798 37365
rect -4629 37363 -4553 37396
rect -4629 37317 -4618 37363
rect -4564 37317 -4553 37363
rect -4445 37363 -4369 37396
rect -4445 37317 -4434 37363
rect -4380 37317 -4369 37363
rect -4261 37363 -4185 37396
rect -4261 37317 -4250 37363
rect -4196 37317 -4185 37363
rect -4016 37354 -3970 37365
rect -4706 37271 -4660 37282
rect -4723 37244 -4706 37246
rect -4522 37271 -4476 37282
rect -4660 37244 -4643 37246
rect -4798 37124 -4711 37244
rect -4655 37124 -4643 37244
rect -4723 37122 -4706 37124
rect -4798 36824 -4706 36944
rect -4660 37122 -4643 37124
rect -4539 36944 -4522 36946
rect -4338 37271 -4292 37282
rect -4355 37244 -4338 37246
rect -4154 37271 -4108 37282
rect -4292 37244 -4275 37246
rect -4355 37124 -4343 37244
rect -4287 37124 -4275 37244
rect -4355 37122 -4338 37124
rect -4476 36944 -4459 36946
rect -4539 36824 -4527 36944
rect -4471 36824 -4459 36944
rect -4539 36822 -4522 36824
rect -4706 36786 -4660 36797
rect -4476 36822 -4459 36824
rect -4522 36786 -4476 36797
rect -4292 37122 -4275 37124
rect -4171 36944 -4154 36946
rect -4033 37244 -4016 37246
rect -3970 37244 -3953 37246
rect -4033 37123 -4021 37244
rect -3965 37123 -3953 37244
rect -4033 37121 -4016 37123
rect -4108 36944 -4091 36946
rect -4171 36824 -4159 36944
rect -4103 36824 -4091 36944
rect -4171 36822 -4154 36824
rect -4338 36786 -4292 36797
rect -4108 36822 -4091 36824
rect -4154 36786 -4108 36797
rect -4629 36748 -4618 36751
rect -4564 36748 -4553 36751
rect -4445 36748 -4434 36751
rect -4380 36748 -4369 36751
rect -4261 36748 -4250 36751
rect -4196 36748 -4185 36751
rect -4844 36703 -4798 36714
rect -4631 36692 -4619 36748
rect -4563 36692 -4551 36748
rect -4631 36678 -4551 36692
rect -4447 36692 -4435 36748
rect -4379 36692 -4367 36748
rect -4447 36678 -4367 36692
rect -4263 36692 -4251 36748
rect -4195 36692 -4183 36748
rect -3970 37121 -3953 37123
rect -4016 36703 -3970 36714
rect -4263 36678 -4183 36692
rect -4631 36598 -4551 36600
rect -5521 36542 -5507 36598
rect -5451 36542 -4619 36598
rect -4563 36542 -4551 36598
rect -5521 36530 -5433 36542
rect -4631 36540 -4551 36542
rect -5303 36482 -5233 36494
rect -4447 36482 -4367 36484
rect -5303 36426 -5291 36482
rect -5235 36426 -4435 36482
rect -4379 36426 -4367 36482
rect -5303 36414 -5233 36426
rect -4447 36424 -4367 36426
rect -4118 36482 -4038 36484
rect -3851 36482 -3781 36494
rect -4118 36426 -4106 36482
rect -4050 36426 -3849 36482
rect -3793 36426 -3781 36482
rect -4118 36424 -4038 36426
rect -3851 36416 -3781 36426
rect -4263 36366 -4183 36368
rect -5019 36310 -4251 36366
rect -4195 36310 -4183 36366
rect -5019 35579 -4963 36310
rect -4263 36308 -4183 36310
rect -4631 36216 -4551 36230
rect -4844 36194 -4798 36205
rect -4631 36160 -4619 36216
rect -4563 36160 -4551 36216
rect -4447 36216 -4367 36230
rect -4447 36160 -4435 36216
rect -4379 36160 -4367 36216
rect -4263 36216 -4183 36230
rect -4263 36160 -4251 36216
rect -4195 36160 -4183 36216
rect -4016 36194 -3970 36205
rect -4629 36157 -4618 36160
rect -4564 36157 -4553 36160
rect -4445 36157 -4434 36160
rect -4380 36157 -4369 36160
rect -4261 36157 -4250 36160
rect -4196 36157 -4185 36160
rect -4706 36111 -4660 36122
rect -4798 35937 -4706 36111
rect -4706 35926 -4660 35937
rect -4522 36111 -4476 36122
rect -4522 35926 -4476 35937
rect -4338 36111 -4292 36122
rect -4154 36111 -4108 36122
rect -4171 36084 -4154 36086
rect -4108 36084 -4091 36086
rect -4171 35964 -4159 36084
rect -4103 35964 -4091 36084
rect -4171 35962 -4154 35964
rect -4338 35926 -4292 35937
rect -4108 35962 -4091 35964
rect -4154 35926 -4108 35937
rect -4844 35709 -4798 35854
rect -4629 35845 -4618 35891
rect -4564 35845 -4553 35891
rect -4629 35812 -4553 35845
rect -4445 35845 -4434 35891
rect -4380 35845 -4369 35891
rect -4445 35812 -4369 35845
rect -4261 35845 -4250 35891
rect -4196 35845 -4185 35891
rect -4261 35812 -4185 35845
rect -4016 35709 -3970 35854
rect -4856 35697 -4776 35709
rect -4856 35641 -4844 35697
rect -4788 35641 -4776 35697
rect -4856 35629 -4776 35641
rect -4038 35697 -3958 35709
rect -4038 35641 -4026 35697
rect -3970 35641 -3958 35697
rect -4038 35629 -3958 35641
rect -3685 35579 -3605 35589
rect -5019 35523 -3673 35579
rect -3617 35523 -3605 35579
rect -3685 35521 -3605 35523
rect -3851 35470 -3781 35472
rect -5019 35469 -3781 35470
rect -5019 35415 -3849 35469
rect -3793 35415 -3781 35469
rect -5019 35414 -3781 35415
rect -5019 34393 -4963 35414
rect -3851 35406 -3781 35414
rect -4355 35362 -4269 35366
rect -4355 35306 -4343 35362
rect -4287 35306 -4269 35362
rect -4355 35294 -4269 35306
rect -4844 35149 -4798 35160
rect -4629 35158 -4553 35191
rect -4629 35112 -4618 35158
rect -4564 35112 -4553 35158
rect -4445 35158 -4369 35191
rect -4445 35112 -4434 35158
rect -4380 35112 -4369 35158
rect -4261 35158 -4185 35191
rect -4261 35112 -4250 35158
rect -4196 35112 -4185 35158
rect -4016 35149 -3970 35160
rect -4706 35066 -4660 35077
rect -4723 35039 -4706 35041
rect -4522 35066 -4476 35077
rect -4660 35039 -4643 35041
rect -4798 34919 -4711 35039
rect -4655 34919 -4643 35039
rect -4723 34917 -4706 34919
rect -4798 34619 -4706 34739
rect -4660 34917 -4643 34919
rect -4539 34739 -4522 34741
rect -4338 35066 -4292 35077
rect -4355 35039 -4338 35041
rect -4154 35066 -4108 35077
rect -4292 35039 -4275 35041
rect -4355 34919 -4343 35039
rect -4287 34919 -4275 35039
rect -4355 34917 -4338 34919
rect -4476 34739 -4459 34741
rect -4539 34619 -4527 34739
rect -4471 34619 -4459 34739
rect -4539 34617 -4522 34619
rect -4706 34581 -4660 34592
rect -4476 34617 -4459 34619
rect -4522 34581 -4476 34592
rect -4292 34917 -4275 34919
rect -4171 34739 -4154 34741
rect -4033 35039 -4016 35041
rect -3970 35039 -3953 35041
rect -4033 34918 -4021 35039
rect -3965 34918 -3953 35039
rect -4033 34916 -4016 34918
rect -4108 34739 -4091 34741
rect -4171 34619 -4159 34739
rect -4103 34619 -4091 34739
rect -4171 34617 -4154 34619
rect -4338 34581 -4292 34592
rect -4108 34617 -4091 34619
rect -4154 34581 -4108 34592
rect -4629 34543 -4618 34546
rect -4564 34543 -4553 34546
rect -4445 34543 -4434 34546
rect -4380 34543 -4369 34546
rect -4261 34543 -4250 34546
rect -4196 34543 -4185 34546
rect -4844 34498 -4798 34509
rect -4631 34487 -4619 34543
rect -4563 34487 -4551 34543
rect -4631 34473 -4551 34487
rect -4447 34487 -4435 34543
rect -4379 34487 -4367 34543
rect -4447 34473 -4367 34487
rect -4263 34487 -4251 34543
rect -4195 34487 -4183 34543
rect -3970 34916 -3953 34918
rect -4016 34498 -3970 34509
rect -4263 34473 -4183 34487
rect -4631 34393 -4551 34395
rect -5019 34337 -4619 34393
rect -4563 34337 -4551 34393
rect -3533 34393 -3477 37619
rect 4448 37619 5995 37675
rect 3951 36598 4039 36610
rect 4448 36598 4504 37619
rect 5117 37567 5203 37571
rect 5117 37511 5129 37567
rect 5185 37511 5203 37567
rect 5117 37499 5203 37511
rect 4628 37354 4674 37365
rect 4843 37363 4919 37396
rect 4843 37317 4854 37363
rect 4908 37317 4919 37363
rect 5027 37363 5103 37396
rect 5027 37317 5038 37363
rect 5092 37317 5103 37363
rect 5211 37363 5287 37396
rect 5211 37317 5222 37363
rect 5276 37317 5287 37363
rect 5456 37354 5502 37365
rect 4766 37271 4812 37282
rect 4749 37244 4766 37246
rect 4950 37271 4996 37282
rect 4812 37244 4829 37246
rect 4674 37124 4761 37244
rect 4817 37124 4829 37244
rect 4749 37122 4766 37124
rect 4674 36824 4766 36944
rect 4812 37122 4829 37124
rect 4933 36944 4950 36946
rect 5134 37271 5180 37282
rect 5117 37244 5134 37246
rect 5318 37271 5364 37282
rect 5180 37244 5197 37246
rect 5117 37124 5129 37244
rect 5185 37124 5197 37244
rect 5117 37122 5134 37124
rect 4996 36944 5013 36946
rect 4933 36824 4945 36944
rect 5001 36824 5013 36944
rect 4933 36822 4950 36824
rect 4766 36786 4812 36797
rect 4996 36822 5013 36824
rect 4950 36786 4996 36797
rect 5180 37122 5197 37124
rect 5301 36944 5318 36946
rect 5439 37244 5456 37246
rect 5502 37244 5519 37246
rect 5439 37123 5451 37244
rect 5507 37123 5519 37244
rect 5439 37121 5456 37123
rect 5364 36944 5381 36946
rect 5301 36824 5313 36944
rect 5369 36824 5381 36944
rect 5301 36822 5318 36824
rect 5134 36786 5180 36797
rect 5364 36822 5381 36824
rect 5318 36786 5364 36797
rect 4843 36748 4854 36751
rect 4908 36748 4919 36751
rect 5027 36748 5038 36751
rect 5092 36748 5103 36751
rect 5211 36748 5222 36751
rect 5276 36748 5287 36751
rect 4628 36703 4674 36714
rect 4841 36692 4853 36748
rect 4909 36692 4921 36748
rect 4841 36678 4921 36692
rect 5025 36692 5037 36748
rect 5093 36692 5105 36748
rect 5025 36678 5105 36692
rect 5209 36692 5221 36748
rect 5277 36692 5289 36748
rect 5502 37121 5519 37123
rect 5456 36703 5502 36714
rect 5209 36678 5289 36692
rect 4841 36598 4921 36600
rect 3951 36542 3965 36598
rect 4021 36542 4853 36598
rect 4909 36542 4921 36598
rect 3951 36530 4039 36542
rect 4841 36540 4921 36542
rect 4169 36482 4239 36494
rect 5025 36482 5105 36484
rect 4169 36426 4181 36482
rect 4237 36426 5037 36482
rect 5093 36426 5105 36482
rect 4169 36414 4239 36426
rect 5025 36424 5105 36426
rect 5354 36482 5434 36484
rect 5621 36482 5691 36494
rect 5354 36426 5366 36482
rect 5422 36426 5623 36482
rect 5679 36426 5691 36482
rect 5354 36424 5434 36426
rect 5621 36416 5691 36426
rect 5209 36366 5289 36368
rect 4453 36310 5221 36366
rect 5277 36310 5289 36366
rect 4453 35579 4509 36310
rect 5209 36308 5289 36310
rect 4841 36216 4921 36230
rect 4628 36194 4674 36205
rect 4841 36160 4853 36216
rect 4909 36160 4921 36216
rect 5025 36216 5105 36230
rect 5025 36160 5037 36216
rect 5093 36160 5105 36216
rect 5209 36216 5289 36230
rect 5209 36160 5221 36216
rect 5277 36160 5289 36216
rect 5456 36194 5502 36205
rect 4843 36157 4854 36160
rect 4908 36157 4919 36160
rect 5027 36157 5038 36160
rect 5092 36157 5103 36160
rect 5211 36157 5222 36160
rect 5276 36157 5287 36160
rect 4766 36111 4812 36122
rect 4674 35937 4766 36111
rect 4766 35926 4812 35937
rect 4950 36111 4996 36122
rect 4950 35926 4996 35937
rect 5134 36111 5180 36122
rect 5318 36111 5364 36122
rect 5301 36084 5318 36086
rect 5364 36084 5381 36086
rect 5301 35964 5313 36084
rect 5369 35964 5381 36084
rect 5301 35962 5318 35964
rect 5134 35926 5180 35937
rect 5364 35962 5381 35964
rect 5318 35926 5364 35937
rect 4628 35709 4674 35854
rect 4843 35845 4854 35891
rect 4908 35845 4919 35891
rect 4843 35812 4919 35845
rect 5027 35845 5038 35891
rect 5092 35845 5103 35891
rect 5027 35812 5103 35845
rect 5211 35845 5222 35891
rect 5276 35845 5287 35891
rect 5211 35812 5287 35845
rect 5456 35709 5502 35854
rect 4616 35697 4696 35709
rect 4616 35641 4628 35697
rect 4684 35641 4696 35697
rect 4616 35629 4696 35641
rect 5434 35697 5514 35709
rect 5434 35641 5446 35697
rect 5502 35641 5514 35697
rect 5434 35629 5514 35641
rect 5787 35579 5867 35589
rect 4453 35523 5799 35579
rect 5855 35523 5867 35579
rect 5787 35521 5867 35523
rect 5621 35470 5691 35472
rect 4453 35469 5691 35470
rect 4453 35415 5623 35469
rect 5679 35415 5691 35469
rect 4453 35414 5691 35415
rect -2869 35362 -2783 35366
rect -2869 35306 -2857 35362
rect -2801 35306 -2783 35362
rect -2869 35294 -2783 35306
rect -3358 35149 -3312 35160
rect -3143 35158 -3067 35191
rect -3143 35112 -3132 35158
rect -3078 35112 -3067 35158
rect -2959 35158 -2883 35191
rect -2959 35112 -2948 35158
rect -2894 35112 -2883 35158
rect -2775 35158 -2699 35191
rect -2775 35112 -2764 35158
rect -2710 35112 -2699 35158
rect -2530 35149 -2484 35160
rect -3220 35066 -3174 35077
rect -3237 35039 -3220 35041
rect -3036 35066 -2990 35077
rect -3174 35039 -3157 35041
rect -3312 34919 -3225 35039
rect -3169 34919 -3157 35039
rect -3237 34917 -3220 34919
rect -3312 34619 -3220 34739
rect -3174 34917 -3157 34919
rect -3053 34739 -3036 34741
rect -2852 35066 -2806 35077
rect -2869 35039 -2852 35041
rect -2668 35066 -2622 35077
rect -2806 35039 -2789 35041
rect -2869 34919 -2857 35039
rect -2801 34919 -2789 35039
rect -2869 34917 -2852 34919
rect -2990 34739 -2973 34741
rect -3053 34619 -3041 34739
rect -2985 34619 -2973 34739
rect -3053 34617 -3036 34619
rect -3220 34581 -3174 34592
rect -2990 34617 -2973 34619
rect -3036 34581 -2990 34592
rect -2806 34917 -2789 34919
rect -2685 34739 -2668 34741
rect -2547 35039 -2530 35041
rect -2484 35039 -2467 35041
rect -2547 34918 -2535 35039
rect -2479 34918 -2467 35039
rect -2547 34916 -2530 34918
rect -2622 34739 -2605 34741
rect -2685 34619 -2673 34739
rect -2617 34619 -2605 34739
rect -2685 34617 -2668 34619
rect -2852 34581 -2806 34592
rect -2622 34617 -2605 34619
rect -2668 34581 -2622 34592
rect -3143 34543 -3132 34546
rect -3078 34543 -3067 34546
rect -2959 34543 -2948 34546
rect -2894 34543 -2883 34546
rect -2775 34543 -2764 34546
rect -2710 34543 -2699 34546
rect -3358 34498 -3312 34509
rect -3145 34487 -3133 34543
rect -3077 34487 -3065 34543
rect -3145 34473 -3065 34487
rect -2961 34487 -2949 34543
rect -2893 34487 -2881 34543
rect -2961 34473 -2881 34487
rect -2777 34487 -2765 34543
rect -2709 34487 -2697 34543
rect -2484 34916 -2467 34918
rect -2530 34498 -2484 34509
rect -2777 34473 -2697 34487
rect -3145 34393 -3065 34395
rect -3533 34337 -3133 34393
rect -3077 34337 -3065 34393
rect 4453 34393 4509 35414
rect 5621 35406 5691 35414
rect 5117 35362 5203 35366
rect 5117 35306 5129 35362
rect 5185 35306 5203 35362
rect 5117 35294 5203 35306
rect 4628 35149 4674 35160
rect 4843 35158 4919 35191
rect 4843 35112 4854 35158
rect 4908 35112 4919 35158
rect 5027 35158 5103 35191
rect 5027 35112 5038 35158
rect 5092 35112 5103 35158
rect 5211 35158 5287 35191
rect 5211 35112 5222 35158
rect 5276 35112 5287 35158
rect 5456 35149 5502 35160
rect 4766 35066 4812 35077
rect 4749 35039 4766 35041
rect 4950 35066 4996 35077
rect 4812 35039 4829 35041
rect 4674 34919 4761 35039
rect 4817 34919 4829 35039
rect 4749 34917 4766 34919
rect 4674 34619 4766 34739
rect 4812 34917 4829 34919
rect 4933 34739 4950 34741
rect 5134 35066 5180 35077
rect 5117 35039 5134 35041
rect 5318 35066 5364 35077
rect 5180 35039 5197 35041
rect 5117 34919 5129 35039
rect 5185 34919 5197 35039
rect 5117 34917 5134 34919
rect 4996 34739 5013 34741
rect 4933 34619 4945 34739
rect 5001 34619 5013 34739
rect 4933 34617 4950 34619
rect 4766 34581 4812 34592
rect 4996 34617 5013 34619
rect 4950 34581 4996 34592
rect 5180 34917 5197 34919
rect 5301 34739 5318 34741
rect 5439 35039 5456 35041
rect 5502 35039 5519 35041
rect 5439 34918 5451 35039
rect 5507 34918 5519 35039
rect 5439 34916 5456 34918
rect 5364 34739 5381 34741
rect 5301 34619 5313 34739
rect 5369 34619 5381 34739
rect 5301 34617 5318 34619
rect 5134 34581 5180 34592
rect 5364 34617 5381 34619
rect 5318 34581 5364 34592
rect 4843 34543 4854 34546
rect 4908 34543 4919 34546
rect 5027 34543 5038 34546
rect 5092 34543 5103 34546
rect 5211 34543 5222 34546
rect 5276 34543 5287 34546
rect 4628 34498 4674 34509
rect 4841 34487 4853 34543
rect 4909 34487 4921 34543
rect 4841 34473 4921 34487
rect 5025 34487 5037 34543
rect 5093 34487 5105 34543
rect 5025 34473 5105 34487
rect 5209 34487 5221 34543
rect 5277 34487 5289 34543
rect 5502 34916 5519 34918
rect 5456 34498 5502 34509
rect 5209 34473 5289 34487
rect 4841 34393 4921 34395
rect 4453 34337 4853 34393
rect 4909 34337 4921 34393
rect 5939 34393 5995 37619
rect 13920 37620 15467 37676
rect 13423 36599 13511 36611
rect 13920 36599 13976 37620
rect 14589 37568 14675 37572
rect 14589 37512 14601 37568
rect 14657 37512 14675 37568
rect 14589 37500 14675 37512
rect 14100 37355 14146 37366
rect 14315 37364 14391 37397
rect 14315 37318 14326 37364
rect 14380 37318 14391 37364
rect 14499 37364 14575 37397
rect 14499 37318 14510 37364
rect 14564 37318 14575 37364
rect 14683 37364 14759 37397
rect 14683 37318 14694 37364
rect 14748 37318 14759 37364
rect 14928 37355 14974 37366
rect 14238 37272 14284 37283
rect 14221 37245 14238 37247
rect 14422 37272 14468 37283
rect 14284 37245 14301 37247
rect 14146 37125 14233 37245
rect 14289 37125 14301 37245
rect 14221 37123 14238 37125
rect 14146 36825 14238 36945
rect 14284 37123 14301 37125
rect 14405 36945 14422 36947
rect 14606 37272 14652 37283
rect 14589 37245 14606 37247
rect 14790 37272 14836 37283
rect 14652 37245 14669 37247
rect 14589 37125 14601 37245
rect 14657 37125 14669 37245
rect 14589 37123 14606 37125
rect 14468 36945 14485 36947
rect 14405 36825 14417 36945
rect 14473 36825 14485 36945
rect 14405 36823 14422 36825
rect 14238 36787 14284 36798
rect 14468 36823 14485 36825
rect 14422 36787 14468 36798
rect 14652 37123 14669 37125
rect 14773 36945 14790 36947
rect 14911 37245 14928 37247
rect 14974 37245 14991 37247
rect 14911 37124 14923 37245
rect 14979 37124 14991 37245
rect 14911 37122 14928 37124
rect 14836 36945 14853 36947
rect 14773 36825 14785 36945
rect 14841 36825 14853 36945
rect 14773 36823 14790 36825
rect 14606 36787 14652 36798
rect 14836 36823 14853 36825
rect 14790 36787 14836 36798
rect 14315 36749 14326 36752
rect 14380 36749 14391 36752
rect 14499 36749 14510 36752
rect 14564 36749 14575 36752
rect 14683 36749 14694 36752
rect 14748 36749 14759 36752
rect 14100 36704 14146 36715
rect 14313 36693 14325 36749
rect 14381 36693 14393 36749
rect 14313 36679 14393 36693
rect 14497 36693 14509 36749
rect 14565 36693 14577 36749
rect 14497 36679 14577 36693
rect 14681 36693 14693 36749
rect 14749 36693 14761 36749
rect 14974 37122 14991 37124
rect 14928 36704 14974 36715
rect 14681 36679 14761 36693
rect 14313 36599 14393 36601
rect 13423 36543 13437 36599
rect 13493 36543 14325 36599
rect 14381 36543 14393 36599
rect 13423 36531 13511 36543
rect 14313 36541 14393 36543
rect 13641 36483 13711 36495
rect 14497 36483 14577 36485
rect 13641 36427 13653 36483
rect 13709 36427 14509 36483
rect 14565 36427 14577 36483
rect 13641 36415 13711 36427
rect 14497 36425 14577 36427
rect 14826 36483 14906 36485
rect 15093 36483 15163 36495
rect 14826 36427 14838 36483
rect 14894 36427 15095 36483
rect 15151 36427 15163 36483
rect 14826 36425 14906 36427
rect 15093 36417 15163 36427
rect 14681 36367 14761 36369
rect 13925 36311 14693 36367
rect 14749 36311 14761 36367
rect 13925 35580 13981 36311
rect 14681 36309 14761 36311
rect 14313 36217 14393 36231
rect 14100 36195 14146 36206
rect 14313 36161 14325 36217
rect 14381 36161 14393 36217
rect 14497 36217 14577 36231
rect 14497 36161 14509 36217
rect 14565 36161 14577 36217
rect 14681 36217 14761 36231
rect 14681 36161 14693 36217
rect 14749 36161 14761 36217
rect 14928 36195 14974 36206
rect 14315 36158 14326 36161
rect 14380 36158 14391 36161
rect 14499 36158 14510 36161
rect 14564 36158 14575 36161
rect 14683 36158 14694 36161
rect 14748 36158 14759 36161
rect 14238 36112 14284 36123
rect 14146 35938 14238 36112
rect 14238 35927 14284 35938
rect 14422 36112 14468 36123
rect 14422 35927 14468 35938
rect 14606 36112 14652 36123
rect 14790 36112 14836 36123
rect 14773 36085 14790 36087
rect 14836 36085 14853 36087
rect 14773 35965 14785 36085
rect 14841 35965 14853 36085
rect 14773 35963 14790 35965
rect 14606 35927 14652 35938
rect 14836 35963 14853 35965
rect 14790 35927 14836 35938
rect 14100 35710 14146 35855
rect 14315 35846 14326 35892
rect 14380 35846 14391 35892
rect 14315 35813 14391 35846
rect 14499 35846 14510 35892
rect 14564 35846 14575 35892
rect 14499 35813 14575 35846
rect 14683 35846 14694 35892
rect 14748 35846 14759 35892
rect 14683 35813 14759 35846
rect 14928 35710 14974 35855
rect 14088 35698 14168 35710
rect 14088 35642 14100 35698
rect 14156 35642 14168 35698
rect 14088 35630 14168 35642
rect 14906 35698 14986 35710
rect 14906 35642 14918 35698
rect 14974 35642 14986 35698
rect 14906 35630 14986 35642
rect 15259 35580 15339 35590
rect 13925 35524 15271 35580
rect 15327 35524 15339 35580
rect 15259 35522 15339 35524
rect 15093 35471 15163 35473
rect 13925 35470 15163 35471
rect 13925 35416 15095 35470
rect 15151 35416 15163 35470
rect 13925 35415 15163 35416
rect 6603 35362 6689 35366
rect 6603 35306 6615 35362
rect 6671 35306 6689 35362
rect 6603 35294 6689 35306
rect 6114 35149 6160 35160
rect 6329 35158 6405 35191
rect 6329 35112 6340 35158
rect 6394 35112 6405 35158
rect 6513 35158 6589 35191
rect 6513 35112 6524 35158
rect 6578 35112 6589 35158
rect 6697 35158 6773 35191
rect 6697 35112 6708 35158
rect 6762 35112 6773 35158
rect 6942 35149 6988 35160
rect 6252 35066 6298 35077
rect 6235 35039 6252 35041
rect 6436 35066 6482 35077
rect 6298 35039 6315 35041
rect 6160 34919 6247 35039
rect 6303 34919 6315 35039
rect 6235 34917 6252 34919
rect 6160 34619 6252 34739
rect 6298 34917 6315 34919
rect 6419 34739 6436 34741
rect 6620 35066 6666 35077
rect 6603 35039 6620 35041
rect 6804 35066 6850 35077
rect 6666 35039 6683 35041
rect 6603 34919 6615 35039
rect 6671 34919 6683 35039
rect 6603 34917 6620 34919
rect 6482 34739 6499 34741
rect 6419 34619 6431 34739
rect 6487 34619 6499 34739
rect 6419 34617 6436 34619
rect 6252 34581 6298 34592
rect 6482 34617 6499 34619
rect 6436 34581 6482 34592
rect 6666 34917 6683 34919
rect 6787 34739 6804 34741
rect 6925 35039 6942 35041
rect 6988 35039 7005 35041
rect 6925 34918 6937 35039
rect 6993 34918 7005 35039
rect 6925 34916 6942 34918
rect 6850 34739 6867 34741
rect 6787 34619 6799 34739
rect 6855 34619 6867 34739
rect 6787 34617 6804 34619
rect 6620 34581 6666 34592
rect 6850 34617 6867 34619
rect 6804 34581 6850 34592
rect 6329 34543 6340 34546
rect 6394 34543 6405 34546
rect 6513 34543 6524 34546
rect 6578 34543 6589 34546
rect 6697 34543 6708 34546
rect 6762 34543 6773 34546
rect 6114 34498 6160 34509
rect 6327 34487 6339 34543
rect 6395 34487 6407 34543
rect 6327 34473 6407 34487
rect 6511 34487 6523 34543
rect 6579 34487 6591 34543
rect 6511 34473 6591 34487
rect 6695 34487 6707 34543
rect 6763 34487 6775 34543
rect 6988 34916 7005 34918
rect 6942 34498 6988 34509
rect 6695 34473 6775 34487
rect 6327 34393 6407 34395
rect 5939 34337 6339 34393
rect 6395 34337 6407 34393
rect 13925 34394 13981 35415
rect 15093 35407 15163 35415
rect 14589 35363 14675 35367
rect 14589 35307 14601 35363
rect 14657 35307 14675 35363
rect 14589 35295 14675 35307
rect 14100 35150 14146 35161
rect 14315 35159 14391 35192
rect 14315 35113 14326 35159
rect 14380 35113 14391 35159
rect 14499 35159 14575 35192
rect 14499 35113 14510 35159
rect 14564 35113 14575 35159
rect 14683 35159 14759 35192
rect 14683 35113 14694 35159
rect 14748 35113 14759 35159
rect 14928 35150 14974 35161
rect 14238 35067 14284 35078
rect 14221 35040 14238 35042
rect 14422 35067 14468 35078
rect 14284 35040 14301 35042
rect 14146 34920 14233 35040
rect 14289 34920 14301 35040
rect 14221 34918 14238 34920
rect 14146 34620 14238 34740
rect 14284 34918 14301 34920
rect 14405 34740 14422 34742
rect 14606 35067 14652 35078
rect 14589 35040 14606 35042
rect 14790 35067 14836 35078
rect 14652 35040 14669 35042
rect 14589 34920 14601 35040
rect 14657 34920 14669 35040
rect 14589 34918 14606 34920
rect 14468 34740 14485 34742
rect 14405 34620 14417 34740
rect 14473 34620 14485 34740
rect 14405 34618 14422 34620
rect 14238 34582 14284 34593
rect 14468 34618 14485 34620
rect 14422 34582 14468 34593
rect 14652 34918 14669 34920
rect 14773 34740 14790 34742
rect 14911 35040 14928 35042
rect 14974 35040 14991 35042
rect 14911 34919 14923 35040
rect 14979 34919 14991 35040
rect 14911 34917 14928 34919
rect 14836 34740 14853 34742
rect 14773 34620 14785 34740
rect 14841 34620 14853 34740
rect 14773 34618 14790 34620
rect 14606 34582 14652 34593
rect 14836 34618 14853 34620
rect 14790 34582 14836 34593
rect 14315 34544 14326 34547
rect 14380 34544 14391 34547
rect 14499 34544 14510 34547
rect 14564 34544 14575 34547
rect 14683 34544 14694 34547
rect 14748 34544 14759 34547
rect 14100 34499 14146 34510
rect 14313 34488 14325 34544
rect 14381 34488 14393 34544
rect 14313 34474 14393 34488
rect 14497 34488 14509 34544
rect 14565 34488 14577 34544
rect 14497 34474 14577 34488
rect 14681 34488 14693 34544
rect 14749 34488 14761 34544
rect 14974 34917 14991 34919
rect 14928 34499 14974 34510
rect 14681 34474 14761 34488
rect 14313 34394 14393 34396
rect 13925 34338 14325 34394
rect 14381 34338 14393 34394
rect 15411 34394 15467 37620
rect 23392 37620 24939 37676
rect 22895 36599 22983 36611
rect 23392 36599 23448 37620
rect 24061 37568 24147 37572
rect 24061 37512 24073 37568
rect 24129 37512 24147 37568
rect 24061 37500 24147 37512
rect 23572 37355 23618 37366
rect 23787 37364 23863 37397
rect 23787 37318 23798 37364
rect 23852 37318 23863 37364
rect 23971 37364 24047 37397
rect 23971 37318 23982 37364
rect 24036 37318 24047 37364
rect 24155 37364 24231 37397
rect 24155 37318 24166 37364
rect 24220 37318 24231 37364
rect 24400 37355 24446 37366
rect 23710 37272 23756 37283
rect 23693 37245 23710 37247
rect 23894 37272 23940 37283
rect 23756 37245 23773 37247
rect 23618 37125 23705 37245
rect 23761 37125 23773 37245
rect 23693 37123 23710 37125
rect 23618 36825 23710 36945
rect 23756 37123 23773 37125
rect 23877 36945 23894 36947
rect 24078 37272 24124 37283
rect 24061 37245 24078 37247
rect 24262 37272 24308 37283
rect 24124 37245 24141 37247
rect 24061 37125 24073 37245
rect 24129 37125 24141 37245
rect 24061 37123 24078 37125
rect 23940 36945 23957 36947
rect 23877 36825 23889 36945
rect 23945 36825 23957 36945
rect 23877 36823 23894 36825
rect 23710 36787 23756 36798
rect 23940 36823 23957 36825
rect 23894 36787 23940 36798
rect 24124 37123 24141 37125
rect 24245 36945 24262 36947
rect 24383 37245 24400 37247
rect 24446 37245 24463 37247
rect 24383 37124 24395 37245
rect 24451 37124 24463 37245
rect 24383 37122 24400 37124
rect 24308 36945 24325 36947
rect 24245 36825 24257 36945
rect 24313 36825 24325 36945
rect 24245 36823 24262 36825
rect 24078 36787 24124 36798
rect 24308 36823 24325 36825
rect 24262 36787 24308 36798
rect 23787 36749 23798 36752
rect 23852 36749 23863 36752
rect 23971 36749 23982 36752
rect 24036 36749 24047 36752
rect 24155 36749 24166 36752
rect 24220 36749 24231 36752
rect 23572 36704 23618 36715
rect 23785 36693 23797 36749
rect 23853 36693 23865 36749
rect 23785 36679 23865 36693
rect 23969 36693 23981 36749
rect 24037 36693 24049 36749
rect 23969 36679 24049 36693
rect 24153 36693 24165 36749
rect 24221 36693 24233 36749
rect 24446 37122 24463 37124
rect 24400 36704 24446 36715
rect 24153 36679 24233 36693
rect 23785 36599 23865 36601
rect 22895 36543 22909 36599
rect 22965 36543 23797 36599
rect 23853 36543 23865 36599
rect 22895 36531 22983 36543
rect 23785 36541 23865 36543
rect 23113 36483 23183 36495
rect 23969 36483 24049 36485
rect 23113 36427 23125 36483
rect 23181 36427 23981 36483
rect 24037 36427 24049 36483
rect 23113 36415 23183 36427
rect 23969 36425 24049 36427
rect 24298 36483 24378 36485
rect 24565 36483 24635 36495
rect 24298 36427 24310 36483
rect 24366 36427 24567 36483
rect 24623 36427 24635 36483
rect 24298 36425 24378 36427
rect 24565 36417 24635 36427
rect 24153 36367 24233 36369
rect 23397 36311 24165 36367
rect 24221 36311 24233 36367
rect 23397 35580 23453 36311
rect 24153 36309 24233 36311
rect 23785 36217 23865 36231
rect 23572 36195 23618 36206
rect 23785 36161 23797 36217
rect 23853 36161 23865 36217
rect 23969 36217 24049 36231
rect 23969 36161 23981 36217
rect 24037 36161 24049 36217
rect 24153 36217 24233 36231
rect 24153 36161 24165 36217
rect 24221 36161 24233 36217
rect 24400 36195 24446 36206
rect 23787 36158 23798 36161
rect 23852 36158 23863 36161
rect 23971 36158 23982 36161
rect 24036 36158 24047 36161
rect 24155 36158 24166 36161
rect 24220 36158 24231 36161
rect 23710 36112 23756 36123
rect 23618 35938 23710 36112
rect 23710 35927 23756 35938
rect 23894 36112 23940 36123
rect 23894 35927 23940 35938
rect 24078 36112 24124 36123
rect 24262 36112 24308 36123
rect 24245 36085 24262 36087
rect 24308 36085 24325 36087
rect 24245 35965 24257 36085
rect 24313 35965 24325 36085
rect 24245 35963 24262 35965
rect 24078 35927 24124 35938
rect 24308 35963 24325 35965
rect 24262 35927 24308 35938
rect 23572 35710 23618 35855
rect 23787 35846 23798 35892
rect 23852 35846 23863 35892
rect 23787 35813 23863 35846
rect 23971 35846 23982 35892
rect 24036 35846 24047 35892
rect 23971 35813 24047 35846
rect 24155 35846 24166 35892
rect 24220 35846 24231 35892
rect 24155 35813 24231 35846
rect 24400 35710 24446 35855
rect 23560 35698 23640 35710
rect 23560 35642 23572 35698
rect 23628 35642 23640 35698
rect 23560 35630 23640 35642
rect 24378 35698 24458 35710
rect 24378 35642 24390 35698
rect 24446 35642 24458 35698
rect 24378 35630 24458 35642
rect 24731 35580 24811 35590
rect 23397 35524 24743 35580
rect 24799 35524 24811 35580
rect 24731 35522 24811 35524
rect 24565 35471 24635 35473
rect 23397 35470 24635 35471
rect 23397 35416 24567 35470
rect 24623 35416 24635 35470
rect 23397 35415 24635 35416
rect 16075 35363 16161 35367
rect 16075 35307 16087 35363
rect 16143 35307 16161 35363
rect 16075 35295 16161 35307
rect 15586 35150 15632 35161
rect 15801 35159 15877 35192
rect 15801 35113 15812 35159
rect 15866 35113 15877 35159
rect 15985 35159 16061 35192
rect 15985 35113 15996 35159
rect 16050 35113 16061 35159
rect 16169 35159 16245 35192
rect 16169 35113 16180 35159
rect 16234 35113 16245 35159
rect 16414 35150 16460 35161
rect 15724 35067 15770 35078
rect 15707 35040 15724 35042
rect 15908 35067 15954 35078
rect 15770 35040 15787 35042
rect 15632 34920 15719 35040
rect 15775 34920 15787 35040
rect 15707 34918 15724 34920
rect 15632 34620 15724 34740
rect 15770 34918 15787 34920
rect 15891 34740 15908 34742
rect 16092 35067 16138 35078
rect 16075 35040 16092 35042
rect 16276 35067 16322 35078
rect 16138 35040 16155 35042
rect 16075 34920 16087 35040
rect 16143 34920 16155 35040
rect 16075 34918 16092 34920
rect 15954 34740 15971 34742
rect 15891 34620 15903 34740
rect 15959 34620 15971 34740
rect 15891 34618 15908 34620
rect 15724 34582 15770 34593
rect 15954 34618 15971 34620
rect 15908 34582 15954 34593
rect 16138 34918 16155 34920
rect 16259 34740 16276 34742
rect 16397 35040 16414 35042
rect 16460 35040 16477 35042
rect 16397 34919 16409 35040
rect 16465 34919 16477 35040
rect 16397 34917 16414 34919
rect 16322 34740 16339 34742
rect 16259 34620 16271 34740
rect 16327 34620 16339 34740
rect 16259 34618 16276 34620
rect 16092 34582 16138 34593
rect 16322 34618 16339 34620
rect 16276 34582 16322 34593
rect 15801 34544 15812 34547
rect 15866 34544 15877 34547
rect 15985 34544 15996 34547
rect 16050 34544 16061 34547
rect 16169 34544 16180 34547
rect 16234 34544 16245 34547
rect 15586 34499 15632 34510
rect 15799 34488 15811 34544
rect 15867 34488 15879 34544
rect 15799 34474 15879 34488
rect 15983 34488 15995 34544
rect 16051 34488 16063 34544
rect 15983 34474 16063 34488
rect 16167 34488 16179 34544
rect 16235 34488 16247 34544
rect 16460 34917 16477 34919
rect 16414 34499 16460 34510
rect 16167 34474 16247 34488
rect 15799 34394 15879 34396
rect 15411 34338 15811 34394
rect 15867 34338 15879 34394
rect 23397 34394 23453 35415
rect 24565 35407 24635 35415
rect 24061 35363 24147 35367
rect 24061 35307 24073 35363
rect 24129 35307 24147 35363
rect 24061 35295 24147 35307
rect 23572 35150 23618 35161
rect 23787 35159 23863 35192
rect 23787 35113 23798 35159
rect 23852 35113 23863 35159
rect 23971 35159 24047 35192
rect 23971 35113 23982 35159
rect 24036 35113 24047 35159
rect 24155 35159 24231 35192
rect 24155 35113 24166 35159
rect 24220 35113 24231 35159
rect 24400 35150 24446 35161
rect 23710 35067 23756 35078
rect 23693 35040 23710 35042
rect 23894 35067 23940 35078
rect 23756 35040 23773 35042
rect 23618 34920 23705 35040
rect 23761 34920 23773 35040
rect 23693 34918 23710 34920
rect 23618 34620 23710 34740
rect 23756 34918 23773 34920
rect 23877 34740 23894 34742
rect 24078 35067 24124 35078
rect 24061 35040 24078 35042
rect 24262 35067 24308 35078
rect 24124 35040 24141 35042
rect 24061 34920 24073 35040
rect 24129 34920 24141 35040
rect 24061 34918 24078 34920
rect 23940 34740 23957 34742
rect 23877 34620 23889 34740
rect 23945 34620 23957 34740
rect 23877 34618 23894 34620
rect 23710 34582 23756 34593
rect 23940 34618 23957 34620
rect 23894 34582 23940 34593
rect 24124 34918 24141 34920
rect 24245 34740 24262 34742
rect 24383 35040 24400 35042
rect 24446 35040 24463 35042
rect 24383 34919 24395 35040
rect 24451 34919 24463 35040
rect 24383 34917 24400 34919
rect 24308 34740 24325 34742
rect 24245 34620 24257 34740
rect 24313 34620 24325 34740
rect 24245 34618 24262 34620
rect 24078 34582 24124 34593
rect 24308 34618 24325 34620
rect 24262 34582 24308 34593
rect 23787 34544 23798 34547
rect 23852 34544 23863 34547
rect 23971 34544 23982 34547
rect 24036 34544 24047 34547
rect 24155 34544 24166 34547
rect 24220 34544 24231 34547
rect 23572 34499 23618 34510
rect 23785 34488 23797 34544
rect 23853 34488 23865 34544
rect 23785 34474 23865 34488
rect 23969 34488 23981 34544
rect 24037 34488 24049 34544
rect 23969 34474 24049 34488
rect 24153 34488 24165 34544
rect 24221 34488 24233 34544
rect 24446 34917 24463 34919
rect 24400 34499 24446 34510
rect 24153 34474 24233 34488
rect 23785 34394 23865 34396
rect 23397 34338 23797 34394
rect 23853 34338 23865 34394
rect 24883 34394 24939 37620
rect 32864 37620 34411 37676
rect 32367 36599 32455 36611
rect 32864 36599 32920 37620
rect 33533 37568 33619 37572
rect 33533 37512 33545 37568
rect 33601 37512 33619 37568
rect 33533 37500 33619 37512
rect 33044 37355 33090 37366
rect 33259 37364 33335 37397
rect 33259 37318 33270 37364
rect 33324 37318 33335 37364
rect 33443 37364 33519 37397
rect 33443 37318 33454 37364
rect 33508 37318 33519 37364
rect 33627 37364 33703 37397
rect 33627 37318 33638 37364
rect 33692 37318 33703 37364
rect 33872 37355 33918 37366
rect 33182 37272 33228 37283
rect 33165 37245 33182 37247
rect 33366 37272 33412 37283
rect 33228 37245 33245 37247
rect 33090 37125 33177 37245
rect 33233 37125 33245 37245
rect 33165 37123 33182 37125
rect 33090 36825 33182 36945
rect 33228 37123 33245 37125
rect 33349 36945 33366 36947
rect 33550 37272 33596 37283
rect 33533 37245 33550 37247
rect 33734 37272 33780 37283
rect 33596 37245 33613 37247
rect 33533 37125 33545 37245
rect 33601 37125 33613 37245
rect 33533 37123 33550 37125
rect 33412 36945 33429 36947
rect 33349 36825 33361 36945
rect 33417 36825 33429 36945
rect 33349 36823 33366 36825
rect 33182 36787 33228 36798
rect 33412 36823 33429 36825
rect 33366 36787 33412 36798
rect 33596 37123 33613 37125
rect 33717 36945 33734 36947
rect 33855 37245 33872 37247
rect 33918 37245 33935 37247
rect 33855 37124 33867 37245
rect 33923 37124 33935 37245
rect 33855 37122 33872 37124
rect 33780 36945 33797 36947
rect 33717 36825 33729 36945
rect 33785 36825 33797 36945
rect 33717 36823 33734 36825
rect 33550 36787 33596 36798
rect 33780 36823 33797 36825
rect 33734 36787 33780 36798
rect 33259 36749 33270 36752
rect 33324 36749 33335 36752
rect 33443 36749 33454 36752
rect 33508 36749 33519 36752
rect 33627 36749 33638 36752
rect 33692 36749 33703 36752
rect 33044 36704 33090 36715
rect 33257 36693 33269 36749
rect 33325 36693 33337 36749
rect 33257 36679 33337 36693
rect 33441 36693 33453 36749
rect 33509 36693 33521 36749
rect 33441 36679 33521 36693
rect 33625 36693 33637 36749
rect 33693 36693 33705 36749
rect 33918 37122 33935 37124
rect 33872 36704 33918 36715
rect 33625 36679 33705 36693
rect 33257 36599 33337 36601
rect 32367 36543 32381 36599
rect 32437 36543 33269 36599
rect 33325 36543 33337 36599
rect 32367 36531 32455 36543
rect 33257 36541 33337 36543
rect 32585 36483 32655 36495
rect 33441 36483 33521 36485
rect 32585 36427 32597 36483
rect 32653 36427 33453 36483
rect 33509 36427 33521 36483
rect 32585 36415 32655 36427
rect 33441 36425 33521 36427
rect 33770 36483 33850 36485
rect 34037 36483 34107 36495
rect 33770 36427 33782 36483
rect 33838 36427 34039 36483
rect 34095 36427 34107 36483
rect 33770 36425 33850 36427
rect 34037 36417 34107 36427
rect 33625 36367 33705 36369
rect 32869 36311 33637 36367
rect 33693 36311 33705 36367
rect 32869 35580 32925 36311
rect 33625 36309 33705 36311
rect 33257 36217 33337 36231
rect 33044 36195 33090 36206
rect 33257 36161 33269 36217
rect 33325 36161 33337 36217
rect 33441 36217 33521 36231
rect 33441 36161 33453 36217
rect 33509 36161 33521 36217
rect 33625 36217 33705 36231
rect 33625 36161 33637 36217
rect 33693 36161 33705 36217
rect 33872 36195 33918 36206
rect 33259 36158 33270 36161
rect 33324 36158 33335 36161
rect 33443 36158 33454 36161
rect 33508 36158 33519 36161
rect 33627 36158 33638 36161
rect 33692 36158 33703 36161
rect 33182 36112 33228 36123
rect 33090 35938 33182 36112
rect 33182 35927 33228 35938
rect 33366 36112 33412 36123
rect 33366 35927 33412 35938
rect 33550 36112 33596 36123
rect 33734 36112 33780 36123
rect 33717 36085 33734 36087
rect 33780 36085 33797 36087
rect 33717 35965 33729 36085
rect 33785 35965 33797 36085
rect 33717 35963 33734 35965
rect 33550 35927 33596 35938
rect 33780 35963 33797 35965
rect 33734 35927 33780 35938
rect 33044 35710 33090 35855
rect 33259 35846 33270 35892
rect 33324 35846 33335 35892
rect 33259 35813 33335 35846
rect 33443 35846 33454 35892
rect 33508 35846 33519 35892
rect 33443 35813 33519 35846
rect 33627 35846 33638 35892
rect 33692 35846 33703 35892
rect 33627 35813 33703 35846
rect 33872 35710 33918 35855
rect 33032 35698 33112 35710
rect 33032 35642 33044 35698
rect 33100 35642 33112 35698
rect 33032 35630 33112 35642
rect 33850 35698 33930 35710
rect 33850 35642 33862 35698
rect 33918 35642 33930 35698
rect 33850 35630 33930 35642
rect 34203 35580 34283 35590
rect 32869 35524 34215 35580
rect 34271 35524 34283 35580
rect 34203 35522 34283 35524
rect 34037 35471 34107 35473
rect 32869 35470 34107 35471
rect 32869 35416 34039 35470
rect 34095 35416 34107 35470
rect 32869 35415 34107 35416
rect 25547 35363 25633 35367
rect 25547 35307 25559 35363
rect 25615 35307 25633 35363
rect 25547 35295 25633 35307
rect 25058 35150 25104 35161
rect 25273 35159 25349 35192
rect 25273 35113 25284 35159
rect 25338 35113 25349 35159
rect 25457 35159 25533 35192
rect 25457 35113 25468 35159
rect 25522 35113 25533 35159
rect 25641 35159 25717 35192
rect 25641 35113 25652 35159
rect 25706 35113 25717 35159
rect 25886 35150 25932 35161
rect 25196 35067 25242 35078
rect 25179 35040 25196 35042
rect 25380 35067 25426 35078
rect 25242 35040 25259 35042
rect 25104 34920 25191 35040
rect 25247 34920 25259 35040
rect 25179 34918 25196 34920
rect 25104 34620 25196 34740
rect 25242 34918 25259 34920
rect 25363 34740 25380 34742
rect 25564 35067 25610 35078
rect 25547 35040 25564 35042
rect 25748 35067 25794 35078
rect 25610 35040 25627 35042
rect 25547 34920 25559 35040
rect 25615 34920 25627 35040
rect 25547 34918 25564 34920
rect 25426 34740 25443 34742
rect 25363 34620 25375 34740
rect 25431 34620 25443 34740
rect 25363 34618 25380 34620
rect 25196 34582 25242 34593
rect 25426 34618 25443 34620
rect 25380 34582 25426 34593
rect 25610 34918 25627 34920
rect 25731 34740 25748 34742
rect 25869 35040 25886 35042
rect 25932 35040 25949 35042
rect 25869 34919 25881 35040
rect 25937 34919 25949 35040
rect 25869 34917 25886 34919
rect 25794 34740 25811 34742
rect 25731 34620 25743 34740
rect 25799 34620 25811 34740
rect 25731 34618 25748 34620
rect 25564 34582 25610 34593
rect 25794 34618 25811 34620
rect 25748 34582 25794 34593
rect 25273 34544 25284 34547
rect 25338 34544 25349 34547
rect 25457 34544 25468 34547
rect 25522 34544 25533 34547
rect 25641 34544 25652 34547
rect 25706 34544 25717 34547
rect 25058 34499 25104 34510
rect 25271 34488 25283 34544
rect 25339 34488 25351 34544
rect 25271 34474 25351 34488
rect 25455 34488 25467 34544
rect 25523 34488 25535 34544
rect 25455 34474 25535 34488
rect 25639 34488 25651 34544
rect 25707 34488 25719 34544
rect 25932 34917 25949 34919
rect 25886 34499 25932 34510
rect 25639 34474 25719 34488
rect 25271 34394 25351 34396
rect 24883 34338 25283 34394
rect 25339 34338 25351 34394
rect 32869 34394 32925 35415
rect 34037 35407 34107 35415
rect 33533 35363 33619 35367
rect 33533 35307 33545 35363
rect 33601 35307 33619 35363
rect 33533 35295 33619 35307
rect 33044 35150 33090 35161
rect 33259 35159 33335 35192
rect 33259 35113 33270 35159
rect 33324 35113 33335 35159
rect 33443 35159 33519 35192
rect 33443 35113 33454 35159
rect 33508 35113 33519 35159
rect 33627 35159 33703 35192
rect 33627 35113 33638 35159
rect 33692 35113 33703 35159
rect 33872 35150 33918 35161
rect 33182 35067 33228 35078
rect 33165 35040 33182 35042
rect 33366 35067 33412 35078
rect 33228 35040 33245 35042
rect 33090 34920 33177 35040
rect 33233 34920 33245 35040
rect 33165 34918 33182 34920
rect 33090 34620 33182 34740
rect 33228 34918 33245 34920
rect 33349 34740 33366 34742
rect 33550 35067 33596 35078
rect 33533 35040 33550 35042
rect 33734 35067 33780 35078
rect 33596 35040 33613 35042
rect 33533 34920 33545 35040
rect 33601 34920 33613 35040
rect 33533 34918 33550 34920
rect 33412 34740 33429 34742
rect 33349 34620 33361 34740
rect 33417 34620 33429 34740
rect 33349 34618 33366 34620
rect 33182 34582 33228 34593
rect 33412 34618 33429 34620
rect 33366 34582 33412 34593
rect 33596 34918 33613 34920
rect 33717 34740 33734 34742
rect 33855 35040 33872 35042
rect 33918 35040 33935 35042
rect 33855 34919 33867 35040
rect 33923 34919 33935 35040
rect 33855 34917 33872 34919
rect 33780 34740 33797 34742
rect 33717 34620 33729 34740
rect 33785 34620 33797 34740
rect 33717 34618 33734 34620
rect 33550 34582 33596 34593
rect 33780 34618 33797 34620
rect 33734 34582 33780 34593
rect 33259 34544 33270 34547
rect 33324 34544 33335 34547
rect 33443 34544 33454 34547
rect 33508 34544 33519 34547
rect 33627 34544 33638 34547
rect 33692 34544 33703 34547
rect 33044 34499 33090 34510
rect 33257 34488 33269 34544
rect 33325 34488 33337 34544
rect 33257 34474 33337 34488
rect 33441 34488 33453 34544
rect 33509 34488 33521 34544
rect 33441 34474 33521 34488
rect 33625 34488 33637 34544
rect 33693 34488 33705 34544
rect 33918 34917 33935 34919
rect 33872 34499 33918 34510
rect 33625 34474 33705 34488
rect 33257 34394 33337 34396
rect 32869 34338 33269 34394
rect 33325 34338 33337 34394
rect 34355 34394 34411 37620
rect 42336 37620 43883 37676
rect 41839 36599 41927 36611
rect 42336 36599 42392 37620
rect 43005 37568 43091 37572
rect 43005 37512 43017 37568
rect 43073 37512 43091 37568
rect 43005 37500 43091 37512
rect 42516 37355 42562 37366
rect 42731 37364 42807 37397
rect 42731 37318 42742 37364
rect 42796 37318 42807 37364
rect 42915 37364 42991 37397
rect 42915 37318 42926 37364
rect 42980 37318 42991 37364
rect 43099 37364 43175 37397
rect 43099 37318 43110 37364
rect 43164 37318 43175 37364
rect 43344 37355 43390 37366
rect 42654 37272 42700 37283
rect 42637 37245 42654 37247
rect 42838 37272 42884 37283
rect 42700 37245 42717 37247
rect 42562 37125 42649 37245
rect 42705 37125 42717 37245
rect 42637 37123 42654 37125
rect 42562 36825 42654 36945
rect 42700 37123 42717 37125
rect 42821 36945 42838 36947
rect 43022 37272 43068 37283
rect 43005 37245 43022 37247
rect 43206 37272 43252 37283
rect 43068 37245 43085 37247
rect 43005 37125 43017 37245
rect 43073 37125 43085 37245
rect 43005 37123 43022 37125
rect 42884 36945 42901 36947
rect 42821 36825 42833 36945
rect 42889 36825 42901 36945
rect 42821 36823 42838 36825
rect 42654 36787 42700 36798
rect 42884 36823 42901 36825
rect 42838 36787 42884 36798
rect 43068 37123 43085 37125
rect 43189 36945 43206 36947
rect 43327 37245 43344 37247
rect 43390 37245 43407 37247
rect 43327 37124 43339 37245
rect 43395 37124 43407 37245
rect 43327 37122 43344 37124
rect 43252 36945 43269 36947
rect 43189 36825 43201 36945
rect 43257 36825 43269 36945
rect 43189 36823 43206 36825
rect 43022 36787 43068 36798
rect 43252 36823 43269 36825
rect 43206 36787 43252 36798
rect 42731 36749 42742 36752
rect 42796 36749 42807 36752
rect 42915 36749 42926 36752
rect 42980 36749 42991 36752
rect 43099 36749 43110 36752
rect 43164 36749 43175 36752
rect 42516 36704 42562 36715
rect 42729 36693 42741 36749
rect 42797 36693 42809 36749
rect 42729 36679 42809 36693
rect 42913 36693 42925 36749
rect 42981 36693 42993 36749
rect 42913 36679 42993 36693
rect 43097 36693 43109 36749
rect 43165 36693 43177 36749
rect 43390 37122 43407 37124
rect 43344 36704 43390 36715
rect 43097 36679 43177 36693
rect 42729 36599 42809 36601
rect 41839 36543 41853 36599
rect 41909 36543 42741 36599
rect 42797 36543 42809 36599
rect 41839 36531 41927 36543
rect 42729 36541 42809 36543
rect 42057 36483 42127 36495
rect 42913 36483 42993 36485
rect 42057 36427 42069 36483
rect 42125 36427 42925 36483
rect 42981 36427 42993 36483
rect 42057 36415 42127 36427
rect 42913 36425 42993 36427
rect 43242 36483 43322 36485
rect 43509 36483 43579 36495
rect 43242 36427 43254 36483
rect 43310 36427 43511 36483
rect 43567 36427 43579 36483
rect 43242 36425 43322 36427
rect 43509 36417 43579 36427
rect 43097 36367 43177 36369
rect 42341 36311 43109 36367
rect 43165 36311 43177 36367
rect 42341 35580 42397 36311
rect 43097 36309 43177 36311
rect 42729 36217 42809 36231
rect 42516 36195 42562 36206
rect 42729 36161 42741 36217
rect 42797 36161 42809 36217
rect 42913 36217 42993 36231
rect 42913 36161 42925 36217
rect 42981 36161 42993 36217
rect 43097 36217 43177 36231
rect 43097 36161 43109 36217
rect 43165 36161 43177 36217
rect 43344 36195 43390 36206
rect 42731 36158 42742 36161
rect 42796 36158 42807 36161
rect 42915 36158 42926 36161
rect 42980 36158 42991 36161
rect 43099 36158 43110 36161
rect 43164 36158 43175 36161
rect 42654 36112 42700 36123
rect 42562 35938 42654 36112
rect 42654 35927 42700 35938
rect 42838 36112 42884 36123
rect 42838 35927 42884 35938
rect 43022 36112 43068 36123
rect 43206 36112 43252 36123
rect 43189 36085 43206 36087
rect 43252 36085 43269 36087
rect 43189 35965 43201 36085
rect 43257 35965 43269 36085
rect 43189 35963 43206 35965
rect 43022 35927 43068 35938
rect 43252 35963 43269 35965
rect 43206 35927 43252 35938
rect 42516 35710 42562 35855
rect 42731 35846 42742 35892
rect 42796 35846 42807 35892
rect 42731 35813 42807 35846
rect 42915 35846 42926 35892
rect 42980 35846 42991 35892
rect 42915 35813 42991 35846
rect 43099 35846 43110 35892
rect 43164 35846 43175 35892
rect 43099 35813 43175 35846
rect 43344 35710 43390 35855
rect 42504 35698 42584 35710
rect 42504 35642 42516 35698
rect 42572 35642 42584 35698
rect 42504 35630 42584 35642
rect 43322 35698 43402 35710
rect 43322 35642 43334 35698
rect 43390 35642 43402 35698
rect 43322 35630 43402 35642
rect 43675 35580 43755 35590
rect 42341 35524 43687 35580
rect 43743 35524 43755 35580
rect 43675 35522 43755 35524
rect 43509 35471 43579 35473
rect 42341 35470 43579 35471
rect 42341 35416 43511 35470
rect 43567 35416 43579 35470
rect 42341 35415 43579 35416
rect 35019 35363 35105 35367
rect 35019 35307 35031 35363
rect 35087 35307 35105 35363
rect 35019 35295 35105 35307
rect 34530 35150 34576 35161
rect 34745 35159 34821 35192
rect 34745 35113 34756 35159
rect 34810 35113 34821 35159
rect 34929 35159 35005 35192
rect 34929 35113 34940 35159
rect 34994 35113 35005 35159
rect 35113 35159 35189 35192
rect 35113 35113 35124 35159
rect 35178 35113 35189 35159
rect 35358 35150 35404 35161
rect 34668 35067 34714 35078
rect 34651 35040 34668 35042
rect 34852 35067 34898 35078
rect 34714 35040 34731 35042
rect 34576 34920 34663 35040
rect 34719 34920 34731 35040
rect 34651 34918 34668 34920
rect 34576 34620 34668 34740
rect 34714 34918 34731 34920
rect 34835 34740 34852 34742
rect 35036 35067 35082 35078
rect 35019 35040 35036 35042
rect 35220 35067 35266 35078
rect 35082 35040 35099 35042
rect 35019 34920 35031 35040
rect 35087 34920 35099 35040
rect 35019 34918 35036 34920
rect 34898 34740 34915 34742
rect 34835 34620 34847 34740
rect 34903 34620 34915 34740
rect 34835 34618 34852 34620
rect 34668 34582 34714 34593
rect 34898 34618 34915 34620
rect 34852 34582 34898 34593
rect 35082 34918 35099 34920
rect 35203 34740 35220 34742
rect 35341 35040 35358 35042
rect 35404 35040 35421 35042
rect 35341 34919 35353 35040
rect 35409 34919 35421 35040
rect 35341 34917 35358 34919
rect 35266 34740 35283 34742
rect 35203 34620 35215 34740
rect 35271 34620 35283 34740
rect 35203 34618 35220 34620
rect 35036 34582 35082 34593
rect 35266 34618 35283 34620
rect 35220 34582 35266 34593
rect 34745 34544 34756 34547
rect 34810 34544 34821 34547
rect 34929 34544 34940 34547
rect 34994 34544 35005 34547
rect 35113 34544 35124 34547
rect 35178 34544 35189 34547
rect 34530 34499 34576 34510
rect 34743 34488 34755 34544
rect 34811 34488 34823 34544
rect 34743 34474 34823 34488
rect 34927 34488 34939 34544
rect 34995 34488 35007 34544
rect 34927 34474 35007 34488
rect 35111 34488 35123 34544
rect 35179 34488 35191 34544
rect 35404 34917 35421 34919
rect 35358 34499 35404 34510
rect 35111 34474 35191 34488
rect 34743 34394 34823 34396
rect 34355 34338 34755 34394
rect 34811 34338 34823 34394
rect 42341 34394 42397 35415
rect 43509 35407 43579 35415
rect 43005 35363 43091 35367
rect 43005 35307 43017 35363
rect 43073 35307 43091 35363
rect 43005 35295 43091 35307
rect 42516 35150 42562 35161
rect 42731 35159 42807 35192
rect 42731 35113 42742 35159
rect 42796 35113 42807 35159
rect 42915 35159 42991 35192
rect 42915 35113 42926 35159
rect 42980 35113 42991 35159
rect 43099 35159 43175 35192
rect 43099 35113 43110 35159
rect 43164 35113 43175 35159
rect 43344 35150 43390 35161
rect 42654 35067 42700 35078
rect 42637 35040 42654 35042
rect 42838 35067 42884 35078
rect 42700 35040 42717 35042
rect 42562 34920 42649 35040
rect 42705 34920 42717 35040
rect 42637 34918 42654 34920
rect 42562 34620 42654 34740
rect 42700 34918 42717 34920
rect 42821 34740 42838 34742
rect 43022 35067 43068 35078
rect 43005 35040 43022 35042
rect 43206 35067 43252 35078
rect 43068 35040 43085 35042
rect 43005 34920 43017 35040
rect 43073 34920 43085 35040
rect 43005 34918 43022 34920
rect 42884 34740 42901 34742
rect 42821 34620 42833 34740
rect 42889 34620 42901 34740
rect 42821 34618 42838 34620
rect 42654 34582 42700 34593
rect 42884 34618 42901 34620
rect 42838 34582 42884 34593
rect 43068 34918 43085 34920
rect 43189 34740 43206 34742
rect 43327 35040 43344 35042
rect 43390 35040 43407 35042
rect 43327 34919 43339 35040
rect 43395 34919 43407 35040
rect 43327 34917 43344 34919
rect 43252 34740 43269 34742
rect 43189 34620 43201 34740
rect 43257 34620 43269 34740
rect 43189 34618 43206 34620
rect 43022 34582 43068 34593
rect 43252 34618 43269 34620
rect 43206 34582 43252 34593
rect 42731 34544 42742 34547
rect 42796 34544 42807 34547
rect 42915 34544 42926 34547
rect 42980 34544 42991 34547
rect 43099 34544 43110 34547
rect 43164 34544 43175 34547
rect 42516 34499 42562 34510
rect 42729 34488 42741 34544
rect 42797 34488 42809 34544
rect 42729 34474 42809 34488
rect 42913 34488 42925 34544
rect 42981 34488 42993 34544
rect 42913 34474 42993 34488
rect 43097 34488 43109 34544
rect 43165 34488 43177 34544
rect 43390 34917 43407 34919
rect 43344 34499 43390 34510
rect 43097 34474 43177 34488
rect 42729 34394 42809 34396
rect 42341 34338 42741 34394
rect 42797 34338 42809 34394
rect 43827 34394 43883 37620
rect 44491 35363 44577 35367
rect 44491 35307 44503 35363
rect 44559 35307 44577 35363
rect 44491 35295 44577 35307
rect 44002 35150 44048 35161
rect 44217 35159 44293 35192
rect 44217 35113 44228 35159
rect 44282 35113 44293 35159
rect 44401 35159 44477 35192
rect 44401 35113 44412 35159
rect 44466 35113 44477 35159
rect 44585 35159 44661 35192
rect 44585 35113 44596 35159
rect 44650 35113 44661 35159
rect 44830 35150 44876 35161
rect 44140 35067 44186 35078
rect 44123 35040 44140 35042
rect 44324 35067 44370 35078
rect 44186 35040 44203 35042
rect 44048 34920 44135 35040
rect 44191 34920 44203 35040
rect 44123 34918 44140 34920
rect 44048 34620 44140 34740
rect 44186 34918 44203 34920
rect 44307 34740 44324 34742
rect 44508 35067 44554 35078
rect 44491 35040 44508 35042
rect 44692 35067 44738 35078
rect 44554 35040 44571 35042
rect 44491 34920 44503 35040
rect 44559 34920 44571 35040
rect 44491 34918 44508 34920
rect 44370 34740 44387 34742
rect 44307 34620 44319 34740
rect 44375 34620 44387 34740
rect 44307 34618 44324 34620
rect 44140 34582 44186 34593
rect 44370 34618 44387 34620
rect 44324 34582 44370 34593
rect 44554 34918 44571 34920
rect 44675 34740 44692 34742
rect 44813 35040 44830 35042
rect 44876 35040 44893 35042
rect 44813 34919 44825 35040
rect 44881 34919 44893 35040
rect 44813 34917 44830 34919
rect 44738 34740 44755 34742
rect 44675 34620 44687 34740
rect 44743 34620 44755 34740
rect 44675 34618 44692 34620
rect 44508 34582 44554 34593
rect 44738 34618 44755 34620
rect 44692 34582 44738 34593
rect 44217 34544 44228 34547
rect 44282 34544 44293 34547
rect 44401 34544 44412 34547
rect 44466 34544 44477 34547
rect 44585 34544 44596 34547
rect 44650 34544 44661 34547
rect 44002 34499 44048 34510
rect 44215 34488 44227 34544
rect 44283 34488 44295 34544
rect 44215 34474 44295 34488
rect 44399 34488 44411 34544
rect 44467 34488 44479 34544
rect 44399 34474 44479 34488
rect 44583 34488 44595 34544
rect 44651 34488 44663 34544
rect 44876 34917 44893 34919
rect 44830 34499 44876 34510
rect 44583 34474 44663 34488
rect 44215 34394 44295 34396
rect 43827 34338 44227 34394
rect 44283 34338 44295 34394
rect -4631 34335 -4551 34337
rect -3145 34335 -3065 34337
rect 4841 34335 4921 34337
rect 6327 34335 6407 34337
rect 14313 34336 14393 34338
rect 15799 34336 15879 34338
rect 23785 34336 23865 34338
rect 25271 34336 25351 34338
rect 33257 34336 33337 34338
rect 34743 34336 34823 34338
rect 42729 34336 42809 34338
rect 44215 34336 44295 34338
rect -5439 34277 -5369 34291
rect -4447 34277 -4367 34279
rect -5439 34221 -5427 34277
rect -5371 34221 -4435 34277
rect -4379 34221 -4367 34277
rect -5439 34209 -5369 34221
rect -4447 34219 -4367 34221
rect -4118 34277 -4038 34279
rect -3675 34277 -3615 34287
rect -2961 34277 -2881 34279
rect -4118 34221 -4106 34277
rect -4050 34221 -3673 34277
rect -3617 34221 -2949 34277
rect -2893 34221 -2881 34277
rect -4118 34219 -4038 34221
rect -3675 34209 -3615 34221
rect -2961 34219 -2881 34221
rect -2632 34277 -2552 34279
rect -2365 34277 -2295 34289
rect -2632 34221 -2620 34277
rect -2564 34221 -2363 34277
rect -2307 34221 -2295 34277
rect -2632 34219 -2552 34221
rect -2365 34211 -2295 34221
rect 4033 34277 4103 34291
rect 5025 34277 5105 34279
rect 4033 34221 4045 34277
rect 4101 34221 5037 34277
rect 5093 34221 5105 34277
rect 4033 34209 4103 34221
rect 5025 34219 5105 34221
rect 5354 34277 5434 34279
rect 5797 34277 5857 34287
rect 6511 34277 6591 34279
rect 5354 34221 5366 34277
rect 5422 34221 5799 34277
rect 5855 34221 6523 34277
rect 6579 34221 6591 34277
rect 5354 34219 5434 34221
rect 5797 34209 5857 34221
rect 6511 34219 6591 34221
rect 6840 34277 6920 34279
rect 7107 34277 7177 34289
rect 6840 34221 6852 34277
rect 6908 34221 7109 34277
rect 7165 34221 7177 34277
rect 6840 34219 6920 34221
rect 7107 34211 7177 34221
rect 13505 34278 13575 34292
rect 14497 34278 14577 34280
rect 13505 34222 13517 34278
rect 13573 34222 14509 34278
rect 14565 34222 14577 34278
rect 13505 34210 13575 34222
rect 14497 34220 14577 34222
rect 14826 34278 14906 34280
rect 15269 34278 15329 34288
rect 15983 34278 16063 34280
rect 14826 34222 14838 34278
rect 14894 34222 15271 34278
rect 15327 34222 15995 34278
rect 16051 34222 16063 34278
rect 14826 34220 14906 34222
rect 15269 34210 15329 34222
rect 15983 34220 16063 34222
rect 16312 34278 16392 34280
rect 16579 34278 16649 34290
rect 16312 34222 16324 34278
rect 16380 34222 16581 34278
rect 16637 34222 16649 34278
rect 16312 34220 16392 34222
rect 16579 34212 16649 34222
rect 22977 34278 23047 34292
rect 23969 34278 24049 34280
rect 22977 34222 22989 34278
rect 23045 34222 23981 34278
rect 24037 34222 24049 34278
rect 22977 34210 23047 34222
rect 23969 34220 24049 34222
rect 24298 34278 24378 34280
rect 24741 34278 24801 34288
rect 25455 34278 25535 34280
rect 24298 34222 24310 34278
rect 24366 34222 24743 34278
rect 24799 34222 25467 34278
rect 25523 34222 25535 34278
rect 24298 34220 24378 34222
rect 24741 34210 24801 34222
rect 25455 34220 25535 34222
rect 25784 34278 25864 34280
rect 26051 34278 26121 34290
rect 25784 34222 25796 34278
rect 25852 34222 26053 34278
rect 26109 34222 26121 34278
rect 25784 34220 25864 34222
rect 26051 34212 26121 34222
rect 32449 34278 32519 34292
rect 33441 34278 33521 34280
rect 32449 34222 32461 34278
rect 32517 34222 33453 34278
rect 33509 34222 33521 34278
rect 32449 34210 32519 34222
rect 33441 34220 33521 34222
rect 33770 34278 33850 34280
rect 34213 34278 34273 34288
rect 34927 34278 35007 34280
rect 33770 34222 33782 34278
rect 33838 34222 34215 34278
rect 34271 34222 34939 34278
rect 34995 34222 35007 34278
rect 33770 34220 33850 34222
rect 34213 34210 34273 34222
rect 34927 34220 35007 34222
rect 35256 34278 35336 34280
rect 35523 34278 35593 34290
rect 35256 34222 35268 34278
rect 35324 34222 35525 34278
rect 35581 34222 35593 34278
rect 35256 34220 35336 34222
rect 35523 34212 35593 34222
rect 41921 34278 41991 34292
rect 42913 34278 42993 34280
rect 41921 34222 41933 34278
rect 41989 34222 42925 34278
rect 42981 34222 42993 34278
rect 41921 34210 41991 34222
rect 42913 34220 42993 34222
rect 43242 34278 43322 34280
rect 43685 34278 43745 34288
rect 44399 34278 44479 34280
rect 43242 34222 43254 34278
rect 43310 34222 43687 34278
rect 43743 34222 44411 34278
rect 44467 34222 44479 34278
rect 43242 34220 43322 34222
rect 43685 34210 43745 34222
rect 44399 34220 44479 34222
rect 44728 34278 44808 34280
rect 44995 34278 45065 34290
rect 44728 34222 44740 34278
rect 44796 34222 44997 34278
rect 45053 34222 45065 34278
rect 44728 34220 44808 34222
rect 44995 34212 45065 34222
rect -4263 34161 -4183 34163
rect -2777 34161 -2697 34163
rect 5209 34161 5289 34163
rect 6695 34161 6775 34163
rect 14681 34162 14761 34164
rect 16167 34162 16247 34164
rect 24153 34162 24233 34164
rect 25639 34162 25719 34164
rect 33625 34162 33705 34164
rect 35111 34162 35191 34164
rect 43097 34162 43177 34164
rect 44583 34162 44663 34164
rect -5155 34105 -4251 34161
rect -4195 34105 -4183 34161
rect -5721 33375 -5639 33387
rect -5155 33375 -5099 34105
rect -4263 34103 -4183 34105
rect -3533 34105 -2765 34161
rect -2709 34105 -2697 34161
rect -4631 34011 -4551 34025
rect -4844 33989 -4798 34000
rect -4631 33955 -4619 34011
rect -4563 33955 -4551 34011
rect -4447 34011 -4367 34025
rect -4447 33955 -4435 34011
rect -4379 33955 -4367 34011
rect -4263 34011 -4183 34025
rect -4263 33955 -4251 34011
rect -4195 33955 -4183 34011
rect -4016 33989 -3970 34000
rect -4629 33952 -4618 33955
rect -4564 33952 -4553 33955
rect -4445 33952 -4434 33955
rect -4380 33952 -4369 33955
rect -4261 33952 -4250 33955
rect -4196 33952 -4185 33955
rect -4706 33906 -4660 33917
rect -4798 33732 -4706 33906
rect -4706 33721 -4660 33732
rect -4522 33906 -4476 33917
rect -4522 33721 -4476 33732
rect -4338 33906 -4292 33917
rect -4154 33906 -4108 33917
rect -4171 33879 -4154 33881
rect -4108 33879 -4091 33881
rect -4171 33759 -4159 33879
rect -4103 33759 -4091 33879
rect -4171 33757 -4154 33759
rect -4338 33721 -4292 33732
rect -4108 33757 -4091 33759
rect -4154 33721 -4108 33732
rect -4844 33504 -4798 33649
rect -4629 33640 -4618 33686
rect -4564 33640 -4553 33686
rect -4629 33607 -4553 33640
rect -4445 33640 -4434 33686
rect -4380 33640 -4369 33686
rect -4445 33607 -4369 33640
rect -4261 33640 -4250 33686
rect -4196 33640 -4185 33686
rect -4261 33607 -4185 33640
rect -4016 33504 -3970 33649
rect -4856 33492 -4776 33504
rect -4856 33436 -4844 33492
rect -4788 33436 -4776 33492
rect -4856 33424 -4776 33436
rect -4038 33492 -3960 33504
rect -4038 33436 -4026 33492
rect -3970 33436 -3960 33492
rect -4038 33424 -3960 33436
rect -5721 33319 -5707 33375
rect -5651 33319 -5099 33375
rect -3533 33375 -3477 34105
rect -2777 34103 -2697 34105
rect 4317 34105 5221 34161
rect 5277 34105 5289 34161
rect -3145 34011 -3065 34025
rect -3358 33989 -3312 34000
rect -3145 33955 -3133 34011
rect -3077 33955 -3065 34011
rect -2961 34011 -2881 34025
rect -2961 33955 -2949 34011
rect -2893 33955 -2881 34011
rect -2777 34011 -2697 34025
rect -2777 33955 -2765 34011
rect -2709 33955 -2697 34011
rect -2530 33989 -2484 34000
rect -3143 33952 -3132 33955
rect -3078 33952 -3067 33955
rect -2959 33952 -2948 33955
rect -2894 33952 -2883 33955
rect -2775 33952 -2764 33955
rect -2710 33952 -2699 33955
rect -3220 33906 -3174 33917
rect -3312 33732 -3220 33906
rect -3220 33721 -3174 33732
rect -3036 33906 -2990 33917
rect -3036 33721 -2990 33732
rect -2852 33906 -2806 33917
rect -2668 33906 -2622 33917
rect -2685 33879 -2668 33881
rect -2622 33879 -2605 33881
rect -2685 33759 -2673 33879
rect -2617 33759 -2605 33879
rect -2685 33757 -2668 33759
rect -2852 33721 -2806 33732
rect -2622 33757 -2605 33759
rect -2668 33721 -2622 33732
rect -3358 33504 -3312 33649
rect -3143 33640 -3132 33686
rect -3078 33640 -3067 33686
rect -3143 33607 -3067 33640
rect -2959 33640 -2948 33686
rect -2894 33640 -2883 33686
rect -2959 33607 -2883 33640
rect -2775 33640 -2764 33686
rect -2710 33640 -2699 33686
rect -2775 33607 -2699 33640
rect -2530 33504 -2484 33649
rect -3370 33492 -3290 33504
rect -3370 33436 -3358 33492
rect -3302 33436 -3290 33492
rect -3370 33424 -3290 33436
rect -2552 33492 -2474 33504
rect -2552 33436 -2540 33492
rect -2484 33436 -2474 33492
rect -2552 33424 -2474 33436
rect -2199 33375 -2119 33385
rect -3533 33319 -2187 33375
rect -2131 33319 -2119 33375
rect -5721 33307 -5639 33319
rect -10921 31969 -5827 32169
rect -5155 32072 -5099 33319
rect -2199 33317 -2119 33319
rect 3751 33375 3833 33387
rect 4317 33375 4373 34105
rect 5209 34103 5289 34105
rect 5939 34105 6707 34161
rect 6763 34105 6775 34161
rect 4841 34011 4921 34025
rect 4628 33989 4674 34000
rect 4841 33955 4853 34011
rect 4909 33955 4921 34011
rect 5025 34011 5105 34025
rect 5025 33955 5037 34011
rect 5093 33955 5105 34011
rect 5209 34011 5289 34025
rect 5209 33955 5221 34011
rect 5277 33955 5289 34011
rect 5456 33989 5502 34000
rect 4843 33952 4854 33955
rect 4908 33952 4919 33955
rect 5027 33952 5038 33955
rect 5092 33952 5103 33955
rect 5211 33952 5222 33955
rect 5276 33952 5287 33955
rect 4766 33906 4812 33917
rect 4674 33732 4766 33906
rect 4766 33721 4812 33732
rect 4950 33906 4996 33917
rect 4950 33721 4996 33732
rect 5134 33906 5180 33917
rect 5318 33906 5364 33917
rect 5301 33879 5318 33881
rect 5364 33879 5381 33881
rect 5301 33759 5313 33879
rect 5369 33759 5381 33879
rect 5301 33757 5318 33759
rect 5134 33721 5180 33732
rect 5364 33757 5381 33759
rect 5318 33721 5364 33732
rect 4628 33504 4674 33649
rect 4843 33640 4854 33686
rect 4908 33640 4919 33686
rect 4843 33607 4919 33640
rect 5027 33640 5038 33686
rect 5092 33640 5103 33686
rect 5027 33607 5103 33640
rect 5211 33640 5222 33686
rect 5276 33640 5287 33686
rect 5211 33607 5287 33640
rect 5456 33504 5502 33649
rect 4616 33492 4696 33504
rect 4616 33436 4628 33492
rect 4684 33436 4696 33492
rect 4616 33424 4696 33436
rect 5434 33492 5512 33504
rect 5434 33436 5446 33492
rect 5502 33436 5512 33492
rect 5434 33424 5512 33436
rect 3751 33319 3765 33375
rect 3821 33319 4373 33375
rect 5939 33375 5995 34105
rect 6695 34103 6775 34105
rect 13789 34106 14693 34162
rect 14749 34106 14761 34162
rect 6327 34011 6407 34025
rect 6114 33989 6160 34000
rect 6327 33955 6339 34011
rect 6395 33955 6407 34011
rect 6511 34011 6591 34025
rect 6511 33955 6523 34011
rect 6579 33955 6591 34011
rect 6695 34011 6775 34025
rect 6695 33955 6707 34011
rect 6763 33955 6775 34011
rect 6942 33989 6988 34000
rect 6329 33952 6340 33955
rect 6394 33952 6405 33955
rect 6513 33952 6524 33955
rect 6578 33952 6589 33955
rect 6697 33952 6708 33955
rect 6762 33952 6773 33955
rect 6252 33906 6298 33917
rect 6160 33732 6252 33906
rect 6252 33721 6298 33732
rect 6436 33906 6482 33917
rect 6436 33721 6482 33732
rect 6620 33906 6666 33917
rect 6804 33906 6850 33917
rect 6787 33879 6804 33881
rect 6850 33879 6867 33881
rect 6787 33759 6799 33879
rect 6855 33759 6867 33879
rect 6787 33757 6804 33759
rect 6620 33721 6666 33732
rect 6850 33757 6867 33759
rect 6804 33721 6850 33732
rect 6114 33504 6160 33649
rect 6329 33640 6340 33686
rect 6394 33640 6405 33686
rect 6329 33607 6405 33640
rect 6513 33640 6524 33686
rect 6578 33640 6589 33686
rect 6513 33607 6589 33640
rect 6697 33640 6708 33686
rect 6762 33640 6773 33686
rect 6697 33607 6773 33640
rect 6942 33504 6988 33649
rect 6102 33492 6182 33504
rect 6102 33436 6114 33492
rect 6170 33436 6182 33492
rect 6102 33424 6182 33436
rect 6920 33492 6998 33504
rect 6920 33436 6932 33492
rect 6988 33436 6998 33492
rect 6920 33424 6998 33436
rect 7273 33375 7353 33385
rect 5939 33319 7285 33375
rect 7341 33319 7353 33375
rect 3751 33307 3833 33319
rect -3675 33264 -3605 33266
rect -2375 33265 -2295 33267
rect -5019 33208 -3673 33264
rect -3617 33208 -3605 33264
rect -5019 32188 -4963 33208
rect -3675 33196 -3605 33208
rect -3533 33209 -2363 33265
rect -2307 33209 -2295 33265
rect -4355 33157 -4269 33161
rect -4355 33101 -4343 33157
rect -4287 33101 -4269 33157
rect -4355 33089 -4269 33101
rect -4844 32944 -4798 32955
rect -4629 32953 -4553 32986
rect -4629 32907 -4618 32953
rect -4564 32907 -4553 32953
rect -4445 32953 -4369 32986
rect -4445 32907 -4434 32953
rect -4380 32907 -4369 32953
rect -4261 32953 -4185 32986
rect -4261 32907 -4250 32953
rect -4196 32907 -4185 32953
rect -4016 32944 -3970 32955
rect -4706 32861 -4660 32872
rect -4723 32834 -4706 32836
rect -4522 32861 -4476 32872
rect -4660 32834 -4643 32836
rect -4798 32714 -4711 32834
rect -4655 32714 -4643 32834
rect -4723 32712 -4706 32714
rect -4798 32414 -4706 32534
rect -4660 32712 -4643 32714
rect -4539 32534 -4522 32536
rect -4338 32861 -4292 32872
rect -4355 32834 -4338 32836
rect -4154 32861 -4108 32872
rect -4292 32834 -4275 32836
rect -4355 32714 -4343 32834
rect -4287 32714 -4275 32834
rect -4355 32712 -4338 32714
rect -4476 32534 -4459 32536
rect -4539 32414 -4527 32534
rect -4471 32414 -4459 32534
rect -4539 32412 -4522 32414
rect -4706 32376 -4660 32387
rect -4476 32412 -4459 32414
rect -4522 32376 -4476 32387
rect -4292 32712 -4275 32714
rect -4171 32534 -4154 32536
rect -4033 32834 -4016 32836
rect -3970 32834 -3953 32836
rect -4033 32713 -4021 32834
rect -3965 32713 -3953 32834
rect -4033 32711 -4016 32713
rect -4108 32534 -4091 32536
rect -4171 32414 -4159 32534
rect -4103 32414 -4091 32534
rect -4171 32412 -4154 32414
rect -4338 32376 -4292 32387
rect -4108 32412 -4091 32414
rect -4154 32376 -4108 32387
rect -4629 32338 -4618 32341
rect -4564 32338 -4553 32341
rect -4445 32338 -4434 32341
rect -4380 32338 -4369 32341
rect -4261 32338 -4250 32341
rect -4196 32338 -4185 32341
rect -4844 32293 -4798 32304
rect -4631 32282 -4619 32338
rect -4563 32282 -4551 32338
rect -4631 32268 -4551 32282
rect -4447 32282 -4435 32338
rect -4379 32282 -4367 32338
rect -4447 32268 -4367 32282
rect -4263 32282 -4251 32338
rect -4195 32282 -4183 32338
rect -3970 32711 -3953 32713
rect -4016 32293 -3970 32304
rect -4263 32268 -4183 32282
rect -4631 32188 -4551 32190
rect -5019 32132 -4619 32188
rect -4563 32132 -4551 32188
rect -3533 32189 -3477 33209
rect -2375 33197 -2295 33209
rect -2869 33158 -2783 33162
rect -2869 33102 -2857 33158
rect -2801 33102 -2783 33158
rect -2869 33090 -2783 33102
rect -3358 32945 -3312 32956
rect -3143 32954 -3067 32987
rect -3143 32908 -3132 32954
rect -3078 32908 -3067 32954
rect -2959 32954 -2883 32987
rect -2959 32908 -2948 32954
rect -2894 32908 -2883 32954
rect -2775 32954 -2699 32987
rect -2775 32908 -2764 32954
rect -2710 32908 -2699 32954
rect -2530 32945 -2484 32956
rect -3220 32862 -3174 32873
rect -3237 32835 -3220 32837
rect -3036 32862 -2990 32873
rect -3174 32835 -3157 32837
rect -3312 32715 -3225 32835
rect -3169 32715 -3157 32835
rect -3237 32713 -3220 32715
rect -3312 32415 -3220 32535
rect -3174 32713 -3157 32715
rect -3053 32535 -3036 32537
rect -2852 32862 -2806 32873
rect -2869 32835 -2852 32837
rect -2668 32862 -2622 32873
rect -2806 32835 -2789 32837
rect -2869 32715 -2857 32835
rect -2801 32715 -2789 32835
rect -2869 32713 -2852 32715
rect -2990 32535 -2973 32537
rect -3053 32415 -3041 32535
rect -2985 32415 -2973 32535
rect -3053 32413 -3036 32415
rect -3220 32377 -3174 32388
rect -2990 32413 -2973 32415
rect -3036 32377 -2990 32388
rect -2806 32713 -2789 32715
rect -2685 32535 -2668 32537
rect -2547 32835 -2530 32837
rect -2484 32835 -2467 32837
rect -2547 32714 -2535 32835
rect -2479 32714 -2467 32835
rect -2547 32712 -2530 32714
rect -2622 32535 -2605 32537
rect -2685 32415 -2673 32535
rect -2617 32415 -2605 32535
rect -2685 32413 -2668 32415
rect -2852 32377 -2806 32388
rect -2622 32413 -2605 32415
rect -2668 32377 -2622 32388
rect -3143 32339 -3132 32342
rect -3078 32339 -3067 32342
rect -2959 32339 -2948 32342
rect -2894 32339 -2883 32342
rect -2775 32339 -2764 32342
rect -2710 32339 -2699 32342
rect -3358 32294 -3312 32305
rect -3145 32283 -3133 32339
rect -3077 32283 -3065 32339
rect -3145 32269 -3065 32283
rect -2961 32283 -2949 32339
rect -2893 32283 -2881 32339
rect -2961 32269 -2881 32283
rect -2777 32283 -2765 32339
rect -2709 32283 -2697 32339
rect -2484 32712 -2467 32714
rect -2530 32294 -2484 32305
rect -2777 32269 -2697 32283
rect -3145 32189 -3065 32191
rect -3533 32133 -3133 32189
rect -3077 32133 -3065 32189
rect -4631 32130 -4551 32132
rect -3145 32131 -3065 32133
rect -4447 32072 -4367 32074
rect -5155 32016 -4435 32072
rect -4379 32016 -4367 32072
rect -4447 32014 -4367 32016
rect -4118 32072 -4038 32074
rect -3851 32073 -3781 32084
rect -2961 32073 -2881 32075
rect -3851 32072 -2949 32073
rect -4118 32016 -4106 32072
rect -4050 32016 -3849 32072
rect -3793 32017 -2949 32072
rect -2893 32017 -2881 32073
rect -3793 32016 -3533 32017
rect -4118 32014 -4038 32016
rect -3851 32006 -3781 32016
rect -2961 32015 -2881 32017
rect -2632 32073 -2552 32075
rect -2189 32073 -2119 32083
rect -2632 32017 -2620 32073
rect -2564 32017 -2187 32073
rect -2131 32017 -2119 32073
rect -2632 32015 -2552 32017
rect -2189 32005 -2119 32017
rect -10921 31362 -10317 31969
rect -12288 31114 -10317 31362
rect -12288 28819 -12030 31114
rect -10921 30549 -10317 31114
rect -9986 31829 -9940 31840
rect -9771 31838 -9675 31869
rect -9771 31792 -9760 31838
rect -9686 31792 -9675 31838
rect -9506 31829 -9052 31969
rect -9848 31746 -9802 31757
rect -9865 31462 -9848 31472
rect -9644 31746 -9506 31757
rect -9802 31462 -9785 31472
rect -9865 31222 -9853 31462
rect -9797 31222 -9785 31462
rect -9865 31212 -9848 31222
rect -9802 31212 -9785 31222
rect -9848 31161 -9802 31172
rect -9598 31172 -9506 31746
rect -9644 31161 -9506 31172
rect -9986 31078 -9940 31089
rect -9771 31080 -9760 31126
rect -9686 31080 -9675 31126
rect -10211 31005 -10131 31015
rect -10211 30949 -10199 31005
rect -10143 30949 -10131 31005
rect -10211 30939 -10131 30949
rect -9771 31005 -9675 31080
rect -9460 31161 -9098 31829
rect -9506 31078 -9460 31089
rect -8883 31838 -8787 31869
rect -8883 31792 -8872 31838
rect -8798 31792 -8787 31838
rect -8618 31829 -8572 31969
rect -9052 31746 -8914 31757
rect -9052 31172 -8960 31746
rect -8756 31746 -8710 31757
rect -8773 31462 -8756 31472
rect -8710 31462 -8693 31472
rect -8773 31222 -8761 31462
rect -8705 31222 -8693 31462
rect -8773 31212 -8756 31222
rect -9052 31161 -8914 31172
rect -8710 31212 -8693 31222
rect -8756 31161 -8710 31172
rect -9098 31078 -9052 31089
rect -8883 31080 -8872 31126
rect -8798 31080 -8787 31126
rect -9771 30949 -9751 31005
rect -9695 30949 -9675 31005
rect -9771 30731 -9675 30949
rect -8883 30861 -8787 31080
rect -8403 31838 -8307 31869
rect -8403 31792 -8392 31838
rect -8318 31792 -8307 31838
rect -8138 31829 -8092 31969
rect -8572 31746 -8434 31757
rect -8572 31172 -8480 31746
rect -8276 31746 -8230 31757
rect -8293 31462 -8276 31472
rect -8230 31462 -8213 31472
rect -8293 31222 -8281 31462
rect -8225 31222 -8213 31462
rect -8293 31212 -8276 31222
rect -8572 31161 -8434 31172
rect -8230 31212 -8213 31222
rect -8276 31161 -8230 31172
rect -8618 31078 -8572 31089
rect -8403 31080 -8392 31126
rect -8318 31080 -8307 31126
rect -8403 30939 -8307 31080
rect -8138 31078 -8092 31089
rect -7795 31169 -6327 31969
rect -6027 31169 -5827 31969
rect -1445 31969 3645 32169
rect 4317 32072 4373 33319
rect 7273 33317 7353 33319
rect 13223 33376 13305 33388
rect 13789 33376 13845 34106
rect 14681 34104 14761 34106
rect 15411 34106 16179 34162
rect 16235 34106 16247 34162
rect 14313 34012 14393 34026
rect 14100 33990 14146 34001
rect 14313 33956 14325 34012
rect 14381 33956 14393 34012
rect 14497 34012 14577 34026
rect 14497 33956 14509 34012
rect 14565 33956 14577 34012
rect 14681 34012 14761 34026
rect 14681 33956 14693 34012
rect 14749 33956 14761 34012
rect 14928 33990 14974 34001
rect 14315 33953 14326 33956
rect 14380 33953 14391 33956
rect 14499 33953 14510 33956
rect 14564 33953 14575 33956
rect 14683 33953 14694 33956
rect 14748 33953 14759 33956
rect 14238 33907 14284 33918
rect 14146 33733 14238 33907
rect 14238 33722 14284 33733
rect 14422 33907 14468 33918
rect 14422 33722 14468 33733
rect 14606 33907 14652 33918
rect 14790 33907 14836 33918
rect 14773 33880 14790 33882
rect 14836 33880 14853 33882
rect 14773 33760 14785 33880
rect 14841 33760 14853 33880
rect 14773 33758 14790 33760
rect 14606 33722 14652 33733
rect 14836 33758 14853 33760
rect 14790 33722 14836 33733
rect 14100 33505 14146 33650
rect 14315 33641 14326 33687
rect 14380 33641 14391 33687
rect 14315 33608 14391 33641
rect 14499 33641 14510 33687
rect 14564 33641 14575 33687
rect 14499 33608 14575 33641
rect 14683 33641 14694 33687
rect 14748 33641 14759 33687
rect 14683 33608 14759 33641
rect 14928 33505 14974 33650
rect 14088 33493 14168 33505
rect 14088 33437 14100 33493
rect 14156 33437 14168 33493
rect 14088 33425 14168 33437
rect 14906 33493 14984 33505
rect 14906 33437 14918 33493
rect 14974 33437 14984 33493
rect 14906 33425 14984 33437
rect 13223 33320 13237 33376
rect 13293 33320 13845 33376
rect 15411 33376 15467 34106
rect 16167 34104 16247 34106
rect 23261 34106 24165 34162
rect 24221 34106 24233 34162
rect 15799 34012 15879 34026
rect 15586 33990 15632 34001
rect 15799 33956 15811 34012
rect 15867 33956 15879 34012
rect 15983 34012 16063 34026
rect 15983 33956 15995 34012
rect 16051 33956 16063 34012
rect 16167 34012 16247 34026
rect 16167 33956 16179 34012
rect 16235 33956 16247 34012
rect 16414 33990 16460 34001
rect 15801 33953 15812 33956
rect 15866 33953 15877 33956
rect 15985 33953 15996 33956
rect 16050 33953 16061 33956
rect 16169 33953 16180 33956
rect 16234 33953 16245 33956
rect 15724 33907 15770 33918
rect 15632 33733 15724 33907
rect 15724 33722 15770 33733
rect 15908 33907 15954 33918
rect 15908 33722 15954 33733
rect 16092 33907 16138 33918
rect 16276 33907 16322 33918
rect 16259 33880 16276 33882
rect 16322 33880 16339 33882
rect 16259 33760 16271 33880
rect 16327 33760 16339 33880
rect 16259 33758 16276 33760
rect 16092 33722 16138 33733
rect 16322 33758 16339 33760
rect 16276 33722 16322 33733
rect 15586 33505 15632 33650
rect 15801 33641 15812 33687
rect 15866 33641 15877 33687
rect 15801 33608 15877 33641
rect 15985 33641 15996 33687
rect 16050 33641 16061 33687
rect 15985 33608 16061 33641
rect 16169 33641 16180 33687
rect 16234 33641 16245 33687
rect 16169 33608 16245 33641
rect 16414 33505 16460 33650
rect 15574 33493 15654 33505
rect 15574 33437 15586 33493
rect 15642 33437 15654 33493
rect 15574 33425 15654 33437
rect 16392 33493 16470 33505
rect 16392 33437 16404 33493
rect 16460 33437 16470 33493
rect 16392 33425 16470 33437
rect 16745 33376 16825 33386
rect 15411 33320 16757 33376
rect 16813 33320 16825 33376
rect 13223 33308 13305 33320
rect 5797 33264 5867 33266
rect 7097 33265 7177 33267
rect 4453 33208 5799 33264
rect 5855 33208 5867 33264
rect 4453 32188 4509 33208
rect 5797 33196 5867 33208
rect 5939 33209 7109 33265
rect 7165 33209 7177 33265
rect 5117 33157 5203 33161
rect 5117 33101 5129 33157
rect 5185 33101 5203 33157
rect 5117 33089 5203 33101
rect 4628 32944 4674 32955
rect 4843 32953 4919 32986
rect 4843 32907 4854 32953
rect 4908 32907 4919 32953
rect 5027 32953 5103 32986
rect 5027 32907 5038 32953
rect 5092 32907 5103 32953
rect 5211 32953 5287 32986
rect 5211 32907 5222 32953
rect 5276 32907 5287 32953
rect 5456 32944 5502 32955
rect 4766 32861 4812 32872
rect 4749 32834 4766 32836
rect 4950 32861 4996 32872
rect 4812 32834 4829 32836
rect 4674 32714 4761 32834
rect 4817 32714 4829 32834
rect 4749 32712 4766 32714
rect 4674 32414 4766 32534
rect 4812 32712 4829 32714
rect 4933 32534 4950 32536
rect 5134 32861 5180 32872
rect 5117 32834 5134 32836
rect 5318 32861 5364 32872
rect 5180 32834 5197 32836
rect 5117 32714 5129 32834
rect 5185 32714 5197 32834
rect 5117 32712 5134 32714
rect 4996 32534 5013 32536
rect 4933 32414 4945 32534
rect 5001 32414 5013 32534
rect 4933 32412 4950 32414
rect 4766 32376 4812 32387
rect 4996 32412 5013 32414
rect 4950 32376 4996 32387
rect 5180 32712 5197 32714
rect 5301 32534 5318 32536
rect 5439 32834 5456 32836
rect 5502 32834 5519 32836
rect 5439 32713 5451 32834
rect 5507 32713 5519 32834
rect 5439 32711 5456 32713
rect 5364 32534 5381 32536
rect 5301 32414 5313 32534
rect 5369 32414 5381 32534
rect 5301 32412 5318 32414
rect 5134 32376 5180 32387
rect 5364 32412 5381 32414
rect 5318 32376 5364 32387
rect 4843 32338 4854 32341
rect 4908 32338 4919 32341
rect 5027 32338 5038 32341
rect 5092 32338 5103 32341
rect 5211 32338 5222 32341
rect 5276 32338 5287 32341
rect 4628 32293 4674 32304
rect 4841 32282 4853 32338
rect 4909 32282 4921 32338
rect 4841 32268 4921 32282
rect 5025 32282 5037 32338
rect 5093 32282 5105 32338
rect 5025 32268 5105 32282
rect 5209 32282 5221 32338
rect 5277 32282 5289 32338
rect 5502 32711 5519 32713
rect 5456 32293 5502 32304
rect 5209 32268 5289 32282
rect 4841 32188 4921 32190
rect 4453 32132 4853 32188
rect 4909 32132 4921 32188
rect 5939 32189 5995 33209
rect 7097 33197 7177 33209
rect 6603 33158 6689 33162
rect 6603 33102 6615 33158
rect 6671 33102 6689 33158
rect 6603 33090 6689 33102
rect 6114 32945 6160 32956
rect 6329 32954 6405 32987
rect 6329 32908 6340 32954
rect 6394 32908 6405 32954
rect 6513 32954 6589 32987
rect 6513 32908 6524 32954
rect 6578 32908 6589 32954
rect 6697 32954 6773 32987
rect 6697 32908 6708 32954
rect 6762 32908 6773 32954
rect 6942 32945 6988 32956
rect 6252 32862 6298 32873
rect 6235 32835 6252 32837
rect 6436 32862 6482 32873
rect 6298 32835 6315 32837
rect 6160 32715 6247 32835
rect 6303 32715 6315 32835
rect 6235 32713 6252 32715
rect 6160 32415 6252 32535
rect 6298 32713 6315 32715
rect 6419 32535 6436 32537
rect 6620 32862 6666 32873
rect 6603 32835 6620 32837
rect 6804 32862 6850 32873
rect 6666 32835 6683 32837
rect 6603 32715 6615 32835
rect 6671 32715 6683 32835
rect 6603 32713 6620 32715
rect 6482 32535 6499 32537
rect 6419 32415 6431 32535
rect 6487 32415 6499 32535
rect 6419 32413 6436 32415
rect 6252 32377 6298 32388
rect 6482 32413 6499 32415
rect 6436 32377 6482 32388
rect 6666 32713 6683 32715
rect 6787 32535 6804 32537
rect 6925 32835 6942 32837
rect 6988 32835 7005 32837
rect 6925 32714 6937 32835
rect 6993 32714 7005 32835
rect 6925 32712 6942 32714
rect 6850 32535 6867 32537
rect 6787 32415 6799 32535
rect 6855 32415 6867 32535
rect 6787 32413 6804 32415
rect 6620 32377 6666 32388
rect 6850 32413 6867 32415
rect 6804 32377 6850 32388
rect 6329 32339 6340 32342
rect 6394 32339 6405 32342
rect 6513 32339 6524 32342
rect 6578 32339 6589 32342
rect 6697 32339 6708 32342
rect 6762 32339 6773 32342
rect 6114 32294 6160 32305
rect 6327 32283 6339 32339
rect 6395 32283 6407 32339
rect 6327 32269 6407 32283
rect 6511 32283 6523 32339
rect 6579 32283 6591 32339
rect 6511 32269 6591 32283
rect 6695 32283 6707 32339
rect 6763 32283 6775 32339
rect 6988 32712 7005 32714
rect 6942 32294 6988 32305
rect 6695 32269 6775 32283
rect 6327 32189 6407 32191
rect 5939 32133 6339 32189
rect 6395 32133 6407 32189
rect 4841 32130 4921 32132
rect 6327 32131 6407 32133
rect 5025 32072 5105 32074
rect 4317 32016 5037 32072
rect 5093 32016 5105 32072
rect 5025 32014 5105 32016
rect 5354 32072 5434 32074
rect 5621 32073 5691 32084
rect 6511 32073 6591 32075
rect 5621 32072 6523 32073
rect 5354 32016 5366 32072
rect 5422 32016 5623 32072
rect 5679 32017 6523 32072
rect 6579 32017 6591 32073
rect 5679 32016 5939 32017
rect 5354 32014 5434 32016
rect 5621 32006 5691 32016
rect 6511 32015 6591 32017
rect 6840 32073 6920 32075
rect 7283 32073 7353 32083
rect 6840 32017 6852 32073
rect 6908 32017 7285 32073
rect 7341 32017 7353 32073
rect 6840 32015 6920 32017
rect 7283 32005 7353 32017
rect -5303 31956 -5233 31968
rect -4263 31956 -4183 31958
rect -2777 31957 -2697 31959
rect -5303 31900 -5291 31956
rect -5235 31900 -4251 31956
rect -4195 31900 -4183 31956
rect -5303 31888 -5233 31900
rect -8951 30849 -8787 30861
rect -8471 30927 -8307 30939
rect -8471 30871 -8459 30927
rect -8403 30871 -8307 30927
rect -8471 30859 -8307 30871
rect -8951 30793 -8939 30849
rect -8883 30793 -8787 30849
rect -8951 30781 -8787 30793
rect -8883 30731 -8787 30781
rect -9986 30709 -9940 30720
rect -10880 30409 -10834 30549
rect -10665 30418 -10569 30449
rect -10665 30372 -10654 30418
rect -10580 30372 -10569 30418
rect -10400 30409 -10354 30549
rect -10834 30326 -10696 30337
rect -10834 29752 -10742 30326
rect -10538 30326 -10492 30337
rect -10555 30042 -10538 30052
rect -10492 30042 -10475 30052
rect -10555 29802 -10543 30042
rect -10487 29802 -10475 30042
rect -10555 29792 -10538 29802
rect -10834 29741 -10696 29752
rect -10492 29792 -10475 29802
rect -10538 29741 -10492 29752
rect -10880 29658 -10834 29669
rect -10665 29660 -10654 29706
rect -10580 29660 -10569 29706
rect -10665 29519 -10569 29660
rect -9771 30718 -9471 30731
rect -9771 30672 -9760 30718
rect -9686 30685 -9556 30718
rect -9686 30672 -9675 30685
rect -9567 30672 -9556 30685
rect -9482 30672 -9471 30718
rect -9302 30709 -9256 30720
rect -9940 30626 -9802 30637
rect -9940 30452 -9848 30626
rect -9644 30626 -9598 30637
rect -9661 30567 -9644 30577
rect -9440 30626 -9302 30637
rect -9598 30567 -9581 30577
rect -9661 30511 -9649 30567
rect -9593 30511 -9581 30567
rect -9661 30501 -9644 30511
rect -9940 30441 -9802 30452
rect -9598 30501 -9581 30511
rect -9644 30441 -9598 30452
rect -9394 30452 -9302 30626
rect -9440 30441 -9302 30452
rect -9986 30229 -9940 30369
rect -9771 30360 -9760 30406
rect -9686 30360 -9675 30406
rect -9771 30329 -9675 30360
rect -9567 30360 -9556 30406
rect -9482 30360 -9471 30406
rect -9567 30329 -9471 30360
rect -9087 30718 -8787 30731
rect -9087 30672 -9076 30718
rect -9002 30685 -8872 30718
rect -9002 30672 -8991 30685
rect -8883 30672 -8872 30685
rect -8798 30672 -8787 30718
rect -8618 30709 -8572 30720
rect -9164 30626 -9118 30637
rect -9181 30567 -9164 30577
rect -8960 30626 -8914 30637
rect -9118 30567 -9101 30577
rect -9181 30511 -9169 30567
rect -9113 30511 -9101 30567
rect -9181 30501 -9164 30511
rect -9118 30501 -9101 30511
rect -8977 30567 -8960 30577
rect -8756 30626 -8710 30637
rect -8914 30567 -8897 30577
rect -8977 30511 -8965 30567
rect -8909 30511 -8897 30567
rect -8977 30501 -8960 30511
rect -9164 30441 -9118 30452
rect -8914 30501 -8897 30511
rect -8773 30567 -8756 30577
rect -8710 30567 -8693 30577
rect -8773 30511 -8761 30567
rect -8705 30511 -8693 30567
rect -8773 30501 -8756 30511
rect -8960 30441 -8914 30452
rect -8710 30501 -8693 30511
rect -8756 30441 -8710 30452
rect -9302 30229 -9256 30369
rect -9087 30360 -9076 30406
rect -9002 30360 -8991 30406
rect -9087 30329 -8991 30360
rect -8883 30360 -8872 30406
rect -8798 30360 -8787 30406
rect -8883 30329 -8787 30360
rect -8403 30718 -8307 30859
rect -7795 30973 -5827 31169
rect -5019 31169 -4963 31900
rect -4263 31898 -4183 31900
rect -3533 31901 -2765 31957
rect -2709 31901 -2697 31957
rect -4631 31806 -4551 31820
rect -4844 31784 -4798 31795
rect -4631 31750 -4619 31806
rect -4563 31750 -4551 31806
rect -4447 31806 -4367 31820
rect -4447 31750 -4435 31806
rect -4379 31750 -4367 31806
rect -4263 31806 -4183 31820
rect -4263 31750 -4251 31806
rect -4195 31750 -4183 31806
rect -4016 31784 -3970 31795
rect -4629 31747 -4618 31750
rect -4564 31747 -4553 31750
rect -4445 31747 -4434 31750
rect -4380 31747 -4369 31750
rect -4261 31747 -4250 31750
rect -4196 31747 -4185 31750
rect -4706 31701 -4660 31712
rect -4798 31527 -4706 31701
rect -4706 31516 -4660 31527
rect -4522 31701 -4476 31712
rect -4522 31516 -4476 31527
rect -4338 31701 -4292 31712
rect -4154 31701 -4108 31712
rect -4171 31674 -4154 31676
rect -4108 31674 -4091 31676
rect -4171 31554 -4159 31674
rect -4103 31554 -4091 31674
rect -4171 31552 -4154 31554
rect -4338 31516 -4292 31527
rect -4108 31552 -4091 31554
rect -4154 31516 -4108 31527
rect -4844 31299 -4798 31444
rect -4629 31435 -4618 31481
rect -4564 31435 -4553 31481
rect -4629 31402 -4553 31435
rect -4445 31435 -4434 31481
rect -4380 31435 -4369 31481
rect -4445 31402 -4369 31435
rect -4261 31435 -4250 31481
rect -4196 31435 -4185 31481
rect -4261 31402 -4185 31435
rect -4016 31299 -3970 31444
rect -4856 31287 -4776 31299
rect -4856 31231 -4844 31287
rect -4788 31231 -4776 31287
rect -4856 31219 -4776 31231
rect -4038 31287 -3960 31299
rect -4038 31231 -4026 31287
rect -3970 31231 -3960 31287
rect -4038 31219 -3960 31231
rect -3685 31169 -3605 31179
rect -5019 31113 -3673 31169
rect -3617 31113 -3605 31169
rect -3685 31111 -3605 31113
rect -3851 31060 -3781 31062
rect -7795 30833 -7695 30973
rect -5927 30833 -5827 30973
rect -7795 30793 -5827 30833
rect -5019 31059 -3781 31060
rect -5019 31005 -3849 31059
rect -3793 31005 -3781 31059
rect -5019 31004 -3781 31005
rect -8403 30672 -8392 30718
rect -8318 30672 -8307 30718
rect -8138 30709 -8092 30720
rect -8572 30626 -8434 30637
rect -8572 30452 -8480 30626
rect -8276 30626 -8230 30637
rect -8293 30567 -8276 30577
rect -8230 30567 -8213 30577
rect -8293 30511 -8281 30567
rect -8225 30511 -8213 30567
rect -8293 30501 -8276 30511
rect -8572 30441 -8434 30452
rect -8230 30501 -8213 30511
rect -8276 30441 -8230 30452
rect -8618 30229 -8572 30369
rect -8403 30360 -8392 30406
rect -8318 30360 -8307 30406
rect -8403 30329 -8307 30360
rect -8138 30229 -8092 30369
rect -7758 30653 -7712 30793
rect -10023 30199 -8055 30229
rect -10023 30166 -8755 30199
rect -10023 30090 -9985 30166
rect -9905 30090 -8755 30166
rect -10023 30059 -8755 30090
rect -8155 30059 -8055 30199
rect -10023 30029 -8055 30059
rect -7543 30662 -7447 30693
rect -7543 30616 -7532 30662
rect -7458 30616 -7447 30662
rect -7339 30662 -7243 30693
rect -7339 30616 -7328 30662
rect -7254 30616 -7243 30662
rect -7074 30653 -7028 30793
rect -7712 30570 -7574 30581
rect -7416 30570 -7370 30581
rect -7212 30570 -7074 30581
rect -7712 29996 -7620 30570
rect -7433 30330 -7421 30570
rect -7365 30330 -7353 30570
rect -7712 29985 -7574 29996
rect -7416 29985 -7370 29996
rect -7166 29996 -7074 30570
rect -7212 29985 -7074 29996
rect -7758 29902 -7712 29913
rect -7543 29904 -7532 29950
rect -7458 29930 -7447 29950
rect -7339 29930 -7328 29950
rect -7458 29904 -7328 29930
rect -7254 29904 -7243 29950
rect -7543 29877 -7243 29904
rect -6859 30662 -6763 30693
rect -6859 30616 -6848 30662
rect -6774 30616 -6763 30662
rect -6655 30662 -6559 30693
rect -6655 30616 -6644 30662
rect -6570 30616 -6559 30662
rect -6390 30653 -6344 30793
rect -6936 30570 -6890 30581
rect -6732 30570 -6686 30581
rect -6528 30570 -6482 30581
rect -6749 30330 -6737 30570
rect -6681 30330 -6669 30570
rect -6953 29996 -6941 30236
rect -6885 29996 -6873 30236
rect -6545 29996 -6533 30236
rect -6477 29996 -6465 30236
rect -6936 29985 -6890 29996
rect -6732 29985 -6686 29996
rect -6528 29985 -6482 29996
rect -7074 29902 -7028 29913
rect -6859 29904 -6848 29950
rect -6774 29930 -6763 29950
rect -6655 29930 -6644 29950
rect -6774 29904 -6644 29930
rect -6570 29904 -6559 29950
rect -6859 29877 -6559 29904
rect -6175 30662 -6079 30693
rect -6175 30616 -6164 30662
rect -6090 30616 -6079 30662
rect -5910 30653 -5864 30793
rect -6344 30570 -6206 30581
rect -6344 29996 -6252 30570
rect -6048 30570 -6002 30581
rect -6065 30286 -6048 30296
rect -6002 30286 -5985 30296
rect -6065 30046 -6053 30286
rect -5997 30046 -5985 30286
rect -6065 30036 -6048 30046
rect -6344 29985 -6206 29996
rect -6002 30036 -5985 30046
rect -6048 29985 -6002 29996
rect -6390 29902 -6344 29913
rect -6175 29904 -6164 29950
rect -6090 29904 -6079 29950
rect -7543 29829 -7447 29877
rect -10400 29658 -10354 29669
rect -10023 29799 -8055 29829
rect -10023 29659 -8755 29799
rect -8155 29659 -8055 29799
rect -10023 29629 -8055 29659
rect -7543 29773 -7523 29829
rect -7467 29773 -7447 29829
rect -10733 29507 -10569 29519
rect -10733 29451 -10721 29507
rect -10665 29451 -10569 29507
rect -10733 29439 -10569 29451
rect -12630 28619 -12030 28819
rect -10880 29289 -10834 29300
rect -10665 29298 -10569 29439
rect -9986 29489 -9940 29500
rect -10665 29252 -10654 29298
rect -10580 29252 -10569 29298
rect -10400 29289 -10354 29300
rect -10834 29206 -10696 29217
rect -10834 29032 -10742 29206
rect -10538 29206 -10492 29217
rect -10555 29147 -10538 29157
rect -10492 29147 -10475 29157
rect -10555 29091 -10543 29147
rect -10487 29091 -10475 29147
rect -10555 29081 -10538 29091
rect -10834 29021 -10696 29032
rect -10492 29081 -10475 29091
rect -10538 29021 -10492 29032
rect -10880 28809 -10834 28949
rect -10665 28940 -10654 28986
rect -10580 28940 -10569 28986
rect -10665 28909 -10569 28940
rect -10400 28809 -10354 28949
rect -12593 28479 -12547 28619
rect -12378 28488 -12282 28519
rect -12378 28442 -12367 28488
rect -12293 28442 -12282 28488
rect -12113 28479 -12067 28619
rect -12547 28396 -12409 28407
rect -12547 27822 -12455 28396
rect -12251 28396 -12205 28407
rect -12268 28112 -12251 28122
rect -12205 28112 -12188 28122
rect -12268 27872 -12256 28112
rect -12200 27872 -12188 28112
rect -12268 27862 -12251 27872
rect -12547 27811 -12409 27822
rect -12205 27862 -12188 27872
rect -12251 27811 -12205 27822
rect -12593 27728 -12547 27739
rect -12378 27730 -12367 27776
rect -12293 27730 -12282 27776
rect -12378 27589 -12282 27730
rect -12113 27728 -12067 27739
rect -10921 27889 -10317 28809
rect -9771 29498 -9675 29529
rect -9771 29452 -9760 29498
rect -9686 29452 -9675 29498
rect -9506 29489 -9052 29629
rect -9848 29406 -9802 29417
rect -9865 29122 -9848 29132
rect -9644 29406 -9506 29417
rect -9802 29122 -9785 29132
rect -9865 28882 -9853 29122
rect -9797 28882 -9785 29122
rect -9865 28872 -9848 28882
rect -9802 28872 -9785 28882
rect -9848 28821 -9802 28832
rect -9598 28832 -9506 29406
rect -9644 28821 -9506 28832
rect -9986 28738 -9940 28749
rect -9771 28740 -9760 28786
rect -9686 28740 -9675 28786
rect -9771 28665 -9675 28740
rect -9460 28821 -9098 29489
rect -9506 28738 -9460 28749
rect -8883 29498 -8787 29529
rect -8883 29452 -8872 29498
rect -8798 29452 -8787 29498
rect -8618 29489 -8572 29629
rect -9052 29406 -8914 29417
rect -9052 28832 -8960 29406
rect -8756 29406 -8710 29417
rect -8773 29122 -8756 29132
rect -8710 29122 -8693 29132
rect -8773 28882 -8761 29122
rect -8705 28882 -8693 29122
rect -8773 28872 -8756 28882
rect -9052 28821 -8914 28832
rect -8710 28872 -8693 28882
rect -8756 28821 -8710 28832
rect -9098 28738 -9052 28749
rect -8883 28740 -8872 28786
rect -8798 28740 -8787 28786
rect -9771 28609 -9751 28665
rect -9695 28609 -9675 28665
rect -9771 28391 -9675 28609
rect -8883 28521 -8787 28740
rect -8403 29498 -8307 29529
rect -8403 29452 -8392 29498
rect -8318 29452 -8307 29498
rect -8138 29489 -8092 29629
rect -8572 29406 -8434 29417
rect -8572 28832 -8480 29406
rect -8276 29406 -8230 29417
rect -8293 29122 -8276 29132
rect -8230 29122 -8213 29132
rect -8293 28882 -8281 29122
rect -8225 28882 -8213 29122
rect -8293 28872 -8276 28882
rect -8572 28821 -8434 28832
rect -8230 28872 -8213 28882
rect -8276 28821 -8230 28832
rect -8618 28738 -8572 28749
rect -8403 28740 -8392 28786
rect -8318 28740 -8307 28786
rect -8403 28599 -8307 28740
rect -7758 29533 -7712 29544
rect -7543 29542 -7447 29773
rect -6859 29673 -6763 29877
rect -6175 29763 -6079 29904
rect -5019 29983 -4963 31004
rect -3851 30996 -3781 31004
rect -4355 30952 -4269 30956
rect -4355 30896 -4343 30952
rect -4287 30896 -4269 30952
rect -4355 30884 -4269 30896
rect -4844 30739 -4798 30750
rect -4629 30748 -4553 30781
rect -4629 30702 -4618 30748
rect -4564 30702 -4553 30748
rect -4445 30748 -4369 30781
rect -4445 30702 -4434 30748
rect -4380 30702 -4369 30748
rect -4261 30748 -4185 30781
rect -4261 30702 -4250 30748
rect -4196 30702 -4185 30748
rect -4016 30739 -3970 30750
rect -4706 30656 -4660 30667
rect -4723 30629 -4706 30631
rect -4522 30656 -4476 30667
rect -4660 30629 -4643 30631
rect -4798 30509 -4711 30629
rect -4655 30509 -4643 30629
rect -4723 30507 -4706 30509
rect -4798 30209 -4706 30329
rect -4660 30507 -4643 30509
rect -4539 30329 -4522 30331
rect -4338 30656 -4292 30667
rect -4355 30629 -4338 30631
rect -4154 30656 -4108 30667
rect -4292 30629 -4275 30631
rect -4355 30509 -4343 30629
rect -4287 30509 -4275 30629
rect -4355 30507 -4338 30509
rect -4476 30329 -4459 30331
rect -4539 30209 -4527 30329
rect -4471 30209 -4459 30329
rect -4539 30207 -4522 30209
rect -4706 30171 -4660 30182
rect -4476 30207 -4459 30209
rect -4522 30171 -4476 30182
rect -4292 30507 -4275 30509
rect -4171 30329 -4154 30331
rect -4033 30629 -4016 30631
rect -3970 30629 -3953 30631
rect -4033 30508 -4021 30629
rect -3965 30508 -3953 30629
rect -4033 30506 -4016 30508
rect -4108 30329 -4091 30331
rect -4171 30209 -4159 30329
rect -4103 30209 -4091 30329
rect -4171 30207 -4154 30209
rect -4338 30171 -4292 30182
rect -4108 30207 -4091 30209
rect -4154 30171 -4108 30182
rect -4629 30133 -4618 30136
rect -4564 30133 -4553 30136
rect -4445 30133 -4434 30136
rect -4380 30133 -4369 30136
rect -4261 30133 -4250 30136
rect -4196 30133 -4185 30136
rect -4844 30088 -4798 30099
rect -4631 30077 -4619 30133
rect -4563 30077 -4551 30133
rect -4631 30063 -4551 30077
rect -4447 30077 -4435 30133
rect -4379 30077 -4367 30133
rect -4447 30063 -4367 30077
rect -4263 30077 -4251 30133
rect -4195 30077 -4183 30133
rect -3970 30506 -3953 30508
rect -4016 30088 -3970 30099
rect -4263 30063 -4183 30077
rect -4631 29983 -4551 29985
rect -5019 29927 -4619 29983
rect -4563 29927 -4551 29983
rect -4631 29925 -4551 29927
rect -5910 29902 -5864 29913
rect -5439 29867 -5369 29881
rect -4447 29867 -4367 29869
rect -5439 29811 -5427 29867
rect -5371 29811 -4435 29867
rect -4379 29811 -4367 29867
rect -5439 29799 -5369 29811
rect -4447 29809 -4367 29811
rect -4118 29867 -4038 29869
rect -3675 29867 -3615 29879
rect -4118 29811 -4106 29867
rect -4050 29811 -3673 29867
rect -3617 29811 -3615 29867
rect -4118 29809 -4038 29811
rect -3675 29799 -3615 29811
rect -6243 29751 -6079 29763
rect -6243 29695 -6231 29751
rect -6175 29695 -6079 29751
rect -6243 29683 -6079 29695
rect -5673 29751 -5595 29762
rect -4263 29751 -4183 29753
rect -5673 29750 -4251 29751
rect -5673 29696 -5661 29750
rect -5607 29696 -4251 29750
rect -5673 29695 -4251 29696
rect -4195 29695 -4183 29751
rect -5673 29684 -5595 29695
rect -4263 29693 -4183 29695
rect -6859 29617 -6839 29673
rect -6783 29617 -6763 29673
rect -7543 29496 -7532 29542
rect -7458 29496 -7447 29542
rect -7278 29533 -7028 29544
rect -7620 29450 -7574 29461
rect -7637 29391 -7620 29401
rect -7416 29450 -7278 29461
rect -7574 29391 -7557 29401
rect -7637 29335 -7625 29391
rect -7569 29335 -7557 29391
rect -7637 29325 -7620 29335
rect -7574 29325 -7557 29335
rect -7620 29265 -7574 29276
rect -7370 29276 -7278 29450
rect -7416 29265 -7278 29276
rect -7758 29053 -7712 29193
rect -7543 29184 -7532 29230
rect -7458 29184 -7447 29230
rect -7543 29153 -7447 29184
rect -7232 29193 -7074 29533
rect -6859 29542 -6763 29617
rect -6859 29496 -6848 29542
rect -6774 29496 -6763 29542
rect -6594 29533 -6548 29544
rect -7028 29450 -6890 29461
rect -7028 29276 -6936 29450
rect -6732 29450 -6686 29461
rect -6749 29391 -6732 29401
rect -6686 29391 -6669 29401
rect -6749 29335 -6737 29391
rect -6681 29335 -6669 29391
rect -6749 29325 -6732 29335
rect -7028 29265 -6890 29276
rect -6686 29325 -6669 29335
rect -6732 29265 -6686 29276
rect -7278 29182 -7028 29193
rect -6859 29184 -6848 29230
rect -6774 29184 -6763 29230
rect -7232 29053 -7074 29182
rect -6859 29153 -6763 29184
rect -6594 29053 -6548 29193
rect -6390 29533 -6344 29544
rect -6175 29542 -6079 29683
rect -4631 29601 -4551 29615
rect -4844 29579 -4798 29590
rect -6175 29496 -6164 29542
rect -6090 29496 -6079 29542
rect -5910 29533 -5864 29544
rect -6344 29450 -6206 29461
rect -6344 29276 -6252 29450
rect -6048 29450 -6002 29461
rect -6065 29391 -6048 29401
rect -6002 29391 -5985 29401
rect -6065 29335 -6053 29391
rect -5997 29335 -5985 29391
rect -6065 29325 -6048 29335
rect -6344 29265 -6206 29276
rect -6002 29325 -5985 29335
rect -6048 29265 -6002 29276
rect -6390 29053 -6344 29193
rect -6175 29184 -6164 29230
rect -6090 29184 -6079 29230
rect -6175 29153 -6079 29184
rect -5910 29053 -5864 29193
rect -4631 29545 -4619 29601
rect -4563 29545 -4551 29601
rect -4447 29601 -4367 29615
rect -4447 29545 -4435 29601
rect -4379 29545 -4367 29601
rect -4263 29601 -4183 29615
rect -4263 29545 -4251 29601
rect -4195 29545 -4183 29601
rect -4016 29579 -3970 29590
rect -4629 29542 -4618 29545
rect -4564 29542 -4553 29545
rect -4445 29542 -4434 29545
rect -4380 29542 -4369 29545
rect -4261 29542 -4250 29545
rect -4196 29542 -4185 29545
rect -4706 29496 -4660 29507
rect -4798 29322 -4706 29496
rect -4706 29311 -4660 29322
rect -4522 29496 -4476 29507
rect -4522 29311 -4476 29322
rect -4338 29496 -4292 29507
rect -4154 29496 -4108 29507
rect -4171 29469 -4154 29471
rect -4108 29469 -4091 29471
rect -4171 29349 -4159 29469
rect -4103 29349 -4091 29469
rect -4171 29347 -4154 29349
rect -4338 29311 -4292 29322
rect -4108 29347 -4091 29349
rect -4154 29311 -4108 29322
rect -4844 29094 -4798 29239
rect -4629 29230 -4618 29276
rect -4564 29230 -4553 29276
rect -4629 29197 -4553 29230
rect -4445 29230 -4434 29276
rect -4380 29230 -4369 29276
rect -4445 29197 -4369 29230
rect -4261 29230 -4250 29276
rect -4196 29230 -4185 29276
rect -4261 29197 -4185 29230
rect -4016 29094 -3970 29239
rect -4856 29082 -4776 29094
rect -8138 28738 -8092 28749
rect -7795 29013 -5827 29053
rect -4856 29026 -4844 29082
rect -4788 29026 -4776 29082
rect -4856 29014 -4776 29026
rect -4038 29082 -3958 29094
rect -4038 29026 -4026 29082
rect -3970 29026 -3958 29082
rect -4038 29014 -3958 29026
rect -7795 28873 -7695 29013
rect -5927 28873 -5827 29013
rect -5622 28964 -5536 28976
rect -5429 28964 -5369 28968
rect -3533 28964 -3477 31901
rect -2777 31899 -2697 31901
rect -3145 31807 -3065 31821
rect -3358 31785 -3312 31796
rect -3145 31751 -3133 31807
rect -3077 31751 -3065 31807
rect -2961 31807 -2881 31821
rect -2961 31751 -2949 31807
rect -2893 31751 -2881 31807
rect -2777 31807 -2697 31821
rect -2777 31751 -2765 31807
rect -2709 31751 -2697 31807
rect -2530 31785 -2484 31796
rect -3143 31748 -3132 31751
rect -3078 31748 -3067 31751
rect -2959 31748 -2948 31751
rect -2894 31748 -2883 31751
rect -2775 31748 -2764 31751
rect -2710 31748 -2699 31751
rect -3220 31702 -3174 31713
rect -3312 31528 -3220 31702
rect -3220 31517 -3174 31528
rect -3036 31702 -2990 31713
rect -3036 31517 -2990 31528
rect -2852 31702 -2806 31713
rect -2668 31702 -2622 31713
rect -2685 31675 -2668 31677
rect -2622 31675 -2605 31677
rect -2685 31555 -2673 31675
rect -2617 31555 -2605 31675
rect -2685 31553 -2668 31555
rect -2852 31517 -2806 31528
rect -2622 31553 -2605 31555
rect -2668 31517 -2622 31528
rect -3358 31300 -3312 31445
rect -3143 31436 -3132 31482
rect -3078 31436 -3067 31482
rect -3143 31403 -3067 31436
rect -2959 31436 -2948 31482
rect -2894 31436 -2883 31482
rect -2959 31403 -2883 31436
rect -2775 31436 -2764 31482
rect -2710 31436 -2699 31482
rect -2775 31403 -2699 31436
rect -2530 31300 -2484 31445
rect -3370 31288 -3290 31300
rect -3370 31232 -3358 31288
rect -3302 31232 -3290 31288
rect -3370 31220 -3290 31232
rect -2552 31288 -2474 31300
rect -2552 31232 -2540 31288
rect -2484 31232 -2474 31288
rect -2552 31220 -2474 31232
rect -1445 31169 -1245 31969
rect -1045 31169 -845 31969
rect -1445 30549 -845 31169
rect -514 31829 -468 31840
rect -299 31838 -203 31869
rect -299 31792 -288 31838
rect -214 31792 -203 31838
rect -34 31829 420 31969
rect -376 31746 -330 31757
rect -393 31462 -376 31472
rect -172 31746 -34 31757
rect -330 31462 -313 31472
rect -393 31222 -381 31462
rect -325 31222 -313 31462
rect -393 31212 -376 31222
rect -330 31212 -313 31222
rect -376 31161 -330 31172
rect -126 31172 -34 31746
rect -172 31161 -34 31172
rect -514 31078 -468 31089
rect -299 31080 -288 31126
rect -214 31080 -203 31126
rect -299 31005 -203 31080
rect 12 31161 374 31829
rect -34 31078 12 31089
rect 589 31838 685 31869
rect 589 31792 600 31838
rect 674 31792 685 31838
rect 854 31829 900 31969
rect 420 31746 558 31757
rect 420 31172 512 31746
rect 716 31746 762 31757
rect 699 31462 716 31472
rect 762 31462 779 31472
rect 699 31222 711 31462
rect 767 31222 779 31462
rect 699 31212 716 31222
rect 420 31161 558 31172
rect 762 31212 779 31222
rect 716 31161 762 31172
rect 374 31078 420 31089
rect 589 31080 600 31126
rect 674 31080 685 31126
rect -299 30949 -279 31005
rect -223 30949 -203 31005
rect -299 30731 -203 30949
rect 589 30861 685 31080
rect 1069 31838 1165 31869
rect 1069 31792 1080 31838
rect 1154 31792 1165 31838
rect 1334 31829 1380 31969
rect 900 31746 1038 31757
rect 900 31172 992 31746
rect 1196 31746 1242 31757
rect 1179 31462 1196 31472
rect 1242 31462 1259 31472
rect 1179 31222 1191 31462
rect 1247 31222 1259 31462
rect 1179 31212 1196 31222
rect 900 31161 1038 31172
rect 1242 31212 1259 31222
rect 1196 31161 1242 31172
rect 854 31078 900 31089
rect 1069 31080 1080 31126
rect 1154 31080 1165 31126
rect 1069 30939 1165 31080
rect 1334 31078 1380 31089
rect 1677 31169 3145 31969
rect 3445 31169 3645 31969
rect 8027 31970 13117 32170
rect 13789 32073 13845 33320
rect 16745 33318 16825 33320
rect 22695 33376 22777 33388
rect 23261 33376 23317 34106
rect 24153 34104 24233 34106
rect 24883 34106 25651 34162
rect 25707 34106 25719 34162
rect 23785 34012 23865 34026
rect 23572 33990 23618 34001
rect 23785 33956 23797 34012
rect 23853 33956 23865 34012
rect 23969 34012 24049 34026
rect 23969 33956 23981 34012
rect 24037 33956 24049 34012
rect 24153 34012 24233 34026
rect 24153 33956 24165 34012
rect 24221 33956 24233 34012
rect 24400 33990 24446 34001
rect 23787 33953 23798 33956
rect 23852 33953 23863 33956
rect 23971 33953 23982 33956
rect 24036 33953 24047 33956
rect 24155 33953 24166 33956
rect 24220 33953 24231 33956
rect 23710 33907 23756 33918
rect 23618 33733 23710 33907
rect 23710 33722 23756 33733
rect 23894 33907 23940 33918
rect 23894 33722 23940 33733
rect 24078 33907 24124 33918
rect 24262 33907 24308 33918
rect 24245 33880 24262 33882
rect 24308 33880 24325 33882
rect 24245 33760 24257 33880
rect 24313 33760 24325 33880
rect 24245 33758 24262 33760
rect 24078 33722 24124 33733
rect 24308 33758 24325 33760
rect 24262 33722 24308 33733
rect 23572 33505 23618 33650
rect 23787 33641 23798 33687
rect 23852 33641 23863 33687
rect 23787 33608 23863 33641
rect 23971 33641 23982 33687
rect 24036 33641 24047 33687
rect 23971 33608 24047 33641
rect 24155 33641 24166 33687
rect 24220 33641 24231 33687
rect 24155 33608 24231 33641
rect 24400 33505 24446 33650
rect 23560 33493 23640 33505
rect 23560 33437 23572 33493
rect 23628 33437 23640 33493
rect 23560 33425 23640 33437
rect 24378 33493 24456 33505
rect 24378 33437 24390 33493
rect 24446 33437 24456 33493
rect 24378 33425 24456 33437
rect 22695 33320 22709 33376
rect 22765 33320 23317 33376
rect 24883 33376 24939 34106
rect 25639 34104 25719 34106
rect 32733 34106 33637 34162
rect 33693 34106 33705 34162
rect 25271 34012 25351 34026
rect 25058 33990 25104 34001
rect 25271 33956 25283 34012
rect 25339 33956 25351 34012
rect 25455 34012 25535 34026
rect 25455 33956 25467 34012
rect 25523 33956 25535 34012
rect 25639 34012 25719 34026
rect 25639 33956 25651 34012
rect 25707 33956 25719 34012
rect 25886 33990 25932 34001
rect 25273 33953 25284 33956
rect 25338 33953 25349 33956
rect 25457 33953 25468 33956
rect 25522 33953 25533 33956
rect 25641 33953 25652 33956
rect 25706 33953 25717 33956
rect 25196 33907 25242 33918
rect 25104 33733 25196 33907
rect 25196 33722 25242 33733
rect 25380 33907 25426 33918
rect 25380 33722 25426 33733
rect 25564 33907 25610 33918
rect 25748 33907 25794 33918
rect 25731 33880 25748 33882
rect 25794 33880 25811 33882
rect 25731 33760 25743 33880
rect 25799 33760 25811 33880
rect 25731 33758 25748 33760
rect 25564 33722 25610 33733
rect 25794 33758 25811 33760
rect 25748 33722 25794 33733
rect 25058 33505 25104 33650
rect 25273 33641 25284 33687
rect 25338 33641 25349 33687
rect 25273 33608 25349 33641
rect 25457 33641 25468 33687
rect 25522 33641 25533 33687
rect 25457 33608 25533 33641
rect 25641 33641 25652 33687
rect 25706 33641 25717 33687
rect 25641 33608 25717 33641
rect 25886 33505 25932 33650
rect 25046 33493 25126 33505
rect 25046 33437 25058 33493
rect 25114 33437 25126 33493
rect 25046 33425 25126 33437
rect 25864 33493 25942 33505
rect 25864 33437 25876 33493
rect 25932 33437 25942 33493
rect 25864 33425 25942 33437
rect 26217 33376 26297 33386
rect 24883 33320 26229 33376
rect 26285 33320 26297 33376
rect 22695 33308 22777 33320
rect 15269 33265 15339 33267
rect 16569 33266 16649 33268
rect 13925 33209 15271 33265
rect 15327 33209 15339 33265
rect 13925 32189 13981 33209
rect 15269 33197 15339 33209
rect 15411 33210 16581 33266
rect 16637 33210 16649 33266
rect 14589 33158 14675 33162
rect 14589 33102 14601 33158
rect 14657 33102 14675 33158
rect 14589 33090 14675 33102
rect 14100 32945 14146 32956
rect 14315 32954 14391 32987
rect 14315 32908 14326 32954
rect 14380 32908 14391 32954
rect 14499 32954 14575 32987
rect 14499 32908 14510 32954
rect 14564 32908 14575 32954
rect 14683 32954 14759 32987
rect 14683 32908 14694 32954
rect 14748 32908 14759 32954
rect 14928 32945 14974 32956
rect 14238 32862 14284 32873
rect 14221 32835 14238 32837
rect 14422 32862 14468 32873
rect 14284 32835 14301 32837
rect 14146 32715 14233 32835
rect 14289 32715 14301 32835
rect 14221 32713 14238 32715
rect 14146 32415 14238 32535
rect 14284 32713 14301 32715
rect 14405 32535 14422 32537
rect 14606 32862 14652 32873
rect 14589 32835 14606 32837
rect 14790 32862 14836 32873
rect 14652 32835 14669 32837
rect 14589 32715 14601 32835
rect 14657 32715 14669 32835
rect 14589 32713 14606 32715
rect 14468 32535 14485 32537
rect 14405 32415 14417 32535
rect 14473 32415 14485 32535
rect 14405 32413 14422 32415
rect 14238 32377 14284 32388
rect 14468 32413 14485 32415
rect 14422 32377 14468 32388
rect 14652 32713 14669 32715
rect 14773 32535 14790 32537
rect 14911 32835 14928 32837
rect 14974 32835 14991 32837
rect 14911 32714 14923 32835
rect 14979 32714 14991 32835
rect 14911 32712 14928 32714
rect 14836 32535 14853 32537
rect 14773 32415 14785 32535
rect 14841 32415 14853 32535
rect 14773 32413 14790 32415
rect 14606 32377 14652 32388
rect 14836 32413 14853 32415
rect 14790 32377 14836 32388
rect 14315 32339 14326 32342
rect 14380 32339 14391 32342
rect 14499 32339 14510 32342
rect 14564 32339 14575 32342
rect 14683 32339 14694 32342
rect 14748 32339 14759 32342
rect 14100 32294 14146 32305
rect 14313 32283 14325 32339
rect 14381 32283 14393 32339
rect 14313 32269 14393 32283
rect 14497 32283 14509 32339
rect 14565 32283 14577 32339
rect 14497 32269 14577 32283
rect 14681 32283 14693 32339
rect 14749 32283 14761 32339
rect 14974 32712 14991 32714
rect 14928 32294 14974 32305
rect 14681 32269 14761 32283
rect 14313 32189 14393 32191
rect 13925 32133 14325 32189
rect 14381 32133 14393 32189
rect 15411 32190 15467 33210
rect 16569 33198 16649 33210
rect 16075 33159 16161 33163
rect 16075 33103 16087 33159
rect 16143 33103 16161 33159
rect 16075 33091 16161 33103
rect 15586 32946 15632 32957
rect 15801 32955 15877 32988
rect 15801 32909 15812 32955
rect 15866 32909 15877 32955
rect 15985 32955 16061 32988
rect 15985 32909 15996 32955
rect 16050 32909 16061 32955
rect 16169 32955 16245 32988
rect 16169 32909 16180 32955
rect 16234 32909 16245 32955
rect 16414 32946 16460 32957
rect 15724 32863 15770 32874
rect 15707 32836 15724 32838
rect 15908 32863 15954 32874
rect 15770 32836 15787 32838
rect 15632 32716 15719 32836
rect 15775 32716 15787 32836
rect 15707 32714 15724 32716
rect 15632 32416 15724 32536
rect 15770 32714 15787 32716
rect 15891 32536 15908 32538
rect 16092 32863 16138 32874
rect 16075 32836 16092 32838
rect 16276 32863 16322 32874
rect 16138 32836 16155 32838
rect 16075 32716 16087 32836
rect 16143 32716 16155 32836
rect 16075 32714 16092 32716
rect 15954 32536 15971 32538
rect 15891 32416 15903 32536
rect 15959 32416 15971 32536
rect 15891 32414 15908 32416
rect 15724 32378 15770 32389
rect 15954 32414 15971 32416
rect 15908 32378 15954 32389
rect 16138 32714 16155 32716
rect 16259 32536 16276 32538
rect 16397 32836 16414 32838
rect 16460 32836 16477 32838
rect 16397 32715 16409 32836
rect 16465 32715 16477 32836
rect 16397 32713 16414 32715
rect 16322 32536 16339 32538
rect 16259 32416 16271 32536
rect 16327 32416 16339 32536
rect 16259 32414 16276 32416
rect 16092 32378 16138 32389
rect 16322 32414 16339 32416
rect 16276 32378 16322 32389
rect 15801 32340 15812 32343
rect 15866 32340 15877 32343
rect 15985 32340 15996 32343
rect 16050 32340 16061 32343
rect 16169 32340 16180 32343
rect 16234 32340 16245 32343
rect 15586 32295 15632 32306
rect 15799 32284 15811 32340
rect 15867 32284 15879 32340
rect 15799 32270 15879 32284
rect 15983 32284 15995 32340
rect 16051 32284 16063 32340
rect 15983 32270 16063 32284
rect 16167 32284 16179 32340
rect 16235 32284 16247 32340
rect 16460 32713 16477 32715
rect 16414 32295 16460 32306
rect 16167 32270 16247 32284
rect 15799 32190 15879 32192
rect 15411 32134 15811 32190
rect 15867 32134 15879 32190
rect 14313 32131 14393 32133
rect 15799 32132 15879 32134
rect 14497 32073 14577 32075
rect 13789 32017 14509 32073
rect 14565 32017 14577 32073
rect 14497 32015 14577 32017
rect 14826 32073 14906 32075
rect 15093 32074 15163 32085
rect 15983 32074 16063 32076
rect 15093 32073 15995 32074
rect 14826 32017 14838 32073
rect 14894 32017 15095 32073
rect 15151 32018 15995 32073
rect 16051 32018 16063 32074
rect 15151 32017 15411 32018
rect 14826 32015 14906 32017
rect 15093 32007 15163 32017
rect 15983 32016 16063 32018
rect 16312 32074 16392 32076
rect 16755 32074 16825 32084
rect 16312 32018 16324 32074
rect 16380 32018 16757 32074
rect 16813 32018 16825 32074
rect 16312 32016 16392 32018
rect 16755 32006 16825 32018
rect 4169 31956 4239 31968
rect 5209 31956 5289 31958
rect 6695 31957 6775 31959
rect 4169 31900 4181 31956
rect 4237 31900 5221 31956
rect 5277 31900 5289 31956
rect 4169 31888 4239 31900
rect 521 30849 685 30861
rect 1001 30927 1165 30939
rect 1001 30871 1013 30927
rect 1069 30871 1165 30927
rect 1001 30859 1165 30871
rect 521 30793 533 30849
rect 589 30793 685 30849
rect 521 30781 685 30793
rect 589 30731 685 30781
rect -514 30709 -468 30720
rect -1408 30409 -1362 30549
rect -1193 30418 -1097 30449
rect -1193 30372 -1182 30418
rect -1108 30372 -1097 30418
rect -928 30409 -882 30549
rect -1362 30326 -1224 30337
rect -1362 29752 -1270 30326
rect -1066 30326 -1020 30337
rect -1083 30042 -1066 30052
rect -1020 30042 -1003 30052
rect -1083 29802 -1071 30042
rect -1015 29802 -1003 30042
rect -1083 29792 -1066 29802
rect -1362 29741 -1224 29752
rect -1020 29792 -1003 29802
rect -1066 29741 -1020 29752
rect -1408 29658 -1362 29669
rect -1193 29660 -1182 29706
rect -1108 29660 -1097 29706
rect -1193 29519 -1097 29660
rect -299 30718 1 30731
rect -299 30672 -288 30718
rect -214 30685 -84 30718
rect -214 30672 -203 30685
rect -95 30672 -84 30685
rect -10 30672 1 30718
rect 170 30709 216 30720
rect -468 30626 -330 30637
rect -468 30452 -376 30626
rect -172 30626 -126 30637
rect -189 30567 -172 30577
rect 32 30626 170 30637
rect -126 30567 -109 30577
rect -189 30511 -177 30567
rect -121 30511 -109 30567
rect -189 30501 -172 30511
rect -468 30441 -330 30452
rect -126 30501 -109 30511
rect -172 30441 -126 30452
rect 78 30452 170 30626
rect 32 30441 170 30452
rect -514 30229 -468 30369
rect -299 30360 -288 30406
rect -214 30360 -203 30406
rect -299 30329 -203 30360
rect -95 30360 -84 30406
rect -10 30360 1 30406
rect -95 30329 1 30360
rect 385 30718 685 30731
rect 385 30672 396 30718
rect 470 30685 600 30718
rect 470 30672 481 30685
rect 589 30672 600 30685
rect 674 30672 685 30718
rect 854 30709 900 30720
rect 308 30626 354 30637
rect 291 30567 308 30577
rect 512 30626 558 30637
rect 354 30567 371 30577
rect 291 30511 303 30567
rect 359 30511 371 30567
rect 291 30501 308 30511
rect 354 30501 371 30511
rect 495 30567 512 30577
rect 716 30626 762 30637
rect 558 30567 575 30577
rect 495 30511 507 30567
rect 563 30511 575 30567
rect 495 30501 512 30511
rect 308 30441 354 30452
rect 558 30501 575 30511
rect 699 30567 716 30577
rect 762 30567 779 30577
rect 699 30511 711 30567
rect 767 30511 779 30567
rect 699 30501 716 30511
rect 512 30441 558 30452
rect 762 30501 779 30511
rect 716 30441 762 30452
rect 170 30229 216 30369
rect 385 30360 396 30406
rect 470 30360 481 30406
rect 385 30329 481 30360
rect 589 30360 600 30406
rect 674 30360 685 30406
rect 589 30329 685 30360
rect 1069 30718 1165 30859
rect 1677 30973 3645 31169
rect 4453 31169 4509 31900
rect 5209 31898 5289 31900
rect 5939 31901 6707 31957
rect 6763 31901 6775 31957
rect 4841 31806 4921 31820
rect 4628 31784 4674 31795
rect 4841 31750 4853 31806
rect 4909 31750 4921 31806
rect 5025 31806 5105 31820
rect 5025 31750 5037 31806
rect 5093 31750 5105 31806
rect 5209 31806 5289 31820
rect 5209 31750 5221 31806
rect 5277 31750 5289 31806
rect 5456 31784 5502 31795
rect 4843 31747 4854 31750
rect 4908 31747 4919 31750
rect 5027 31747 5038 31750
rect 5092 31747 5103 31750
rect 5211 31747 5222 31750
rect 5276 31747 5287 31750
rect 4766 31701 4812 31712
rect 4674 31527 4766 31701
rect 4766 31516 4812 31527
rect 4950 31701 4996 31712
rect 4950 31516 4996 31527
rect 5134 31701 5180 31712
rect 5318 31701 5364 31712
rect 5301 31674 5318 31676
rect 5364 31674 5381 31676
rect 5301 31554 5313 31674
rect 5369 31554 5381 31674
rect 5301 31552 5318 31554
rect 5134 31516 5180 31527
rect 5364 31552 5381 31554
rect 5318 31516 5364 31527
rect 4628 31299 4674 31444
rect 4843 31435 4854 31481
rect 4908 31435 4919 31481
rect 4843 31402 4919 31435
rect 5027 31435 5038 31481
rect 5092 31435 5103 31481
rect 5027 31402 5103 31435
rect 5211 31435 5222 31481
rect 5276 31435 5287 31481
rect 5211 31402 5287 31435
rect 5456 31299 5502 31444
rect 4616 31287 4696 31299
rect 4616 31231 4628 31287
rect 4684 31231 4696 31287
rect 4616 31219 4696 31231
rect 5434 31287 5512 31299
rect 5434 31231 5446 31287
rect 5502 31231 5512 31287
rect 5434 31219 5512 31231
rect 5787 31169 5867 31179
rect 4453 31113 5799 31169
rect 5855 31113 5867 31169
rect 5787 31111 5867 31113
rect 5621 31060 5691 31062
rect 1677 30833 1777 30973
rect 3545 30833 3645 30973
rect 1677 30793 3645 30833
rect 4453 31059 5691 31060
rect 4453 31005 5623 31059
rect 5679 31005 5691 31059
rect 4453 31004 5691 31005
rect 1069 30672 1080 30718
rect 1154 30672 1165 30718
rect 1334 30709 1380 30720
rect 900 30626 1038 30637
rect 900 30452 992 30626
rect 1196 30626 1242 30637
rect 1179 30567 1196 30577
rect 1242 30567 1259 30577
rect 1179 30511 1191 30567
rect 1247 30511 1259 30567
rect 1179 30501 1196 30511
rect 900 30441 1038 30452
rect 1242 30501 1259 30511
rect 1196 30441 1242 30452
rect 854 30229 900 30369
rect 1069 30360 1080 30406
rect 1154 30360 1165 30406
rect 1069 30329 1165 30360
rect 1334 30229 1380 30369
rect 1714 30653 1760 30793
rect -551 30199 1417 30229
rect -551 30059 717 30199
rect 1317 30059 1417 30199
rect -551 30029 1417 30059
rect 1929 30662 2025 30693
rect 1929 30616 1940 30662
rect 2014 30616 2025 30662
rect 2133 30662 2229 30693
rect 2133 30616 2144 30662
rect 2218 30616 2229 30662
rect 2398 30653 2444 30793
rect 1760 30570 1898 30581
rect 2056 30570 2102 30581
rect 2260 30570 2398 30581
rect 1760 29996 1852 30570
rect 2039 30330 2051 30570
rect 2107 30330 2119 30570
rect 1760 29985 1898 29996
rect 2056 29985 2102 29996
rect 2306 29996 2398 30570
rect 2260 29985 2398 29996
rect 1714 29902 1760 29913
rect 1929 29904 1940 29950
rect 2014 29930 2025 29950
rect 2133 29930 2144 29950
rect 2014 29904 2144 29930
rect 2218 29904 2229 29950
rect 1929 29877 2229 29904
rect 2613 30662 2709 30693
rect 2613 30616 2624 30662
rect 2698 30616 2709 30662
rect 2817 30662 2913 30693
rect 2817 30616 2828 30662
rect 2902 30616 2913 30662
rect 3082 30653 3128 30793
rect 2536 30570 2582 30581
rect 2740 30570 2786 30581
rect 2944 30570 2990 30581
rect 2723 30330 2735 30570
rect 2791 30330 2803 30570
rect 2519 29996 2531 30236
rect 2587 29996 2599 30236
rect 2927 29996 2939 30236
rect 2995 29996 3007 30236
rect 2536 29985 2582 29996
rect 2740 29985 2786 29996
rect 2944 29985 2990 29996
rect 2398 29902 2444 29913
rect 2613 29904 2624 29950
rect 2698 29930 2709 29950
rect 2817 29930 2828 29950
rect 2698 29904 2828 29930
rect 2902 29904 2913 29950
rect 2613 29877 2913 29904
rect 3297 30662 3393 30693
rect 3297 30616 3308 30662
rect 3382 30616 3393 30662
rect 3562 30653 3608 30793
rect 3128 30570 3266 30581
rect 3128 29996 3220 30570
rect 3424 30570 3470 30581
rect 3407 30286 3424 30296
rect 3470 30286 3487 30296
rect 3407 30046 3419 30286
rect 3475 30046 3487 30286
rect 3407 30036 3424 30046
rect 3128 29985 3266 29996
rect 3470 30036 3487 30046
rect 3424 29985 3470 29996
rect 3082 29902 3128 29913
rect 3297 29904 3308 29950
rect 3382 29904 3393 29950
rect 1929 29829 2025 29877
rect -928 29658 -882 29669
rect -551 29799 1417 29829
rect -551 29659 717 29799
rect 1317 29659 1417 29799
rect -551 29629 1417 29659
rect 1929 29773 1949 29829
rect 2005 29773 2025 29829
rect -1261 29507 -1097 29519
rect -1261 29451 -1249 29507
rect -1193 29451 -1097 29507
rect -1261 29439 -1097 29451
rect -5622 28908 -5610 28964
rect -5554 28908 -5427 28964
rect -5371 28908 -3477 28964
rect -1408 29289 -1362 29300
rect -1193 29298 -1097 29439
rect -514 29489 -468 29500
rect -1193 29252 -1182 29298
rect -1108 29252 -1097 29298
rect -928 29289 -882 29300
rect -1362 29206 -1224 29217
rect -1362 29032 -1270 29206
rect -1066 29206 -1020 29217
rect -1083 29147 -1066 29157
rect -1020 29147 -1003 29157
rect -1083 29091 -1071 29147
rect -1015 29091 -1003 29147
rect -1083 29081 -1066 29091
rect -1362 29021 -1224 29032
rect -1020 29081 -1003 29091
rect -1066 29021 -1020 29032
rect -5622 28896 -5536 28908
rect -5429 28896 -5369 28908
rect -8951 28509 -8787 28521
rect -8471 28587 -8307 28599
rect -8471 28531 -8459 28587
rect -8403 28531 -8307 28587
rect -8471 28519 -8307 28531
rect -8951 28453 -8939 28509
rect -8883 28453 -8787 28509
rect -8951 28441 -8787 28453
rect -8883 28391 -8787 28441
rect -9986 28369 -9940 28380
rect -9771 28378 -9471 28391
rect -9771 28332 -9760 28378
rect -9686 28345 -9556 28378
rect -9686 28332 -9675 28345
rect -9567 28332 -9556 28345
rect -9482 28332 -9471 28378
rect -9302 28369 -9256 28380
rect -9940 28286 -9802 28297
rect -9940 28112 -9848 28286
rect -9644 28286 -9598 28297
rect -9661 28227 -9644 28237
rect -9440 28286 -9302 28297
rect -9598 28227 -9581 28237
rect -9661 28171 -9649 28227
rect -9593 28171 -9581 28227
rect -9661 28161 -9644 28171
rect -9940 28101 -9802 28112
rect -9598 28161 -9581 28171
rect -9644 28101 -9598 28112
rect -9394 28112 -9302 28286
rect -9440 28101 -9302 28112
rect -9986 27889 -9940 28029
rect -9771 28020 -9760 28066
rect -9686 28020 -9675 28066
rect -9771 27989 -9675 28020
rect -9567 28020 -9556 28066
rect -9482 28020 -9471 28066
rect -9567 27989 -9471 28020
rect -9087 28378 -8787 28391
rect -9087 28332 -9076 28378
rect -9002 28345 -8872 28378
rect -9002 28332 -8991 28345
rect -8883 28332 -8872 28345
rect -8798 28332 -8787 28378
rect -8618 28369 -8572 28380
rect -9164 28286 -9118 28297
rect -9181 28227 -9164 28237
rect -8960 28286 -8914 28297
rect -9118 28227 -9101 28237
rect -9181 28171 -9169 28227
rect -9113 28171 -9101 28227
rect -9181 28161 -9164 28171
rect -9118 28161 -9101 28171
rect -8977 28227 -8960 28237
rect -8756 28286 -8710 28297
rect -8914 28227 -8897 28237
rect -8977 28171 -8965 28227
rect -8909 28171 -8897 28227
rect -8977 28161 -8960 28171
rect -9164 28101 -9118 28112
rect -8914 28161 -8897 28171
rect -8773 28227 -8756 28237
rect -8710 28227 -8693 28237
rect -8773 28171 -8761 28227
rect -8705 28171 -8693 28227
rect -8773 28161 -8756 28171
rect -8960 28101 -8914 28112
rect -8710 28161 -8693 28171
rect -8756 28101 -8710 28112
rect -9302 27889 -9256 28029
rect -9087 28020 -9076 28066
rect -9002 28020 -8991 28066
rect -9087 27989 -8991 28020
rect -8883 28020 -8872 28066
rect -8798 28020 -8787 28066
rect -8883 27989 -8787 28020
rect -8403 28378 -8307 28519
rect -7795 28689 -5827 28873
rect -1408 28809 -1362 28949
rect -1193 28940 -1182 28986
rect -1108 28940 -1097 28986
rect -1193 28909 -1097 28940
rect -928 28809 -882 28949
rect -8403 28332 -8392 28378
rect -8318 28332 -8307 28378
rect -8138 28369 -8092 28380
rect -8572 28286 -8434 28297
rect -8572 28112 -8480 28286
rect -8276 28286 -8230 28297
rect -8293 28227 -8276 28237
rect -8230 28227 -8213 28237
rect -8293 28171 -8281 28227
rect -8225 28171 -8213 28227
rect -8293 28161 -8276 28171
rect -8572 28101 -8434 28112
rect -8230 28161 -8213 28171
rect -8276 28101 -8230 28112
rect -8618 27889 -8572 28029
rect -8403 28020 -8392 28066
rect -8318 28020 -8307 28066
rect -8403 27989 -8307 28020
rect -8138 27889 -8092 28029
rect -7795 27889 -6327 28689
rect -6027 28089 -5827 28689
rect -1445 28089 -845 28809
rect -299 29498 -203 29529
rect -299 29452 -288 29498
rect -214 29452 -203 29498
rect -34 29489 420 29629
rect -376 29406 -330 29417
rect -393 29122 -376 29132
rect -172 29406 -34 29417
rect -330 29122 -313 29132
rect -393 28882 -381 29122
rect -325 28882 -313 29122
rect -393 28872 -376 28882
rect -330 28872 -313 28882
rect -376 28821 -330 28832
rect -126 28832 -34 29406
rect -172 28821 -34 28832
rect -514 28738 -468 28749
rect -299 28740 -288 28786
rect -214 28740 -203 28786
rect -299 28665 -203 28740
rect 12 28821 374 29489
rect -34 28738 12 28749
rect 589 29498 685 29529
rect 589 29452 600 29498
rect 674 29452 685 29498
rect 854 29489 900 29629
rect 420 29406 558 29417
rect 420 28832 512 29406
rect 716 29406 762 29417
rect 699 29122 716 29132
rect 762 29122 779 29132
rect 699 28882 711 29122
rect 767 28882 779 29122
rect 699 28872 716 28882
rect 420 28821 558 28832
rect 762 28872 779 28882
rect 716 28821 762 28832
rect 374 28738 420 28749
rect 589 28740 600 28786
rect 674 28740 685 28786
rect -299 28609 -279 28665
rect -223 28609 -203 28665
rect -299 28391 -203 28609
rect 589 28521 685 28740
rect 1069 29498 1165 29529
rect 1069 29452 1080 29498
rect 1154 29452 1165 29498
rect 1334 29489 1380 29629
rect 900 29406 1038 29417
rect 900 28832 992 29406
rect 1196 29406 1242 29417
rect 1179 29122 1196 29132
rect 1242 29122 1259 29132
rect 1179 28882 1191 29122
rect 1247 28882 1259 29122
rect 1179 28872 1196 28882
rect 900 28821 1038 28832
rect 1242 28872 1259 28882
rect 1196 28821 1242 28832
rect 854 28738 900 28749
rect 1069 28740 1080 28786
rect 1154 28740 1165 28786
rect 1069 28599 1165 28740
rect 1714 29533 1760 29544
rect 1929 29542 2025 29773
rect 2613 29673 2709 29877
rect 3297 29763 3393 29904
rect 4453 29983 4509 31004
rect 5621 30996 5691 31004
rect 5117 30952 5203 30956
rect 5117 30896 5129 30952
rect 5185 30896 5203 30952
rect 5117 30884 5203 30896
rect 4628 30739 4674 30750
rect 4843 30748 4919 30781
rect 4843 30702 4854 30748
rect 4908 30702 4919 30748
rect 5027 30748 5103 30781
rect 5027 30702 5038 30748
rect 5092 30702 5103 30748
rect 5211 30748 5287 30781
rect 5211 30702 5222 30748
rect 5276 30702 5287 30748
rect 5456 30739 5502 30750
rect 4766 30656 4812 30667
rect 4749 30629 4766 30631
rect 4950 30656 4996 30667
rect 4812 30629 4829 30631
rect 4674 30509 4761 30629
rect 4817 30509 4829 30629
rect 4749 30507 4766 30509
rect 4674 30209 4766 30329
rect 4812 30507 4829 30509
rect 4933 30329 4950 30331
rect 5134 30656 5180 30667
rect 5117 30629 5134 30631
rect 5318 30656 5364 30667
rect 5180 30629 5197 30631
rect 5117 30509 5129 30629
rect 5185 30509 5197 30629
rect 5117 30507 5134 30509
rect 4996 30329 5013 30331
rect 4933 30209 4945 30329
rect 5001 30209 5013 30329
rect 4933 30207 4950 30209
rect 4766 30171 4812 30182
rect 4996 30207 5013 30209
rect 4950 30171 4996 30182
rect 5180 30507 5197 30509
rect 5301 30329 5318 30331
rect 5439 30629 5456 30631
rect 5502 30629 5519 30631
rect 5439 30508 5451 30629
rect 5507 30508 5519 30629
rect 5439 30506 5456 30508
rect 5364 30329 5381 30331
rect 5301 30209 5313 30329
rect 5369 30209 5381 30329
rect 5301 30207 5318 30209
rect 5134 30171 5180 30182
rect 5364 30207 5381 30209
rect 5318 30171 5364 30182
rect 4843 30133 4854 30136
rect 4908 30133 4919 30136
rect 5027 30133 5038 30136
rect 5092 30133 5103 30136
rect 5211 30133 5222 30136
rect 5276 30133 5287 30136
rect 4628 30088 4674 30099
rect 4841 30077 4853 30133
rect 4909 30077 4921 30133
rect 4841 30063 4921 30077
rect 5025 30077 5037 30133
rect 5093 30077 5105 30133
rect 5025 30063 5105 30077
rect 5209 30077 5221 30133
rect 5277 30077 5289 30133
rect 5502 30506 5519 30508
rect 5456 30088 5502 30099
rect 5209 30063 5289 30077
rect 4841 29983 4921 29985
rect 4453 29927 4853 29983
rect 4909 29927 4921 29983
rect 4841 29925 4921 29927
rect 3562 29902 3608 29913
rect 4033 29867 4103 29881
rect 5025 29867 5105 29869
rect 4033 29811 4045 29867
rect 4101 29811 5037 29867
rect 5093 29811 5105 29867
rect 4033 29799 4103 29811
rect 5025 29809 5105 29811
rect 5354 29867 5434 29869
rect 5797 29867 5857 29879
rect 5354 29811 5366 29867
rect 5422 29811 5799 29867
rect 5855 29811 5857 29867
rect 5354 29809 5434 29811
rect 5797 29799 5857 29811
rect 3229 29751 3393 29763
rect 3229 29695 3241 29751
rect 3297 29695 3393 29751
rect 3229 29683 3393 29695
rect 3799 29751 3877 29762
rect 5209 29751 5289 29753
rect 3799 29750 5221 29751
rect 3799 29696 3811 29750
rect 3865 29696 5221 29750
rect 3799 29695 5221 29696
rect 5277 29695 5289 29751
rect 3799 29684 3877 29695
rect 5209 29693 5289 29695
rect 2613 29617 2633 29673
rect 2689 29617 2709 29673
rect 1929 29496 1940 29542
rect 2014 29496 2025 29542
rect 2194 29533 2444 29544
rect 1852 29450 1898 29461
rect 1835 29391 1852 29401
rect 2056 29450 2194 29461
rect 1898 29391 1915 29401
rect 1835 29335 1847 29391
rect 1903 29335 1915 29391
rect 1835 29325 1852 29335
rect 1898 29325 1915 29335
rect 1852 29265 1898 29276
rect 2102 29276 2194 29450
rect 2056 29265 2194 29276
rect 1714 29053 1760 29193
rect 1929 29184 1940 29230
rect 2014 29184 2025 29230
rect 1929 29153 2025 29184
rect 2240 29193 2398 29533
rect 2613 29542 2709 29617
rect 2613 29496 2624 29542
rect 2698 29496 2709 29542
rect 2878 29533 2924 29544
rect 2444 29450 2582 29461
rect 2444 29276 2536 29450
rect 2740 29450 2786 29461
rect 2723 29391 2740 29401
rect 2786 29391 2803 29401
rect 2723 29335 2735 29391
rect 2791 29335 2803 29391
rect 2723 29325 2740 29335
rect 2444 29265 2582 29276
rect 2786 29325 2803 29335
rect 2740 29265 2786 29276
rect 2194 29182 2444 29193
rect 2613 29184 2624 29230
rect 2698 29184 2709 29230
rect 2240 29053 2398 29182
rect 2613 29153 2709 29184
rect 2878 29053 2924 29193
rect 3082 29533 3128 29544
rect 3297 29542 3393 29683
rect 4841 29601 4921 29615
rect 4628 29579 4674 29590
rect 3297 29496 3308 29542
rect 3382 29496 3393 29542
rect 3562 29533 3608 29544
rect 3128 29450 3266 29461
rect 3128 29276 3220 29450
rect 3424 29450 3470 29461
rect 3407 29391 3424 29401
rect 3470 29391 3487 29401
rect 3407 29335 3419 29391
rect 3475 29335 3487 29391
rect 3407 29325 3424 29335
rect 3128 29265 3266 29276
rect 3470 29325 3487 29335
rect 3424 29265 3470 29276
rect 3082 29053 3128 29193
rect 3297 29184 3308 29230
rect 3382 29184 3393 29230
rect 3297 29153 3393 29184
rect 3562 29053 3608 29193
rect 4841 29545 4853 29601
rect 4909 29545 4921 29601
rect 5025 29601 5105 29615
rect 5025 29545 5037 29601
rect 5093 29545 5105 29601
rect 5209 29601 5289 29615
rect 5209 29545 5221 29601
rect 5277 29545 5289 29601
rect 5456 29579 5502 29590
rect 4843 29542 4854 29545
rect 4908 29542 4919 29545
rect 5027 29542 5038 29545
rect 5092 29542 5103 29545
rect 5211 29542 5222 29545
rect 5276 29542 5287 29545
rect 4766 29496 4812 29507
rect 4674 29322 4766 29496
rect 4766 29311 4812 29322
rect 4950 29496 4996 29507
rect 4950 29311 4996 29322
rect 5134 29496 5180 29507
rect 5318 29496 5364 29507
rect 5301 29469 5318 29471
rect 5364 29469 5381 29471
rect 5301 29349 5313 29469
rect 5369 29349 5381 29469
rect 5301 29347 5318 29349
rect 5134 29311 5180 29322
rect 5364 29347 5381 29349
rect 5318 29311 5364 29322
rect 4628 29094 4674 29239
rect 4843 29230 4854 29276
rect 4908 29230 4919 29276
rect 4843 29197 4919 29230
rect 5027 29230 5038 29276
rect 5092 29230 5103 29276
rect 5027 29197 5103 29230
rect 5211 29230 5222 29276
rect 5276 29230 5287 29276
rect 5211 29197 5287 29230
rect 5456 29094 5502 29239
rect 4616 29082 4696 29094
rect 1334 28738 1380 28749
rect 1677 29013 3645 29053
rect 4616 29026 4628 29082
rect 4684 29026 4696 29082
rect 4616 29014 4696 29026
rect 5434 29082 5514 29094
rect 5434 29026 5446 29082
rect 5502 29026 5514 29082
rect 5434 29014 5514 29026
rect 1677 28873 1777 29013
rect 3545 28873 3645 29013
rect 3850 28964 3936 28976
rect 4043 28964 4103 28968
rect 5939 28964 5995 31901
rect 6695 31899 6775 31901
rect 6327 31807 6407 31821
rect 6114 31785 6160 31796
rect 6327 31751 6339 31807
rect 6395 31751 6407 31807
rect 6511 31807 6591 31821
rect 6511 31751 6523 31807
rect 6579 31751 6591 31807
rect 6695 31807 6775 31821
rect 6695 31751 6707 31807
rect 6763 31751 6775 31807
rect 6942 31785 6988 31796
rect 6329 31748 6340 31751
rect 6394 31748 6405 31751
rect 6513 31748 6524 31751
rect 6578 31748 6589 31751
rect 6697 31748 6708 31751
rect 6762 31748 6773 31751
rect 6252 31702 6298 31713
rect 6160 31528 6252 31702
rect 6252 31517 6298 31528
rect 6436 31702 6482 31713
rect 6436 31517 6482 31528
rect 6620 31702 6666 31713
rect 6804 31702 6850 31713
rect 6787 31675 6804 31677
rect 6850 31675 6867 31677
rect 6787 31555 6799 31675
rect 6855 31555 6867 31675
rect 6787 31553 6804 31555
rect 6620 31517 6666 31528
rect 6850 31553 6867 31555
rect 6804 31517 6850 31528
rect 6114 31300 6160 31445
rect 6329 31436 6340 31482
rect 6394 31436 6405 31482
rect 6329 31403 6405 31436
rect 6513 31436 6524 31482
rect 6578 31436 6589 31482
rect 6513 31403 6589 31436
rect 6697 31436 6708 31482
rect 6762 31436 6773 31482
rect 6697 31403 6773 31436
rect 6942 31300 6988 31445
rect 6102 31288 6182 31300
rect 6102 31232 6114 31288
rect 6170 31232 6182 31288
rect 6102 31220 6182 31232
rect 6920 31288 6998 31300
rect 6920 31232 6932 31288
rect 6988 31232 6998 31288
rect 6920 31220 6998 31232
rect 8027 31170 8227 31970
rect 8427 31170 8627 31970
rect 8027 30550 8627 31170
rect 8958 31830 9004 31841
rect 9173 31839 9269 31870
rect 9173 31793 9184 31839
rect 9258 31793 9269 31839
rect 9438 31830 9892 31970
rect 9096 31747 9142 31758
rect 9079 31463 9096 31473
rect 9300 31747 9438 31758
rect 9142 31463 9159 31473
rect 9079 31223 9091 31463
rect 9147 31223 9159 31463
rect 9079 31213 9096 31223
rect 9142 31213 9159 31223
rect 9096 31162 9142 31173
rect 9346 31173 9438 31747
rect 9300 31162 9438 31173
rect 8958 31079 9004 31090
rect 9173 31081 9184 31127
rect 9258 31081 9269 31127
rect 9173 31006 9269 31081
rect 9484 31162 9846 31830
rect 9438 31079 9484 31090
rect 10061 31839 10157 31870
rect 10061 31793 10072 31839
rect 10146 31793 10157 31839
rect 10326 31830 10372 31970
rect 9892 31747 10030 31758
rect 9892 31173 9984 31747
rect 10188 31747 10234 31758
rect 10171 31463 10188 31473
rect 10234 31463 10251 31473
rect 10171 31223 10183 31463
rect 10239 31223 10251 31463
rect 10171 31213 10188 31223
rect 9892 31162 10030 31173
rect 10234 31213 10251 31223
rect 10188 31162 10234 31173
rect 9846 31079 9892 31090
rect 10061 31081 10072 31127
rect 10146 31081 10157 31127
rect 9173 30950 9193 31006
rect 9249 30950 9269 31006
rect 9173 30732 9269 30950
rect 10061 30862 10157 31081
rect 10541 31839 10637 31870
rect 10541 31793 10552 31839
rect 10626 31793 10637 31839
rect 10806 31830 10852 31970
rect 10372 31747 10510 31758
rect 10372 31173 10464 31747
rect 10668 31747 10714 31758
rect 10651 31463 10668 31473
rect 10714 31463 10731 31473
rect 10651 31223 10663 31463
rect 10719 31223 10731 31463
rect 10651 31213 10668 31223
rect 10372 31162 10510 31173
rect 10714 31213 10731 31223
rect 10668 31162 10714 31173
rect 10326 31079 10372 31090
rect 10541 31081 10552 31127
rect 10626 31081 10637 31127
rect 10541 30940 10637 31081
rect 10806 31079 10852 31090
rect 11149 31170 12617 31970
rect 12917 31170 13117 31970
rect 17499 31970 22589 32170
rect 23261 32073 23317 33320
rect 26217 33318 26297 33320
rect 32167 33376 32249 33388
rect 32733 33376 32789 34106
rect 33625 34104 33705 34106
rect 34355 34106 35123 34162
rect 35179 34106 35191 34162
rect 33257 34012 33337 34026
rect 33044 33990 33090 34001
rect 33257 33956 33269 34012
rect 33325 33956 33337 34012
rect 33441 34012 33521 34026
rect 33441 33956 33453 34012
rect 33509 33956 33521 34012
rect 33625 34012 33705 34026
rect 33625 33956 33637 34012
rect 33693 33956 33705 34012
rect 33872 33990 33918 34001
rect 33259 33953 33270 33956
rect 33324 33953 33335 33956
rect 33443 33953 33454 33956
rect 33508 33953 33519 33956
rect 33627 33953 33638 33956
rect 33692 33953 33703 33956
rect 33182 33907 33228 33918
rect 33090 33733 33182 33907
rect 33182 33722 33228 33733
rect 33366 33907 33412 33918
rect 33366 33722 33412 33733
rect 33550 33907 33596 33918
rect 33734 33907 33780 33918
rect 33717 33880 33734 33882
rect 33780 33880 33797 33882
rect 33717 33760 33729 33880
rect 33785 33760 33797 33880
rect 33717 33758 33734 33760
rect 33550 33722 33596 33733
rect 33780 33758 33797 33760
rect 33734 33722 33780 33733
rect 33044 33505 33090 33650
rect 33259 33641 33270 33687
rect 33324 33641 33335 33687
rect 33259 33608 33335 33641
rect 33443 33641 33454 33687
rect 33508 33641 33519 33687
rect 33443 33608 33519 33641
rect 33627 33641 33638 33687
rect 33692 33641 33703 33687
rect 33627 33608 33703 33641
rect 33872 33505 33918 33650
rect 33032 33493 33112 33505
rect 33032 33437 33044 33493
rect 33100 33437 33112 33493
rect 33032 33425 33112 33437
rect 33850 33493 33928 33505
rect 33850 33437 33862 33493
rect 33918 33437 33928 33493
rect 33850 33425 33928 33437
rect 32167 33320 32181 33376
rect 32237 33320 32789 33376
rect 34355 33376 34411 34106
rect 35111 34104 35191 34106
rect 42205 34106 43109 34162
rect 43165 34106 43177 34162
rect 34743 34012 34823 34026
rect 34530 33990 34576 34001
rect 34743 33956 34755 34012
rect 34811 33956 34823 34012
rect 34927 34012 35007 34026
rect 34927 33956 34939 34012
rect 34995 33956 35007 34012
rect 35111 34012 35191 34026
rect 35111 33956 35123 34012
rect 35179 33956 35191 34012
rect 35358 33990 35404 34001
rect 34745 33953 34756 33956
rect 34810 33953 34821 33956
rect 34929 33953 34940 33956
rect 34994 33953 35005 33956
rect 35113 33953 35124 33956
rect 35178 33953 35189 33956
rect 34668 33907 34714 33918
rect 34576 33733 34668 33907
rect 34668 33722 34714 33733
rect 34852 33907 34898 33918
rect 34852 33722 34898 33733
rect 35036 33907 35082 33918
rect 35220 33907 35266 33918
rect 35203 33880 35220 33882
rect 35266 33880 35283 33882
rect 35203 33760 35215 33880
rect 35271 33760 35283 33880
rect 35203 33758 35220 33760
rect 35036 33722 35082 33733
rect 35266 33758 35283 33760
rect 35220 33722 35266 33733
rect 34530 33505 34576 33650
rect 34745 33641 34756 33687
rect 34810 33641 34821 33687
rect 34745 33608 34821 33641
rect 34929 33641 34940 33687
rect 34994 33641 35005 33687
rect 34929 33608 35005 33641
rect 35113 33641 35124 33687
rect 35178 33641 35189 33687
rect 35113 33608 35189 33641
rect 35358 33505 35404 33650
rect 34518 33493 34598 33505
rect 34518 33437 34530 33493
rect 34586 33437 34598 33493
rect 34518 33425 34598 33437
rect 35336 33493 35414 33505
rect 35336 33437 35348 33493
rect 35404 33437 35414 33493
rect 35336 33425 35414 33437
rect 35689 33376 35769 33386
rect 34355 33320 35701 33376
rect 35757 33320 35769 33376
rect 32167 33308 32249 33320
rect 24741 33265 24811 33267
rect 26041 33266 26121 33268
rect 23397 33209 24743 33265
rect 24799 33209 24811 33265
rect 23397 32189 23453 33209
rect 24741 33197 24811 33209
rect 24883 33210 26053 33266
rect 26109 33210 26121 33266
rect 24061 33158 24147 33162
rect 24061 33102 24073 33158
rect 24129 33102 24147 33158
rect 24061 33090 24147 33102
rect 23572 32945 23618 32956
rect 23787 32954 23863 32987
rect 23787 32908 23798 32954
rect 23852 32908 23863 32954
rect 23971 32954 24047 32987
rect 23971 32908 23982 32954
rect 24036 32908 24047 32954
rect 24155 32954 24231 32987
rect 24155 32908 24166 32954
rect 24220 32908 24231 32954
rect 24400 32945 24446 32956
rect 23710 32862 23756 32873
rect 23693 32835 23710 32837
rect 23894 32862 23940 32873
rect 23756 32835 23773 32837
rect 23618 32715 23705 32835
rect 23761 32715 23773 32835
rect 23693 32713 23710 32715
rect 23618 32415 23710 32535
rect 23756 32713 23773 32715
rect 23877 32535 23894 32537
rect 24078 32862 24124 32873
rect 24061 32835 24078 32837
rect 24262 32862 24308 32873
rect 24124 32835 24141 32837
rect 24061 32715 24073 32835
rect 24129 32715 24141 32835
rect 24061 32713 24078 32715
rect 23940 32535 23957 32537
rect 23877 32415 23889 32535
rect 23945 32415 23957 32535
rect 23877 32413 23894 32415
rect 23710 32377 23756 32388
rect 23940 32413 23957 32415
rect 23894 32377 23940 32388
rect 24124 32713 24141 32715
rect 24245 32535 24262 32537
rect 24383 32835 24400 32837
rect 24446 32835 24463 32837
rect 24383 32714 24395 32835
rect 24451 32714 24463 32835
rect 24383 32712 24400 32714
rect 24308 32535 24325 32537
rect 24245 32415 24257 32535
rect 24313 32415 24325 32535
rect 24245 32413 24262 32415
rect 24078 32377 24124 32388
rect 24308 32413 24325 32415
rect 24262 32377 24308 32388
rect 23787 32339 23798 32342
rect 23852 32339 23863 32342
rect 23971 32339 23982 32342
rect 24036 32339 24047 32342
rect 24155 32339 24166 32342
rect 24220 32339 24231 32342
rect 23572 32294 23618 32305
rect 23785 32283 23797 32339
rect 23853 32283 23865 32339
rect 23785 32269 23865 32283
rect 23969 32283 23981 32339
rect 24037 32283 24049 32339
rect 23969 32269 24049 32283
rect 24153 32283 24165 32339
rect 24221 32283 24233 32339
rect 24446 32712 24463 32714
rect 24400 32294 24446 32305
rect 24153 32269 24233 32283
rect 23785 32189 23865 32191
rect 23397 32133 23797 32189
rect 23853 32133 23865 32189
rect 24883 32190 24939 33210
rect 26041 33198 26121 33210
rect 25547 33159 25633 33163
rect 25547 33103 25559 33159
rect 25615 33103 25633 33159
rect 25547 33091 25633 33103
rect 25058 32946 25104 32957
rect 25273 32955 25349 32988
rect 25273 32909 25284 32955
rect 25338 32909 25349 32955
rect 25457 32955 25533 32988
rect 25457 32909 25468 32955
rect 25522 32909 25533 32955
rect 25641 32955 25717 32988
rect 25641 32909 25652 32955
rect 25706 32909 25717 32955
rect 25886 32946 25932 32957
rect 25196 32863 25242 32874
rect 25179 32836 25196 32838
rect 25380 32863 25426 32874
rect 25242 32836 25259 32838
rect 25104 32716 25191 32836
rect 25247 32716 25259 32836
rect 25179 32714 25196 32716
rect 25104 32416 25196 32536
rect 25242 32714 25259 32716
rect 25363 32536 25380 32538
rect 25564 32863 25610 32874
rect 25547 32836 25564 32838
rect 25748 32863 25794 32874
rect 25610 32836 25627 32838
rect 25547 32716 25559 32836
rect 25615 32716 25627 32836
rect 25547 32714 25564 32716
rect 25426 32536 25443 32538
rect 25363 32416 25375 32536
rect 25431 32416 25443 32536
rect 25363 32414 25380 32416
rect 25196 32378 25242 32389
rect 25426 32414 25443 32416
rect 25380 32378 25426 32389
rect 25610 32714 25627 32716
rect 25731 32536 25748 32538
rect 25869 32836 25886 32838
rect 25932 32836 25949 32838
rect 25869 32715 25881 32836
rect 25937 32715 25949 32836
rect 25869 32713 25886 32715
rect 25794 32536 25811 32538
rect 25731 32416 25743 32536
rect 25799 32416 25811 32536
rect 25731 32414 25748 32416
rect 25564 32378 25610 32389
rect 25794 32414 25811 32416
rect 25748 32378 25794 32389
rect 25273 32340 25284 32343
rect 25338 32340 25349 32343
rect 25457 32340 25468 32343
rect 25522 32340 25533 32343
rect 25641 32340 25652 32343
rect 25706 32340 25717 32343
rect 25058 32295 25104 32306
rect 25271 32284 25283 32340
rect 25339 32284 25351 32340
rect 25271 32270 25351 32284
rect 25455 32284 25467 32340
rect 25523 32284 25535 32340
rect 25455 32270 25535 32284
rect 25639 32284 25651 32340
rect 25707 32284 25719 32340
rect 25932 32713 25949 32715
rect 25886 32295 25932 32306
rect 25639 32270 25719 32284
rect 25271 32190 25351 32192
rect 24883 32134 25283 32190
rect 25339 32134 25351 32190
rect 23785 32131 23865 32133
rect 25271 32132 25351 32134
rect 23969 32073 24049 32075
rect 23261 32017 23981 32073
rect 24037 32017 24049 32073
rect 23969 32015 24049 32017
rect 24298 32073 24378 32075
rect 24565 32074 24635 32085
rect 25455 32074 25535 32076
rect 24565 32073 25467 32074
rect 24298 32017 24310 32073
rect 24366 32017 24567 32073
rect 24623 32018 25467 32073
rect 25523 32018 25535 32074
rect 24623 32017 24883 32018
rect 24298 32015 24378 32017
rect 24565 32007 24635 32017
rect 25455 32016 25535 32018
rect 25784 32074 25864 32076
rect 26227 32074 26297 32084
rect 25784 32018 25796 32074
rect 25852 32018 26229 32074
rect 26285 32018 26297 32074
rect 25784 32016 25864 32018
rect 26227 32006 26297 32018
rect 13641 31957 13711 31969
rect 14681 31957 14761 31959
rect 16167 31958 16247 31960
rect 13641 31901 13653 31957
rect 13709 31901 14693 31957
rect 14749 31901 14761 31957
rect 13641 31889 13711 31901
rect 9993 30850 10157 30862
rect 10473 30928 10637 30940
rect 10473 30872 10485 30928
rect 10541 30872 10637 30928
rect 10473 30860 10637 30872
rect 9993 30794 10005 30850
rect 10061 30794 10157 30850
rect 9993 30782 10157 30794
rect 10061 30732 10157 30782
rect 8958 30710 9004 30721
rect 8064 30410 8110 30550
rect 8279 30419 8375 30450
rect 8279 30373 8290 30419
rect 8364 30373 8375 30419
rect 8544 30410 8590 30550
rect 8110 30327 8248 30338
rect 8110 29753 8202 30327
rect 8406 30327 8452 30338
rect 8389 30043 8406 30053
rect 8452 30043 8469 30053
rect 8389 29803 8401 30043
rect 8457 29803 8469 30043
rect 8389 29793 8406 29803
rect 8110 29742 8248 29753
rect 8452 29793 8469 29803
rect 8406 29742 8452 29753
rect 8064 29659 8110 29670
rect 8279 29661 8290 29707
rect 8364 29661 8375 29707
rect 8279 29520 8375 29661
rect 9173 30719 9473 30732
rect 9173 30673 9184 30719
rect 9258 30686 9388 30719
rect 9258 30673 9269 30686
rect 9377 30673 9388 30686
rect 9462 30673 9473 30719
rect 9642 30710 9688 30721
rect 9004 30627 9142 30638
rect 9004 30453 9096 30627
rect 9300 30627 9346 30638
rect 9283 30568 9300 30578
rect 9504 30627 9642 30638
rect 9346 30568 9363 30578
rect 9283 30512 9295 30568
rect 9351 30512 9363 30568
rect 9283 30502 9300 30512
rect 9004 30442 9142 30453
rect 9346 30502 9363 30512
rect 9300 30442 9346 30453
rect 9550 30453 9642 30627
rect 9504 30442 9642 30453
rect 8958 30230 9004 30370
rect 9173 30361 9184 30407
rect 9258 30361 9269 30407
rect 9173 30330 9269 30361
rect 9377 30361 9388 30407
rect 9462 30361 9473 30407
rect 9377 30330 9473 30361
rect 9857 30719 10157 30732
rect 9857 30673 9868 30719
rect 9942 30686 10072 30719
rect 9942 30673 9953 30686
rect 10061 30673 10072 30686
rect 10146 30673 10157 30719
rect 10326 30710 10372 30721
rect 9780 30627 9826 30638
rect 9763 30568 9780 30578
rect 9984 30627 10030 30638
rect 9826 30568 9843 30578
rect 9763 30512 9775 30568
rect 9831 30512 9843 30568
rect 9763 30502 9780 30512
rect 9826 30502 9843 30512
rect 9967 30568 9984 30578
rect 10188 30627 10234 30638
rect 10030 30568 10047 30578
rect 9967 30512 9979 30568
rect 10035 30512 10047 30568
rect 9967 30502 9984 30512
rect 9780 30442 9826 30453
rect 10030 30502 10047 30512
rect 10171 30568 10188 30578
rect 10234 30568 10251 30578
rect 10171 30512 10183 30568
rect 10239 30512 10251 30568
rect 10171 30502 10188 30512
rect 9984 30442 10030 30453
rect 10234 30502 10251 30512
rect 10188 30442 10234 30453
rect 9642 30230 9688 30370
rect 9857 30361 9868 30407
rect 9942 30361 9953 30407
rect 9857 30330 9953 30361
rect 10061 30361 10072 30407
rect 10146 30361 10157 30407
rect 10061 30330 10157 30361
rect 10541 30719 10637 30860
rect 11149 30974 13117 31170
rect 13925 31170 13981 31901
rect 14681 31899 14761 31901
rect 15411 31902 16179 31958
rect 16235 31902 16247 31958
rect 14313 31807 14393 31821
rect 14100 31785 14146 31796
rect 14313 31751 14325 31807
rect 14381 31751 14393 31807
rect 14497 31807 14577 31821
rect 14497 31751 14509 31807
rect 14565 31751 14577 31807
rect 14681 31807 14761 31821
rect 14681 31751 14693 31807
rect 14749 31751 14761 31807
rect 14928 31785 14974 31796
rect 14315 31748 14326 31751
rect 14380 31748 14391 31751
rect 14499 31748 14510 31751
rect 14564 31748 14575 31751
rect 14683 31748 14694 31751
rect 14748 31748 14759 31751
rect 14238 31702 14284 31713
rect 14146 31528 14238 31702
rect 14238 31517 14284 31528
rect 14422 31702 14468 31713
rect 14422 31517 14468 31528
rect 14606 31702 14652 31713
rect 14790 31702 14836 31713
rect 14773 31675 14790 31677
rect 14836 31675 14853 31677
rect 14773 31555 14785 31675
rect 14841 31555 14853 31675
rect 14773 31553 14790 31555
rect 14606 31517 14652 31528
rect 14836 31553 14853 31555
rect 14790 31517 14836 31528
rect 14100 31300 14146 31445
rect 14315 31436 14326 31482
rect 14380 31436 14391 31482
rect 14315 31403 14391 31436
rect 14499 31436 14510 31482
rect 14564 31436 14575 31482
rect 14499 31403 14575 31436
rect 14683 31436 14694 31482
rect 14748 31436 14759 31482
rect 14683 31403 14759 31436
rect 14928 31300 14974 31445
rect 14088 31288 14168 31300
rect 14088 31232 14100 31288
rect 14156 31232 14168 31288
rect 14088 31220 14168 31232
rect 14906 31288 14984 31300
rect 14906 31232 14918 31288
rect 14974 31232 14984 31288
rect 14906 31220 14984 31232
rect 15259 31170 15339 31180
rect 13925 31114 15271 31170
rect 15327 31114 15339 31170
rect 15259 31112 15339 31114
rect 15093 31061 15163 31063
rect 11149 30834 11249 30974
rect 13017 30834 13117 30974
rect 11149 30794 13117 30834
rect 13925 31060 15163 31061
rect 13925 31006 15095 31060
rect 15151 31006 15163 31060
rect 13925 31005 15163 31006
rect 10541 30673 10552 30719
rect 10626 30673 10637 30719
rect 10806 30710 10852 30721
rect 10372 30627 10510 30638
rect 10372 30453 10464 30627
rect 10668 30627 10714 30638
rect 10651 30568 10668 30578
rect 10714 30568 10731 30578
rect 10651 30512 10663 30568
rect 10719 30512 10731 30568
rect 10651 30502 10668 30512
rect 10372 30442 10510 30453
rect 10714 30502 10731 30512
rect 10668 30442 10714 30453
rect 10326 30230 10372 30370
rect 10541 30361 10552 30407
rect 10626 30361 10637 30407
rect 10541 30330 10637 30361
rect 10806 30230 10852 30370
rect 11186 30654 11232 30794
rect 8921 30200 10889 30230
rect 8921 30060 10189 30200
rect 10789 30060 10889 30200
rect 8921 30030 10889 30060
rect 11401 30663 11497 30694
rect 11401 30617 11412 30663
rect 11486 30617 11497 30663
rect 11605 30663 11701 30694
rect 11605 30617 11616 30663
rect 11690 30617 11701 30663
rect 11870 30654 11916 30794
rect 11232 30571 11370 30582
rect 11528 30571 11574 30582
rect 11732 30571 11870 30582
rect 11232 29997 11324 30571
rect 11511 30331 11523 30571
rect 11579 30331 11591 30571
rect 11232 29986 11370 29997
rect 11528 29986 11574 29997
rect 11778 29997 11870 30571
rect 11732 29986 11870 29997
rect 11186 29903 11232 29914
rect 11401 29905 11412 29951
rect 11486 29931 11497 29951
rect 11605 29931 11616 29951
rect 11486 29905 11616 29931
rect 11690 29905 11701 29951
rect 11401 29878 11701 29905
rect 12085 30663 12181 30694
rect 12085 30617 12096 30663
rect 12170 30617 12181 30663
rect 12289 30663 12385 30694
rect 12289 30617 12300 30663
rect 12374 30617 12385 30663
rect 12554 30654 12600 30794
rect 12008 30571 12054 30582
rect 12212 30571 12258 30582
rect 12416 30571 12462 30582
rect 12195 30331 12207 30571
rect 12263 30331 12275 30571
rect 11991 29997 12003 30237
rect 12059 29997 12071 30237
rect 12399 29997 12411 30237
rect 12467 29997 12479 30237
rect 12008 29986 12054 29997
rect 12212 29986 12258 29997
rect 12416 29986 12462 29997
rect 11870 29903 11916 29914
rect 12085 29905 12096 29951
rect 12170 29931 12181 29951
rect 12289 29931 12300 29951
rect 12170 29905 12300 29931
rect 12374 29905 12385 29951
rect 12085 29878 12385 29905
rect 12769 30663 12865 30694
rect 12769 30617 12780 30663
rect 12854 30617 12865 30663
rect 13034 30654 13080 30794
rect 12600 30571 12738 30582
rect 12600 29997 12692 30571
rect 12896 30571 12942 30582
rect 12879 30287 12896 30297
rect 12942 30287 12959 30297
rect 12879 30047 12891 30287
rect 12947 30047 12959 30287
rect 12879 30037 12896 30047
rect 12600 29986 12738 29997
rect 12942 30037 12959 30047
rect 12896 29986 12942 29997
rect 12554 29903 12600 29914
rect 12769 29905 12780 29951
rect 12854 29905 12865 29951
rect 11401 29830 11497 29878
rect 8544 29659 8590 29670
rect 8921 29800 10889 29830
rect 8921 29660 10189 29800
rect 10789 29660 10889 29800
rect 8921 29630 10889 29660
rect 11401 29774 11421 29830
rect 11477 29774 11497 29830
rect 8211 29508 8375 29520
rect 8211 29452 8223 29508
rect 8279 29452 8375 29508
rect 8211 29440 8375 29452
rect 3850 28908 3862 28964
rect 3918 28908 4045 28964
rect 4101 28908 5995 28964
rect 8064 29290 8110 29301
rect 8279 29299 8375 29440
rect 8958 29490 9004 29501
rect 8279 29253 8290 29299
rect 8364 29253 8375 29299
rect 8544 29290 8590 29301
rect 8110 29207 8248 29218
rect 8110 29033 8202 29207
rect 8406 29207 8452 29218
rect 8389 29148 8406 29158
rect 8452 29148 8469 29158
rect 8389 29092 8401 29148
rect 8457 29092 8469 29148
rect 8389 29082 8406 29092
rect 8110 29022 8248 29033
rect 8452 29082 8469 29092
rect 8406 29022 8452 29033
rect 3850 28896 3936 28908
rect 4043 28896 4103 28908
rect 521 28509 685 28521
rect 1001 28587 1165 28599
rect 1001 28531 1013 28587
rect 1069 28531 1165 28587
rect 1001 28519 1165 28531
rect 521 28453 533 28509
rect 589 28453 685 28509
rect 521 28441 685 28453
rect 589 28391 685 28441
rect -6027 27889 -845 28089
rect -514 28369 -468 28380
rect -299 28378 1 28391
rect -299 28332 -288 28378
rect -214 28345 -84 28378
rect -214 28332 -203 28345
rect -95 28332 -84 28345
rect -10 28332 1 28378
rect 170 28369 216 28380
rect -468 28286 -330 28297
rect -468 28112 -376 28286
rect -172 28286 -126 28297
rect -189 28227 -172 28237
rect 32 28286 170 28297
rect -126 28227 -109 28237
rect -189 28171 -177 28227
rect -121 28171 -109 28227
rect -189 28161 -172 28171
rect -468 28101 -330 28112
rect -126 28161 -109 28171
rect -172 28101 -126 28112
rect 78 28112 170 28286
rect 32 28101 170 28112
rect -514 27889 -468 28029
rect -299 28020 -288 28066
rect -214 28020 -203 28066
rect -299 27989 -203 28020
rect -95 28020 -84 28066
rect -10 28020 1 28066
rect -95 27989 1 28020
rect 385 28378 685 28391
rect 385 28332 396 28378
rect 470 28345 600 28378
rect 470 28332 481 28345
rect 589 28332 600 28345
rect 674 28332 685 28378
rect 854 28369 900 28380
rect 308 28286 354 28297
rect 291 28227 308 28237
rect 512 28286 558 28297
rect 354 28227 371 28237
rect 291 28171 303 28227
rect 359 28171 371 28227
rect 291 28161 308 28171
rect 354 28161 371 28171
rect 495 28227 512 28237
rect 716 28286 762 28297
rect 558 28227 575 28237
rect 495 28171 507 28227
rect 563 28171 575 28227
rect 495 28161 512 28171
rect 308 28101 354 28112
rect 558 28161 575 28171
rect 699 28227 716 28237
rect 762 28227 779 28237
rect 699 28171 711 28227
rect 767 28171 779 28227
rect 699 28161 716 28171
rect 512 28101 558 28112
rect 762 28161 779 28171
rect 716 28101 762 28112
rect 170 27889 216 28029
rect 385 28020 396 28066
rect 470 28020 481 28066
rect 385 27989 481 28020
rect 589 28020 600 28066
rect 674 28020 685 28066
rect 589 27989 685 28020
rect 1069 28378 1165 28519
rect 1677 28689 3645 28873
rect 8064 28810 8110 28950
rect 8279 28941 8290 28987
rect 8364 28941 8375 28987
rect 8279 28910 8375 28941
rect 8544 28810 8590 28950
rect 1069 28332 1080 28378
rect 1154 28332 1165 28378
rect 1334 28369 1380 28380
rect 900 28286 1038 28297
rect 900 28112 992 28286
rect 1196 28286 1242 28297
rect 1179 28227 1196 28237
rect 1242 28227 1259 28237
rect 1179 28171 1191 28227
rect 1247 28171 1259 28227
rect 1179 28161 1196 28171
rect 900 28101 1038 28112
rect 1242 28161 1259 28171
rect 1196 28101 1242 28112
rect 854 27889 900 28029
rect 1069 28020 1080 28066
rect 1154 28020 1165 28066
rect 1069 27989 1165 28020
rect 1334 27889 1380 28029
rect 1677 27889 3145 28689
rect 3445 28089 3645 28689
rect 8027 28089 8627 28810
rect 9173 29499 9269 29530
rect 9173 29453 9184 29499
rect 9258 29453 9269 29499
rect 9438 29490 9892 29630
rect 9096 29407 9142 29418
rect 9079 29123 9096 29133
rect 9300 29407 9438 29418
rect 9142 29123 9159 29133
rect 9079 28883 9091 29123
rect 9147 28883 9159 29123
rect 9079 28873 9096 28883
rect 9142 28873 9159 28883
rect 9096 28822 9142 28833
rect 9346 28833 9438 29407
rect 9300 28822 9438 28833
rect 8958 28739 9004 28750
rect 9173 28741 9184 28787
rect 9258 28741 9269 28787
rect 9173 28666 9269 28741
rect 9484 28822 9846 29490
rect 9438 28739 9484 28750
rect 10061 29499 10157 29530
rect 10061 29453 10072 29499
rect 10146 29453 10157 29499
rect 10326 29490 10372 29630
rect 9892 29407 10030 29418
rect 9892 28833 9984 29407
rect 10188 29407 10234 29418
rect 10171 29123 10188 29133
rect 10234 29123 10251 29133
rect 10171 28883 10183 29123
rect 10239 28883 10251 29123
rect 10171 28873 10188 28883
rect 9892 28822 10030 28833
rect 10234 28873 10251 28883
rect 10188 28822 10234 28833
rect 9846 28739 9892 28750
rect 10061 28741 10072 28787
rect 10146 28741 10157 28787
rect 9173 28610 9193 28666
rect 9249 28610 9269 28666
rect 9173 28392 9269 28610
rect 10061 28522 10157 28741
rect 10541 29499 10637 29530
rect 10541 29453 10552 29499
rect 10626 29453 10637 29499
rect 10806 29490 10852 29630
rect 10372 29407 10510 29418
rect 10372 28833 10464 29407
rect 10668 29407 10714 29418
rect 10651 29123 10668 29133
rect 10714 29123 10731 29133
rect 10651 28883 10663 29123
rect 10719 28883 10731 29123
rect 10651 28873 10668 28883
rect 10372 28822 10510 28833
rect 10714 28873 10731 28883
rect 10668 28822 10714 28833
rect 10326 28739 10372 28750
rect 10541 28741 10552 28787
rect 10626 28741 10637 28787
rect 10541 28600 10637 28741
rect 11186 29534 11232 29545
rect 11401 29543 11497 29774
rect 12085 29674 12181 29878
rect 12769 29764 12865 29905
rect 13925 29984 13981 31005
rect 15093 30997 15163 31005
rect 14589 30953 14675 30957
rect 14589 30897 14601 30953
rect 14657 30897 14675 30953
rect 14589 30885 14675 30897
rect 14100 30740 14146 30751
rect 14315 30749 14391 30782
rect 14315 30703 14326 30749
rect 14380 30703 14391 30749
rect 14499 30749 14575 30782
rect 14499 30703 14510 30749
rect 14564 30703 14575 30749
rect 14683 30749 14759 30782
rect 14683 30703 14694 30749
rect 14748 30703 14759 30749
rect 14928 30740 14974 30751
rect 14238 30657 14284 30668
rect 14221 30630 14238 30632
rect 14422 30657 14468 30668
rect 14284 30630 14301 30632
rect 14146 30510 14233 30630
rect 14289 30510 14301 30630
rect 14221 30508 14238 30510
rect 14146 30210 14238 30330
rect 14284 30508 14301 30510
rect 14405 30330 14422 30332
rect 14606 30657 14652 30668
rect 14589 30630 14606 30632
rect 14790 30657 14836 30668
rect 14652 30630 14669 30632
rect 14589 30510 14601 30630
rect 14657 30510 14669 30630
rect 14589 30508 14606 30510
rect 14468 30330 14485 30332
rect 14405 30210 14417 30330
rect 14473 30210 14485 30330
rect 14405 30208 14422 30210
rect 14238 30172 14284 30183
rect 14468 30208 14485 30210
rect 14422 30172 14468 30183
rect 14652 30508 14669 30510
rect 14773 30330 14790 30332
rect 14911 30630 14928 30632
rect 14974 30630 14991 30632
rect 14911 30509 14923 30630
rect 14979 30509 14991 30630
rect 14911 30507 14928 30509
rect 14836 30330 14853 30332
rect 14773 30210 14785 30330
rect 14841 30210 14853 30330
rect 14773 30208 14790 30210
rect 14606 30172 14652 30183
rect 14836 30208 14853 30210
rect 14790 30172 14836 30183
rect 14315 30134 14326 30137
rect 14380 30134 14391 30137
rect 14499 30134 14510 30137
rect 14564 30134 14575 30137
rect 14683 30134 14694 30137
rect 14748 30134 14759 30137
rect 14100 30089 14146 30100
rect 14313 30078 14325 30134
rect 14381 30078 14393 30134
rect 14313 30064 14393 30078
rect 14497 30078 14509 30134
rect 14565 30078 14577 30134
rect 14497 30064 14577 30078
rect 14681 30078 14693 30134
rect 14749 30078 14761 30134
rect 14974 30507 14991 30509
rect 14928 30089 14974 30100
rect 14681 30064 14761 30078
rect 14313 29984 14393 29986
rect 13925 29928 14325 29984
rect 14381 29928 14393 29984
rect 14313 29926 14393 29928
rect 13034 29903 13080 29914
rect 13505 29868 13575 29882
rect 14497 29868 14577 29870
rect 13505 29812 13517 29868
rect 13573 29812 14509 29868
rect 14565 29812 14577 29868
rect 13505 29800 13575 29812
rect 14497 29810 14577 29812
rect 14826 29868 14906 29870
rect 15269 29868 15329 29880
rect 14826 29812 14838 29868
rect 14894 29812 15271 29868
rect 15327 29812 15329 29868
rect 14826 29810 14906 29812
rect 15269 29800 15329 29812
rect 12701 29752 12865 29764
rect 12701 29696 12713 29752
rect 12769 29696 12865 29752
rect 12701 29684 12865 29696
rect 13271 29752 13349 29763
rect 14681 29752 14761 29754
rect 13271 29751 14693 29752
rect 13271 29697 13283 29751
rect 13337 29697 14693 29751
rect 13271 29696 14693 29697
rect 14749 29696 14761 29752
rect 13271 29685 13349 29696
rect 14681 29694 14761 29696
rect 12085 29618 12105 29674
rect 12161 29618 12181 29674
rect 11401 29497 11412 29543
rect 11486 29497 11497 29543
rect 11666 29534 11916 29545
rect 11324 29451 11370 29462
rect 11307 29392 11324 29402
rect 11528 29451 11666 29462
rect 11370 29392 11387 29402
rect 11307 29336 11319 29392
rect 11375 29336 11387 29392
rect 11307 29326 11324 29336
rect 11370 29326 11387 29336
rect 11324 29266 11370 29277
rect 11574 29277 11666 29451
rect 11528 29266 11666 29277
rect 11186 29054 11232 29194
rect 11401 29185 11412 29231
rect 11486 29185 11497 29231
rect 11401 29154 11497 29185
rect 11712 29194 11870 29534
rect 12085 29543 12181 29618
rect 12085 29497 12096 29543
rect 12170 29497 12181 29543
rect 12350 29534 12396 29545
rect 11916 29451 12054 29462
rect 11916 29277 12008 29451
rect 12212 29451 12258 29462
rect 12195 29392 12212 29402
rect 12258 29392 12275 29402
rect 12195 29336 12207 29392
rect 12263 29336 12275 29392
rect 12195 29326 12212 29336
rect 11916 29266 12054 29277
rect 12258 29326 12275 29336
rect 12212 29266 12258 29277
rect 11666 29183 11916 29194
rect 12085 29185 12096 29231
rect 12170 29185 12181 29231
rect 11712 29054 11870 29183
rect 12085 29154 12181 29185
rect 12350 29054 12396 29194
rect 12554 29534 12600 29545
rect 12769 29543 12865 29684
rect 14313 29602 14393 29616
rect 14100 29580 14146 29591
rect 12769 29497 12780 29543
rect 12854 29497 12865 29543
rect 13034 29534 13080 29545
rect 12600 29451 12738 29462
rect 12600 29277 12692 29451
rect 12896 29451 12942 29462
rect 12879 29392 12896 29402
rect 12942 29392 12959 29402
rect 12879 29336 12891 29392
rect 12947 29336 12959 29392
rect 12879 29326 12896 29336
rect 12600 29266 12738 29277
rect 12942 29326 12959 29336
rect 12896 29266 12942 29277
rect 12554 29054 12600 29194
rect 12769 29185 12780 29231
rect 12854 29185 12865 29231
rect 12769 29154 12865 29185
rect 13034 29054 13080 29194
rect 14313 29546 14325 29602
rect 14381 29546 14393 29602
rect 14497 29602 14577 29616
rect 14497 29546 14509 29602
rect 14565 29546 14577 29602
rect 14681 29602 14761 29616
rect 14681 29546 14693 29602
rect 14749 29546 14761 29602
rect 14928 29580 14974 29591
rect 14315 29543 14326 29546
rect 14380 29543 14391 29546
rect 14499 29543 14510 29546
rect 14564 29543 14575 29546
rect 14683 29543 14694 29546
rect 14748 29543 14759 29546
rect 14238 29497 14284 29508
rect 14146 29323 14238 29497
rect 14238 29312 14284 29323
rect 14422 29497 14468 29508
rect 14422 29312 14468 29323
rect 14606 29497 14652 29508
rect 14790 29497 14836 29508
rect 14773 29470 14790 29472
rect 14836 29470 14853 29472
rect 14773 29350 14785 29470
rect 14841 29350 14853 29470
rect 14773 29348 14790 29350
rect 14606 29312 14652 29323
rect 14836 29348 14853 29350
rect 14790 29312 14836 29323
rect 14100 29095 14146 29240
rect 14315 29231 14326 29277
rect 14380 29231 14391 29277
rect 14315 29198 14391 29231
rect 14499 29231 14510 29277
rect 14564 29231 14575 29277
rect 14499 29198 14575 29231
rect 14683 29231 14694 29277
rect 14748 29231 14759 29277
rect 14683 29198 14759 29231
rect 14928 29095 14974 29240
rect 14088 29083 14168 29095
rect 10806 28739 10852 28750
rect 11149 29014 13117 29054
rect 14088 29027 14100 29083
rect 14156 29027 14168 29083
rect 14088 29015 14168 29027
rect 14906 29083 14986 29095
rect 14906 29027 14918 29083
rect 14974 29027 14986 29083
rect 14906 29015 14986 29027
rect 11149 28874 11249 29014
rect 13017 28874 13117 29014
rect 13322 28965 13408 28977
rect 13515 28965 13575 28969
rect 15411 28965 15467 31902
rect 16167 31900 16247 31902
rect 15799 31808 15879 31822
rect 15586 31786 15632 31797
rect 15799 31752 15811 31808
rect 15867 31752 15879 31808
rect 15983 31808 16063 31822
rect 15983 31752 15995 31808
rect 16051 31752 16063 31808
rect 16167 31808 16247 31822
rect 16167 31752 16179 31808
rect 16235 31752 16247 31808
rect 16414 31786 16460 31797
rect 15801 31749 15812 31752
rect 15866 31749 15877 31752
rect 15985 31749 15996 31752
rect 16050 31749 16061 31752
rect 16169 31749 16180 31752
rect 16234 31749 16245 31752
rect 15724 31703 15770 31714
rect 15632 31529 15724 31703
rect 15724 31518 15770 31529
rect 15908 31703 15954 31714
rect 15908 31518 15954 31529
rect 16092 31703 16138 31714
rect 16276 31703 16322 31714
rect 16259 31676 16276 31678
rect 16322 31676 16339 31678
rect 16259 31556 16271 31676
rect 16327 31556 16339 31676
rect 16259 31554 16276 31556
rect 16092 31518 16138 31529
rect 16322 31554 16339 31556
rect 16276 31518 16322 31529
rect 15586 31301 15632 31446
rect 15801 31437 15812 31483
rect 15866 31437 15877 31483
rect 15801 31404 15877 31437
rect 15985 31437 15996 31483
rect 16050 31437 16061 31483
rect 15985 31404 16061 31437
rect 16169 31437 16180 31483
rect 16234 31437 16245 31483
rect 16169 31404 16245 31437
rect 16414 31301 16460 31446
rect 15574 31289 15654 31301
rect 15574 31233 15586 31289
rect 15642 31233 15654 31289
rect 15574 31221 15654 31233
rect 16392 31289 16470 31301
rect 16392 31233 16404 31289
rect 16460 31233 16470 31289
rect 16392 31221 16470 31233
rect 17499 31170 17699 31970
rect 17899 31170 18099 31970
rect 17499 30550 18099 31170
rect 18430 31830 18476 31841
rect 18645 31839 18741 31870
rect 18645 31793 18656 31839
rect 18730 31793 18741 31839
rect 18910 31830 19364 31970
rect 18568 31747 18614 31758
rect 18551 31463 18568 31473
rect 18772 31747 18910 31758
rect 18614 31463 18631 31473
rect 18551 31223 18563 31463
rect 18619 31223 18631 31463
rect 18551 31213 18568 31223
rect 18614 31213 18631 31223
rect 18568 31162 18614 31173
rect 18818 31173 18910 31747
rect 18772 31162 18910 31173
rect 18430 31079 18476 31090
rect 18645 31081 18656 31127
rect 18730 31081 18741 31127
rect 18645 31006 18741 31081
rect 18956 31162 19318 31830
rect 18910 31079 18956 31090
rect 19533 31839 19629 31870
rect 19533 31793 19544 31839
rect 19618 31793 19629 31839
rect 19798 31830 19844 31970
rect 19364 31747 19502 31758
rect 19364 31173 19456 31747
rect 19660 31747 19706 31758
rect 19643 31463 19660 31473
rect 19706 31463 19723 31473
rect 19643 31223 19655 31463
rect 19711 31223 19723 31463
rect 19643 31213 19660 31223
rect 19364 31162 19502 31173
rect 19706 31213 19723 31223
rect 19660 31162 19706 31173
rect 19318 31079 19364 31090
rect 19533 31081 19544 31127
rect 19618 31081 19629 31127
rect 18645 30950 18665 31006
rect 18721 30950 18741 31006
rect 18645 30732 18741 30950
rect 19533 30862 19629 31081
rect 20013 31839 20109 31870
rect 20013 31793 20024 31839
rect 20098 31793 20109 31839
rect 20278 31830 20324 31970
rect 19844 31747 19982 31758
rect 19844 31173 19936 31747
rect 20140 31747 20186 31758
rect 20123 31463 20140 31473
rect 20186 31463 20203 31473
rect 20123 31223 20135 31463
rect 20191 31223 20203 31463
rect 20123 31213 20140 31223
rect 19844 31162 19982 31173
rect 20186 31213 20203 31223
rect 20140 31162 20186 31173
rect 19798 31079 19844 31090
rect 20013 31081 20024 31127
rect 20098 31081 20109 31127
rect 20013 30940 20109 31081
rect 20278 31079 20324 31090
rect 20621 31170 22089 31970
rect 22389 31170 22589 31970
rect 26971 31970 32061 32170
rect 32733 32073 32789 33320
rect 35689 33318 35769 33320
rect 41639 33376 41721 33388
rect 42205 33376 42261 34106
rect 43097 34104 43177 34106
rect 43827 34106 44595 34162
rect 44651 34106 44663 34162
rect 42729 34012 42809 34026
rect 42516 33990 42562 34001
rect 42729 33956 42741 34012
rect 42797 33956 42809 34012
rect 42913 34012 42993 34026
rect 42913 33956 42925 34012
rect 42981 33956 42993 34012
rect 43097 34012 43177 34026
rect 43097 33956 43109 34012
rect 43165 33956 43177 34012
rect 43344 33990 43390 34001
rect 42731 33953 42742 33956
rect 42796 33953 42807 33956
rect 42915 33953 42926 33956
rect 42980 33953 42991 33956
rect 43099 33953 43110 33956
rect 43164 33953 43175 33956
rect 42654 33907 42700 33918
rect 42562 33733 42654 33907
rect 42654 33722 42700 33733
rect 42838 33907 42884 33918
rect 42838 33722 42884 33733
rect 43022 33907 43068 33918
rect 43206 33907 43252 33918
rect 43189 33880 43206 33882
rect 43252 33880 43269 33882
rect 43189 33760 43201 33880
rect 43257 33760 43269 33880
rect 43189 33758 43206 33760
rect 43022 33722 43068 33733
rect 43252 33758 43269 33760
rect 43206 33722 43252 33733
rect 42516 33505 42562 33650
rect 42731 33641 42742 33687
rect 42796 33641 42807 33687
rect 42731 33608 42807 33641
rect 42915 33641 42926 33687
rect 42980 33641 42991 33687
rect 42915 33608 42991 33641
rect 43099 33641 43110 33687
rect 43164 33641 43175 33687
rect 43099 33608 43175 33641
rect 43344 33505 43390 33650
rect 42504 33493 42584 33505
rect 42504 33437 42516 33493
rect 42572 33437 42584 33493
rect 42504 33425 42584 33437
rect 43322 33493 43400 33505
rect 43322 33437 43334 33493
rect 43390 33437 43400 33493
rect 43322 33425 43400 33437
rect 41639 33320 41653 33376
rect 41709 33320 42261 33376
rect 43827 33376 43883 34106
rect 44583 34104 44663 34106
rect 44215 34012 44295 34026
rect 44002 33990 44048 34001
rect 44215 33956 44227 34012
rect 44283 33956 44295 34012
rect 44399 34012 44479 34026
rect 44399 33956 44411 34012
rect 44467 33956 44479 34012
rect 44583 34012 44663 34026
rect 44583 33956 44595 34012
rect 44651 33956 44663 34012
rect 44830 33990 44876 34001
rect 44217 33953 44228 33956
rect 44282 33953 44293 33956
rect 44401 33953 44412 33956
rect 44466 33953 44477 33956
rect 44585 33953 44596 33956
rect 44650 33953 44661 33956
rect 44140 33907 44186 33918
rect 44048 33733 44140 33907
rect 44140 33722 44186 33733
rect 44324 33907 44370 33918
rect 44324 33722 44370 33733
rect 44508 33907 44554 33918
rect 44692 33907 44738 33918
rect 44675 33880 44692 33882
rect 44738 33880 44755 33882
rect 44675 33760 44687 33880
rect 44743 33760 44755 33880
rect 44675 33758 44692 33760
rect 44508 33722 44554 33733
rect 44738 33758 44755 33760
rect 44692 33722 44738 33733
rect 44002 33505 44048 33650
rect 44217 33641 44228 33687
rect 44282 33641 44293 33687
rect 44217 33608 44293 33641
rect 44401 33641 44412 33687
rect 44466 33641 44477 33687
rect 44401 33608 44477 33641
rect 44585 33641 44596 33687
rect 44650 33641 44661 33687
rect 44585 33608 44661 33641
rect 44830 33505 44876 33650
rect 43990 33493 44070 33505
rect 43990 33437 44002 33493
rect 44058 33437 44070 33493
rect 43990 33425 44070 33437
rect 44808 33493 44886 33505
rect 44808 33437 44820 33493
rect 44876 33437 44886 33493
rect 44808 33425 44886 33437
rect 45161 33376 45241 33386
rect 43827 33320 45173 33376
rect 45229 33320 45241 33376
rect 41639 33308 41721 33320
rect 34213 33265 34283 33267
rect 35513 33266 35593 33268
rect 32869 33209 34215 33265
rect 34271 33209 34283 33265
rect 32869 32189 32925 33209
rect 34213 33197 34283 33209
rect 34355 33210 35525 33266
rect 35581 33210 35593 33266
rect 33533 33158 33619 33162
rect 33533 33102 33545 33158
rect 33601 33102 33619 33158
rect 33533 33090 33619 33102
rect 33044 32945 33090 32956
rect 33259 32954 33335 32987
rect 33259 32908 33270 32954
rect 33324 32908 33335 32954
rect 33443 32954 33519 32987
rect 33443 32908 33454 32954
rect 33508 32908 33519 32954
rect 33627 32954 33703 32987
rect 33627 32908 33638 32954
rect 33692 32908 33703 32954
rect 33872 32945 33918 32956
rect 33182 32862 33228 32873
rect 33165 32835 33182 32837
rect 33366 32862 33412 32873
rect 33228 32835 33245 32837
rect 33090 32715 33177 32835
rect 33233 32715 33245 32835
rect 33165 32713 33182 32715
rect 33090 32415 33182 32535
rect 33228 32713 33245 32715
rect 33349 32535 33366 32537
rect 33550 32862 33596 32873
rect 33533 32835 33550 32837
rect 33734 32862 33780 32873
rect 33596 32835 33613 32837
rect 33533 32715 33545 32835
rect 33601 32715 33613 32835
rect 33533 32713 33550 32715
rect 33412 32535 33429 32537
rect 33349 32415 33361 32535
rect 33417 32415 33429 32535
rect 33349 32413 33366 32415
rect 33182 32377 33228 32388
rect 33412 32413 33429 32415
rect 33366 32377 33412 32388
rect 33596 32713 33613 32715
rect 33717 32535 33734 32537
rect 33855 32835 33872 32837
rect 33918 32835 33935 32837
rect 33855 32714 33867 32835
rect 33923 32714 33935 32835
rect 33855 32712 33872 32714
rect 33780 32535 33797 32537
rect 33717 32415 33729 32535
rect 33785 32415 33797 32535
rect 33717 32413 33734 32415
rect 33550 32377 33596 32388
rect 33780 32413 33797 32415
rect 33734 32377 33780 32388
rect 33259 32339 33270 32342
rect 33324 32339 33335 32342
rect 33443 32339 33454 32342
rect 33508 32339 33519 32342
rect 33627 32339 33638 32342
rect 33692 32339 33703 32342
rect 33044 32294 33090 32305
rect 33257 32283 33269 32339
rect 33325 32283 33337 32339
rect 33257 32269 33337 32283
rect 33441 32283 33453 32339
rect 33509 32283 33521 32339
rect 33441 32269 33521 32283
rect 33625 32283 33637 32339
rect 33693 32283 33705 32339
rect 33918 32712 33935 32714
rect 33872 32294 33918 32305
rect 33625 32269 33705 32283
rect 33257 32189 33337 32191
rect 32869 32133 33269 32189
rect 33325 32133 33337 32189
rect 34355 32190 34411 33210
rect 35513 33198 35593 33210
rect 35019 33159 35105 33163
rect 35019 33103 35031 33159
rect 35087 33103 35105 33159
rect 35019 33091 35105 33103
rect 34530 32946 34576 32957
rect 34745 32955 34821 32988
rect 34745 32909 34756 32955
rect 34810 32909 34821 32955
rect 34929 32955 35005 32988
rect 34929 32909 34940 32955
rect 34994 32909 35005 32955
rect 35113 32955 35189 32988
rect 35113 32909 35124 32955
rect 35178 32909 35189 32955
rect 35358 32946 35404 32957
rect 34668 32863 34714 32874
rect 34651 32836 34668 32838
rect 34852 32863 34898 32874
rect 34714 32836 34731 32838
rect 34576 32716 34663 32836
rect 34719 32716 34731 32836
rect 34651 32714 34668 32716
rect 34576 32416 34668 32536
rect 34714 32714 34731 32716
rect 34835 32536 34852 32538
rect 35036 32863 35082 32874
rect 35019 32836 35036 32838
rect 35220 32863 35266 32874
rect 35082 32836 35099 32838
rect 35019 32716 35031 32836
rect 35087 32716 35099 32836
rect 35019 32714 35036 32716
rect 34898 32536 34915 32538
rect 34835 32416 34847 32536
rect 34903 32416 34915 32536
rect 34835 32414 34852 32416
rect 34668 32378 34714 32389
rect 34898 32414 34915 32416
rect 34852 32378 34898 32389
rect 35082 32714 35099 32716
rect 35203 32536 35220 32538
rect 35341 32836 35358 32838
rect 35404 32836 35421 32838
rect 35341 32715 35353 32836
rect 35409 32715 35421 32836
rect 35341 32713 35358 32715
rect 35266 32536 35283 32538
rect 35203 32416 35215 32536
rect 35271 32416 35283 32536
rect 35203 32414 35220 32416
rect 35036 32378 35082 32389
rect 35266 32414 35283 32416
rect 35220 32378 35266 32389
rect 34745 32340 34756 32343
rect 34810 32340 34821 32343
rect 34929 32340 34940 32343
rect 34994 32340 35005 32343
rect 35113 32340 35124 32343
rect 35178 32340 35189 32343
rect 34530 32295 34576 32306
rect 34743 32284 34755 32340
rect 34811 32284 34823 32340
rect 34743 32270 34823 32284
rect 34927 32284 34939 32340
rect 34995 32284 35007 32340
rect 34927 32270 35007 32284
rect 35111 32284 35123 32340
rect 35179 32284 35191 32340
rect 35404 32713 35421 32715
rect 35358 32295 35404 32306
rect 35111 32270 35191 32284
rect 34743 32190 34823 32192
rect 34355 32134 34755 32190
rect 34811 32134 34823 32190
rect 33257 32131 33337 32133
rect 34743 32132 34823 32134
rect 33441 32073 33521 32075
rect 32733 32017 33453 32073
rect 33509 32017 33521 32073
rect 33441 32015 33521 32017
rect 33770 32073 33850 32075
rect 34037 32074 34107 32085
rect 34927 32074 35007 32076
rect 34037 32073 34939 32074
rect 33770 32017 33782 32073
rect 33838 32017 34039 32073
rect 34095 32018 34939 32073
rect 34995 32018 35007 32074
rect 34095 32017 34355 32018
rect 33770 32015 33850 32017
rect 34037 32007 34107 32017
rect 34927 32016 35007 32018
rect 35256 32074 35336 32076
rect 35699 32074 35769 32084
rect 35256 32018 35268 32074
rect 35324 32018 35701 32074
rect 35757 32018 35769 32074
rect 35256 32016 35336 32018
rect 35699 32006 35769 32018
rect 23113 31957 23183 31969
rect 24153 31957 24233 31959
rect 25639 31958 25719 31960
rect 23113 31901 23125 31957
rect 23181 31901 24165 31957
rect 24221 31901 24233 31957
rect 23113 31889 23183 31901
rect 19465 30850 19629 30862
rect 19945 30928 20109 30940
rect 19945 30872 19957 30928
rect 20013 30872 20109 30928
rect 19945 30860 20109 30872
rect 19465 30794 19477 30850
rect 19533 30794 19629 30850
rect 19465 30782 19629 30794
rect 19533 30732 19629 30782
rect 18430 30710 18476 30721
rect 17536 30410 17582 30550
rect 17751 30419 17847 30450
rect 17751 30373 17762 30419
rect 17836 30373 17847 30419
rect 18016 30410 18062 30550
rect 17582 30327 17720 30338
rect 17582 29753 17674 30327
rect 17878 30327 17924 30338
rect 17861 30043 17878 30053
rect 17924 30043 17941 30053
rect 17861 29803 17873 30043
rect 17929 29803 17941 30043
rect 17861 29793 17878 29803
rect 17582 29742 17720 29753
rect 17924 29793 17941 29803
rect 17878 29742 17924 29753
rect 17536 29659 17582 29670
rect 17751 29661 17762 29707
rect 17836 29661 17847 29707
rect 17751 29520 17847 29661
rect 18645 30719 18945 30732
rect 18645 30673 18656 30719
rect 18730 30686 18860 30719
rect 18730 30673 18741 30686
rect 18849 30673 18860 30686
rect 18934 30673 18945 30719
rect 19114 30710 19160 30721
rect 18476 30627 18614 30638
rect 18476 30453 18568 30627
rect 18772 30627 18818 30638
rect 18755 30568 18772 30578
rect 18976 30627 19114 30638
rect 18818 30568 18835 30578
rect 18755 30512 18767 30568
rect 18823 30512 18835 30568
rect 18755 30502 18772 30512
rect 18476 30442 18614 30453
rect 18818 30502 18835 30512
rect 18772 30442 18818 30453
rect 19022 30453 19114 30627
rect 18976 30442 19114 30453
rect 18430 30230 18476 30370
rect 18645 30361 18656 30407
rect 18730 30361 18741 30407
rect 18645 30330 18741 30361
rect 18849 30361 18860 30407
rect 18934 30361 18945 30407
rect 18849 30330 18945 30361
rect 19329 30719 19629 30732
rect 19329 30673 19340 30719
rect 19414 30686 19544 30719
rect 19414 30673 19425 30686
rect 19533 30673 19544 30686
rect 19618 30673 19629 30719
rect 19798 30710 19844 30721
rect 19252 30627 19298 30638
rect 19235 30568 19252 30578
rect 19456 30627 19502 30638
rect 19298 30568 19315 30578
rect 19235 30512 19247 30568
rect 19303 30512 19315 30568
rect 19235 30502 19252 30512
rect 19298 30502 19315 30512
rect 19439 30568 19456 30578
rect 19660 30627 19706 30638
rect 19502 30568 19519 30578
rect 19439 30512 19451 30568
rect 19507 30512 19519 30568
rect 19439 30502 19456 30512
rect 19252 30442 19298 30453
rect 19502 30502 19519 30512
rect 19643 30568 19660 30578
rect 19706 30568 19723 30578
rect 19643 30512 19655 30568
rect 19711 30512 19723 30568
rect 19643 30502 19660 30512
rect 19456 30442 19502 30453
rect 19706 30502 19723 30512
rect 19660 30442 19706 30453
rect 19114 30230 19160 30370
rect 19329 30361 19340 30407
rect 19414 30361 19425 30407
rect 19329 30330 19425 30361
rect 19533 30361 19544 30407
rect 19618 30361 19629 30407
rect 19533 30330 19629 30361
rect 20013 30719 20109 30860
rect 20621 30974 22589 31170
rect 23397 31170 23453 31901
rect 24153 31899 24233 31901
rect 24883 31902 25651 31958
rect 25707 31902 25719 31958
rect 23785 31807 23865 31821
rect 23572 31785 23618 31796
rect 23785 31751 23797 31807
rect 23853 31751 23865 31807
rect 23969 31807 24049 31821
rect 23969 31751 23981 31807
rect 24037 31751 24049 31807
rect 24153 31807 24233 31821
rect 24153 31751 24165 31807
rect 24221 31751 24233 31807
rect 24400 31785 24446 31796
rect 23787 31748 23798 31751
rect 23852 31748 23863 31751
rect 23971 31748 23982 31751
rect 24036 31748 24047 31751
rect 24155 31748 24166 31751
rect 24220 31748 24231 31751
rect 23710 31702 23756 31713
rect 23618 31528 23710 31702
rect 23710 31517 23756 31528
rect 23894 31702 23940 31713
rect 23894 31517 23940 31528
rect 24078 31702 24124 31713
rect 24262 31702 24308 31713
rect 24245 31675 24262 31677
rect 24308 31675 24325 31677
rect 24245 31555 24257 31675
rect 24313 31555 24325 31675
rect 24245 31553 24262 31555
rect 24078 31517 24124 31528
rect 24308 31553 24325 31555
rect 24262 31517 24308 31528
rect 23572 31300 23618 31445
rect 23787 31436 23798 31482
rect 23852 31436 23863 31482
rect 23787 31403 23863 31436
rect 23971 31436 23982 31482
rect 24036 31436 24047 31482
rect 23971 31403 24047 31436
rect 24155 31436 24166 31482
rect 24220 31436 24231 31482
rect 24155 31403 24231 31436
rect 24400 31300 24446 31445
rect 23560 31288 23640 31300
rect 23560 31232 23572 31288
rect 23628 31232 23640 31288
rect 23560 31220 23640 31232
rect 24378 31288 24456 31300
rect 24378 31232 24390 31288
rect 24446 31232 24456 31288
rect 24378 31220 24456 31232
rect 24731 31170 24811 31180
rect 23397 31114 24743 31170
rect 24799 31114 24811 31170
rect 24731 31112 24811 31114
rect 24565 31061 24635 31063
rect 20621 30834 20721 30974
rect 22489 30834 22589 30974
rect 20621 30794 22589 30834
rect 23397 31060 24635 31061
rect 23397 31006 24567 31060
rect 24623 31006 24635 31060
rect 23397 31005 24635 31006
rect 20013 30673 20024 30719
rect 20098 30673 20109 30719
rect 20278 30710 20324 30721
rect 19844 30627 19982 30638
rect 19844 30453 19936 30627
rect 20140 30627 20186 30638
rect 20123 30568 20140 30578
rect 20186 30568 20203 30578
rect 20123 30512 20135 30568
rect 20191 30512 20203 30568
rect 20123 30502 20140 30512
rect 19844 30442 19982 30453
rect 20186 30502 20203 30512
rect 20140 30442 20186 30453
rect 19798 30230 19844 30370
rect 20013 30361 20024 30407
rect 20098 30361 20109 30407
rect 20013 30330 20109 30361
rect 20278 30230 20324 30370
rect 20658 30654 20704 30794
rect 18393 30200 20361 30230
rect 18393 30060 19661 30200
rect 20261 30060 20361 30200
rect 18393 30030 20361 30060
rect 20873 30663 20969 30694
rect 20873 30617 20884 30663
rect 20958 30617 20969 30663
rect 21077 30663 21173 30694
rect 21077 30617 21088 30663
rect 21162 30617 21173 30663
rect 21342 30654 21388 30794
rect 20704 30571 20842 30582
rect 21000 30571 21046 30582
rect 21204 30571 21342 30582
rect 20704 29997 20796 30571
rect 20983 30331 20995 30571
rect 21051 30331 21063 30571
rect 20704 29986 20842 29997
rect 21000 29986 21046 29997
rect 21250 29997 21342 30571
rect 21204 29986 21342 29997
rect 20658 29903 20704 29914
rect 20873 29905 20884 29951
rect 20958 29931 20969 29951
rect 21077 29931 21088 29951
rect 20958 29905 21088 29931
rect 21162 29905 21173 29951
rect 20873 29878 21173 29905
rect 21557 30663 21653 30694
rect 21557 30617 21568 30663
rect 21642 30617 21653 30663
rect 21761 30663 21857 30694
rect 21761 30617 21772 30663
rect 21846 30617 21857 30663
rect 22026 30654 22072 30794
rect 21480 30571 21526 30582
rect 21684 30571 21730 30582
rect 21888 30571 21934 30582
rect 21667 30331 21679 30571
rect 21735 30331 21747 30571
rect 21463 29997 21475 30237
rect 21531 29997 21543 30237
rect 21871 29997 21883 30237
rect 21939 29997 21951 30237
rect 21480 29986 21526 29997
rect 21684 29986 21730 29997
rect 21888 29986 21934 29997
rect 21342 29903 21388 29914
rect 21557 29905 21568 29951
rect 21642 29931 21653 29951
rect 21761 29931 21772 29951
rect 21642 29905 21772 29931
rect 21846 29905 21857 29951
rect 21557 29878 21857 29905
rect 22241 30663 22337 30694
rect 22241 30617 22252 30663
rect 22326 30617 22337 30663
rect 22506 30654 22552 30794
rect 22072 30571 22210 30582
rect 22072 29997 22164 30571
rect 22368 30571 22414 30582
rect 22351 30287 22368 30297
rect 22414 30287 22431 30297
rect 22351 30047 22363 30287
rect 22419 30047 22431 30287
rect 22351 30037 22368 30047
rect 22072 29986 22210 29997
rect 22414 30037 22431 30047
rect 22368 29986 22414 29997
rect 22026 29903 22072 29914
rect 22241 29905 22252 29951
rect 22326 29905 22337 29951
rect 20873 29830 20969 29878
rect 18016 29659 18062 29670
rect 18393 29800 20361 29830
rect 18393 29660 19661 29800
rect 20261 29660 20361 29800
rect 18393 29630 20361 29660
rect 20873 29774 20893 29830
rect 20949 29774 20969 29830
rect 17683 29508 17847 29520
rect 17683 29452 17695 29508
rect 17751 29452 17847 29508
rect 17683 29440 17847 29452
rect 13322 28909 13334 28965
rect 13390 28909 13517 28965
rect 13573 28909 15467 28965
rect 17536 29290 17582 29301
rect 17751 29299 17847 29440
rect 18430 29490 18476 29501
rect 17751 29253 17762 29299
rect 17836 29253 17847 29299
rect 18016 29290 18062 29301
rect 17582 29207 17720 29218
rect 17582 29033 17674 29207
rect 17878 29207 17924 29218
rect 17861 29148 17878 29158
rect 17924 29148 17941 29158
rect 17861 29092 17873 29148
rect 17929 29092 17941 29148
rect 17861 29082 17878 29092
rect 17582 29022 17720 29033
rect 17924 29082 17941 29092
rect 17878 29022 17924 29033
rect 13322 28897 13408 28909
rect 13515 28897 13575 28909
rect 9993 28510 10157 28522
rect 10473 28588 10637 28600
rect 10473 28532 10485 28588
rect 10541 28532 10637 28588
rect 10473 28520 10637 28532
rect 9993 28454 10005 28510
rect 10061 28454 10157 28510
rect 9993 28442 10157 28454
rect 10061 28392 10157 28442
rect 3445 27890 8627 28089
rect 8958 28370 9004 28381
rect 9173 28379 9473 28392
rect 9173 28333 9184 28379
rect 9258 28346 9388 28379
rect 9258 28333 9269 28346
rect 9377 28333 9388 28346
rect 9462 28333 9473 28379
rect 9642 28370 9688 28381
rect 9004 28287 9142 28298
rect 9004 28113 9096 28287
rect 9300 28287 9346 28298
rect 9283 28228 9300 28238
rect 9504 28287 9642 28298
rect 9346 28228 9363 28238
rect 9283 28172 9295 28228
rect 9351 28172 9363 28228
rect 9283 28162 9300 28172
rect 9004 28102 9142 28113
rect 9346 28162 9363 28172
rect 9300 28102 9346 28113
rect 9550 28113 9642 28287
rect 9504 28102 9642 28113
rect 8958 27890 9004 28030
rect 9173 28021 9184 28067
rect 9258 28021 9269 28067
rect 9173 27990 9269 28021
rect 9377 28021 9388 28067
rect 9462 28021 9473 28067
rect 9377 27990 9473 28021
rect 9857 28379 10157 28392
rect 9857 28333 9868 28379
rect 9942 28346 10072 28379
rect 9942 28333 9953 28346
rect 10061 28333 10072 28346
rect 10146 28333 10157 28379
rect 10326 28370 10372 28381
rect 9780 28287 9826 28298
rect 9763 28228 9780 28238
rect 9984 28287 10030 28298
rect 9826 28228 9843 28238
rect 9763 28172 9775 28228
rect 9831 28172 9843 28228
rect 9763 28162 9780 28172
rect 9826 28162 9843 28172
rect 9967 28228 9984 28238
rect 10188 28287 10234 28298
rect 10030 28228 10047 28238
rect 9967 28172 9979 28228
rect 10035 28172 10047 28228
rect 9967 28162 9984 28172
rect 9780 28102 9826 28113
rect 10030 28162 10047 28172
rect 10171 28228 10188 28238
rect 10234 28228 10251 28238
rect 10171 28172 10183 28228
rect 10239 28172 10251 28228
rect 10171 28162 10188 28172
rect 9984 28102 10030 28113
rect 10234 28162 10251 28172
rect 10188 28102 10234 28113
rect 9642 27890 9688 28030
rect 9857 28021 9868 28067
rect 9942 28021 9953 28067
rect 9857 27990 9953 28021
rect 10061 28021 10072 28067
rect 10146 28021 10157 28067
rect 10061 27990 10157 28021
rect 10541 28379 10637 28520
rect 11149 28690 13117 28874
rect 17536 28810 17582 28950
rect 17751 28941 17762 28987
rect 17836 28941 17847 28987
rect 17751 28910 17847 28941
rect 18016 28810 18062 28950
rect 10541 28333 10552 28379
rect 10626 28333 10637 28379
rect 10806 28370 10852 28381
rect 10372 28287 10510 28298
rect 10372 28113 10464 28287
rect 10668 28287 10714 28298
rect 10651 28228 10668 28238
rect 10714 28228 10731 28238
rect 10651 28172 10663 28228
rect 10719 28172 10731 28228
rect 10651 28162 10668 28172
rect 10372 28102 10510 28113
rect 10714 28162 10731 28172
rect 10668 28102 10714 28113
rect 10326 27890 10372 28030
rect 10541 28021 10552 28067
rect 10626 28021 10637 28067
rect 10541 27990 10637 28021
rect 10806 27890 10852 28030
rect 11149 27890 12617 28690
rect 12917 28090 13117 28690
rect 17499 28090 18099 28810
rect 18645 29499 18741 29530
rect 18645 29453 18656 29499
rect 18730 29453 18741 29499
rect 18910 29490 19364 29630
rect 18568 29407 18614 29418
rect 18551 29123 18568 29133
rect 18772 29407 18910 29418
rect 18614 29123 18631 29133
rect 18551 28883 18563 29123
rect 18619 28883 18631 29123
rect 18551 28873 18568 28883
rect 18614 28873 18631 28883
rect 18568 28822 18614 28833
rect 18818 28833 18910 29407
rect 18772 28822 18910 28833
rect 18430 28739 18476 28750
rect 18645 28741 18656 28787
rect 18730 28741 18741 28787
rect 18645 28666 18741 28741
rect 18956 28822 19318 29490
rect 18910 28739 18956 28750
rect 19533 29499 19629 29530
rect 19533 29453 19544 29499
rect 19618 29453 19629 29499
rect 19798 29490 19844 29630
rect 19364 29407 19502 29418
rect 19364 28833 19456 29407
rect 19660 29407 19706 29418
rect 19643 29123 19660 29133
rect 19706 29123 19723 29133
rect 19643 28883 19655 29123
rect 19711 28883 19723 29123
rect 19643 28873 19660 28883
rect 19364 28822 19502 28833
rect 19706 28873 19723 28883
rect 19660 28822 19706 28833
rect 19318 28739 19364 28750
rect 19533 28741 19544 28787
rect 19618 28741 19629 28787
rect 18645 28610 18665 28666
rect 18721 28610 18741 28666
rect 18645 28392 18741 28610
rect 19533 28522 19629 28741
rect 20013 29499 20109 29530
rect 20013 29453 20024 29499
rect 20098 29453 20109 29499
rect 20278 29490 20324 29630
rect 19844 29407 19982 29418
rect 19844 28833 19936 29407
rect 20140 29407 20186 29418
rect 20123 29123 20140 29133
rect 20186 29123 20203 29133
rect 20123 28883 20135 29123
rect 20191 28883 20203 29123
rect 20123 28873 20140 28883
rect 19844 28822 19982 28833
rect 20186 28873 20203 28883
rect 20140 28822 20186 28833
rect 19798 28739 19844 28750
rect 20013 28741 20024 28787
rect 20098 28741 20109 28787
rect 20013 28600 20109 28741
rect 20658 29534 20704 29545
rect 20873 29543 20969 29774
rect 21557 29674 21653 29878
rect 22241 29764 22337 29905
rect 23397 29984 23453 31005
rect 24565 30997 24635 31005
rect 24061 30953 24147 30957
rect 24061 30897 24073 30953
rect 24129 30897 24147 30953
rect 24061 30885 24147 30897
rect 23572 30740 23618 30751
rect 23787 30749 23863 30782
rect 23787 30703 23798 30749
rect 23852 30703 23863 30749
rect 23971 30749 24047 30782
rect 23971 30703 23982 30749
rect 24036 30703 24047 30749
rect 24155 30749 24231 30782
rect 24155 30703 24166 30749
rect 24220 30703 24231 30749
rect 24400 30740 24446 30751
rect 23710 30657 23756 30668
rect 23693 30630 23710 30632
rect 23894 30657 23940 30668
rect 23756 30630 23773 30632
rect 23618 30510 23705 30630
rect 23761 30510 23773 30630
rect 23693 30508 23710 30510
rect 23618 30210 23710 30330
rect 23756 30508 23773 30510
rect 23877 30330 23894 30332
rect 24078 30657 24124 30668
rect 24061 30630 24078 30632
rect 24262 30657 24308 30668
rect 24124 30630 24141 30632
rect 24061 30510 24073 30630
rect 24129 30510 24141 30630
rect 24061 30508 24078 30510
rect 23940 30330 23957 30332
rect 23877 30210 23889 30330
rect 23945 30210 23957 30330
rect 23877 30208 23894 30210
rect 23710 30172 23756 30183
rect 23940 30208 23957 30210
rect 23894 30172 23940 30183
rect 24124 30508 24141 30510
rect 24245 30330 24262 30332
rect 24383 30630 24400 30632
rect 24446 30630 24463 30632
rect 24383 30509 24395 30630
rect 24451 30509 24463 30630
rect 24383 30507 24400 30509
rect 24308 30330 24325 30332
rect 24245 30210 24257 30330
rect 24313 30210 24325 30330
rect 24245 30208 24262 30210
rect 24078 30172 24124 30183
rect 24308 30208 24325 30210
rect 24262 30172 24308 30183
rect 23787 30134 23798 30137
rect 23852 30134 23863 30137
rect 23971 30134 23982 30137
rect 24036 30134 24047 30137
rect 24155 30134 24166 30137
rect 24220 30134 24231 30137
rect 23572 30089 23618 30100
rect 23785 30078 23797 30134
rect 23853 30078 23865 30134
rect 23785 30064 23865 30078
rect 23969 30078 23981 30134
rect 24037 30078 24049 30134
rect 23969 30064 24049 30078
rect 24153 30078 24165 30134
rect 24221 30078 24233 30134
rect 24446 30507 24463 30509
rect 24400 30089 24446 30100
rect 24153 30064 24233 30078
rect 23785 29984 23865 29986
rect 23397 29928 23797 29984
rect 23853 29928 23865 29984
rect 23785 29926 23865 29928
rect 22506 29903 22552 29914
rect 22977 29868 23047 29882
rect 23969 29868 24049 29870
rect 22977 29812 22989 29868
rect 23045 29812 23981 29868
rect 24037 29812 24049 29868
rect 22977 29800 23047 29812
rect 23969 29810 24049 29812
rect 24298 29868 24378 29870
rect 24741 29868 24801 29880
rect 24298 29812 24310 29868
rect 24366 29812 24743 29868
rect 24799 29812 24801 29868
rect 24298 29810 24378 29812
rect 24741 29800 24801 29812
rect 22173 29752 22337 29764
rect 22173 29696 22185 29752
rect 22241 29696 22337 29752
rect 22173 29684 22337 29696
rect 22743 29752 22821 29763
rect 24153 29752 24233 29754
rect 22743 29751 24165 29752
rect 22743 29697 22755 29751
rect 22809 29697 24165 29751
rect 22743 29696 24165 29697
rect 24221 29696 24233 29752
rect 22743 29685 22821 29696
rect 24153 29694 24233 29696
rect 21557 29618 21577 29674
rect 21633 29618 21653 29674
rect 20873 29497 20884 29543
rect 20958 29497 20969 29543
rect 21138 29534 21388 29545
rect 20796 29451 20842 29462
rect 20779 29392 20796 29402
rect 21000 29451 21138 29462
rect 20842 29392 20859 29402
rect 20779 29336 20791 29392
rect 20847 29336 20859 29392
rect 20779 29326 20796 29336
rect 20842 29326 20859 29336
rect 20796 29266 20842 29277
rect 21046 29277 21138 29451
rect 21000 29266 21138 29277
rect 20658 29054 20704 29194
rect 20873 29185 20884 29231
rect 20958 29185 20969 29231
rect 20873 29154 20969 29185
rect 21184 29194 21342 29534
rect 21557 29543 21653 29618
rect 21557 29497 21568 29543
rect 21642 29497 21653 29543
rect 21822 29534 21868 29545
rect 21388 29451 21526 29462
rect 21388 29277 21480 29451
rect 21684 29451 21730 29462
rect 21667 29392 21684 29402
rect 21730 29392 21747 29402
rect 21667 29336 21679 29392
rect 21735 29336 21747 29392
rect 21667 29326 21684 29336
rect 21388 29266 21526 29277
rect 21730 29326 21747 29336
rect 21684 29266 21730 29277
rect 21138 29183 21388 29194
rect 21557 29185 21568 29231
rect 21642 29185 21653 29231
rect 21184 29054 21342 29183
rect 21557 29154 21653 29185
rect 21822 29054 21868 29194
rect 22026 29534 22072 29545
rect 22241 29543 22337 29684
rect 23785 29602 23865 29616
rect 23572 29580 23618 29591
rect 22241 29497 22252 29543
rect 22326 29497 22337 29543
rect 22506 29534 22552 29545
rect 22072 29451 22210 29462
rect 22072 29277 22164 29451
rect 22368 29451 22414 29462
rect 22351 29392 22368 29402
rect 22414 29392 22431 29402
rect 22351 29336 22363 29392
rect 22419 29336 22431 29392
rect 22351 29326 22368 29336
rect 22072 29266 22210 29277
rect 22414 29326 22431 29336
rect 22368 29266 22414 29277
rect 22026 29054 22072 29194
rect 22241 29185 22252 29231
rect 22326 29185 22337 29231
rect 22241 29154 22337 29185
rect 22506 29054 22552 29194
rect 23785 29546 23797 29602
rect 23853 29546 23865 29602
rect 23969 29602 24049 29616
rect 23969 29546 23981 29602
rect 24037 29546 24049 29602
rect 24153 29602 24233 29616
rect 24153 29546 24165 29602
rect 24221 29546 24233 29602
rect 24400 29580 24446 29591
rect 23787 29543 23798 29546
rect 23852 29543 23863 29546
rect 23971 29543 23982 29546
rect 24036 29543 24047 29546
rect 24155 29543 24166 29546
rect 24220 29543 24231 29546
rect 23710 29497 23756 29508
rect 23618 29323 23710 29497
rect 23710 29312 23756 29323
rect 23894 29497 23940 29508
rect 23894 29312 23940 29323
rect 24078 29497 24124 29508
rect 24262 29497 24308 29508
rect 24245 29470 24262 29472
rect 24308 29470 24325 29472
rect 24245 29350 24257 29470
rect 24313 29350 24325 29470
rect 24245 29348 24262 29350
rect 24078 29312 24124 29323
rect 24308 29348 24325 29350
rect 24262 29312 24308 29323
rect 23572 29095 23618 29240
rect 23787 29231 23798 29277
rect 23852 29231 23863 29277
rect 23787 29198 23863 29231
rect 23971 29231 23982 29277
rect 24036 29231 24047 29277
rect 23971 29198 24047 29231
rect 24155 29231 24166 29277
rect 24220 29231 24231 29277
rect 24155 29198 24231 29231
rect 24400 29095 24446 29240
rect 23560 29083 23640 29095
rect 20278 28739 20324 28750
rect 20621 29014 22589 29054
rect 23560 29027 23572 29083
rect 23628 29027 23640 29083
rect 23560 29015 23640 29027
rect 24378 29083 24458 29095
rect 24378 29027 24390 29083
rect 24446 29027 24458 29083
rect 24378 29015 24458 29027
rect 20621 28874 20721 29014
rect 22489 28874 22589 29014
rect 22794 28965 22880 28977
rect 22987 28965 23047 28969
rect 24883 28965 24939 31902
rect 25639 31900 25719 31902
rect 25271 31808 25351 31822
rect 25058 31786 25104 31797
rect 25271 31752 25283 31808
rect 25339 31752 25351 31808
rect 25455 31808 25535 31822
rect 25455 31752 25467 31808
rect 25523 31752 25535 31808
rect 25639 31808 25719 31822
rect 25639 31752 25651 31808
rect 25707 31752 25719 31808
rect 25886 31786 25932 31797
rect 25273 31749 25284 31752
rect 25338 31749 25349 31752
rect 25457 31749 25468 31752
rect 25522 31749 25533 31752
rect 25641 31749 25652 31752
rect 25706 31749 25717 31752
rect 25196 31703 25242 31714
rect 25104 31529 25196 31703
rect 25196 31518 25242 31529
rect 25380 31703 25426 31714
rect 25380 31518 25426 31529
rect 25564 31703 25610 31714
rect 25748 31703 25794 31714
rect 25731 31676 25748 31678
rect 25794 31676 25811 31678
rect 25731 31556 25743 31676
rect 25799 31556 25811 31676
rect 25731 31554 25748 31556
rect 25564 31518 25610 31529
rect 25794 31554 25811 31556
rect 25748 31518 25794 31529
rect 25058 31301 25104 31446
rect 25273 31437 25284 31483
rect 25338 31437 25349 31483
rect 25273 31404 25349 31437
rect 25457 31437 25468 31483
rect 25522 31437 25533 31483
rect 25457 31404 25533 31437
rect 25641 31437 25652 31483
rect 25706 31437 25717 31483
rect 25641 31404 25717 31437
rect 25886 31301 25932 31446
rect 25046 31289 25126 31301
rect 25046 31233 25058 31289
rect 25114 31233 25126 31289
rect 25046 31221 25126 31233
rect 25864 31289 25942 31301
rect 25864 31233 25876 31289
rect 25932 31233 25942 31289
rect 25864 31221 25942 31233
rect 26971 31170 27171 31970
rect 27371 31170 27571 31970
rect 26971 30550 27571 31170
rect 27902 31830 27948 31841
rect 28117 31839 28213 31870
rect 28117 31793 28128 31839
rect 28202 31793 28213 31839
rect 28382 31830 28836 31970
rect 28040 31747 28086 31758
rect 28023 31463 28040 31473
rect 28244 31747 28382 31758
rect 28086 31463 28103 31473
rect 28023 31223 28035 31463
rect 28091 31223 28103 31463
rect 28023 31213 28040 31223
rect 28086 31213 28103 31223
rect 28040 31162 28086 31173
rect 28290 31173 28382 31747
rect 28244 31162 28382 31173
rect 27902 31079 27948 31090
rect 28117 31081 28128 31127
rect 28202 31081 28213 31127
rect 28117 31006 28213 31081
rect 28428 31162 28790 31830
rect 28382 31079 28428 31090
rect 29005 31839 29101 31870
rect 29005 31793 29016 31839
rect 29090 31793 29101 31839
rect 29270 31830 29316 31970
rect 28836 31747 28974 31758
rect 28836 31173 28928 31747
rect 29132 31747 29178 31758
rect 29115 31463 29132 31473
rect 29178 31463 29195 31473
rect 29115 31223 29127 31463
rect 29183 31223 29195 31463
rect 29115 31213 29132 31223
rect 28836 31162 28974 31173
rect 29178 31213 29195 31223
rect 29132 31162 29178 31173
rect 28790 31079 28836 31090
rect 29005 31081 29016 31127
rect 29090 31081 29101 31127
rect 28117 30950 28137 31006
rect 28193 30950 28213 31006
rect 28117 30732 28213 30950
rect 29005 30862 29101 31081
rect 29485 31839 29581 31870
rect 29485 31793 29496 31839
rect 29570 31793 29581 31839
rect 29750 31830 29796 31970
rect 29316 31747 29454 31758
rect 29316 31173 29408 31747
rect 29612 31747 29658 31758
rect 29595 31463 29612 31473
rect 29658 31463 29675 31473
rect 29595 31223 29607 31463
rect 29663 31223 29675 31463
rect 29595 31213 29612 31223
rect 29316 31162 29454 31173
rect 29658 31213 29675 31223
rect 29612 31162 29658 31173
rect 29270 31079 29316 31090
rect 29485 31081 29496 31127
rect 29570 31081 29581 31127
rect 29485 30940 29581 31081
rect 29750 31079 29796 31090
rect 30093 31170 31561 31970
rect 31861 31170 32061 31970
rect 36443 31970 41533 32170
rect 42205 32073 42261 33320
rect 45161 33318 45241 33320
rect 43685 33265 43755 33267
rect 44985 33266 45065 33268
rect 42341 33209 43687 33265
rect 43743 33209 43755 33265
rect 42341 32189 42397 33209
rect 43685 33197 43755 33209
rect 43827 33210 44997 33266
rect 45053 33210 45065 33266
rect 43005 33158 43091 33162
rect 43005 33102 43017 33158
rect 43073 33102 43091 33158
rect 43005 33090 43091 33102
rect 42516 32945 42562 32956
rect 42731 32954 42807 32987
rect 42731 32908 42742 32954
rect 42796 32908 42807 32954
rect 42915 32954 42991 32987
rect 42915 32908 42926 32954
rect 42980 32908 42991 32954
rect 43099 32954 43175 32987
rect 43099 32908 43110 32954
rect 43164 32908 43175 32954
rect 43344 32945 43390 32956
rect 42654 32862 42700 32873
rect 42637 32835 42654 32837
rect 42838 32862 42884 32873
rect 42700 32835 42717 32837
rect 42562 32715 42649 32835
rect 42705 32715 42717 32835
rect 42637 32713 42654 32715
rect 42562 32415 42654 32535
rect 42700 32713 42717 32715
rect 42821 32535 42838 32537
rect 43022 32862 43068 32873
rect 43005 32835 43022 32837
rect 43206 32862 43252 32873
rect 43068 32835 43085 32837
rect 43005 32715 43017 32835
rect 43073 32715 43085 32835
rect 43005 32713 43022 32715
rect 42884 32535 42901 32537
rect 42821 32415 42833 32535
rect 42889 32415 42901 32535
rect 42821 32413 42838 32415
rect 42654 32377 42700 32388
rect 42884 32413 42901 32415
rect 42838 32377 42884 32388
rect 43068 32713 43085 32715
rect 43189 32535 43206 32537
rect 43327 32835 43344 32837
rect 43390 32835 43407 32837
rect 43327 32714 43339 32835
rect 43395 32714 43407 32835
rect 43327 32712 43344 32714
rect 43252 32535 43269 32537
rect 43189 32415 43201 32535
rect 43257 32415 43269 32535
rect 43189 32413 43206 32415
rect 43022 32377 43068 32388
rect 43252 32413 43269 32415
rect 43206 32377 43252 32388
rect 42731 32339 42742 32342
rect 42796 32339 42807 32342
rect 42915 32339 42926 32342
rect 42980 32339 42991 32342
rect 43099 32339 43110 32342
rect 43164 32339 43175 32342
rect 42516 32294 42562 32305
rect 42729 32283 42741 32339
rect 42797 32283 42809 32339
rect 42729 32269 42809 32283
rect 42913 32283 42925 32339
rect 42981 32283 42993 32339
rect 42913 32269 42993 32283
rect 43097 32283 43109 32339
rect 43165 32283 43177 32339
rect 43390 32712 43407 32714
rect 43344 32294 43390 32305
rect 43097 32269 43177 32283
rect 42729 32189 42809 32191
rect 42341 32133 42741 32189
rect 42797 32133 42809 32189
rect 43827 32190 43883 33210
rect 44985 33198 45065 33210
rect 44491 33159 44577 33163
rect 44491 33103 44503 33159
rect 44559 33103 44577 33159
rect 44491 33091 44577 33103
rect 44002 32946 44048 32957
rect 44217 32955 44293 32988
rect 44217 32909 44228 32955
rect 44282 32909 44293 32955
rect 44401 32955 44477 32988
rect 44401 32909 44412 32955
rect 44466 32909 44477 32955
rect 44585 32955 44661 32988
rect 44585 32909 44596 32955
rect 44650 32909 44661 32955
rect 44830 32946 44876 32957
rect 44140 32863 44186 32874
rect 44123 32836 44140 32838
rect 44324 32863 44370 32874
rect 44186 32836 44203 32838
rect 44048 32716 44135 32836
rect 44191 32716 44203 32836
rect 44123 32714 44140 32716
rect 44048 32416 44140 32536
rect 44186 32714 44203 32716
rect 44307 32536 44324 32538
rect 44508 32863 44554 32874
rect 44491 32836 44508 32838
rect 44692 32863 44738 32874
rect 44554 32836 44571 32838
rect 44491 32716 44503 32836
rect 44559 32716 44571 32836
rect 44491 32714 44508 32716
rect 44370 32536 44387 32538
rect 44307 32416 44319 32536
rect 44375 32416 44387 32536
rect 44307 32414 44324 32416
rect 44140 32378 44186 32389
rect 44370 32414 44387 32416
rect 44324 32378 44370 32389
rect 44554 32714 44571 32716
rect 44675 32536 44692 32538
rect 44813 32836 44830 32838
rect 44876 32836 44893 32838
rect 44813 32715 44825 32836
rect 44881 32715 44893 32836
rect 44813 32713 44830 32715
rect 44738 32536 44755 32538
rect 44675 32416 44687 32536
rect 44743 32416 44755 32536
rect 44675 32414 44692 32416
rect 44508 32378 44554 32389
rect 44738 32414 44755 32416
rect 44692 32378 44738 32389
rect 44217 32340 44228 32343
rect 44282 32340 44293 32343
rect 44401 32340 44412 32343
rect 44466 32340 44477 32343
rect 44585 32340 44596 32343
rect 44650 32340 44661 32343
rect 44002 32295 44048 32306
rect 44215 32284 44227 32340
rect 44283 32284 44295 32340
rect 44215 32270 44295 32284
rect 44399 32284 44411 32340
rect 44467 32284 44479 32340
rect 44399 32270 44479 32284
rect 44583 32284 44595 32340
rect 44651 32284 44663 32340
rect 44876 32713 44893 32715
rect 44830 32295 44876 32306
rect 44583 32270 44663 32284
rect 44215 32190 44295 32192
rect 43827 32134 44227 32190
rect 44283 32134 44295 32190
rect 42729 32131 42809 32133
rect 44215 32132 44295 32134
rect 42913 32073 42993 32075
rect 42205 32017 42925 32073
rect 42981 32017 42993 32073
rect 42913 32015 42993 32017
rect 43242 32073 43322 32075
rect 43509 32074 43579 32085
rect 44399 32074 44479 32076
rect 43509 32073 44411 32074
rect 43242 32017 43254 32073
rect 43310 32017 43511 32073
rect 43567 32018 44411 32073
rect 44467 32018 44479 32074
rect 43567 32017 43827 32018
rect 43242 32015 43322 32017
rect 43509 32007 43579 32017
rect 44399 32016 44479 32018
rect 44728 32074 44808 32076
rect 45171 32074 45241 32084
rect 44728 32018 44740 32074
rect 44796 32018 45173 32074
rect 45229 32018 45241 32074
rect 44728 32016 44808 32018
rect 45171 32006 45241 32018
rect 32585 31957 32655 31969
rect 33625 31957 33705 31959
rect 35111 31958 35191 31960
rect 32585 31901 32597 31957
rect 32653 31901 33637 31957
rect 33693 31901 33705 31957
rect 32585 31889 32655 31901
rect 28937 30850 29101 30862
rect 29417 30928 29581 30940
rect 29417 30872 29429 30928
rect 29485 30872 29581 30928
rect 29417 30860 29581 30872
rect 28937 30794 28949 30850
rect 29005 30794 29101 30850
rect 28937 30782 29101 30794
rect 29005 30732 29101 30782
rect 27902 30710 27948 30721
rect 27008 30410 27054 30550
rect 27223 30419 27319 30450
rect 27223 30373 27234 30419
rect 27308 30373 27319 30419
rect 27488 30410 27534 30550
rect 27054 30327 27192 30338
rect 27054 29753 27146 30327
rect 27350 30327 27396 30338
rect 27333 30043 27350 30053
rect 27396 30043 27413 30053
rect 27333 29803 27345 30043
rect 27401 29803 27413 30043
rect 27333 29793 27350 29803
rect 27054 29742 27192 29753
rect 27396 29793 27413 29803
rect 27350 29742 27396 29753
rect 27008 29659 27054 29670
rect 27223 29661 27234 29707
rect 27308 29661 27319 29707
rect 27223 29520 27319 29661
rect 28117 30719 28417 30732
rect 28117 30673 28128 30719
rect 28202 30686 28332 30719
rect 28202 30673 28213 30686
rect 28321 30673 28332 30686
rect 28406 30673 28417 30719
rect 28586 30710 28632 30721
rect 27948 30627 28086 30638
rect 27948 30453 28040 30627
rect 28244 30627 28290 30638
rect 28227 30568 28244 30578
rect 28448 30627 28586 30638
rect 28290 30568 28307 30578
rect 28227 30512 28239 30568
rect 28295 30512 28307 30568
rect 28227 30502 28244 30512
rect 27948 30442 28086 30453
rect 28290 30502 28307 30512
rect 28244 30442 28290 30453
rect 28494 30453 28586 30627
rect 28448 30442 28586 30453
rect 27902 30230 27948 30370
rect 28117 30361 28128 30407
rect 28202 30361 28213 30407
rect 28117 30330 28213 30361
rect 28321 30361 28332 30407
rect 28406 30361 28417 30407
rect 28321 30330 28417 30361
rect 28801 30719 29101 30732
rect 28801 30673 28812 30719
rect 28886 30686 29016 30719
rect 28886 30673 28897 30686
rect 29005 30673 29016 30686
rect 29090 30673 29101 30719
rect 29270 30710 29316 30721
rect 28724 30627 28770 30638
rect 28707 30568 28724 30578
rect 28928 30627 28974 30638
rect 28770 30568 28787 30578
rect 28707 30512 28719 30568
rect 28775 30512 28787 30568
rect 28707 30502 28724 30512
rect 28770 30502 28787 30512
rect 28911 30568 28928 30578
rect 29132 30627 29178 30638
rect 28974 30568 28991 30578
rect 28911 30512 28923 30568
rect 28979 30512 28991 30568
rect 28911 30502 28928 30512
rect 28724 30442 28770 30453
rect 28974 30502 28991 30512
rect 29115 30568 29132 30578
rect 29178 30568 29195 30578
rect 29115 30512 29127 30568
rect 29183 30512 29195 30568
rect 29115 30502 29132 30512
rect 28928 30442 28974 30453
rect 29178 30502 29195 30512
rect 29132 30442 29178 30453
rect 28586 30230 28632 30370
rect 28801 30361 28812 30407
rect 28886 30361 28897 30407
rect 28801 30330 28897 30361
rect 29005 30361 29016 30407
rect 29090 30361 29101 30407
rect 29005 30330 29101 30361
rect 29485 30719 29581 30860
rect 30093 30974 32061 31170
rect 32869 31170 32925 31901
rect 33625 31899 33705 31901
rect 34355 31902 35123 31958
rect 35179 31902 35191 31958
rect 33257 31807 33337 31821
rect 33044 31785 33090 31796
rect 33257 31751 33269 31807
rect 33325 31751 33337 31807
rect 33441 31807 33521 31821
rect 33441 31751 33453 31807
rect 33509 31751 33521 31807
rect 33625 31807 33705 31821
rect 33625 31751 33637 31807
rect 33693 31751 33705 31807
rect 33872 31785 33918 31796
rect 33259 31748 33270 31751
rect 33324 31748 33335 31751
rect 33443 31748 33454 31751
rect 33508 31748 33519 31751
rect 33627 31748 33638 31751
rect 33692 31748 33703 31751
rect 33182 31702 33228 31713
rect 33090 31528 33182 31702
rect 33182 31517 33228 31528
rect 33366 31702 33412 31713
rect 33366 31517 33412 31528
rect 33550 31702 33596 31713
rect 33734 31702 33780 31713
rect 33717 31675 33734 31677
rect 33780 31675 33797 31677
rect 33717 31555 33729 31675
rect 33785 31555 33797 31675
rect 33717 31553 33734 31555
rect 33550 31517 33596 31528
rect 33780 31553 33797 31555
rect 33734 31517 33780 31528
rect 33044 31300 33090 31445
rect 33259 31436 33270 31482
rect 33324 31436 33335 31482
rect 33259 31403 33335 31436
rect 33443 31436 33454 31482
rect 33508 31436 33519 31482
rect 33443 31403 33519 31436
rect 33627 31436 33638 31482
rect 33692 31436 33703 31482
rect 33627 31403 33703 31436
rect 33872 31300 33918 31445
rect 33032 31288 33112 31300
rect 33032 31232 33044 31288
rect 33100 31232 33112 31288
rect 33032 31220 33112 31232
rect 33850 31288 33928 31300
rect 33850 31232 33862 31288
rect 33918 31232 33928 31288
rect 33850 31220 33928 31232
rect 34203 31170 34283 31180
rect 32869 31114 34215 31170
rect 34271 31114 34283 31170
rect 34203 31112 34283 31114
rect 34037 31061 34107 31063
rect 30093 30834 30193 30974
rect 31961 30834 32061 30974
rect 30093 30794 32061 30834
rect 32869 31060 34107 31061
rect 32869 31006 34039 31060
rect 34095 31006 34107 31060
rect 32869 31005 34107 31006
rect 29485 30673 29496 30719
rect 29570 30673 29581 30719
rect 29750 30710 29796 30721
rect 29316 30627 29454 30638
rect 29316 30453 29408 30627
rect 29612 30627 29658 30638
rect 29595 30568 29612 30578
rect 29658 30568 29675 30578
rect 29595 30512 29607 30568
rect 29663 30512 29675 30568
rect 29595 30502 29612 30512
rect 29316 30442 29454 30453
rect 29658 30502 29675 30512
rect 29612 30442 29658 30453
rect 29270 30230 29316 30370
rect 29485 30361 29496 30407
rect 29570 30361 29581 30407
rect 29485 30330 29581 30361
rect 29750 30230 29796 30370
rect 30130 30654 30176 30794
rect 27865 30200 29833 30230
rect 27865 30060 29133 30200
rect 29733 30060 29833 30200
rect 27865 30030 29833 30060
rect 30345 30663 30441 30694
rect 30345 30617 30356 30663
rect 30430 30617 30441 30663
rect 30549 30663 30645 30694
rect 30549 30617 30560 30663
rect 30634 30617 30645 30663
rect 30814 30654 30860 30794
rect 30176 30571 30314 30582
rect 30472 30571 30518 30582
rect 30676 30571 30814 30582
rect 30176 29997 30268 30571
rect 30455 30331 30467 30571
rect 30523 30331 30535 30571
rect 30176 29986 30314 29997
rect 30472 29986 30518 29997
rect 30722 29997 30814 30571
rect 30676 29986 30814 29997
rect 30130 29903 30176 29914
rect 30345 29905 30356 29951
rect 30430 29931 30441 29951
rect 30549 29931 30560 29951
rect 30430 29905 30560 29931
rect 30634 29905 30645 29951
rect 30345 29878 30645 29905
rect 31029 30663 31125 30694
rect 31029 30617 31040 30663
rect 31114 30617 31125 30663
rect 31233 30663 31329 30694
rect 31233 30617 31244 30663
rect 31318 30617 31329 30663
rect 31498 30654 31544 30794
rect 30952 30571 30998 30582
rect 31156 30571 31202 30582
rect 31360 30571 31406 30582
rect 31139 30331 31151 30571
rect 31207 30331 31219 30571
rect 30935 29997 30947 30237
rect 31003 29997 31015 30237
rect 31343 29997 31355 30237
rect 31411 29997 31423 30237
rect 30952 29986 30998 29997
rect 31156 29986 31202 29997
rect 31360 29986 31406 29997
rect 30814 29903 30860 29914
rect 31029 29905 31040 29951
rect 31114 29931 31125 29951
rect 31233 29931 31244 29951
rect 31114 29905 31244 29931
rect 31318 29905 31329 29951
rect 31029 29878 31329 29905
rect 31713 30663 31809 30694
rect 31713 30617 31724 30663
rect 31798 30617 31809 30663
rect 31978 30654 32024 30794
rect 31544 30571 31682 30582
rect 31544 29997 31636 30571
rect 31840 30571 31886 30582
rect 31823 30287 31840 30297
rect 31886 30287 31903 30297
rect 31823 30047 31835 30287
rect 31891 30047 31903 30287
rect 31823 30037 31840 30047
rect 31544 29986 31682 29997
rect 31886 30037 31903 30047
rect 31840 29986 31886 29997
rect 31498 29903 31544 29914
rect 31713 29905 31724 29951
rect 31798 29905 31809 29951
rect 30345 29830 30441 29878
rect 27488 29659 27534 29670
rect 27865 29800 29833 29830
rect 27865 29660 29133 29800
rect 29733 29660 29833 29800
rect 27865 29630 29833 29660
rect 30345 29774 30365 29830
rect 30421 29774 30441 29830
rect 27155 29508 27319 29520
rect 27155 29452 27167 29508
rect 27223 29452 27319 29508
rect 27155 29440 27319 29452
rect 22794 28909 22806 28965
rect 22862 28909 22989 28965
rect 23045 28909 24939 28965
rect 27008 29290 27054 29301
rect 27223 29299 27319 29440
rect 27902 29490 27948 29501
rect 27223 29253 27234 29299
rect 27308 29253 27319 29299
rect 27488 29290 27534 29301
rect 27054 29207 27192 29218
rect 27054 29033 27146 29207
rect 27350 29207 27396 29218
rect 27333 29148 27350 29158
rect 27396 29148 27413 29158
rect 27333 29092 27345 29148
rect 27401 29092 27413 29148
rect 27333 29082 27350 29092
rect 27054 29022 27192 29033
rect 27396 29082 27413 29092
rect 27350 29022 27396 29033
rect 22794 28897 22880 28909
rect 22987 28897 23047 28909
rect 19465 28510 19629 28522
rect 19945 28588 20109 28600
rect 19945 28532 19957 28588
rect 20013 28532 20109 28588
rect 19945 28520 20109 28532
rect 19465 28454 19477 28510
rect 19533 28454 19629 28510
rect 19465 28442 19629 28454
rect 19533 28392 19629 28442
rect 12917 27890 18099 28090
rect 18430 28370 18476 28381
rect 18645 28379 18945 28392
rect 18645 28333 18656 28379
rect 18730 28346 18860 28379
rect 18730 28333 18741 28346
rect 18849 28333 18860 28346
rect 18934 28333 18945 28379
rect 19114 28370 19160 28381
rect 18476 28287 18614 28298
rect 18476 28113 18568 28287
rect 18772 28287 18818 28298
rect 18755 28228 18772 28238
rect 18976 28287 19114 28298
rect 18818 28228 18835 28238
rect 18755 28172 18767 28228
rect 18823 28172 18835 28228
rect 18755 28162 18772 28172
rect 18476 28102 18614 28113
rect 18818 28162 18835 28172
rect 18772 28102 18818 28113
rect 19022 28113 19114 28287
rect 18976 28102 19114 28113
rect 18430 27890 18476 28030
rect 18645 28021 18656 28067
rect 18730 28021 18741 28067
rect 18645 27990 18741 28021
rect 18849 28021 18860 28067
rect 18934 28021 18945 28067
rect 18849 27990 18945 28021
rect 19329 28379 19629 28392
rect 19329 28333 19340 28379
rect 19414 28346 19544 28379
rect 19414 28333 19425 28346
rect 19533 28333 19544 28346
rect 19618 28333 19629 28379
rect 19798 28370 19844 28381
rect 19252 28287 19298 28298
rect 19235 28228 19252 28238
rect 19456 28287 19502 28298
rect 19298 28228 19315 28238
rect 19235 28172 19247 28228
rect 19303 28172 19315 28228
rect 19235 28162 19252 28172
rect 19298 28162 19315 28172
rect 19439 28228 19456 28238
rect 19660 28287 19706 28298
rect 19502 28228 19519 28238
rect 19439 28172 19451 28228
rect 19507 28172 19519 28228
rect 19439 28162 19456 28172
rect 19252 28102 19298 28113
rect 19502 28162 19519 28172
rect 19643 28228 19660 28238
rect 19706 28228 19723 28238
rect 19643 28172 19655 28228
rect 19711 28172 19723 28228
rect 19643 28162 19660 28172
rect 19456 28102 19502 28113
rect 19706 28162 19723 28172
rect 19660 28102 19706 28113
rect 19114 27890 19160 28030
rect 19329 28021 19340 28067
rect 19414 28021 19425 28067
rect 19329 27990 19425 28021
rect 19533 28021 19544 28067
rect 19618 28021 19629 28067
rect 19533 27990 19629 28021
rect 20013 28379 20109 28520
rect 20621 28690 22589 28874
rect 27008 28810 27054 28950
rect 27223 28941 27234 28987
rect 27308 28941 27319 28987
rect 27223 28910 27319 28941
rect 27488 28810 27534 28950
rect 20013 28333 20024 28379
rect 20098 28333 20109 28379
rect 20278 28370 20324 28381
rect 19844 28287 19982 28298
rect 19844 28113 19936 28287
rect 20140 28287 20186 28298
rect 20123 28228 20140 28238
rect 20186 28228 20203 28238
rect 20123 28172 20135 28228
rect 20191 28172 20203 28228
rect 20123 28162 20140 28172
rect 19844 28102 19982 28113
rect 20186 28162 20203 28172
rect 20140 28102 20186 28113
rect 19798 27890 19844 28030
rect 20013 28021 20024 28067
rect 20098 28021 20109 28067
rect 20013 27990 20109 28021
rect 20278 27890 20324 28030
rect 20621 27890 22089 28690
rect 22389 28090 22589 28690
rect 26971 28090 27571 28810
rect 28117 29499 28213 29530
rect 28117 29453 28128 29499
rect 28202 29453 28213 29499
rect 28382 29490 28836 29630
rect 28040 29407 28086 29418
rect 28023 29123 28040 29133
rect 28244 29407 28382 29418
rect 28086 29123 28103 29133
rect 28023 28883 28035 29123
rect 28091 28883 28103 29123
rect 28023 28873 28040 28883
rect 28086 28873 28103 28883
rect 28040 28822 28086 28833
rect 28290 28833 28382 29407
rect 28244 28822 28382 28833
rect 27902 28739 27948 28750
rect 28117 28741 28128 28787
rect 28202 28741 28213 28787
rect 28117 28666 28213 28741
rect 28428 28822 28790 29490
rect 28382 28739 28428 28750
rect 29005 29499 29101 29530
rect 29005 29453 29016 29499
rect 29090 29453 29101 29499
rect 29270 29490 29316 29630
rect 28836 29407 28974 29418
rect 28836 28833 28928 29407
rect 29132 29407 29178 29418
rect 29115 29123 29132 29133
rect 29178 29123 29195 29133
rect 29115 28883 29127 29123
rect 29183 28883 29195 29123
rect 29115 28873 29132 28883
rect 28836 28822 28974 28833
rect 29178 28873 29195 28883
rect 29132 28822 29178 28833
rect 28790 28739 28836 28750
rect 29005 28741 29016 28787
rect 29090 28741 29101 28787
rect 28117 28610 28137 28666
rect 28193 28610 28213 28666
rect 28117 28392 28213 28610
rect 29005 28522 29101 28741
rect 29485 29499 29581 29530
rect 29485 29453 29496 29499
rect 29570 29453 29581 29499
rect 29750 29490 29796 29630
rect 29316 29407 29454 29418
rect 29316 28833 29408 29407
rect 29612 29407 29658 29418
rect 29595 29123 29612 29133
rect 29658 29123 29675 29133
rect 29595 28883 29607 29123
rect 29663 28883 29675 29123
rect 29595 28873 29612 28883
rect 29316 28822 29454 28833
rect 29658 28873 29675 28883
rect 29612 28822 29658 28833
rect 29270 28739 29316 28750
rect 29485 28741 29496 28787
rect 29570 28741 29581 28787
rect 29485 28600 29581 28741
rect 30130 29534 30176 29545
rect 30345 29543 30441 29774
rect 31029 29674 31125 29878
rect 31713 29764 31809 29905
rect 32869 29984 32925 31005
rect 34037 30997 34107 31005
rect 33533 30953 33619 30957
rect 33533 30897 33545 30953
rect 33601 30897 33619 30953
rect 33533 30885 33619 30897
rect 33044 30740 33090 30751
rect 33259 30749 33335 30782
rect 33259 30703 33270 30749
rect 33324 30703 33335 30749
rect 33443 30749 33519 30782
rect 33443 30703 33454 30749
rect 33508 30703 33519 30749
rect 33627 30749 33703 30782
rect 33627 30703 33638 30749
rect 33692 30703 33703 30749
rect 33872 30740 33918 30751
rect 33182 30657 33228 30668
rect 33165 30630 33182 30632
rect 33366 30657 33412 30668
rect 33228 30630 33245 30632
rect 33090 30510 33177 30630
rect 33233 30510 33245 30630
rect 33165 30508 33182 30510
rect 33090 30210 33182 30330
rect 33228 30508 33245 30510
rect 33349 30330 33366 30332
rect 33550 30657 33596 30668
rect 33533 30630 33550 30632
rect 33734 30657 33780 30668
rect 33596 30630 33613 30632
rect 33533 30510 33545 30630
rect 33601 30510 33613 30630
rect 33533 30508 33550 30510
rect 33412 30330 33429 30332
rect 33349 30210 33361 30330
rect 33417 30210 33429 30330
rect 33349 30208 33366 30210
rect 33182 30172 33228 30183
rect 33412 30208 33429 30210
rect 33366 30172 33412 30183
rect 33596 30508 33613 30510
rect 33717 30330 33734 30332
rect 33855 30630 33872 30632
rect 33918 30630 33935 30632
rect 33855 30509 33867 30630
rect 33923 30509 33935 30630
rect 33855 30507 33872 30509
rect 33780 30330 33797 30332
rect 33717 30210 33729 30330
rect 33785 30210 33797 30330
rect 33717 30208 33734 30210
rect 33550 30172 33596 30183
rect 33780 30208 33797 30210
rect 33734 30172 33780 30183
rect 33259 30134 33270 30137
rect 33324 30134 33335 30137
rect 33443 30134 33454 30137
rect 33508 30134 33519 30137
rect 33627 30134 33638 30137
rect 33692 30134 33703 30137
rect 33044 30089 33090 30100
rect 33257 30078 33269 30134
rect 33325 30078 33337 30134
rect 33257 30064 33337 30078
rect 33441 30078 33453 30134
rect 33509 30078 33521 30134
rect 33441 30064 33521 30078
rect 33625 30078 33637 30134
rect 33693 30078 33705 30134
rect 33918 30507 33935 30509
rect 33872 30089 33918 30100
rect 33625 30064 33705 30078
rect 33257 29984 33337 29986
rect 32869 29928 33269 29984
rect 33325 29928 33337 29984
rect 33257 29926 33337 29928
rect 31978 29903 32024 29914
rect 32449 29868 32519 29882
rect 33441 29868 33521 29870
rect 32449 29812 32461 29868
rect 32517 29812 33453 29868
rect 33509 29812 33521 29868
rect 32449 29800 32519 29812
rect 33441 29810 33521 29812
rect 33770 29868 33850 29870
rect 34213 29868 34273 29880
rect 33770 29812 33782 29868
rect 33838 29812 34215 29868
rect 34271 29812 34273 29868
rect 33770 29810 33850 29812
rect 34213 29800 34273 29812
rect 31645 29752 31809 29764
rect 31645 29696 31657 29752
rect 31713 29696 31809 29752
rect 31645 29684 31809 29696
rect 32215 29752 32293 29763
rect 33625 29752 33705 29754
rect 32215 29751 33637 29752
rect 32215 29697 32227 29751
rect 32281 29697 33637 29751
rect 32215 29696 33637 29697
rect 33693 29696 33705 29752
rect 32215 29685 32293 29696
rect 33625 29694 33705 29696
rect 31029 29618 31049 29674
rect 31105 29618 31125 29674
rect 30345 29497 30356 29543
rect 30430 29497 30441 29543
rect 30610 29534 30860 29545
rect 30268 29451 30314 29462
rect 30251 29392 30268 29402
rect 30472 29451 30610 29462
rect 30314 29392 30331 29402
rect 30251 29336 30263 29392
rect 30319 29336 30331 29392
rect 30251 29326 30268 29336
rect 30314 29326 30331 29336
rect 30268 29266 30314 29277
rect 30518 29277 30610 29451
rect 30472 29266 30610 29277
rect 30130 29054 30176 29194
rect 30345 29185 30356 29231
rect 30430 29185 30441 29231
rect 30345 29154 30441 29185
rect 30656 29194 30814 29534
rect 31029 29543 31125 29618
rect 31029 29497 31040 29543
rect 31114 29497 31125 29543
rect 31294 29534 31340 29545
rect 30860 29451 30998 29462
rect 30860 29277 30952 29451
rect 31156 29451 31202 29462
rect 31139 29392 31156 29402
rect 31202 29392 31219 29402
rect 31139 29336 31151 29392
rect 31207 29336 31219 29392
rect 31139 29326 31156 29336
rect 30860 29266 30998 29277
rect 31202 29326 31219 29336
rect 31156 29266 31202 29277
rect 30610 29183 30860 29194
rect 31029 29185 31040 29231
rect 31114 29185 31125 29231
rect 30656 29054 30814 29183
rect 31029 29154 31125 29185
rect 31294 29054 31340 29194
rect 31498 29534 31544 29545
rect 31713 29543 31809 29684
rect 33257 29602 33337 29616
rect 33044 29580 33090 29591
rect 31713 29497 31724 29543
rect 31798 29497 31809 29543
rect 31978 29534 32024 29545
rect 31544 29451 31682 29462
rect 31544 29277 31636 29451
rect 31840 29451 31886 29462
rect 31823 29392 31840 29402
rect 31886 29392 31903 29402
rect 31823 29336 31835 29392
rect 31891 29336 31903 29392
rect 31823 29326 31840 29336
rect 31544 29266 31682 29277
rect 31886 29326 31903 29336
rect 31840 29266 31886 29277
rect 31498 29054 31544 29194
rect 31713 29185 31724 29231
rect 31798 29185 31809 29231
rect 31713 29154 31809 29185
rect 31978 29054 32024 29194
rect 33257 29546 33269 29602
rect 33325 29546 33337 29602
rect 33441 29602 33521 29616
rect 33441 29546 33453 29602
rect 33509 29546 33521 29602
rect 33625 29602 33705 29616
rect 33625 29546 33637 29602
rect 33693 29546 33705 29602
rect 33872 29580 33918 29591
rect 33259 29543 33270 29546
rect 33324 29543 33335 29546
rect 33443 29543 33454 29546
rect 33508 29543 33519 29546
rect 33627 29543 33638 29546
rect 33692 29543 33703 29546
rect 33182 29497 33228 29508
rect 33090 29323 33182 29497
rect 33182 29312 33228 29323
rect 33366 29497 33412 29508
rect 33366 29312 33412 29323
rect 33550 29497 33596 29508
rect 33734 29497 33780 29508
rect 33717 29470 33734 29472
rect 33780 29470 33797 29472
rect 33717 29350 33729 29470
rect 33785 29350 33797 29470
rect 33717 29348 33734 29350
rect 33550 29312 33596 29323
rect 33780 29348 33797 29350
rect 33734 29312 33780 29323
rect 33044 29095 33090 29240
rect 33259 29231 33270 29277
rect 33324 29231 33335 29277
rect 33259 29198 33335 29231
rect 33443 29231 33454 29277
rect 33508 29231 33519 29277
rect 33443 29198 33519 29231
rect 33627 29231 33638 29277
rect 33692 29231 33703 29277
rect 33627 29198 33703 29231
rect 33872 29095 33918 29240
rect 33032 29083 33112 29095
rect 29750 28739 29796 28750
rect 30093 29014 32061 29054
rect 33032 29027 33044 29083
rect 33100 29027 33112 29083
rect 33032 29015 33112 29027
rect 33850 29083 33930 29095
rect 33850 29027 33862 29083
rect 33918 29027 33930 29083
rect 33850 29015 33930 29027
rect 30093 28874 30193 29014
rect 31961 28874 32061 29014
rect 32266 28965 32352 28977
rect 32459 28965 32519 28969
rect 34355 28965 34411 31902
rect 35111 31900 35191 31902
rect 34743 31808 34823 31822
rect 34530 31786 34576 31797
rect 34743 31752 34755 31808
rect 34811 31752 34823 31808
rect 34927 31808 35007 31822
rect 34927 31752 34939 31808
rect 34995 31752 35007 31808
rect 35111 31808 35191 31822
rect 35111 31752 35123 31808
rect 35179 31752 35191 31808
rect 35358 31786 35404 31797
rect 34745 31749 34756 31752
rect 34810 31749 34821 31752
rect 34929 31749 34940 31752
rect 34994 31749 35005 31752
rect 35113 31749 35124 31752
rect 35178 31749 35189 31752
rect 34668 31703 34714 31714
rect 34576 31529 34668 31703
rect 34668 31518 34714 31529
rect 34852 31703 34898 31714
rect 34852 31518 34898 31529
rect 35036 31703 35082 31714
rect 35220 31703 35266 31714
rect 35203 31676 35220 31678
rect 35266 31676 35283 31678
rect 35203 31556 35215 31676
rect 35271 31556 35283 31676
rect 35203 31554 35220 31556
rect 35036 31518 35082 31529
rect 35266 31554 35283 31556
rect 35220 31518 35266 31529
rect 34530 31301 34576 31446
rect 34745 31437 34756 31483
rect 34810 31437 34821 31483
rect 34745 31404 34821 31437
rect 34929 31437 34940 31483
rect 34994 31437 35005 31483
rect 34929 31404 35005 31437
rect 35113 31437 35124 31483
rect 35178 31437 35189 31483
rect 35113 31404 35189 31437
rect 35358 31301 35404 31446
rect 34518 31289 34598 31301
rect 34518 31233 34530 31289
rect 34586 31233 34598 31289
rect 34518 31221 34598 31233
rect 35336 31289 35414 31301
rect 35336 31233 35348 31289
rect 35404 31233 35414 31289
rect 35336 31221 35414 31233
rect 36443 31170 36643 31970
rect 36843 31170 37043 31970
rect 36443 30550 37043 31170
rect 37374 31830 37420 31841
rect 37589 31839 37685 31870
rect 37589 31793 37600 31839
rect 37674 31793 37685 31839
rect 37854 31830 38308 31970
rect 37512 31747 37558 31758
rect 37495 31463 37512 31473
rect 37716 31747 37854 31758
rect 37558 31463 37575 31473
rect 37495 31223 37507 31463
rect 37563 31223 37575 31463
rect 37495 31213 37512 31223
rect 37558 31213 37575 31223
rect 37512 31162 37558 31173
rect 37762 31173 37854 31747
rect 37716 31162 37854 31173
rect 37374 31079 37420 31090
rect 37589 31081 37600 31127
rect 37674 31081 37685 31127
rect 37589 31006 37685 31081
rect 37900 31162 38262 31830
rect 37854 31079 37900 31090
rect 38477 31839 38573 31870
rect 38477 31793 38488 31839
rect 38562 31793 38573 31839
rect 38742 31830 38788 31970
rect 38308 31747 38446 31758
rect 38308 31173 38400 31747
rect 38604 31747 38650 31758
rect 38587 31463 38604 31473
rect 38650 31463 38667 31473
rect 38587 31223 38599 31463
rect 38655 31223 38667 31463
rect 38587 31213 38604 31223
rect 38308 31162 38446 31173
rect 38650 31213 38667 31223
rect 38604 31162 38650 31173
rect 38262 31079 38308 31090
rect 38477 31081 38488 31127
rect 38562 31081 38573 31127
rect 37589 30950 37609 31006
rect 37665 30950 37685 31006
rect 37589 30732 37685 30950
rect 38477 30862 38573 31081
rect 38957 31839 39053 31870
rect 38957 31793 38968 31839
rect 39042 31793 39053 31839
rect 39222 31830 39268 31970
rect 38788 31747 38926 31758
rect 38788 31173 38880 31747
rect 39084 31747 39130 31758
rect 39067 31463 39084 31473
rect 39130 31463 39147 31473
rect 39067 31223 39079 31463
rect 39135 31223 39147 31463
rect 39067 31213 39084 31223
rect 38788 31162 38926 31173
rect 39130 31213 39147 31223
rect 39084 31162 39130 31173
rect 38742 31079 38788 31090
rect 38957 31081 38968 31127
rect 39042 31081 39053 31127
rect 38957 30940 39053 31081
rect 39222 31079 39268 31090
rect 39565 31170 41033 31970
rect 41333 31170 41533 31970
rect 42057 31957 42127 31969
rect 43097 31957 43177 31959
rect 44583 31958 44663 31960
rect 42057 31901 42069 31957
rect 42125 31901 43109 31957
rect 43165 31901 43177 31957
rect 42057 31889 42127 31901
rect 38409 30850 38573 30862
rect 38889 30928 39053 30940
rect 38889 30872 38901 30928
rect 38957 30872 39053 30928
rect 38889 30860 39053 30872
rect 38409 30794 38421 30850
rect 38477 30794 38573 30850
rect 38409 30782 38573 30794
rect 38477 30732 38573 30782
rect 37374 30710 37420 30721
rect 36480 30410 36526 30550
rect 36695 30419 36791 30450
rect 36695 30373 36706 30419
rect 36780 30373 36791 30419
rect 36960 30410 37006 30550
rect 36526 30327 36664 30338
rect 36526 29753 36618 30327
rect 36822 30327 36868 30338
rect 36805 30043 36822 30053
rect 36868 30043 36885 30053
rect 36805 29803 36817 30043
rect 36873 29803 36885 30043
rect 36805 29793 36822 29803
rect 36526 29742 36664 29753
rect 36868 29793 36885 29803
rect 36822 29742 36868 29753
rect 36480 29659 36526 29670
rect 36695 29661 36706 29707
rect 36780 29661 36791 29707
rect 36695 29520 36791 29661
rect 37589 30719 37889 30732
rect 37589 30673 37600 30719
rect 37674 30686 37804 30719
rect 37674 30673 37685 30686
rect 37793 30673 37804 30686
rect 37878 30673 37889 30719
rect 38058 30710 38104 30721
rect 37420 30627 37558 30638
rect 37420 30453 37512 30627
rect 37716 30627 37762 30638
rect 37699 30568 37716 30578
rect 37920 30627 38058 30638
rect 37762 30568 37779 30578
rect 37699 30512 37711 30568
rect 37767 30512 37779 30568
rect 37699 30502 37716 30512
rect 37420 30442 37558 30453
rect 37762 30502 37779 30512
rect 37716 30442 37762 30453
rect 37966 30453 38058 30627
rect 37920 30442 38058 30453
rect 37374 30230 37420 30370
rect 37589 30361 37600 30407
rect 37674 30361 37685 30407
rect 37589 30330 37685 30361
rect 37793 30361 37804 30407
rect 37878 30361 37889 30407
rect 37793 30330 37889 30361
rect 38273 30719 38573 30732
rect 38273 30673 38284 30719
rect 38358 30686 38488 30719
rect 38358 30673 38369 30686
rect 38477 30673 38488 30686
rect 38562 30673 38573 30719
rect 38742 30710 38788 30721
rect 38196 30627 38242 30638
rect 38179 30568 38196 30578
rect 38400 30627 38446 30638
rect 38242 30568 38259 30578
rect 38179 30512 38191 30568
rect 38247 30512 38259 30568
rect 38179 30502 38196 30512
rect 38242 30502 38259 30512
rect 38383 30568 38400 30578
rect 38604 30627 38650 30638
rect 38446 30568 38463 30578
rect 38383 30512 38395 30568
rect 38451 30512 38463 30568
rect 38383 30502 38400 30512
rect 38196 30442 38242 30453
rect 38446 30502 38463 30512
rect 38587 30568 38604 30578
rect 38650 30568 38667 30578
rect 38587 30512 38599 30568
rect 38655 30512 38667 30568
rect 38587 30502 38604 30512
rect 38400 30442 38446 30453
rect 38650 30502 38667 30512
rect 38604 30442 38650 30453
rect 38058 30230 38104 30370
rect 38273 30361 38284 30407
rect 38358 30361 38369 30407
rect 38273 30330 38369 30361
rect 38477 30361 38488 30407
rect 38562 30361 38573 30407
rect 38477 30330 38573 30361
rect 38957 30719 39053 30860
rect 39565 30974 41533 31170
rect 42341 31170 42397 31901
rect 43097 31899 43177 31901
rect 43827 31902 44595 31958
rect 44651 31902 44663 31958
rect 42729 31807 42809 31821
rect 42516 31785 42562 31796
rect 42729 31751 42741 31807
rect 42797 31751 42809 31807
rect 42913 31807 42993 31821
rect 42913 31751 42925 31807
rect 42981 31751 42993 31807
rect 43097 31807 43177 31821
rect 43097 31751 43109 31807
rect 43165 31751 43177 31807
rect 43344 31785 43390 31796
rect 42731 31748 42742 31751
rect 42796 31748 42807 31751
rect 42915 31748 42926 31751
rect 42980 31748 42991 31751
rect 43099 31748 43110 31751
rect 43164 31748 43175 31751
rect 42654 31702 42700 31713
rect 42562 31528 42654 31702
rect 42654 31517 42700 31528
rect 42838 31702 42884 31713
rect 42838 31517 42884 31528
rect 43022 31702 43068 31713
rect 43206 31702 43252 31713
rect 43189 31675 43206 31677
rect 43252 31675 43269 31677
rect 43189 31555 43201 31675
rect 43257 31555 43269 31675
rect 43189 31553 43206 31555
rect 43022 31517 43068 31528
rect 43252 31553 43269 31555
rect 43206 31517 43252 31528
rect 42516 31300 42562 31445
rect 42731 31436 42742 31482
rect 42796 31436 42807 31482
rect 42731 31403 42807 31436
rect 42915 31436 42926 31482
rect 42980 31436 42991 31482
rect 42915 31403 42991 31436
rect 43099 31436 43110 31482
rect 43164 31436 43175 31482
rect 43099 31403 43175 31436
rect 43344 31300 43390 31445
rect 42504 31288 42584 31300
rect 42504 31232 42516 31288
rect 42572 31232 42584 31288
rect 42504 31220 42584 31232
rect 43322 31288 43400 31300
rect 43322 31232 43334 31288
rect 43390 31232 43400 31288
rect 43322 31220 43400 31232
rect 43675 31170 43755 31180
rect 42341 31114 43687 31170
rect 43743 31114 43755 31170
rect 43675 31112 43755 31114
rect 43509 31061 43579 31063
rect 39565 30834 39665 30974
rect 41433 30834 41533 30974
rect 39565 30794 41533 30834
rect 42341 31060 43579 31061
rect 42341 31006 43511 31060
rect 43567 31006 43579 31060
rect 42341 31005 43579 31006
rect 38957 30673 38968 30719
rect 39042 30673 39053 30719
rect 39222 30710 39268 30721
rect 38788 30627 38926 30638
rect 38788 30453 38880 30627
rect 39084 30627 39130 30638
rect 39067 30568 39084 30578
rect 39130 30568 39147 30578
rect 39067 30512 39079 30568
rect 39135 30512 39147 30568
rect 39067 30502 39084 30512
rect 38788 30442 38926 30453
rect 39130 30502 39147 30512
rect 39084 30442 39130 30453
rect 38742 30230 38788 30370
rect 38957 30361 38968 30407
rect 39042 30361 39053 30407
rect 38957 30330 39053 30361
rect 39222 30230 39268 30370
rect 39602 30654 39648 30794
rect 37337 30200 39305 30230
rect 37337 30060 38605 30200
rect 39205 30060 39305 30200
rect 37337 30030 39305 30060
rect 39817 30663 39913 30694
rect 39817 30617 39828 30663
rect 39902 30617 39913 30663
rect 40021 30663 40117 30694
rect 40021 30617 40032 30663
rect 40106 30617 40117 30663
rect 40286 30654 40332 30794
rect 39648 30571 39786 30582
rect 39944 30571 39990 30582
rect 40148 30571 40286 30582
rect 39648 29997 39740 30571
rect 39927 30331 39939 30571
rect 39995 30331 40007 30571
rect 39648 29986 39786 29997
rect 39944 29986 39990 29997
rect 40194 29997 40286 30571
rect 40148 29986 40286 29997
rect 39602 29903 39648 29914
rect 39817 29905 39828 29951
rect 39902 29931 39913 29951
rect 40021 29931 40032 29951
rect 39902 29905 40032 29931
rect 40106 29905 40117 29951
rect 39817 29878 40117 29905
rect 40501 30663 40597 30694
rect 40501 30617 40512 30663
rect 40586 30617 40597 30663
rect 40705 30663 40801 30694
rect 40705 30617 40716 30663
rect 40790 30617 40801 30663
rect 40970 30654 41016 30794
rect 40424 30571 40470 30582
rect 40628 30571 40674 30582
rect 40832 30571 40878 30582
rect 40611 30331 40623 30571
rect 40679 30331 40691 30571
rect 40407 29997 40419 30237
rect 40475 29997 40487 30237
rect 40815 29997 40827 30237
rect 40883 29997 40895 30237
rect 40424 29986 40470 29997
rect 40628 29986 40674 29997
rect 40832 29986 40878 29997
rect 40286 29903 40332 29914
rect 40501 29905 40512 29951
rect 40586 29931 40597 29951
rect 40705 29931 40716 29951
rect 40586 29905 40716 29931
rect 40790 29905 40801 29951
rect 40501 29878 40801 29905
rect 41185 30663 41281 30694
rect 41185 30617 41196 30663
rect 41270 30617 41281 30663
rect 41450 30654 41496 30794
rect 41016 30571 41154 30582
rect 41016 29997 41108 30571
rect 41312 30571 41358 30582
rect 41295 30287 41312 30297
rect 41358 30287 41375 30297
rect 41295 30047 41307 30287
rect 41363 30047 41375 30287
rect 41295 30037 41312 30047
rect 41016 29986 41154 29997
rect 41358 30037 41375 30047
rect 41312 29986 41358 29997
rect 40970 29903 41016 29914
rect 41185 29905 41196 29951
rect 41270 29905 41281 29951
rect 39817 29830 39913 29878
rect 36960 29659 37006 29670
rect 37337 29800 39305 29830
rect 37337 29660 38605 29800
rect 39205 29660 39305 29800
rect 37337 29630 39305 29660
rect 39817 29774 39837 29830
rect 39893 29774 39913 29830
rect 36627 29508 36791 29520
rect 36627 29452 36639 29508
rect 36695 29452 36791 29508
rect 36627 29440 36791 29452
rect 32266 28909 32278 28965
rect 32334 28909 32461 28965
rect 32517 28909 34411 28965
rect 36480 29290 36526 29301
rect 36695 29299 36791 29440
rect 37374 29490 37420 29501
rect 36695 29253 36706 29299
rect 36780 29253 36791 29299
rect 36960 29290 37006 29301
rect 36526 29207 36664 29218
rect 36526 29033 36618 29207
rect 36822 29207 36868 29218
rect 36805 29148 36822 29158
rect 36868 29148 36885 29158
rect 36805 29092 36817 29148
rect 36873 29092 36885 29148
rect 36805 29082 36822 29092
rect 36526 29022 36664 29033
rect 36868 29082 36885 29092
rect 36822 29022 36868 29033
rect 32266 28897 32352 28909
rect 32459 28897 32519 28909
rect 28937 28510 29101 28522
rect 29417 28588 29581 28600
rect 29417 28532 29429 28588
rect 29485 28532 29581 28588
rect 29417 28520 29581 28532
rect 28937 28454 28949 28510
rect 29005 28454 29101 28510
rect 28937 28442 29101 28454
rect 29005 28392 29101 28442
rect 22389 27890 27571 28090
rect 27902 28370 27948 28381
rect 28117 28379 28417 28392
rect 28117 28333 28128 28379
rect 28202 28346 28332 28379
rect 28202 28333 28213 28346
rect 28321 28333 28332 28346
rect 28406 28333 28417 28379
rect 28586 28370 28632 28381
rect 27948 28287 28086 28298
rect 27948 28113 28040 28287
rect 28244 28287 28290 28298
rect 28227 28228 28244 28238
rect 28448 28287 28586 28298
rect 28290 28228 28307 28238
rect 28227 28172 28239 28228
rect 28295 28172 28307 28228
rect 28227 28162 28244 28172
rect 27948 28102 28086 28113
rect 28290 28162 28307 28172
rect 28244 28102 28290 28113
rect 28494 28113 28586 28287
rect 28448 28102 28586 28113
rect 27902 27890 27948 28030
rect 28117 28021 28128 28067
rect 28202 28021 28213 28067
rect 28117 27990 28213 28021
rect 28321 28021 28332 28067
rect 28406 28021 28417 28067
rect 28321 27990 28417 28021
rect 28801 28379 29101 28392
rect 28801 28333 28812 28379
rect 28886 28346 29016 28379
rect 28886 28333 28897 28346
rect 29005 28333 29016 28346
rect 29090 28333 29101 28379
rect 29270 28370 29316 28381
rect 28724 28287 28770 28298
rect 28707 28228 28724 28238
rect 28928 28287 28974 28298
rect 28770 28228 28787 28238
rect 28707 28172 28719 28228
rect 28775 28172 28787 28228
rect 28707 28162 28724 28172
rect 28770 28162 28787 28172
rect 28911 28228 28928 28238
rect 29132 28287 29178 28298
rect 28974 28228 28991 28238
rect 28911 28172 28923 28228
rect 28979 28172 28991 28228
rect 28911 28162 28928 28172
rect 28724 28102 28770 28113
rect 28974 28162 28991 28172
rect 29115 28228 29132 28238
rect 29178 28228 29195 28238
rect 29115 28172 29127 28228
rect 29183 28172 29195 28228
rect 29115 28162 29132 28172
rect 28928 28102 28974 28113
rect 29178 28162 29195 28172
rect 29132 28102 29178 28113
rect 28586 27890 28632 28030
rect 28801 28021 28812 28067
rect 28886 28021 28897 28067
rect 28801 27990 28897 28021
rect 29005 28021 29016 28067
rect 29090 28021 29101 28067
rect 29005 27990 29101 28021
rect 29485 28379 29581 28520
rect 30093 28690 32061 28874
rect 36480 28810 36526 28950
rect 36695 28941 36706 28987
rect 36780 28941 36791 28987
rect 36695 28910 36791 28941
rect 36960 28810 37006 28950
rect 29485 28333 29496 28379
rect 29570 28333 29581 28379
rect 29750 28370 29796 28381
rect 29316 28287 29454 28298
rect 29316 28113 29408 28287
rect 29612 28287 29658 28298
rect 29595 28228 29612 28238
rect 29658 28228 29675 28238
rect 29595 28172 29607 28228
rect 29663 28172 29675 28228
rect 29595 28162 29612 28172
rect 29316 28102 29454 28113
rect 29658 28162 29675 28172
rect 29612 28102 29658 28113
rect 29270 27890 29316 28030
rect 29485 28021 29496 28067
rect 29570 28021 29581 28067
rect 29485 27990 29581 28021
rect 29750 27890 29796 28030
rect 30093 27890 31561 28690
rect 31861 28090 32061 28690
rect 36443 28090 37043 28810
rect 37589 29499 37685 29530
rect 37589 29453 37600 29499
rect 37674 29453 37685 29499
rect 37854 29490 38308 29630
rect 37512 29407 37558 29418
rect 37495 29123 37512 29133
rect 37716 29407 37854 29418
rect 37558 29123 37575 29133
rect 37495 28883 37507 29123
rect 37563 28883 37575 29123
rect 37495 28873 37512 28883
rect 37558 28873 37575 28883
rect 37512 28822 37558 28833
rect 37762 28833 37854 29407
rect 37716 28822 37854 28833
rect 37374 28739 37420 28750
rect 37589 28741 37600 28787
rect 37674 28741 37685 28787
rect 37589 28666 37685 28741
rect 37900 28822 38262 29490
rect 37854 28739 37900 28750
rect 38477 29499 38573 29530
rect 38477 29453 38488 29499
rect 38562 29453 38573 29499
rect 38742 29490 38788 29630
rect 38308 29407 38446 29418
rect 38308 28833 38400 29407
rect 38604 29407 38650 29418
rect 38587 29123 38604 29133
rect 38650 29123 38667 29133
rect 38587 28883 38599 29123
rect 38655 28883 38667 29123
rect 38587 28873 38604 28883
rect 38308 28822 38446 28833
rect 38650 28873 38667 28883
rect 38604 28822 38650 28833
rect 38262 28739 38308 28750
rect 38477 28741 38488 28787
rect 38562 28741 38573 28787
rect 37589 28610 37609 28666
rect 37665 28610 37685 28666
rect 37589 28392 37685 28610
rect 38477 28522 38573 28741
rect 38957 29499 39053 29530
rect 38957 29453 38968 29499
rect 39042 29453 39053 29499
rect 39222 29490 39268 29630
rect 38788 29407 38926 29418
rect 38788 28833 38880 29407
rect 39084 29407 39130 29418
rect 39067 29123 39084 29133
rect 39130 29123 39147 29133
rect 39067 28883 39079 29123
rect 39135 28883 39147 29123
rect 39067 28873 39084 28883
rect 38788 28822 38926 28833
rect 39130 28873 39147 28883
rect 39084 28822 39130 28833
rect 38742 28739 38788 28750
rect 38957 28741 38968 28787
rect 39042 28741 39053 28787
rect 38957 28600 39053 28741
rect 39602 29534 39648 29545
rect 39817 29543 39913 29774
rect 40501 29674 40597 29878
rect 41185 29764 41281 29905
rect 42341 29984 42397 31005
rect 43509 30997 43579 31005
rect 43005 30953 43091 30957
rect 43005 30897 43017 30953
rect 43073 30897 43091 30953
rect 43005 30885 43091 30897
rect 42516 30740 42562 30751
rect 42731 30749 42807 30782
rect 42731 30703 42742 30749
rect 42796 30703 42807 30749
rect 42915 30749 42991 30782
rect 42915 30703 42926 30749
rect 42980 30703 42991 30749
rect 43099 30749 43175 30782
rect 43099 30703 43110 30749
rect 43164 30703 43175 30749
rect 43344 30740 43390 30751
rect 42654 30657 42700 30668
rect 42637 30630 42654 30632
rect 42838 30657 42884 30668
rect 42700 30630 42717 30632
rect 42562 30510 42649 30630
rect 42705 30510 42717 30630
rect 42637 30508 42654 30510
rect 42562 30210 42654 30330
rect 42700 30508 42717 30510
rect 42821 30330 42838 30332
rect 43022 30657 43068 30668
rect 43005 30630 43022 30632
rect 43206 30657 43252 30668
rect 43068 30630 43085 30632
rect 43005 30510 43017 30630
rect 43073 30510 43085 30630
rect 43005 30508 43022 30510
rect 42884 30330 42901 30332
rect 42821 30210 42833 30330
rect 42889 30210 42901 30330
rect 42821 30208 42838 30210
rect 42654 30172 42700 30183
rect 42884 30208 42901 30210
rect 42838 30172 42884 30183
rect 43068 30508 43085 30510
rect 43189 30330 43206 30332
rect 43327 30630 43344 30632
rect 43390 30630 43407 30632
rect 43327 30509 43339 30630
rect 43395 30509 43407 30630
rect 43327 30507 43344 30509
rect 43252 30330 43269 30332
rect 43189 30210 43201 30330
rect 43257 30210 43269 30330
rect 43189 30208 43206 30210
rect 43022 30172 43068 30183
rect 43252 30208 43269 30210
rect 43206 30172 43252 30183
rect 42731 30134 42742 30137
rect 42796 30134 42807 30137
rect 42915 30134 42926 30137
rect 42980 30134 42991 30137
rect 43099 30134 43110 30137
rect 43164 30134 43175 30137
rect 42516 30089 42562 30100
rect 42729 30078 42741 30134
rect 42797 30078 42809 30134
rect 42729 30064 42809 30078
rect 42913 30078 42925 30134
rect 42981 30078 42993 30134
rect 42913 30064 42993 30078
rect 43097 30078 43109 30134
rect 43165 30078 43177 30134
rect 43390 30507 43407 30509
rect 43344 30089 43390 30100
rect 43097 30064 43177 30078
rect 42729 29984 42809 29986
rect 42341 29928 42741 29984
rect 42797 29928 42809 29984
rect 42729 29926 42809 29928
rect 41450 29903 41496 29914
rect 41921 29868 41991 29882
rect 42913 29868 42993 29870
rect 41921 29812 41933 29868
rect 41989 29812 42925 29868
rect 42981 29812 42993 29868
rect 41921 29800 41991 29812
rect 42913 29810 42993 29812
rect 43242 29868 43322 29870
rect 43685 29868 43745 29880
rect 43242 29812 43254 29868
rect 43310 29812 43687 29868
rect 43743 29812 43745 29868
rect 43242 29810 43322 29812
rect 43685 29800 43745 29812
rect 41117 29752 41281 29764
rect 41117 29696 41129 29752
rect 41185 29696 41281 29752
rect 41117 29684 41281 29696
rect 41687 29752 41765 29763
rect 43097 29752 43177 29754
rect 41687 29751 43109 29752
rect 41687 29697 41699 29751
rect 41753 29697 43109 29751
rect 41687 29696 43109 29697
rect 43165 29696 43177 29752
rect 41687 29685 41765 29696
rect 43097 29694 43177 29696
rect 40501 29618 40521 29674
rect 40577 29618 40597 29674
rect 39817 29497 39828 29543
rect 39902 29497 39913 29543
rect 40082 29534 40332 29545
rect 39740 29451 39786 29462
rect 39723 29392 39740 29402
rect 39944 29451 40082 29462
rect 39786 29392 39803 29402
rect 39723 29336 39735 29392
rect 39791 29336 39803 29392
rect 39723 29326 39740 29336
rect 39786 29326 39803 29336
rect 39740 29266 39786 29277
rect 39990 29277 40082 29451
rect 39944 29266 40082 29277
rect 39602 29054 39648 29194
rect 39817 29185 39828 29231
rect 39902 29185 39913 29231
rect 39817 29154 39913 29185
rect 40128 29194 40286 29534
rect 40501 29543 40597 29618
rect 40501 29497 40512 29543
rect 40586 29497 40597 29543
rect 40766 29534 40812 29545
rect 40332 29451 40470 29462
rect 40332 29277 40424 29451
rect 40628 29451 40674 29462
rect 40611 29392 40628 29402
rect 40674 29392 40691 29402
rect 40611 29336 40623 29392
rect 40679 29336 40691 29392
rect 40611 29326 40628 29336
rect 40332 29266 40470 29277
rect 40674 29326 40691 29336
rect 40628 29266 40674 29277
rect 40082 29183 40332 29194
rect 40501 29185 40512 29231
rect 40586 29185 40597 29231
rect 40128 29054 40286 29183
rect 40501 29154 40597 29185
rect 40766 29054 40812 29194
rect 40970 29534 41016 29545
rect 41185 29543 41281 29684
rect 42729 29602 42809 29616
rect 42516 29580 42562 29591
rect 41185 29497 41196 29543
rect 41270 29497 41281 29543
rect 41450 29534 41496 29545
rect 41016 29451 41154 29462
rect 41016 29277 41108 29451
rect 41312 29451 41358 29462
rect 41295 29392 41312 29402
rect 41358 29392 41375 29402
rect 41295 29336 41307 29392
rect 41363 29336 41375 29392
rect 41295 29326 41312 29336
rect 41016 29266 41154 29277
rect 41358 29326 41375 29336
rect 41312 29266 41358 29277
rect 40970 29054 41016 29194
rect 41185 29185 41196 29231
rect 41270 29185 41281 29231
rect 41185 29154 41281 29185
rect 41450 29054 41496 29194
rect 42729 29546 42741 29602
rect 42797 29546 42809 29602
rect 42913 29602 42993 29616
rect 42913 29546 42925 29602
rect 42981 29546 42993 29602
rect 43097 29602 43177 29616
rect 43097 29546 43109 29602
rect 43165 29546 43177 29602
rect 43344 29580 43390 29591
rect 42731 29543 42742 29546
rect 42796 29543 42807 29546
rect 42915 29543 42926 29546
rect 42980 29543 42991 29546
rect 43099 29543 43110 29546
rect 43164 29543 43175 29546
rect 42654 29497 42700 29508
rect 42562 29323 42654 29497
rect 42654 29312 42700 29323
rect 42838 29497 42884 29508
rect 42838 29312 42884 29323
rect 43022 29497 43068 29508
rect 43206 29497 43252 29508
rect 43189 29470 43206 29472
rect 43252 29470 43269 29472
rect 43189 29350 43201 29470
rect 43257 29350 43269 29470
rect 43189 29348 43206 29350
rect 43022 29312 43068 29323
rect 43252 29348 43269 29350
rect 43206 29312 43252 29323
rect 42516 29095 42562 29240
rect 42731 29231 42742 29277
rect 42796 29231 42807 29277
rect 42731 29198 42807 29231
rect 42915 29231 42926 29277
rect 42980 29231 42991 29277
rect 42915 29198 42991 29231
rect 43099 29231 43110 29277
rect 43164 29231 43175 29277
rect 43099 29198 43175 29231
rect 43344 29095 43390 29240
rect 42504 29083 42584 29095
rect 39222 28739 39268 28750
rect 39565 29014 41533 29054
rect 42504 29027 42516 29083
rect 42572 29027 42584 29083
rect 42504 29015 42584 29027
rect 43322 29083 43402 29095
rect 43322 29027 43334 29083
rect 43390 29027 43402 29083
rect 43322 29015 43402 29027
rect 39565 28874 39665 29014
rect 41433 28874 41533 29014
rect 41738 28965 41824 28977
rect 41931 28965 41991 28969
rect 43827 28965 43883 31902
rect 44583 31900 44663 31902
rect 44215 31808 44295 31822
rect 44002 31786 44048 31797
rect 44215 31752 44227 31808
rect 44283 31752 44295 31808
rect 44399 31808 44479 31822
rect 44399 31752 44411 31808
rect 44467 31752 44479 31808
rect 44583 31808 44663 31822
rect 44583 31752 44595 31808
rect 44651 31752 44663 31808
rect 44830 31786 44876 31797
rect 44217 31749 44228 31752
rect 44282 31749 44293 31752
rect 44401 31749 44412 31752
rect 44466 31749 44477 31752
rect 44585 31749 44596 31752
rect 44650 31749 44661 31752
rect 44140 31703 44186 31714
rect 44048 31529 44140 31703
rect 44140 31518 44186 31529
rect 44324 31703 44370 31714
rect 44324 31518 44370 31529
rect 44508 31703 44554 31714
rect 44692 31703 44738 31714
rect 44675 31676 44692 31678
rect 44738 31676 44755 31678
rect 44675 31556 44687 31676
rect 44743 31556 44755 31676
rect 44675 31554 44692 31556
rect 44508 31518 44554 31529
rect 44738 31554 44755 31556
rect 44692 31518 44738 31529
rect 44002 31301 44048 31446
rect 44217 31437 44228 31483
rect 44282 31437 44293 31483
rect 44217 31404 44293 31437
rect 44401 31437 44412 31483
rect 44466 31437 44477 31483
rect 44401 31404 44477 31437
rect 44585 31437 44596 31483
rect 44650 31437 44661 31483
rect 44585 31404 44661 31437
rect 44830 31301 44876 31446
rect 43990 31289 44070 31301
rect 43990 31233 44002 31289
rect 44058 31233 44070 31289
rect 43990 31221 44070 31233
rect 44808 31289 44886 31301
rect 44808 31233 44820 31289
rect 44876 31233 44886 31289
rect 44808 31221 44886 31233
rect 41738 28909 41750 28965
rect 41806 28909 41933 28965
rect 41989 28909 43883 28965
rect 41738 28897 41824 28909
rect 41931 28897 41991 28909
rect 38409 28510 38573 28522
rect 38889 28588 39053 28600
rect 38889 28532 38901 28588
rect 38957 28532 39053 28588
rect 38889 28520 39053 28532
rect 38409 28454 38421 28510
rect 38477 28454 38573 28510
rect 38409 28442 38573 28454
rect 38477 28392 38573 28442
rect 31861 27890 37043 28090
rect 37374 28370 37420 28381
rect 37589 28379 37889 28392
rect 37589 28333 37600 28379
rect 37674 28346 37804 28379
rect 37674 28333 37685 28346
rect 37793 28333 37804 28346
rect 37878 28333 37889 28379
rect 38058 28370 38104 28381
rect 37420 28287 37558 28298
rect 37420 28113 37512 28287
rect 37716 28287 37762 28298
rect 37699 28228 37716 28238
rect 37920 28287 38058 28298
rect 37762 28228 37779 28238
rect 37699 28172 37711 28228
rect 37767 28172 37779 28228
rect 37699 28162 37716 28172
rect 37420 28102 37558 28113
rect 37762 28162 37779 28172
rect 37716 28102 37762 28113
rect 37966 28113 38058 28287
rect 37920 28102 38058 28113
rect 37374 27890 37420 28030
rect 37589 28021 37600 28067
rect 37674 28021 37685 28067
rect 37589 27990 37685 28021
rect 37793 28021 37804 28067
rect 37878 28021 37889 28067
rect 37793 27990 37889 28021
rect 38273 28379 38573 28392
rect 38273 28333 38284 28379
rect 38358 28346 38488 28379
rect 38358 28333 38369 28346
rect 38477 28333 38488 28346
rect 38562 28333 38573 28379
rect 38742 28370 38788 28381
rect 38196 28287 38242 28298
rect 38179 28228 38196 28238
rect 38400 28287 38446 28298
rect 38242 28228 38259 28238
rect 38179 28172 38191 28228
rect 38247 28172 38259 28228
rect 38179 28162 38196 28172
rect 38242 28162 38259 28172
rect 38383 28228 38400 28238
rect 38604 28287 38650 28298
rect 38446 28228 38463 28238
rect 38383 28172 38395 28228
rect 38451 28172 38463 28228
rect 38383 28162 38400 28172
rect 38196 28102 38242 28113
rect 38446 28162 38463 28172
rect 38587 28228 38604 28238
rect 38650 28228 38667 28238
rect 38587 28172 38599 28228
rect 38655 28172 38667 28228
rect 38587 28162 38604 28172
rect 38400 28102 38446 28113
rect 38650 28162 38667 28172
rect 38604 28102 38650 28113
rect 38058 27890 38104 28030
rect 38273 28021 38284 28067
rect 38358 28021 38369 28067
rect 38273 27990 38369 28021
rect 38477 28021 38488 28067
rect 38562 28021 38573 28067
rect 38477 27990 38573 28021
rect 38957 28379 39053 28520
rect 39565 28690 41533 28874
rect 38957 28333 38968 28379
rect 39042 28333 39053 28379
rect 39222 28370 39268 28381
rect 38788 28287 38926 28298
rect 38788 28113 38880 28287
rect 39084 28287 39130 28298
rect 39067 28228 39084 28238
rect 39130 28228 39147 28238
rect 39067 28172 39079 28228
rect 39135 28172 39147 28228
rect 39067 28162 39084 28172
rect 38788 28102 38926 28113
rect 39130 28162 39147 28172
rect 39084 28102 39130 28113
rect 38742 27890 38788 28030
rect 38957 28021 38968 28067
rect 39042 28021 39053 28067
rect 38957 27990 39053 28021
rect 39222 27890 39268 28030
rect 39565 27890 41033 28690
rect 41333 27890 41533 28690
rect 3445 27889 41533 27890
rect -12446 27577 -12282 27589
rect -12446 27521 -12434 27577
rect -12378 27521 -12282 27577
rect -12446 27509 -12282 27521
rect -12593 27359 -12547 27370
rect -12378 27368 -12282 27509
rect -10921 27690 41533 27889
rect -10921 27689 8027 27690
rect -12378 27322 -12367 27368
rect -12293 27322 -12282 27368
rect -12113 27359 -12067 27370
rect -12547 27276 -12409 27287
rect -12547 27102 -12455 27276
rect -12251 27276 -12205 27287
rect -12268 27217 -12251 27227
rect -12205 27217 -12188 27227
rect -12268 27161 -12256 27217
rect -12200 27161 -12188 27217
rect -12268 27151 -12251 27161
rect -12547 27091 -12409 27102
rect -12205 27151 -12188 27161
rect -12251 27091 -12205 27102
rect -12593 26879 -12547 27019
rect -12378 27010 -12367 27056
rect -12293 27010 -12282 27056
rect -12378 26979 -12282 27010
rect -12113 26879 -12067 27019
rect -10921 26879 -10568 27689
rect -12630 26679 -10568 26879
rect -749 26074 -679 26086
rect 7109 26074 7179 26076
rect -749 26018 -737 26074
rect -681 26018 7111 26074
rect 7167 26018 7179 26074
rect -749 26016 -679 26018
rect 7109 26016 7179 26018
rect 3293 25898 3363 25910
rect 11151 25898 11221 25900
rect 3293 25842 3305 25898
rect 3361 25842 11153 25898
rect 11209 25842 11221 25898
rect 3293 25840 3363 25842
rect 11151 25840 11221 25842
rect -8887 25722 -8817 25734
rect -1029 25722 -959 25724
rect -8887 25666 -8875 25722
rect -8819 25666 -1027 25722
rect -971 25666 -959 25722
rect -8887 25664 -8817 25666
rect -1029 25664 -959 25666
rect 7335 25722 7405 25734
rect 15193 25722 15263 25724
rect 7335 25666 7347 25722
rect 7403 25666 15195 25722
rect 15251 25666 15263 25722
rect 7335 25664 7405 25666
rect 15193 25664 15263 25666
rect -4791 25546 -4721 25558
rect 3067 25546 3137 25548
rect -4791 25490 -4779 25546
rect -4723 25490 3069 25546
rect 3125 25490 3137 25546
rect -4791 25488 -4721 25490
rect 3067 25488 3137 25490
rect 11377 25546 11447 25558
rect 19235 25546 19305 25558
rect 11377 25490 11389 25546
rect 11445 25490 19237 25546
rect 19293 25490 19305 25546
rect 11377 25488 11447 25490
rect 19235 25488 19305 25490
rect -8282 25317 -6735 25373
rect -9241 24296 -9171 24308
rect -8282 24296 -8226 25317
rect -7613 25265 -7527 25269
rect -7613 25209 -7601 25265
rect -7545 25209 -7527 25265
rect -7613 25197 -7527 25209
rect -8102 25052 -8056 25063
rect -7887 25061 -7811 25094
rect -7887 25015 -7876 25061
rect -7822 25015 -7811 25061
rect -7703 25061 -7627 25094
rect -7703 25015 -7692 25061
rect -7638 25015 -7627 25061
rect -7519 25061 -7443 25094
rect -7519 25015 -7508 25061
rect -7454 25015 -7443 25061
rect -7274 25052 -7228 25063
rect -7964 24969 -7918 24980
rect -7981 24942 -7964 24944
rect -7780 24969 -7734 24980
rect -7918 24942 -7901 24944
rect -8056 24822 -7969 24942
rect -7913 24822 -7901 24942
rect -7981 24820 -7964 24822
rect -8056 24522 -7964 24642
rect -7918 24820 -7901 24822
rect -7797 24642 -7780 24644
rect -7596 24969 -7550 24980
rect -7613 24942 -7596 24944
rect -7412 24969 -7366 24980
rect -7550 24942 -7533 24944
rect -7613 24822 -7601 24942
rect -7545 24822 -7533 24942
rect -7613 24820 -7596 24822
rect -7734 24642 -7717 24644
rect -7797 24522 -7785 24642
rect -7729 24522 -7717 24642
rect -7797 24520 -7780 24522
rect -7964 24484 -7918 24495
rect -7734 24520 -7717 24522
rect -7780 24484 -7734 24495
rect -7550 24820 -7533 24822
rect -7429 24642 -7412 24644
rect -7291 24942 -7274 24944
rect -7228 24942 -7211 24944
rect -7291 24821 -7279 24942
rect -7223 24821 -7211 24942
rect -7291 24819 -7274 24821
rect -7366 24642 -7349 24644
rect -7429 24522 -7417 24642
rect -7361 24522 -7349 24642
rect -7429 24520 -7412 24522
rect -7596 24484 -7550 24495
rect -7366 24520 -7349 24522
rect -7412 24484 -7366 24495
rect -7887 24446 -7876 24449
rect -7822 24446 -7811 24449
rect -7703 24446 -7692 24449
rect -7638 24446 -7627 24449
rect -7519 24446 -7508 24449
rect -7454 24446 -7443 24449
rect -8102 24401 -8056 24412
rect -7889 24390 -7877 24446
rect -7821 24390 -7809 24446
rect -7889 24376 -7809 24390
rect -7705 24390 -7693 24446
rect -7637 24390 -7625 24446
rect -7705 24376 -7625 24390
rect -7521 24390 -7509 24446
rect -7453 24390 -7441 24446
rect -7228 24819 -7211 24821
rect -7274 24401 -7228 24412
rect -7521 24376 -7441 24390
rect -7889 24296 -7809 24298
rect -9241 24240 -9229 24296
rect -9173 24240 -7877 24296
rect -7821 24240 -7809 24296
rect -9241 24238 -9171 24240
rect -7889 24238 -7809 24240
rect -8561 24180 -8491 24192
rect -7705 24180 -7625 24182
rect -8561 24124 -8549 24180
rect -8493 24124 -7693 24180
rect -7637 24124 -7625 24180
rect -8561 24112 -8491 24124
rect -7705 24122 -7625 24124
rect -7376 24180 -7296 24182
rect -7109 24180 -7039 24192
rect -7376 24124 -7364 24180
rect -7308 24124 -7107 24180
rect -7051 24124 -7039 24180
rect -7376 24122 -7296 24124
rect -7109 24114 -7039 24124
rect -7521 24064 -7441 24066
rect -8277 24008 -7509 24064
rect -7453 24008 -7441 24064
rect -8277 23277 -8221 24008
rect -7521 24006 -7441 24008
rect -7889 23914 -7809 23928
rect -8102 23892 -8056 23903
rect -7889 23858 -7877 23914
rect -7821 23858 -7809 23914
rect -7705 23914 -7625 23928
rect -7705 23858 -7693 23914
rect -7637 23858 -7625 23914
rect -7521 23914 -7441 23928
rect -7521 23858 -7509 23914
rect -7453 23858 -7441 23914
rect -7274 23892 -7228 23903
rect -7887 23855 -7876 23858
rect -7822 23855 -7811 23858
rect -7703 23855 -7692 23858
rect -7638 23855 -7627 23858
rect -7519 23855 -7508 23858
rect -7454 23855 -7443 23858
rect -7964 23809 -7918 23820
rect -8056 23635 -7964 23809
rect -7964 23624 -7918 23635
rect -7780 23809 -7734 23820
rect -7780 23624 -7734 23635
rect -7596 23809 -7550 23820
rect -7412 23809 -7366 23820
rect -7429 23782 -7412 23784
rect -7366 23782 -7349 23784
rect -7429 23662 -7417 23782
rect -7361 23662 -7349 23782
rect -7429 23660 -7412 23662
rect -7596 23624 -7550 23635
rect -7366 23660 -7349 23662
rect -7412 23624 -7366 23635
rect -8102 23407 -8056 23552
rect -7887 23543 -7876 23589
rect -7822 23543 -7811 23589
rect -7887 23510 -7811 23543
rect -7703 23543 -7692 23589
rect -7638 23543 -7627 23589
rect -7703 23510 -7627 23543
rect -7519 23543 -7508 23589
rect -7454 23543 -7443 23589
rect -7519 23510 -7443 23543
rect -7274 23407 -7228 23552
rect -8114 23395 -8034 23407
rect -8114 23339 -8102 23395
rect -8046 23339 -8034 23395
rect -8114 23327 -8034 23339
rect -7296 23395 -7216 23407
rect -7296 23339 -7284 23395
rect -7228 23339 -7216 23395
rect -7296 23327 -7216 23339
rect -6943 23277 -6863 23287
rect -8277 23221 -6931 23277
rect -6875 23221 -6863 23277
rect -6943 23219 -6863 23221
rect -7109 23168 -7039 23170
rect -8277 23167 -7039 23168
rect -8277 23113 -7107 23167
rect -7051 23113 -7039 23167
rect -8277 23112 -7039 23113
rect -8277 22091 -8221 23112
rect -7109 23104 -7039 23112
rect -7613 23060 -7527 23064
rect -7613 23004 -7601 23060
rect -7545 23004 -7527 23060
rect -7613 22992 -7527 23004
rect -8102 22847 -8056 22858
rect -7887 22856 -7811 22889
rect -7887 22810 -7876 22856
rect -7822 22810 -7811 22856
rect -7703 22856 -7627 22889
rect -7703 22810 -7692 22856
rect -7638 22810 -7627 22856
rect -7519 22856 -7443 22889
rect -7519 22810 -7508 22856
rect -7454 22810 -7443 22856
rect -7274 22847 -7228 22858
rect -7964 22764 -7918 22775
rect -7981 22737 -7964 22739
rect -7780 22764 -7734 22775
rect -7918 22737 -7901 22739
rect -8056 22617 -7969 22737
rect -7913 22617 -7901 22737
rect -7981 22615 -7964 22617
rect -8056 22317 -7964 22437
rect -7918 22615 -7901 22617
rect -7797 22437 -7780 22439
rect -7596 22764 -7550 22775
rect -7613 22737 -7596 22739
rect -7412 22764 -7366 22775
rect -7550 22737 -7533 22739
rect -7613 22617 -7601 22737
rect -7545 22617 -7533 22737
rect -7613 22615 -7596 22617
rect -7734 22437 -7717 22439
rect -7797 22317 -7785 22437
rect -7729 22317 -7717 22437
rect -7797 22315 -7780 22317
rect -7964 22279 -7918 22290
rect -7734 22315 -7717 22317
rect -7780 22279 -7734 22290
rect -7550 22615 -7533 22617
rect -7429 22437 -7412 22439
rect -7291 22737 -7274 22739
rect -7228 22737 -7211 22739
rect -7291 22616 -7279 22737
rect -7223 22616 -7211 22737
rect -7291 22614 -7274 22616
rect -7366 22437 -7349 22439
rect -7429 22317 -7417 22437
rect -7361 22317 -7349 22437
rect -7429 22315 -7412 22317
rect -7596 22279 -7550 22290
rect -7366 22315 -7349 22317
rect -7412 22279 -7366 22290
rect -7887 22241 -7876 22244
rect -7822 22241 -7811 22244
rect -7703 22241 -7692 22244
rect -7638 22241 -7627 22244
rect -7519 22241 -7508 22244
rect -7454 22241 -7443 22244
rect -8102 22196 -8056 22207
rect -7889 22185 -7877 22241
rect -7821 22185 -7809 22241
rect -7889 22171 -7809 22185
rect -7705 22185 -7693 22241
rect -7637 22185 -7625 22241
rect -7705 22171 -7625 22185
rect -7521 22185 -7509 22241
rect -7453 22185 -7441 22241
rect -7228 22614 -7211 22616
rect -7274 22196 -7228 22207
rect -7521 22171 -7441 22185
rect -7889 22091 -7809 22093
rect -8277 22035 -7877 22091
rect -7821 22035 -7809 22091
rect -6791 22091 -6735 25317
rect -4240 25314 -2693 25370
rect -5229 24293 -5159 24305
rect -4240 24293 -4184 25314
rect -3571 25262 -3485 25266
rect -3571 25206 -3559 25262
rect -3503 25206 -3485 25262
rect -3571 25194 -3485 25206
rect -4060 25049 -4014 25060
rect -3845 25058 -3769 25091
rect -3845 25012 -3834 25058
rect -3780 25012 -3769 25058
rect -3661 25058 -3585 25091
rect -3661 25012 -3650 25058
rect -3596 25012 -3585 25058
rect -3477 25058 -3401 25091
rect -3477 25012 -3466 25058
rect -3412 25012 -3401 25058
rect -3232 25049 -3186 25060
rect -3922 24966 -3876 24977
rect -3939 24939 -3922 24941
rect -3738 24966 -3692 24977
rect -3876 24939 -3859 24941
rect -4014 24819 -3927 24939
rect -3871 24819 -3859 24939
rect -3939 24817 -3922 24819
rect -4014 24519 -3922 24639
rect -3876 24817 -3859 24819
rect -3755 24639 -3738 24641
rect -3554 24966 -3508 24977
rect -3571 24939 -3554 24941
rect -3370 24966 -3324 24977
rect -3508 24939 -3491 24941
rect -3571 24819 -3559 24939
rect -3503 24819 -3491 24939
rect -3571 24817 -3554 24819
rect -3692 24639 -3675 24641
rect -3755 24519 -3743 24639
rect -3687 24519 -3675 24639
rect -3755 24517 -3738 24519
rect -3922 24481 -3876 24492
rect -3692 24517 -3675 24519
rect -3738 24481 -3692 24492
rect -3508 24817 -3491 24819
rect -3387 24639 -3370 24641
rect -3249 24939 -3232 24941
rect -3186 24939 -3169 24941
rect -3249 24818 -3237 24939
rect -3181 24818 -3169 24939
rect -3249 24816 -3232 24818
rect -3324 24639 -3307 24641
rect -3387 24519 -3375 24639
rect -3319 24519 -3307 24639
rect -3387 24517 -3370 24519
rect -3554 24481 -3508 24492
rect -3324 24517 -3307 24519
rect -3370 24481 -3324 24492
rect -3845 24443 -3834 24446
rect -3780 24443 -3769 24446
rect -3661 24443 -3650 24446
rect -3596 24443 -3585 24446
rect -3477 24443 -3466 24446
rect -3412 24443 -3401 24446
rect -4060 24398 -4014 24409
rect -3847 24387 -3835 24443
rect -3779 24387 -3767 24443
rect -3847 24373 -3767 24387
rect -3663 24387 -3651 24443
rect -3595 24387 -3583 24443
rect -3663 24373 -3583 24387
rect -3479 24387 -3467 24443
rect -3411 24387 -3399 24443
rect -3186 24816 -3169 24818
rect -3232 24398 -3186 24409
rect -3479 24373 -3399 24387
rect -3847 24293 -3767 24295
rect -5229 24237 -5217 24293
rect -5161 24237 -3835 24293
rect -3779 24237 -3767 24293
rect -5229 24235 -5159 24237
rect -3847 24235 -3767 24237
rect -4519 24177 -4449 24189
rect -3663 24177 -3583 24179
rect -4519 24121 -4507 24177
rect -4451 24121 -3651 24177
rect -3595 24121 -3583 24177
rect -4519 24109 -4449 24121
rect -3663 24119 -3583 24121
rect -3334 24177 -3254 24179
rect -3067 24177 -2997 24189
rect -3334 24121 -3322 24177
rect -3266 24121 -3065 24177
rect -3009 24121 -2997 24177
rect -3334 24119 -3254 24121
rect -3067 24111 -2997 24121
rect -3479 24061 -3399 24063
rect -4235 24005 -3467 24061
rect -3411 24005 -3399 24061
rect -4235 23274 -4179 24005
rect -3479 24003 -3399 24005
rect -3847 23911 -3767 23925
rect -4060 23889 -4014 23900
rect -3847 23855 -3835 23911
rect -3779 23855 -3767 23911
rect -3663 23911 -3583 23925
rect -3663 23855 -3651 23911
rect -3595 23855 -3583 23911
rect -3479 23911 -3399 23925
rect -3479 23855 -3467 23911
rect -3411 23855 -3399 23911
rect -3232 23889 -3186 23900
rect -3845 23852 -3834 23855
rect -3780 23852 -3769 23855
rect -3661 23852 -3650 23855
rect -3596 23852 -3585 23855
rect -3477 23852 -3466 23855
rect -3412 23852 -3401 23855
rect -3922 23806 -3876 23817
rect -4014 23632 -3922 23806
rect -3922 23621 -3876 23632
rect -3738 23806 -3692 23817
rect -3738 23621 -3692 23632
rect -3554 23806 -3508 23817
rect -3370 23806 -3324 23817
rect -3387 23779 -3370 23781
rect -3324 23779 -3307 23781
rect -3387 23659 -3375 23779
rect -3319 23659 -3307 23779
rect -3387 23657 -3370 23659
rect -3554 23621 -3508 23632
rect -3324 23657 -3307 23659
rect -3370 23621 -3324 23632
rect -4060 23404 -4014 23549
rect -3845 23540 -3834 23586
rect -3780 23540 -3769 23586
rect -3845 23507 -3769 23540
rect -3661 23540 -3650 23586
rect -3596 23540 -3585 23586
rect -3661 23507 -3585 23540
rect -3477 23540 -3466 23586
rect -3412 23540 -3401 23586
rect -3477 23507 -3401 23540
rect -3232 23404 -3186 23549
rect -4072 23392 -3992 23404
rect -4072 23336 -4060 23392
rect -4004 23336 -3992 23392
rect -4072 23324 -3992 23336
rect -3254 23392 -3174 23404
rect -3254 23336 -3242 23392
rect -3186 23336 -3174 23392
rect -3254 23324 -3174 23336
rect -2901 23274 -2821 23284
rect -4235 23218 -2889 23274
rect -2833 23218 -2821 23274
rect -2901 23216 -2821 23218
rect -3067 23165 -2997 23167
rect -4235 23164 -2997 23165
rect -4235 23110 -3065 23164
rect -3009 23110 -2997 23164
rect -4235 23109 -2997 23110
rect -6127 23060 -6041 23064
rect -6127 23004 -6115 23060
rect -6059 23004 -6041 23060
rect -6127 22992 -6041 23004
rect -6616 22847 -6570 22858
rect -6401 22856 -6325 22889
rect -6401 22810 -6390 22856
rect -6336 22810 -6325 22856
rect -6217 22856 -6141 22889
rect -6217 22810 -6206 22856
rect -6152 22810 -6141 22856
rect -6033 22856 -5957 22889
rect -6033 22810 -6022 22856
rect -5968 22810 -5957 22856
rect -5788 22847 -5742 22858
rect -6478 22764 -6432 22775
rect -6495 22737 -6478 22739
rect -6294 22764 -6248 22775
rect -6432 22737 -6415 22739
rect -6570 22617 -6483 22737
rect -6427 22617 -6415 22737
rect -6495 22615 -6478 22617
rect -6570 22317 -6478 22437
rect -6432 22615 -6415 22617
rect -6311 22437 -6294 22439
rect -6110 22764 -6064 22775
rect -6127 22737 -6110 22739
rect -5926 22764 -5880 22775
rect -6064 22737 -6047 22739
rect -6127 22617 -6115 22737
rect -6059 22617 -6047 22737
rect -6127 22615 -6110 22617
rect -6248 22437 -6231 22439
rect -6311 22317 -6299 22437
rect -6243 22317 -6231 22437
rect -6311 22315 -6294 22317
rect -6478 22279 -6432 22290
rect -6248 22315 -6231 22317
rect -6294 22279 -6248 22290
rect -6064 22615 -6047 22617
rect -5943 22437 -5926 22439
rect -5805 22737 -5788 22739
rect -5742 22737 -5725 22739
rect -5805 22616 -5793 22737
rect -5737 22616 -5725 22737
rect -5805 22614 -5788 22616
rect -5880 22437 -5863 22439
rect -5943 22317 -5931 22437
rect -5875 22317 -5863 22437
rect -5943 22315 -5926 22317
rect -6110 22279 -6064 22290
rect -5880 22315 -5863 22317
rect -5926 22279 -5880 22290
rect -6401 22241 -6390 22244
rect -6336 22241 -6325 22244
rect -6217 22241 -6206 22244
rect -6152 22241 -6141 22244
rect -6033 22241 -6022 22244
rect -5968 22241 -5957 22244
rect -6616 22196 -6570 22207
rect -6403 22185 -6391 22241
rect -6335 22185 -6323 22241
rect -6403 22171 -6323 22185
rect -6219 22185 -6207 22241
rect -6151 22185 -6139 22241
rect -6219 22171 -6139 22185
rect -6035 22185 -6023 22241
rect -5967 22185 -5955 22241
rect -5742 22614 -5725 22616
rect -5788 22196 -5742 22207
rect -6035 22171 -5955 22185
rect -6403 22091 -6323 22093
rect -6791 22035 -6391 22091
rect -6335 22035 -6323 22091
rect -7889 22033 -7809 22035
rect -6403 22033 -6323 22035
rect -4235 22088 -4179 23109
rect -3067 23101 -2997 23109
rect -3571 23057 -3485 23061
rect -3571 23001 -3559 23057
rect -3503 23001 -3485 23057
rect -3571 22989 -3485 23001
rect -4060 22844 -4014 22855
rect -3845 22853 -3769 22886
rect -3845 22807 -3834 22853
rect -3780 22807 -3769 22853
rect -3661 22853 -3585 22886
rect -3661 22807 -3650 22853
rect -3596 22807 -3585 22853
rect -3477 22853 -3401 22886
rect -3477 22807 -3466 22853
rect -3412 22807 -3401 22853
rect -3232 22844 -3186 22855
rect -3922 22761 -3876 22772
rect -3939 22734 -3922 22736
rect -3738 22761 -3692 22772
rect -3876 22734 -3859 22736
rect -4014 22614 -3927 22734
rect -3871 22614 -3859 22734
rect -3939 22612 -3922 22614
rect -4014 22314 -3922 22434
rect -3876 22612 -3859 22614
rect -3755 22434 -3738 22436
rect -3554 22761 -3508 22772
rect -3571 22734 -3554 22736
rect -3370 22761 -3324 22772
rect -3508 22734 -3491 22736
rect -3571 22614 -3559 22734
rect -3503 22614 -3491 22734
rect -3571 22612 -3554 22614
rect -3692 22434 -3675 22436
rect -3755 22314 -3743 22434
rect -3687 22314 -3675 22434
rect -3755 22312 -3738 22314
rect -3922 22276 -3876 22287
rect -3692 22312 -3675 22314
rect -3738 22276 -3692 22287
rect -3508 22612 -3491 22614
rect -3387 22434 -3370 22436
rect -3249 22734 -3232 22736
rect -3186 22734 -3169 22736
rect -3249 22613 -3237 22734
rect -3181 22613 -3169 22734
rect -3249 22611 -3232 22613
rect -3324 22434 -3307 22436
rect -3387 22314 -3375 22434
rect -3319 22314 -3307 22434
rect -3387 22312 -3370 22314
rect -3554 22276 -3508 22287
rect -3324 22312 -3307 22314
rect -3370 22276 -3324 22287
rect -3845 22238 -3834 22241
rect -3780 22238 -3769 22241
rect -3661 22238 -3650 22241
rect -3596 22238 -3585 22241
rect -3477 22238 -3466 22241
rect -3412 22238 -3401 22241
rect -4060 22193 -4014 22204
rect -3847 22182 -3835 22238
rect -3779 22182 -3767 22238
rect -3847 22168 -3767 22182
rect -3663 22182 -3651 22238
rect -3595 22182 -3583 22238
rect -3663 22168 -3583 22182
rect -3479 22182 -3467 22238
rect -3411 22182 -3399 22238
rect -3186 22611 -3169 22613
rect -3232 22193 -3186 22204
rect -3479 22168 -3399 22182
rect -3847 22088 -3767 22090
rect -4235 22032 -3835 22088
rect -3779 22032 -3767 22088
rect -2749 22088 -2693 25314
rect -198 25314 1349 25370
rect -1187 24293 -1117 24305
rect -198 24293 -142 25314
rect 471 25262 557 25266
rect 471 25206 483 25262
rect 539 25206 557 25262
rect 471 25194 557 25206
rect -18 25049 28 25060
rect 197 25058 273 25091
rect 197 25012 208 25058
rect 262 25012 273 25058
rect 381 25058 457 25091
rect 381 25012 392 25058
rect 446 25012 457 25058
rect 565 25058 641 25091
rect 565 25012 576 25058
rect 630 25012 641 25058
rect 810 25049 856 25060
rect 120 24966 166 24977
rect 103 24939 120 24941
rect 304 24966 350 24977
rect 166 24939 183 24941
rect 28 24819 115 24939
rect 171 24819 183 24939
rect 103 24817 120 24819
rect 28 24519 120 24639
rect 166 24817 183 24819
rect 287 24639 304 24641
rect 488 24966 534 24977
rect 471 24939 488 24941
rect 672 24966 718 24977
rect 534 24939 551 24941
rect 471 24819 483 24939
rect 539 24819 551 24939
rect 471 24817 488 24819
rect 350 24639 367 24641
rect 287 24519 299 24639
rect 355 24519 367 24639
rect 287 24517 304 24519
rect 120 24481 166 24492
rect 350 24517 367 24519
rect 304 24481 350 24492
rect 534 24817 551 24819
rect 655 24639 672 24641
rect 793 24939 810 24941
rect 856 24939 873 24941
rect 793 24818 805 24939
rect 861 24818 873 24939
rect 793 24816 810 24818
rect 718 24639 735 24641
rect 655 24519 667 24639
rect 723 24519 735 24639
rect 655 24517 672 24519
rect 488 24481 534 24492
rect 718 24517 735 24519
rect 672 24481 718 24492
rect 197 24443 208 24446
rect 262 24443 273 24446
rect 381 24443 392 24446
rect 446 24443 457 24446
rect 565 24443 576 24446
rect 630 24443 641 24446
rect -18 24398 28 24409
rect 195 24387 207 24443
rect 263 24387 275 24443
rect 195 24373 275 24387
rect 379 24387 391 24443
rect 447 24387 459 24443
rect 379 24373 459 24387
rect 563 24387 575 24443
rect 631 24387 643 24443
rect 856 24816 873 24818
rect 810 24398 856 24409
rect 563 24373 643 24387
rect 195 24293 275 24295
rect -1187 24237 -1175 24293
rect -1119 24237 207 24293
rect 263 24237 275 24293
rect -1187 24235 -1117 24237
rect 195 24235 275 24237
rect -477 24177 -407 24189
rect 379 24177 459 24179
rect -477 24121 -465 24177
rect -409 24121 391 24177
rect 447 24121 459 24177
rect -477 24109 -407 24121
rect 379 24119 459 24121
rect 708 24177 788 24179
rect 975 24177 1045 24189
rect 708 24121 720 24177
rect 776 24121 977 24177
rect 1033 24121 1045 24177
rect 708 24119 788 24121
rect 975 24111 1045 24121
rect 563 24061 643 24063
rect -193 24005 575 24061
rect 631 24005 643 24061
rect -193 23274 -137 24005
rect 563 24003 643 24005
rect 195 23911 275 23925
rect -18 23889 28 23900
rect 195 23855 207 23911
rect 263 23855 275 23911
rect 379 23911 459 23925
rect 379 23855 391 23911
rect 447 23855 459 23911
rect 563 23911 643 23925
rect 563 23855 575 23911
rect 631 23855 643 23911
rect 810 23889 856 23900
rect 197 23852 208 23855
rect 262 23852 273 23855
rect 381 23852 392 23855
rect 446 23852 457 23855
rect 565 23852 576 23855
rect 630 23852 641 23855
rect 120 23806 166 23817
rect 28 23632 120 23806
rect 120 23621 166 23632
rect 304 23806 350 23817
rect 304 23621 350 23632
rect 488 23806 534 23817
rect 672 23806 718 23817
rect 655 23779 672 23781
rect 718 23779 735 23781
rect 655 23659 667 23779
rect 723 23659 735 23779
rect 655 23657 672 23659
rect 488 23621 534 23632
rect 718 23657 735 23659
rect 672 23621 718 23632
rect -18 23404 28 23549
rect 197 23540 208 23586
rect 262 23540 273 23586
rect 197 23507 273 23540
rect 381 23540 392 23586
rect 446 23540 457 23586
rect 381 23507 457 23540
rect 565 23540 576 23586
rect 630 23540 641 23586
rect 565 23507 641 23540
rect 810 23404 856 23549
rect -30 23392 50 23404
rect -30 23336 -18 23392
rect 38 23336 50 23392
rect -30 23324 50 23336
rect 788 23392 868 23404
rect 788 23336 800 23392
rect 856 23336 868 23392
rect 788 23324 868 23336
rect 1141 23274 1221 23284
rect -193 23218 1153 23274
rect 1209 23218 1221 23274
rect 1141 23216 1221 23218
rect 975 23165 1045 23167
rect -193 23164 1045 23165
rect -193 23110 977 23164
rect 1033 23110 1045 23164
rect -193 23109 1045 23110
rect -2085 23057 -1999 23061
rect -2085 23001 -2073 23057
rect -2017 23001 -1999 23057
rect -2085 22989 -1999 23001
rect -2574 22844 -2528 22855
rect -2359 22853 -2283 22886
rect -2359 22807 -2348 22853
rect -2294 22807 -2283 22853
rect -2175 22853 -2099 22886
rect -2175 22807 -2164 22853
rect -2110 22807 -2099 22853
rect -1991 22853 -1915 22886
rect -1991 22807 -1980 22853
rect -1926 22807 -1915 22853
rect -1746 22844 -1700 22855
rect -2436 22761 -2390 22772
rect -2453 22734 -2436 22736
rect -2252 22761 -2206 22772
rect -2390 22734 -2373 22736
rect -2528 22614 -2441 22734
rect -2385 22614 -2373 22734
rect -2453 22612 -2436 22614
rect -2528 22314 -2436 22434
rect -2390 22612 -2373 22614
rect -2269 22434 -2252 22436
rect -2068 22761 -2022 22772
rect -2085 22734 -2068 22736
rect -1884 22761 -1838 22772
rect -2022 22734 -2005 22736
rect -2085 22614 -2073 22734
rect -2017 22614 -2005 22734
rect -2085 22612 -2068 22614
rect -2206 22434 -2189 22436
rect -2269 22314 -2257 22434
rect -2201 22314 -2189 22434
rect -2269 22312 -2252 22314
rect -2436 22276 -2390 22287
rect -2206 22312 -2189 22314
rect -2252 22276 -2206 22287
rect -2022 22612 -2005 22614
rect -1901 22434 -1884 22436
rect -1763 22734 -1746 22736
rect -1700 22734 -1683 22736
rect -1763 22613 -1751 22734
rect -1695 22613 -1683 22734
rect -1763 22611 -1746 22613
rect -1838 22434 -1821 22436
rect -1901 22314 -1889 22434
rect -1833 22314 -1821 22434
rect -1901 22312 -1884 22314
rect -2068 22276 -2022 22287
rect -1838 22312 -1821 22314
rect -1884 22276 -1838 22287
rect -2359 22238 -2348 22241
rect -2294 22238 -2283 22241
rect -2175 22238 -2164 22241
rect -2110 22238 -2099 22241
rect -1991 22238 -1980 22241
rect -1926 22238 -1915 22241
rect -2574 22193 -2528 22204
rect -2361 22182 -2349 22238
rect -2293 22182 -2281 22238
rect -2361 22168 -2281 22182
rect -2177 22182 -2165 22238
rect -2109 22182 -2097 22238
rect -2177 22168 -2097 22182
rect -1993 22182 -1981 22238
rect -1925 22182 -1913 22238
rect -1700 22611 -1683 22613
rect -1746 22193 -1700 22204
rect -1993 22168 -1913 22182
rect -2361 22088 -2281 22090
rect -2749 22032 -2349 22088
rect -2293 22032 -2281 22088
rect -193 22088 -137 23109
rect 975 23101 1045 23109
rect 471 23057 557 23061
rect 471 23001 483 23057
rect 539 23001 557 23057
rect 471 22989 557 23001
rect -18 22844 28 22855
rect 197 22853 273 22886
rect 197 22807 208 22853
rect 262 22807 273 22853
rect 381 22853 457 22886
rect 381 22807 392 22853
rect 446 22807 457 22853
rect 565 22853 641 22886
rect 565 22807 576 22853
rect 630 22807 641 22853
rect 810 22844 856 22855
rect 120 22761 166 22772
rect 103 22734 120 22736
rect 304 22761 350 22772
rect 166 22734 183 22736
rect 28 22614 115 22734
rect 171 22614 183 22734
rect 103 22612 120 22614
rect 28 22314 120 22434
rect 166 22612 183 22614
rect 287 22434 304 22436
rect 488 22761 534 22772
rect 471 22734 488 22736
rect 672 22761 718 22772
rect 534 22734 551 22736
rect 471 22614 483 22734
rect 539 22614 551 22734
rect 471 22612 488 22614
rect 350 22434 367 22436
rect 287 22314 299 22434
rect 355 22314 367 22434
rect 287 22312 304 22314
rect 120 22276 166 22287
rect 350 22312 367 22314
rect 304 22276 350 22287
rect 534 22612 551 22614
rect 655 22434 672 22436
rect 793 22734 810 22736
rect 856 22734 873 22736
rect 793 22613 805 22734
rect 861 22613 873 22734
rect 793 22611 810 22613
rect 718 22434 735 22436
rect 655 22314 667 22434
rect 723 22314 735 22434
rect 655 22312 672 22314
rect 488 22276 534 22287
rect 718 22312 735 22314
rect 672 22276 718 22287
rect 197 22238 208 22241
rect 262 22238 273 22241
rect 381 22238 392 22241
rect 446 22238 457 22241
rect 565 22238 576 22241
rect 630 22238 641 22241
rect -18 22193 28 22204
rect 195 22182 207 22238
rect 263 22182 275 22238
rect 195 22168 275 22182
rect 379 22182 391 22238
rect 447 22182 459 22238
rect 379 22168 459 22182
rect 563 22182 575 22238
rect 631 22182 643 22238
rect 856 22611 873 22613
rect 810 22193 856 22204
rect 563 22168 643 22182
rect 195 22088 275 22090
rect -193 22032 207 22088
rect 263 22032 275 22088
rect 1293 22088 1349 25314
rect 3844 25314 5391 25370
rect 2855 24293 2925 24305
rect 3844 24293 3900 25314
rect 4513 25262 4599 25266
rect 4513 25206 4525 25262
rect 4581 25206 4599 25262
rect 4513 25194 4599 25206
rect 4024 25049 4070 25060
rect 4239 25058 4315 25091
rect 4239 25012 4250 25058
rect 4304 25012 4315 25058
rect 4423 25058 4499 25091
rect 4423 25012 4434 25058
rect 4488 25012 4499 25058
rect 4607 25058 4683 25091
rect 4607 25012 4618 25058
rect 4672 25012 4683 25058
rect 4852 25049 4898 25060
rect 4162 24966 4208 24977
rect 4145 24939 4162 24941
rect 4346 24966 4392 24977
rect 4208 24939 4225 24941
rect 4070 24819 4157 24939
rect 4213 24819 4225 24939
rect 4145 24817 4162 24819
rect 4070 24519 4162 24639
rect 4208 24817 4225 24819
rect 4329 24639 4346 24641
rect 4530 24966 4576 24977
rect 4513 24939 4530 24941
rect 4714 24966 4760 24977
rect 4576 24939 4593 24941
rect 4513 24819 4525 24939
rect 4581 24819 4593 24939
rect 4513 24817 4530 24819
rect 4392 24639 4409 24641
rect 4329 24519 4341 24639
rect 4397 24519 4409 24639
rect 4329 24517 4346 24519
rect 4162 24481 4208 24492
rect 4392 24517 4409 24519
rect 4346 24481 4392 24492
rect 4576 24817 4593 24819
rect 4697 24639 4714 24641
rect 4835 24939 4852 24941
rect 4898 24939 4915 24941
rect 4835 24818 4847 24939
rect 4903 24818 4915 24939
rect 4835 24816 4852 24818
rect 4760 24639 4777 24641
rect 4697 24519 4709 24639
rect 4765 24519 4777 24639
rect 4697 24517 4714 24519
rect 4530 24481 4576 24492
rect 4760 24517 4777 24519
rect 4714 24481 4760 24492
rect 4239 24443 4250 24446
rect 4304 24443 4315 24446
rect 4423 24443 4434 24446
rect 4488 24443 4499 24446
rect 4607 24443 4618 24446
rect 4672 24443 4683 24446
rect 4024 24398 4070 24409
rect 4237 24387 4249 24443
rect 4305 24387 4317 24443
rect 4237 24373 4317 24387
rect 4421 24387 4433 24443
rect 4489 24387 4501 24443
rect 4421 24373 4501 24387
rect 4605 24387 4617 24443
rect 4673 24387 4685 24443
rect 4898 24816 4915 24818
rect 4852 24398 4898 24409
rect 4605 24373 4685 24387
rect 4237 24293 4317 24295
rect 2855 24237 2867 24293
rect 2923 24237 4249 24293
rect 4305 24237 4317 24293
rect 2855 24235 2925 24237
rect 4237 24235 4317 24237
rect 3565 24177 3635 24189
rect 4421 24177 4501 24179
rect 3565 24121 3577 24177
rect 3633 24121 4433 24177
rect 4489 24121 4501 24177
rect 3565 24109 3635 24121
rect 4421 24119 4501 24121
rect 4750 24177 4830 24179
rect 5017 24177 5087 24189
rect 4750 24121 4762 24177
rect 4818 24121 5019 24177
rect 5075 24121 5087 24177
rect 4750 24119 4830 24121
rect 5017 24111 5087 24121
rect 4605 24061 4685 24063
rect 3849 24005 4617 24061
rect 4673 24005 4685 24061
rect 3849 23274 3905 24005
rect 4605 24003 4685 24005
rect 4237 23911 4317 23925
rect 4024 23889 4070 23900
rect 4237 23855 4249 23911
rect 4305 23855 4317 23911
rect 4421 23911 4501 23925
rect 4421 23855 4433 23911
rect 4489 23855 4501 23911
rect 4605 23911 4685 23925
rect 4605 23855 4617 23911
rect 4673 23855 4685 23911
rect 4852 23889 4898 23900
rect 4239 23852 4250 23855
rect 4304 23852 4315 23855
rect 4423 23852 4434 23855
rect 4488 23852 4499 23855
rect 4607 23852 4618 23855
rect 4672 23852 4683 23855
rect 4162 23806 4208 23817
rect 4070 23632 4162 23806
rect 4162 23621 4208 23632
rect 4346 23806 4392 23817
rect 4346 23621 4392 23632
rect 4530 23806 4576 23817
rect 4714 23806 4760 23817
rect 4697 23779 4714 23781
rect 4760 23779 4777 23781
rect 4697 23659 4709 23779
rect 4765 23659 4777 23779
rect 4697 23657 4714 23659
rect 4530 23621 4576 23632
rect 4760 23657 4777 23659
rect 4714 23621 4760 23632
rect 4024 23404 4070 23549
rect 4239 23540 4250 23586
rect 4304 23540 4315 23586
rect 4239 23507 4315 23540
rect 4423 23540 4434 23586
rect 4488 23540 4499 23586
rect 4423 23507 4499 23540
rect 4607 23540 4618 23586
rect 4672 23540 4683 23586
rect 4607 23507 4683 23540
rect 4852 23404 4898 23549
rect 4012 23392 4092 23404
rect 4012 23336 4024 23392
rect 4080 23336 4092 23392
rect 4012 23324 4092 23336
rect 4830 23392 4910 23404
rect 4830 23336 4842 23392
rect 4898 23336 4910 23392
rect 4830 23324 4910 23336
rect 5183 23274 5263 23284
rect 3849 23218 5195 23274
rect 5251 23218 5263 23274
rect 5183 23216 5263 23218
rect 5017 23165 5087 23167
rect 3849 23164 5087 23165
rect 3849 23110 5019 23164
rect 5075 23110 5087 23164
rect 3849 23109 5087 23110
rect 1957 23057 2043 23061
rect 1957 23001 1969 23057
rect 2025 23001 2043 23057
rect 1957 22989 2043 23001
rect 1468 22844 1514 22855
rect 1683 22853 1759 22886
rect 1683 22807 1694 22853
rect 1748 22807 1759 22853
rect 1867 22853 1943 22886
rect 1867 22807 1878 22853
rect 1932 22807 1943 22853
rect 2051 22853 2127 22886
rect 2051 22807 2062 22853
rect 2116 22807 2127 22853
rect 2296 22844 2342 22855
rect 1606 22761 1652 22772
rect 1589 22734 1606 22736
rect 1790 22761 1836 22772
rect 1652 22734 1669 22736
rect 1514 22614 1601 22734
rect 1657 22614 1669 22734
rect 1589 22612 1606 22614
rect 1514 22314 1606 22434
rect 1652 22612 1669 22614
rect 1773 22434 1790 22436
rect 1974 22761 2020 22772
rect 1957 22734 1974 22736
rect 2158 22761 2204 22772
rect 2020 22734 2037 22736
rect 1957 22614 1969 22734
rect 2025 22614 2037 22734
rect 1957 22612 1974 22614
rect 1836 22434 1853 22436
rect 1773 22314 1785 22434
rect 1841 22314 1853 22434
rect 1773 22312 1790 22314
rect 1606 22276 1652 22287
rect 1836 22312 1853 22314
rect 1790 22276 1836 22287
rect 2020 22612 2037 22614
rect 2141 22434 2158 22436
rect 2279 22734 2296 22736
rect 2342 22734 2359 22736
rect 2279 22613 2291 22734
rect 2347 22613 2359 22734
rect 2279 22611 2296 22613
rect 2204 22434 2221 22436
rect 2141 22314 2153 22434
rect 2209 22314 2221 22434
rect 2141 22312 2158 22314
rect 1974 22276 2020 22287
rect 2204 22312 2221 22314
rect 2158 22276 2204 22287
rect 1683 22238 1694 22241
rect 1748 22238 1759 22241
rect 1867 22238 1878 22241
rect 1932 22238 1943 22241
rect 2051 22238 2062 22241
rect 2116 22238 2127 22241
rect 1468 22193 1514 22204
rect 1681 22182 1693 22238
rect 1749 22182 1761 22238
rect 1681 22168 1761 22182
rect 1865 22182 1877 22238
rect 1933 22182 1945 22238
rect 1865 22168 1945 22182
rect 2049 22182 2061 22238
rect 2117 22182 2129 22238
rect 2342 22611 2359 22613
rect 2296 22193 2342 22204
rect 2049 22168 2129 22182
rect 1681 22088 1761 22090
rect 1293 22032 1693 22088
rect 1749 22032 1761 22088
rect 3849 22088 3905 23109
rect 5017 23101 5087 23109
rect 4513 23057 4599 23061
rect 4513 23001 4525 23057
rect 4581 23001 4599 23057
rect 4513 22989 4599 23001
rect 4024 22844 4070 22855
rect 4239 22853 4315 22886
rect 4239 22807 4250 22853
rect 4304 22807 4315 22853
rect 4423 22853 4499 22886
rect 4423 22807 4434 22853
rect 4488 22807 4499 22853
rect 4607 22853 4683 22886
rect 4607 22807 4618 22853
rect 4672 22807 4683 22853
rect 4852 22844 4898 22855
rect 4162 22761 4208 22772
rect 4145 22734 4162 22736
rect 4346 22761 4392 22772
rect 4208 22734 4225 22736
rect 4070 22614 4157 22734
rect 4213 22614 4225 22734
rect 4145 22612 4162 22614
rect 4070 22314 4162 22434
rect 4208 22612 4225 22614
rect 4329 22434 4346 22436
rect 4530 22761 4576 22772
rect 4513 22734 4530 22736
rect 4714 22761 4760 22772
rect 4576 22734 4593 22736
rect 4513 22614 4525 22734
rect 4581 22614 4593 22734
rect 4513 22612 4530 22614
rect 4392 22434 4409 22436
rect 4329 22314 4341 22434
rect 4397 22314 4409 22434
rect 4329 22312 4346 22314
rect 4162 22276 4208 22287
rect 4392 22312 4409 22314
rect 4346 22276 4392 22287
rect 4576 22612 4593 22614
rect 4697 22434 4714 22436
rect 4835 22734 4852 22736
rect 4898 22734 4915 22736
rect 4835 22613 4847 22734
rect 4903 22613 4915 22734
rect 4835 22611 4852 22613
rect 4760 22434 4777 22436
rect 4697 22314 4709 22434
rect 4765 22314 4777 22434
rect 4697 22312 4714 22314
rect 4530 22276 4576 22287
rect 4760 22312 4777 22314
rect 4714 22276 4760 22287
rect 4239 22238 4250 22241
rect 4304 22238 4315 22241
rect 4423 22238 4434 22241
rect 4488 22238 4499 22241
rect 4607 22238 4618 22241
rect 4672 22238 4683 22241
rect 4024 22193 4070 22204
rect 4237 22182 4249 22238
rect 4305 22182 4317 22238
rect 4237 22168 4317 22182
rect 4421 22182 4433 22238
rect 4489 22182 4501 22238
rect 4421 22168 4501 22182
rect 4605 22182 4617 22238
rect 4673 22182 4685 22238
rect 4898 22611 4915 22613
rect 4852 22193 4898 22204
rect 4605 22168 4685 22182
rect 4237 22088 4317 22090
rect 3849 22032 4249 22088
rect 4305 22032 4317 22088
rect 5335 22088 5391 25314
rect 7886 25314 9433 25370
rect 6897 24293 6967 24305
rect 7886 24293 7942 25314
rect 8555 25262 8641 25266
rect 8555 25206 8567 25262
rect 8623 25206 8641 25262
rect 8555 25194 8641 25206
rect 8066 25049 8112 25060
rect 8281 25058 8357 25091
rect 8281 25012 8292 25058
rect 8346 25012 8357 25058
rect 8465 25058 8541 25091
rect 8465 25012 8476 25058
rect 8530 25012 8541 25058
rect 8649 25058 8725 25091
rect 8649 25012 8660 25058
rect 8714 25012 8725 25058
rect 8894 25049 8940 25060
rect 8204 24966 8250 24977
rect 8187 24939 8204 24941
rect 8388 24966 8434 24977
rect 8250 24939 8267 24941
rect 8112 24819 8199 24939
rect 8255 24819 8267 24939
rect 8187 24817 8204 24819
rect 8112 24519 8204 24639
rect 8250 24817 8267 24819
rect 8371 24639 8388 24641
rect 8572 24966 8618 24977
rect 8555 24939 8572 24941
rect 8756 24966 8802 24977
rect 8618 24939 8635 24941
rect 8555 24819 8567 24939
rect 8623 24819 8635 24939
rect 8555 24817 8572 24819
rect 8434 24639 8451 24641
rect 8371 24519 8383 24639
rect 8439 24519 8451 24639
rect 8371 24517 8388 24519
rect 8204 24481 8250 24492
rect 8434 24517 8451 24519
rect 8388 24481 8434 24492
rect 8618 24817 8635 24819
rect 8739 24639 8756 24641
rect 8877 24939 8894 24941
rect 8940 24939 8957 24941
rect 8877 24818 8889 24939
rect 8945 24818 8957 24939
rect 8877 24816 8894 24818
rect 8802 24639 8819 24641
rect 8739 24519 8751 24639
rect 8807 24519 8819 24639
rect 8739 24517 8756 24519
rect 8572 24481 8618 24492
rect 8802 24517 8819 24519
rect 8756 24481 8802 24492
rect 8281 24443 8292 24446
rect 8346 24443 8357 24446
rect 8465 24443 8476 24446
rect 8530 24443 8541 24446
rect 8649 24443 8660 24446
rect 8714 24443 8725 24446
rect 8066 24398 8112 24409
rect 8279 24387 8291 24443
rect 8347 24387 8359 24443
rect 8279 24373 8359 24387
rect 8463 24387 8475 24443
rect 8531 24387 8543 24443
rect 8463 24373 8543 24387
rect 8647 24387 8659 24443
rect 8715 24387 8727 24443
rect 8940 24816 8957 24818
rect 8894 24398 8940 24409
rect 8647 24373 8727 24387
rect 8279 24293 8359 24295
rect 6897 24237 6909 24293
rect 6965 24237 8291 24293
rect 8347 24237 8359 24293
rect 6897 24235 6967 24237
rect 8279 24235 8359 24237
rect 7607 24177 7677 24189
rect 8463 24177 8543 24179
rect 7607 24121 7619 24177
rect 7675 24121 8475 24177
rect 8531 24121 8543 24177
rect 7607 24109 7677 24121
rect 8463 24119 8543 24121
rect 8792 24177 8872 24179
rect 9059 24177 9129 24189
rect 8792 24121 8804 24177
rect 8860 24121 9061 24177
rect 9117 24121 9129 24177
rect 8792 24119 8872 24121
rect 9059 24111 9129 24121
rect 8647 24061 8727 24063
rect 7891 24005 8659 24061
rect 8715 24005 8727 24061
rect 7891 23274 7947 24005
rect 8647 24003 8727 24005
rect 8279 23911 8359 23925
rect 8066 23889 8112 23900
rect 8279 23855 8291 23911
rect 8347 23855 8359 23911
rect 8463 23911 8543 23925
rect 8463 23855 8475 23911
rect 8531 23855 8543 23911
rect 8647 23911 8727 23925
rect 8647 23855 8659 23911
rect 8715 23855 8727 23911
rect 8894 23889 8940 23900
rect 8281 23852 8292 23855
rect 8346 23852 8357 23855
rect 8465 23852 8476 23855
rect 8530 23852 8541 23855
rect 8649 23852 8660 23855
rect 8714 23852 8725 23855
rect 8204 23806 8250 23817
rect 8112 23632 8204 23806
rect 8204 23621 8250 23632
rect 8388 23806 8434 23817
rect 8388 23621 8434 23632
rect 8572 23806 8618 23817
rect 8756 23806 8802 23817
rect 8739 23779 8756 23781
rect 8802 23779 8819 23781
rect 8739 23659 8751 23779
rect 8807 23659 8819 23779
rect 8739 23657 8756 23659
rect 8572 23621 8618 23632
rect 8802 23657 8819 23659
rect 8756 23621 8802 23632
rect 8066 23404 8112 23549
rect 8281 23540 8292 23586
rect 8346 23540 8357 23586
rect 8281 23507 8357 23540
rect 8465 23540 8476 23586
rect 8530 23540 8541 23586
rect 8465 23507 8541 23540
rect 8649 23540 8660 23586
rect 8714 23540 8725 23586
rect 8649 23507 8725 23540
rect 8894 23404 8940 23549
rect 8054 23392 8134 23404
rect 8054 23336 8066 23392
rect 8122 23336 8134 23392
rect 8054 23324 8134 23336
rect 8872 23392 8952 23404
rect 8872 23336 8884 23392
rect 8940 23336 8952 23392
rect 8872 23324 8952 23336
rect 9225 23274 9305 23284
rect 7891 23218 9237 23274
rect 9293 23218 9305 23274
rect 9225 23216 9305 23218
rect 9059 23165 9129 23167
rect 7891 23164 9129 23165
rect 7891 23110 9061 23164
rect 9117 23110 9129 23164
rect 7891 23109 9129 23110
rect 5999 23057 6085 23061
rect 5999 23001 6011 23057
rect 6067 23001 6085 23057
rect 5999 22989 6085 23001
rect 5510 22844 5556 22855
rect 5725 22853 5801 22886
rect 5725 22807 5736 22853
rect 5790 22807 5801 22853
rect 5909 22853 5985 22886
rect 5909 22807 5920 22853
rect 5974 22807 5985 22853
rect 6093 22853 6169 22886
rect 6093 22807 6104 22853
rect 6158 22807 6169 22853
rect 6338 22844 6384 22855
rect 5648 22761 5694 22772
rect 5631 22734 5648 22736
rect 5832 22761 5878 22772
rect 5694 22734 5711 22736
rect 5556 22614 5643 22734
rect 5699 22614 5711 22734
rect 5631 22612 5648 22614
rect 5556 22314 5648 22434
rect 5694 22612 5711 22614
rect 5815 22434 5832 22436
rect 6016 22761 6062 22772
rect 5999 22734 6016 22736
rect 6200 22761 6246 22772
rect 6062 22734 6079 22736
rect 5999 22614 6011 22734
rect 6067 22614 6079 22734
rect 5999 22612 6016 22614
rect 5878 22434 5895 22436
rect 5815 22314 5827 22434
rect 5883 22314 5895 22434
rect 5815 22312 5832 22314
rect 5648 22276 5694 22287
rect 5878 22312 5895 22314
rect 5832 22276 5878 22287
rect 6062 22612 6079 22614
rect 6183 22434 6200 22436
rect 6321 22734 6338 22736
rect 6384 22734 6401 22736
rect 6321 22613 6333 22734
rect 6389 22613 6401 22734
rect 6321 22611 6338 22613
rect 6246 22434 6263 22436
rect 6183 22314 6195 22434
rect 6251 22314 6263 22434
rect 6183 22312 6200 22314
rect 6016 22276 6062 22287
rect 6246 22312 6263 22314
rect 6200 22276 6246 22287
rect 5725 22238 5736 22241
rect 5790 22238 5801 22241
rect 5909 22238 5920 22241
rect 5974 22238 5985 22241
rect 6093 22238 6104 22241
rect 6158 22238 6169 22241
rect 5510 22193 5556 22204
rect 5723 22182 5735 22238
rect 5791 22182 5803 22238
rect 5723 22168 5803 22182
rect 5907 22182 5919 22238
rect 5975 22182 5987 22238
rect 5907 22168 5987 22182
rect 6091 22182 6103 22238
rect 6159 22182 6171 22238
rect 6384 22611 6401 22613
rect 6338 22193 6384 22204
rect 6091 22168 6171 22182
rect 5723 22088 5803 22090
rect 5335 22032 5735 22088
rect 5791 22032 5803 22088
rect 7891 22088 7947 23109
rect 9059 23101 9129 23109
rect 8555 23057 8641 23061
rect 8555 23001 8567 23057
rect 8623 23001 8641 23057
rect 8555 22989 8641 23001
rect 8066 22844 8112 22855
rect 8281 22853 8357 22886
rect 8281 22807 8292 22853
rect 8346 22807 8357 22853
rect 8465 22853 8541 22886
rect 8465 22807 8476 22853
rect 8530 22807 8541 22853
rect 8649 22853 8725 22886
rect 8649 22807 8660 22853
rect 8714 22807 8725 22853
rect 8894 22844 8940 22855
rect 8204 22761 8250 22772
rect 8187 22734 8204 22736
rect 8388 22761 8434 22772
rect 8250 22734 8267 22736
rect 8112 22614 8199 22734
rect 8255 22614 8267 22734
rect 8187 22612 8204 22614
rect 8112 22314 8204 22434
rect 8250 22612 8267 22614
rect 8371 22434 8388 22436
rect 8572 22761 8618 22772
rect 8555 22734 8572 22736
rect 8756 22761 8802 22772
rect 8618 22734 8635 22736
rect 8555 22614 8567 22734
rect 8623 22614 8635 22734
rect 8555 22612 8572 22614
rect 8434 22434 8451 22436
rect 8371 22314 8383 22434
rect 8439 22314 8451 22434
rect 8371 22312 8388 22314
rect 8204 22276 8250 22287
rect 8434 22312 8451 22314
rect 8388 22276 8434 22287
rect 8618 22612 8635 22614
rect 8739 22434 8756 22436
rect 8877 22734 8894 22736
rect 8940 22734 8957 22736
rect 8877 22613 8889 22734
rect 8945 22613 8957 22734
rect 8877 22611 8894 22613
rect 8802 22434 8819 22436
rect 8739 22314 8751 22434
rect 8807 22314 8819 22434
rect 8739 22312 8756 22314
rect 8572 22276 8618 22287
rect 8802 22312 8819 22314
rect 8756 22276 8802 22287
rect 8281 22238 8292 22241
rect 8346 22238 8357 22241
rect 8465 22238 8476 22241
rect 8530 22238 8541 22241
rect 8649 22238 8660 22241
rect 8714 22238 8725 22241
rect 8066 22193 8112 22204
rect 8279 22182 8291 22238
rect 8347 22182 8359 22238
rect 8279 22168 8359 22182
rect 8463 22182 8475 22238
rect 8531 22182 8543 22238
rect 8463 22168 8543 22182
rect 8647 22182 8659 22238
rect 8715 22182 8727 22238
rect 8940 22611 8957 22613
rect 8894 22193 8940 22204
rect 8647 22168 8727 22182
rect 8279 22088 8359 22090
rect 7891 22032 8291 22088
rect 8347 22032 8359 22088
rect 9377 22088 9433 25314
rect 11928 25314 13475 25370
rect 10939 24293 11009 24305
rect 11928 24293 11984 25314
rect 12597 25262 12683 25266
rect 12597 25206 12609 25262
rect 12665 25206 12683 25262
rect 12597 25194 12683 25206
rect 12108 25049 12154 25060
rect 12323 25058 12399 25091
rect 12323 25012 12334 25058
rect 12388 25012 12399 25058
rect 12507 25058 12583 25091
rect 12507 25012 12518 25058
rect 12572 25012 12583 25058
rect 12691 25058 12767 25091
rect 12691 25012 12702 25058
rect 12756 25012 12767 25058
rect 12936 25049 12982 25060
rect 12246 24966 12292 24977
rect 12229 24939 12246 24941
rect 12430 24966 12476 24977
rect 12292 24939 12309 24941
rect 12154 24819 12241 24939
rect 12297 24819 12309 24939
rect 12229 24817 12246 24819
rect 12154 24519 12246 24639
rect 12292 24817 12309 24819
rect 12413 24639 12430 24641
rect 12614 24966 12660 24977
rect 12597 24939 12614 24941
rect 12798 24966 12844 24977
rect 12660 24939 12677 24941
rect 12597 24819 12609 24939
rect 12665 24819 12677 24939
rect 12597 24817 12614 24819
rect 12476 24639 12493 24641
rect 12413 24519 12425 24639
rect 12481 24519 12493 24639
rect 12413 24517 12430 24519
rect 12246 24481 12292 24492
rect 12476 24517 12493 24519
rect 12430 24481 12476 24492
rect 12660 24817 12677 24819
rect 12781 24639 12798 24641
rect 12919 24939 12936 24941
rect 12982 24939 12999 24941
rect 12919 24818 12931 24939
rect 12987 24818 12999 24939
rect 12919 24816 12936 24818
rect 12844 24639 12861 24641
rect 12781 24519 12793 24639
rect 12849 24519 12861 24639
rect 12781 24517 12798 24519
rect 12614 24481 12660 24492
rect 12844 24517 12861 24519
rect 12798 24481 12844 24492
rect 12323 24443 12334 24446
rect 12388 24443 12399 24446
rect 12507 24443 12518 24446
rect 12572 24443 12583 24446
rect 12691 24443 12702 24446
rect 12756 24443 12767 24446
rect 12108 24398 12154 24409
rect 12321 24387 12333 24443
rect 12389 24387 12401 24443
rect 12321 24373 12401 24387
rect 12505 24387 12517 24443
rect 12573 24387 12585 24443
rect 12505 24373 12585 24387
rect 12689 24387 12701 24443
rect 12757 24387 12769 24443
rect 12982 24816 12999 24818
rect 12936 24398 12982 24409
rect 12689 24373 12769 24387
rect 12321 24293 12401 24295
rect 10939 24237 10951 24293
rect 11007 24237 12333 24293
rect 12389 24237 12401 24293
rect 10939 24235 11009 24237
rect 12321 24235 12401 24237
rect 11649 24177 11719 24189
rect 12505 24177 12585 24179
rect 11649 24121 11661 24177
rect 11717 24121 12517 24177
rect 12573 24121 12585 24177
rect 11649 24109 11719 24121
rect 12505 24119 12585 24121
rect 12834 24177 12914 24179
rect 13101 24177 13171 24189
rect 12834 24121 12846 24177
rect 12902 24121 13103 24177
rect 13159 24121 13171 24177
rect 12834 24119 12914 24121
rect 13101 24111 13171 24121
rect 12689 24061 12769 24063
rect 11933 24005 12701 24061
rect 12757 24005 12769 24061
rect 11933 23274 11989 24005
rect 12689 24003 12769 24005
rect 12321 23911 12401 23925
rect 12108 23889 12154 23900
rect 12321 23855 12333 23911
rect 12389 23855 12401 23911
rect 12505 23911 12585 23925
rect 12505 23855 12517 23911
rect 12573 23855 12585 23911
rect 12689 23911 12769 23925
rect 12689 23855 12701 23911
rect 12757 23855 12769 23911
rect 12936 23889 12982 23900
rect 12323 23852 12334 23855
rect 12388 23852 12399 23855
rect 12507 23852 12518 23855
rect 12572 23852 12583 23855
rect 12691 23852 12702 23855
rect 12756 23852 12767 23855
rect 12246 23806 12292 23817
rect 12154 23632 12246 23806
rect 12246 23621 12292 23632
rect 12430 23806 12476 23817
rect 12430 23621 12476 23632
rect 12614 23806 12660 23817
rect 12798 23806 12844 23817
rect 12781 23779 12798 23781
rect 12844 23779 12861 23781
rect 12781 23659 12793 23779
rect 12849 23659 12861 23779
rect 12781 23657 12798 23659
rect 12614 23621 12660 23632
rect 12844 23657 12861 23659
rect 12798 23621 12844 23632
rect 12108 23404 12154 23549
rect 12323 23540 12334 23586
rect 12388 23540 12399 23586
rect 12323 23507 12399 23540
rect 12507 23540 12518 23586
rect 12572 23540 12583 23586
rect 12507 23507 12583 23540
rect 12691 23540 12702 23586
rect 12756 23540 12767 23586
rect 12691 23507 12767 23540
rect 12936 23404 12982 23549
rect 12096 23392 12176 23404
rect 12096 23336 12108 23392
rect 12164 23336 12176 23392
rect 12096 23324 12176 23336
rect 12914 23392 12994 23404
rect 12914 23336 12926 23392
rect 12982 23336 12994 23392
rect 12914 23324 12994 23336
rect 13267 23274 13347 23284
rect 11933 23218 13279 23274
rect 13335 23218 13347 23274
rect 13267 23216 13347 23218
rect 13101 23165 13171 23167
rect 11933 23164 13171 23165
rect 11933 23110 13103 23164
rect 13159 23110 13171 23164
rect 11933 23109 13171 23110
rect 10041 23057 10127 23061
rect 10041 23001 10053 23057
rect 10109 23001 10127 23057
rect 10041 22989 10127 23001
rect 9552 22844 9598 22855
rect 9767 22853 9843 22886
rect 9767 22807 9778 22853
rect 9832 22807 9843 22853
rect 9951 22853 10027 22886
rect 9951 22807 9962 22853
rect 10016 22807 10027 22853
rect 10135 22853 10211 22886
rect 10135 22807 10146 22853
rect 10200 22807 10211 22853
rect 10380 22844 10426 22855
rect 9690 22761 9736 22772
rect 9673 22734 9690 22736
rect 9874 22761 9920 22772
rect 9736 22734 9753 22736
rect 9598 22614 9685 22734
rect 9741 22614 9753 22734
rect 9673 22612 9690 22614
rect 9598 22314 9690 22434
rect 9736 22612 9753 22614
rect 9857 22434 9874 22436
rect 10058 22761 10104 22772
rect 10041 22734 10058 22736
rect 10242 22761 10288 22772
rect 10104 22734 10121 22736
rect 10041 22614 10053 22734
rect 10109 22614 10121 22734
rect 10041 22612 10058 22614
rect 9920 22434 9937 22436
rect 9857 22314 9869 22434
rect 9925 22314 9937 22434
rect 9857 22312 9874 22314
rect 9690 22276 9736 22287
rect 9920 22312 9937 22314
rect 9874 22276 9920 22287
rect 10104 22612 10121 22614
rect 10225 22434 10242 22436
rect 10363 22734 10380 22736
rect 10426 22734 10443 22736
rect 10363 22613 10375 22734
rect 10431 22613 10443 22734
rect 10363 22611 10380 22613
rect 10288 22434 10305 22436
rect 10225 22314 10237 22434
rect 10293 22314 10305 22434
rect 10225 22312 10242 22314
rect 10058 22276 10104 22287
rect 10288 22312 10305 22314
rect 10242 22276 10288 22287
rect 9767 22238 9778 22241
rect 9832 22238 9843 22241
rect 9951 22238 9962 22241
rect 10016 22238 10027 22241
rect 10135 22238 10146 22241
rect 10200 22238 10211 22241
rect 9552 22193 9598 22204
rect 9765 22182 9777 22238
rect 9833 22182 9845 22238
rect 9765 22168 9845 22182
rect 9949 22182 9961 22238
rect 10017 22182 10029 22238
rect 9949 22168 10029 22182
rect 10133 22182 10145 22238
rect 10201 22182 10213 22238
rect 10426 22611 10443 22613
rect 10380 22193 10426 22204
rect 10133 22168 10213 22182
rect 9765 22088 9845 22090
rect 9377 22032 9777 22088
rect 9833 22032 9845 22088
rect 11933 22088 11989 23109
rect 13101 23101 13171 23109
rect 12597 23057 12683 23061
rect 12597 23001 12609 23057
rect 12665 23001 12683 23057
rect 12597 22989 12683 23001
rect 12108 22844 12154 22855
rect 12323 22853 12399 22886
rect 12323 22807 12334 22853
rect 12388 22807 12399 22853
rect 12507 22853 12583 22886
rect 12507 22807 12518 22853
rect 12572 22807 12583 22853
rect 12691 22853 12767 22886
rect 12691 22807 12702 22853
rect 12756 22807 12767 22853
rect 12936 22844 12982 22855
rect 12246 22761 12292 22772
rect 12229 22734 12246 22736
rect 12430 22761 12476 22772
rect 12292 22734 12309 22736
rect 12154 22614 12241 22734
rect 12297 22614 12309 22734
rect 12229 22612 12246 22614
rect 12154 22314 12246 22434
rect 12292 22612 12309 22614
rect 12413 22434 12430 22436
rect 12614 22761 12660 22772
rect 12597 22734 12614 22736
rect 12798 22761 12844 22772
rect 12660 22734 12677 22736
rect 12597 22614 12609 22734
rect 12665 22614 12677 22734
rect 12597 22612 12614 22614
rect 12476 22434 12493 22436
rect 12413 22314 12425 22434
rect 12481 22314 12493 22434
rect 12413 22312 12430 22314
rect 12246 22276 12292 22287
rect 12476 22312 12493 22314
rect 12430 22276 12476 22287
rect 12660 22612 12677 22614
rect 12781 22434 12798 22436
rect 12919 22734 12936 22736
rect 12982 22734 12999 22736
rect 12919 22613 12931 22734
rect 12987 22613 12999 22734
rect 12919 22611 12936 22613
rect 12844 22434 12861 22436
rect 12781 22314 12793 22434
rect 12849 22314 12861 22434
rect 12781 22312 12798 22314
rect 12614 22276 12660 22287
rect 12844 22312 12861 22314
rect 12798 22276 12844 22287
rect 12323 22238 12334 22241
rect 12388 22238 12399 22241
rect 12507 22238 12518 22241
rect 12572 22238 12583 22241
rect 12691 22238 12702 22241
rect 12756 22238 12767 22241
rect 12108 22193 12154 22204
rect 12321 22182 12333 22238
rect 12389 22182 12401 22238
rect 12321 22168 12401 22182
rect 12505 22182 12517 22238
rect 12573 22182 12585 22238
rect 12505 22168 12585 22182
rect 12689 22182 12701 22238
rect 12757 22182 12769 22238
rect 12982 22611 12999 22613
rect 12936 22193 12982 22204
rect 12689 22168 12769 22182
rect 12321 22088 12401 22090
rect 11933 22032 12333 22088
rect 12389 22032 12401 22088
rect 13419 22088 13475 25314
rect 15970 25314 17517 25370
rect 14981 24293 15061 24305
rect 15970 24293 16026 25314
rect 16639 25262 16725 25266
rect 16639 25206 16651 25262
rect 16707 25206 16725 25262
rect 16639 25194 16725 25206
rect 16150 25049 16196 25060
rect 16365 25058 16441 25091
rect 16365 25012 16376 25058
rect 16430 25012 16441 25058
rect 16549 25058 16625 25091
rect 16549 25012 16560 25058
rect 16614 25012 16625 25058
rect 16733 25058 16809 25091
rect 16733 25012 16744 25058
rect 16798 25012 16809 25058
rect 16978 25049 17024 25060
rect 16288 24966 16334 24977
rect 16271 24939 16288 24941
rect 16472 24966 16518 24977
rect 16334 24939 16351 24941
rect 16196 24819 16283 24939
rect 16339 24819 16351 24939
rect 16271 24817 16288 24819
rect 16196 24519 16288 24639
rect 16334 24817 16351 24819
rect 16455 24639 16472 24641
rect 16656 24966 16702 24977
rect 16639 24939 16656 24941
rect 16840 24966 16886 24977
rect 16702 24939 16719 24941
rect 16639 24819 16651 24939
rect 16707 24819 16719 24939
rect 16639 24817 16656 24819
rect 16518 24639 16535 24641
rect 16455 24519 16467 24639
rect 16523 24519 16535 24639
rect 16455 24517 16472 24519
rect 16288 24481 16334 24492
rect 16518 24517 16535 24519
rect 16472 24481 16518 24492
rect 16702 24817 16719 24819
rect 16823 24639 16840 24641
rect 16961 24939 16978 24941
rect 17024 24939 17041 24941
rect 16961 24818 16973 24939
rect 17029 24818 17041 24939
rect 16961 24816 16978 24818
rect 16886 24639 16903 24641
rect 16823 24519 16835 24639
rect 16891 24519 16903 24639
rect 16823 24517 16840 24519
rect 16656 24481 16702 24492
rect 16886 24517 16903 24519
rect 16840 24481 16886 24492
rect 16365 24443 16376 24446
rect 16430 24443 16441 24446
rect 16549 24443 16560 24446
rect 16614 24443 16625 24446
rect 16733 24443 16744 24446
rect 16798 24443 16809 24446
rect 16150 24398 16196 24409
rect 16363 24387 16375 24443
rect 16431 24387 16443 24443
rect 16363 24373 16443 24387
rect 16547 24387 16559 24443
rect 16615 24387 16627 24443
rect 16547 24373 16627 24387
rect 16731 24387 16743 24443
rect 16799 24387 16811 24443
rect 17024 24816 17041 24818
rect 16978 24398 17024 24409
rect 16731 24373 16811 24387
rect 16363 24293 16443 24295
rect 14981 24237 14993 24293
rect 15049 24237 16375 24293
rect 16431 24237 16443 24293
rect 14981 24235 15061 24237
rect 16363 24235 16443 24237
rect 15691 24177 15761 24189
rect 16547 24177 16627 24179
rect 15691 24121 15703 24177
rect 15759 24121 16559 24177
rect 16615 24121 16627 24177
rect 15691 24109 15761 24121
rect 16547 24119 16627 24121
rect 16876 24177 16956 24179
rect 17143 24177 17213 24189
rect 16876 24121 16888 24177
rect 16944 24121 17145 24177
rect 17201 24121 17213 24177
rect 16876 24119 16956 24121
rect 17143 24111 17213 24121
rect 16731 24061 16811 24063
rect 15975 24005 16743 24061
rect 16799 24005 16811 24061
rect 15975 23274 16031 24005
rect 16731 24003 16811 24005
rect 16363 23911 16443 23925
rect 16150 23889 16196 23900
rect 16363 23855 16375 23911
rect 16431 23855 16443 23911
rect 16547 23911 16627 23925
rect 16547 23855 16559 23911
rect 16615 23855 16627 23911
rect 16731 23911 16811 23925
rect 16731 23855 16743 23911
rect 16799 23855 16811 23911
rect 16978 23889 17024 23900
rect 16365 23852 16376 23855
rect 16430 23852 16441 23855
rect 16549 23852 16560 23855
rect 16614 23852 16625 23855
rect 16733 23852 16744 23855
rect 16798 23852 16809 23855
rect 16288 23806 16334 23817
rect 16196 23632 16288 23806
rect 16288 23621 16334 23632
rect 16472 23806 16518 23817
rect 16472 23621 16518 23632
rect 16656 23806 16702 23817
rect 16840 23806 16886 23817
rect 16823 23779 16840 23781
rect 16886 23779 16903 23781
rect 16823 23659 16835 23779
rect 16891 23659 16903 23779
rect 16823 23657 16840 23659
rect 16656 23621 16702 23632
rect 16886 23657 16903 23659
rect 16840 23621 16886 23632
rect 16150 23404 16196 23549
rect 16365 23540 16376 23586
rect 16430 23540 16441 23586
rect 16365 23507 16441 23540
rect 16549 23540 16560 23586
rect 16614 23540 16625 23586
rect 16549 23507 16625 23540
rect 16733 23540 16744 23586
rect 16798 23540 16809 23586
rect 16733 23507 16809 23540
rect 16978 23404 17024 23549
rect 16138 23392 16218 23404
rect 16138 23336 16150 23392
rect 16206 23336 16218 23392
rect 16138 23324 16218 23336
rect 16956 23392 17036 23404
rect 16956 23336 16968 23392
rect 17024 23336 17036 23392
rect 16956 23324 17036 23336
rect 17309 23274 17389 23284
rect 15975 23218 17321 23274
rect 17377 23218 17389 23274
rect 17309 23216 17389 23218
rect 17143 23165 17213 23167
rect 15975 23164 17213 23165
rect 15975 23110 17145 23164
rect 17201 23110 17213 23164
rect 15975 23109 17213 23110
rect 14083 23057 14169 23061
rect 14083 23001 14095 23057
rect 14151 23001 14169 23057
rect 14083 22989 14169 23001
rect 13594 22844 13640 22855
rect 13809 22853 13885 22886
rect 13809 22807 13820 22853
rect 13874 22807 13885 22853
rect 13993 22853 14069 22886
rect 13993 22807 14004 22853
rect 14058 22807 14069 22853
rect 14177 22853 14253 22886
rect 14177 22807 14188 22853
rect 14242 22807 14253 22853
rect 14422 22844 14468 22855
rect 13732 22761 13778 22772
rect 13715 22734 13732 22736
rect 13916 22761 13962 22772
rect 13778 22734 13795 22736
rect 13640 22614 13727 22734
rect 13783 22614 13795 22734
rect 13715 22612 13732 22614
rect 13640 22314 13732 22434
rect 13778 22612 13795 22614
rect 13899 22434 13916 22436
rect 14100 22761 14146 22772
rect 14083 22734 14100 22736
rect 14284 22761 14330 22772
rect 14146 22734 14163 22736
rect 14083 22614 14095 22734
rect 14151 22614 14163 22734
rect 14083 22612 14100 22614
rect 13962 22434 13979 22436
rect 13899 22314 13911 22434
rect 13967 22314 13979 22434
rect 13899 22312 13916 22314
rect 13732 22276 13778 22287
rect 13962 22312 13979 22314
rect 13916 22276 13962 22287
rect 14146 22612 14163 22614
rect 14267 22434 14284 22436
rect 14405 22734 14422 22736
rect 14468 22734 14485 22736
rect 14405 22613 14417 22734
rect 14473 22613 14485 22734
rect 14405 22611 14422 22613
rect 14330 22434 14347 22436
rect 14267 22314 14279 22434
rect 14335 22314 14347 22434
rect 14267 22312 14284 22314
rect 14100 22276 14146 22287
rect 14330 22312 14347 22314
rect 14284 22276 14330 22287
rect 13809 22238 13820 22241
rect 13874 22238 13885 22241
rect 13993 22238 14004 22241
rect 14058 22238 14069 22241
rect 14177 22238 14188 22241
rect 14242 22238 14253 22241
rect 13594 22193 13640 22204
rect 13807 22182 13819 22238
rect 13875 22182 13887 22238
rect 13807 22168 13887 22182
rect 13991 22182 14003 22238
rect 14059 22182 14071 22238
rect 13991 22168 14071 22182
rect 14175 22182 14187 22238
rect 14243 22182 14255 22238
rect 14468 22611 14485 22613
rect 14422 22193 14468 22204
rect 14175 22168 14255 22182
rect 13807 22088 13887 22090
rect 13419 22032 13819 22088
rect 13875 22032 13887 22088
rect 15975 22088 16031 23109
rect 17143 23101 17213 23109
rect 16639 23057 16725 23061
rect 16639 23001 16651 23057
rect 16707 23001 16725 23057
rect 16639 22989 16725 23001
rect 16150 22844 16196 22855
rect 16365 22853 16441 22886
rect 16365 22807 16376 22853
rect 16430 22807 16441 22853
rect 16549 22853 16625 22886
rect 16549 22807 16560 22853
rect 16614 22807 16625 22853
rect 16733 22853 16809 22886
rect 16733 22807 16744 22853
rect 16798 22807 16809 22853
rect 16978 22844 17024 22855
rect 16288 22761 16334 22772
rect 16271 22734 16288 22736
rect 16472 22761 16518 22772
rect 16334 22734 16351 22736
rect 16196 22614 16283 22734
rect 16339 22614 16351 22734
rect 16271 22612 16288 22614
rect 16196 22314 16288 22434
rect 16334 22612 16351 22614
rect 16455 22434 16472 22436
rect 16656 22761 16702 22772
rect 16639 22734 16656 22736
rect 16840 22761 16886 22772
rect 16702 22734 16719 22736
rect 16639 22614 16651 22734
rect 16707 22614 16719 22734
rect 16639 22612 16656 22614
rect 16518 22434 16535 22436
rect 16455 22314 16467 22434
rect 16523 22314 16535 22434
rect 16455 22312 16472 22314
rect 16288 22276 16334 22287
rect 16518 22312 16535 22314
rect 16472 22276 16518 22287
rect 16702 22612 16719 22614
rect 16823 22434 16840 22436
rect 16961 22734 16978 22736
rect 17024 22734 17041 22736
rect 16961 22613 16973 22734
rect 17029 22613 17041 22734
rect 16961 22611 16978 22613
rect 16886 22434 16903 22436
rect 16823 22314 16835 22434
rect 16891 22314 16903 22434
rect 16823 22312 16840 22314
rect 16656 22276 16702 22287
rect 16886 22312 16903 22314
rect 16840 22276 16886 22287
rect 16365 22238 16376 22241
rect 16430 22238 16441 22241
rect 16549 22238 16560 22241
rect 16614 22238 16625 22241
rect 16733 22238 16744 22241
rect 16798 22238 16809 22241
rect 16150 22193 16196 22204
rect 16363 22182 16375 22238
rect 16431 22182 16443 22238
rect 16363 22168 16443 22182
rect 16547 22182 16559 22238
rect 16615 22182 16627 22238
rect 16547 22168 16627 22182
rect 16731 22182 16743 22238
rect 16799 22182 16811 22238
rect 17024 22611 17041 22613
rect 16978 22193 17024 22204
rect 16731 22168 16811 22182
rect 16363 22088 16443 22090
rect 15975 22032 16375 22088
rect 16431 22032 16443 22088
rect 17461 22088 17517 25314
rect 18125 23057 18211 23061
rect 18125 23001 18137 23057
rect 18193 23001 18211 23057
rect 18125 22989 18211 23001
rect 17636 22844 17682 22855
rect 17851 22853 17927 22886
rect 17851 22807 17862 22853
rect 17916 22807 17927 22853
rect 18035 22853 18111 22886
rect 18035 22807 18046 22853
rect 18100 22807 18111 22853
rect 18219 22853 18295 22886
rect 18219 22807 18230 22853
rect 18284 22807 18295 22853
rect 18464 22844 18510 22855
rect 17774 22761 17820 22772
rect 17757 22734 17774 22736
rect 17958 22761 18004 22772
rect 17820 22734 17837 22736
rect 17682 22614 17769 22734
rect 17825 22614 17837 22734
rect 17757 22612 17774 22614
rect 17682 22314 17774 22434
rect 17820 22612 17837 22614
rect 17941 22434 17958 22436
rect 18142 22761 18188 22772
rect 18125 22734 18142 22736
rect 18326 22761 18372 22772
rect 18188 22734 18205 22736
rect 18125 22614 18137 22734
rect 18193 22614 18205 22734
rect 18125 22612 18142 22614
rect 18004 22434 18021 22436
rect 17941 22314 17953 22434
rect 18009 22314 18021 22434
rect 17941 22312 17958 22314
rect 17774 22276 17820 22287
rect 18004 22312 18021 22314
rect 17958 22276 18004 22287
rect 18188 22612 18205 22614
rect 18309 22434 18326 22436
rect 18447 22734 18464 22736
rect 18510 22734 18527 22736
rect 18447 22613 18459 22734
rect 18515 22613 18527 22734
rect 18447 22611 18464 22613
rect 18372 22434 18389 22436
rect 18309 22314 18321 22434
rect 18377 22314 18389 22434
rect 18309 22312 18326 22314
rect 18142 22276 18188 22287
rect 18372 22312 18389 22314
rect 18326 22276 18372 22287
rect 17851 22238 17862 22241
rect 17916 22238 17927 22241
rect 18035 22238 18046 22241
rect 18100 22238 18111 22241
rect 18219 22238 18230 22241
rect 18284 22238 18295 22241
rect 17636 22193 17682 22204
rect 17849 22182 17861 22238
rect 17917 22182 17929 22238
rect 17849 22168 17929 22182
rect 18033 22182 18045 22238
rect 18101 22182 18113 22238
rect 18033 22168 18113 22182
rect 18217 22182 18229 22238
rect 18285 22182 18297 22238
rect 18510 22611 18527 22613
rect 18464 22193 18510 22204
rect 18217 22168 18297 22182
rect 17849 22088 17929 22090
rect 17461 22032 17861 22088
rect 17917 22032 17929 22088
rect -3847 22030 -3767 22032
rect -2361 22030 -2281 22032
rect 195 22030 275 22032
rect 1681 22030 1761 22032
rect 4237 22030 4317 22032
rect 5723 22030 5803 22032
rect 8279 22030 8359 22032
rect 9765 22030 9845 22032
rect 12321 22030 12401 22032
rect 13807 22030 13887 22032
rect 16363 22030 16443 22032
rect 17849 22030 17929 22032
rect -8697 21975 -8627 21989
rect -7705 21975 -7625 21977
rect -8697 21919 -8685 21975
rect -8629 21919 -7693 21975
rect -7637 21919 -7625 21975
rect -8697 21907 -8627 21919
rect -7705 21917 -7625 21919
rect -7376 21975 -7296 21977
rect -6933 21975 -6873 21985
rect -6219 21975 -6139 21977
rect -7376 21919 -7364 21975
rect -7308 21919 -6931 21975
rect -6875 21919 -6207 21975
rect -6151 21919 -6139 21975
rect -7376 21917 -7296 21919
rect -6933 21907 -6873 21919
rect -6219 21917 -6139 21919
rect -5890 21975 -5810 21977
rect -5623 21975 -5553 21987
rect -5083 21975 -5013 21977
rect -5890 21919 -5878 21975
rect -5822 21919 -5621 21975
rect -5565 21919 -5081 21975
rect -5025 21919 -5013 21975
rect -5890 21917 -5810 21919
rect -5623 21909 -5553 21919
rect -5083 21907 -5013 21919
rect -4655 21972 -4585 21986
rect -3663 21972 -3583 21974
rect -4655 21916 -4643 21972
rect -4587 21916 -3651 21972
rect -3595 21916 -3583 21972
rect -4655 21904 -4585 21916
rect -3663 21914 -3583 21916
rect -3334 21972 -3254 21974
rect -2891 21972 -2831 21982
rect -2177 21972 -2097 21974
rect -3334 21916 -3322 21972
rect -3266 21916 -2889 21972
rect -2833 21916 -2165 21972
rect -2109 21916 -2097 21972
rect -3334 21914 -3254 21916
rect -2891 21904 -2831 21916
rect -2177 21914 -2097 21916
rect -1848 21972 -1768 21974
rect -1581 21972 -1511 21984
rect -1029 21972 -959 21984
rect -1848 21916 -1836 21972
rect -1780 21916 -1579 21972
rect -1523 21916 -1027 21972
rect -971 21916 -959 21972
rect -1848 21914 -1768 21916
rect -1581 21906 -1511 21916
rect -1029 21904 -959 21916
rect -613 21972 -543 21986
rect 379 21972 459 21974
rect -613 21916 -601 21972
rect -545 21916 391 21972
rect 447 21916 459 21972
rect -613 21904 -543 21916
rect 379 21914 459 21916
rect 708 21972 788 21974
rect 1151 21972 1211 21982
rect 1865 21972 1945 21974
rect 708 21916 720 21972
rect 776 21916 1153 21972
rect 1209 21916 1877 21972
rect 1933 21916 1945 21972
rect 708 21914 788 21916
rect 1151 21904 1211 21916
rect 1865 21914 1945 21916
rect 2194 21972 2274 21974
rect 2461 21972 2531 21984
rect 3067 21972 3137 21984
rect 2194 21916 2206 21972
rect 2262 21916 2463 21972
rect 2519 21916 3069 21972
rect 3125 21916 3137 21972
rect 2194 21914 2274 21916
rect 2461 21906 2531 21916
rect 3067 21904 3137 21916
rect 3429 21972 3499 21986
rect 4421 21972 4501 21974
rect 3429 21916 3441 21972
rect 3497 21916 4433 21972
rect 4489 21916 4501 21972
rect 3429 21904 3499 21916
rect 4421 21914 4501 21916
rect 4750 21972 4830 21974
rect 5193 21972 5253 21982
rect 5907 21972 5987 21974
rect 4750 21916 4762 21972
rect 4818 21916 5195 21972
rect 5251 21916 5919 21972
rect 5975 21916 5987 21972
rect 4750 21914 4830 21916
rect 5193 21904 5253 21916
rect 5907 21914 5987 21916
rect 6236 21972 6316 21974
rect 6503 21972 6573 21984
rect 7109 21972 7179 21984
rect 6236 21916 6248 21972
rect 6304 21916 6505 21972
rect 6561 21916 7111 21972
rect 7167 21916 7179 21972
rect 6236 21914 6316 21916
rect 6503 21906 6573 21916
rect 7109 21904 7179 21916
rect 7471 21972 7541 21986
rect 8463 21972 8543 21974
rect 7471 21916 7483 21972
rect 7539 21916 8475 21972
rect 8531 21916 8543 21972
rect 7471 21904 7541 21916
rect 8463 21914 8543 21916
rect 8792 21972 8872 21974
rect 9235 21972 9295 21982
rect 9949 21972 10029 21974
rect 8792 21916 8804 21972
rect 8860 21916 9237 21972
rect 9293 21916 9961 21972
rect 10017 21916 10029 21972
rect 8792 21914 8872 21916
rect 9235 21904 9295 21916
rect 9949 21914 10029 21916
rect 10278 21972 10358 21974
rect 10545 21972 10615 21984
rect 11151 21972 11221 21984
rect 10278 21916 10290 21972
rect 10346 21916 10547 21972
rect 10603 21916 11153 21972
rect 11209 21916 11221 21972
rect 10278 21914 10358 21916
rect 10545 21906 10615 21916
rect 11151 21904 11221 21916
rect 11513 21972 11583 21986
rect 12505 21972 12585 21974
rect 11513 21916 11525 21972
rect 11581 21916 12517 21972
rect 12573 21916 12585 21972
rect 11513 21904 11583 21916
rect 12505 21914 12585 21916
rect 12834 21972 12914 21974
rect 13277 21972 13337 21982
rect 13991 21972 14071 21974
rect 12834 21916 12846 21972
rect 12902 21916 13279 21972
rect 13335 21916 14003 21972
rect 14059 21916 14071 21972
rect 12834 21914 12914 21916
rect 13277 21904 13337 21916
rect 13991 21914 14071 21916
rect 14320 21972 14400 21974
rect 14587 21972 14657 21984
rect 15193 21972 15263 21984
rect 14320 21916 14332 21972
rect 14388 21916 14589 21972
rect 14645 21916 15195 21972
rect 15251 21916 15263 21972
rect 14320 21914 14400 21916
rect 14587 21906 14657 21916
rect 15193 21904 15263 21916
rect 15555 21972 15625 21986
rect 16547 21972 16627 21974
rect 15555 21916 15567 21972
rect 15623 21916 16559 21972
rect 16615 21916 16627 21972
rect 15555 21904 15625 21916
rect 16547 21914 16627 21916
rect 16876 21972 16956 21974
rect 17319 21972 17379 21982
rect 18033 21972 18113 21974
rect 16876 21916 16888 21972
rect 16944 21916 17321 21972
rect 17377 21916 18045 21972
rect 18101 21916 18113 21972
rect 16876 21914 16956 21916
rect 17319 21904 17379 21916
rect 18033 21914 18113 21916
rect 18362 21972 18442 21974
rect 18629 21972 18699 21984
rect 19235 21972 19305 21984
rect 18362 21916 18374 21972
rect 18430 21916 18631 21972
rect 18687 21916 19237 21972
rect 19293 21916 19305 21972
rect 18362 21914 18442 21916
rect 18629 21906 18699 21916
rect 19235 21904 19305 21916
rect -7521 21859 -7441 21861
rect -6035 21859 -5955 21861
rect -8413 21803 -7509 21859
rect -7453 21803 -7441 21859
rect -8887 21073 -8817 21075
rect -8413 21073 -8357 21803
rect -7521 21801 -7441 21803
rect -6791 21803 -6023 21859
rect -5967 21803 -5955 21859
rect -3479 21856 -3399 21858
rect -1993 21856 -1913 21858
rect 563 21856 643 21858
rect 2049 21856 2129 21858
rect 4605 21856 4685 21858
rect 6091 21856 6171 21858
rect 8647 21856 8727 21858
rect 10133 21856 10213 21858
rect 12689 21856 12769 21858
rect 14175 21856 14255 21858
rect 16731 21856 16811 21858
rect 18217 21856 18297 21858
rect -7889 21709 -7809 21723
rect -8102 21687 -8056 21698
rect -7889 21653 -7877 21709
rect -7821 21653 -7809 21709
rect -7705 21709 -7625 21723
rect -7705 21653 -7693 21709
rect -7637 21653 -7625 21709
rect -7521 21709 -7441 21723
rect -7521 21653 -7509 21709
rect -7453 21653 -7441 21709
rect -7274 21687 -7228 21698
rect -7887 21650 -7876 21653
rect -7822 21650 -7811 21653
rect -7703 21650 -7692 21653
rect -7638 21650 -7627 21653
rect -7519 21650 -7508 21653
rect -7454 21650 -7443 21653
rect -7964 21604 -7918 21615
rect -8056 21430 -7964 21604
rect -7964 21419 -7918 21430
rect -7780 21604 -7734 21615
rect -7780 21419 -7734 21430
rect -7596 21604 -7550 21615
rect -7412 21604 -7366 21615
rect -7429 21577 -7412 21579
rect -7366 21577 -7349 21579
rect -7429 21457 -7417 21577
rect -7361 21457 -7349 21577
rect -7429 21455 -7412 21457
rect -7596 21419 -7550 21430
rect -7366 21455 -7349 21457
rect -7412 21419 -7366 21430
rect -8102 21202 -8056 21347
rect -7887 21338 -7876 21384
rect -7822 21338 -7811 21384
rect -7887 21305 -7811 21338
rect -7703 21338 -7692 21384
rect -7638 21338 -7627 21384
rect -7703 21305 -7627 21338
rect -7519 21338 -7508 21384
rect -7454 21338 -7443 21384
rect -7519 21305 -7443 21338
rect -7274 21202 -7228 21347
rect -8114 21190 -8034 21202
rect -8114 21134 -8102 21190
rect -8046 21134 -8034 21190
rect -8114 21122 -8034 21134
rect -7296 21190 -7218 21202
rect -7296 21134 -7284 21190
rect -7228 21134 -7218 21190
rect -7296 21122 -7218 21134
rect -8887 21017 -8875 21073
rect -8819 21017 -8357 21073
rect -6791 21073 -6735 21803
rect -6035 21801 -5955 21803
rect -4371 21800 -3467 21856
rect -3411 21800 -3399 21856
rect -6403 21709 -6323 21723
rect -6616 21687 -6570 21698
rect -6403 21653 -6391 21709
rect -6335 21653 -6323 21709
rect -6219 21709 -6139 21723
rect -6219 21653 -6207 21709
rect -6151 21653 -6139 21709
rect -6035 21709 -5955 21723
rect -6035 21653 -6023 21709
rect -5967 21653 -5955 21709
rect -5788 21687 -5742 21698
rect -6401 21650 -6390 21653
rect -6336 21650 -6325 21653
rect -6217 21650 -6206 21653
rect -6152 21650 -6141 21653
rect -6033 21650 -6022 21653
rect -5968 21650 -5957 21653
rect -6478 21604 -6432 21615
rect -6570 21430 -6478 21604
rect -6478 21419 -6432 21430
rect -6294 21604 -6248 21615
rect -6294 21419 -6248 21430
rect -6110 21604 -6064 21615
rect -5926 21604 -5880 21615
rect -5943 21577 -5926 21579
rect -5880 21577 -5863 21579
rect -5943 21457 -5931 21577
rect -5875 21457 -5863 21577
rect -5943 21455 -5926 21457
rect -6110 21419 -6064 21430
rect -5880 21455 -5863 21457
rect -5926 21419 -5880 21430
rect -6616 21202 -6570 21347
rect -6401 21338 -6390 21384
rect -6336 21338 -6325 21384
rect -6401 21305 -6325 21338
rect -6217 21338 -6206 21384
rect -6152 21338 -6141 21384
rect -6217 21305 -6141 21338
rect -6033 21338 -6022 21384
rect -5968 21338 -5957 21384
rect -6033 21305 -5957 21338
rect -5788 21202 -5742 21347
rect -6628 21190 -6548 21202
rect -6628 21134 -6616 21190
rect -6560 21134 -6548 21190
rect -6628 21122 -6548 21134
rect -5810 21190 -5732 21202
rect -5810 21134 -5798 21190
rect -5742 21134 -5732 21190
rect -5810 21122 -5732 21134
rect -5457 21073 -5377 21083
rect -6791 21017 -5445 21073
rect -5389 21017 -5377 21073
rect -8887 21005 -8817 21017
rect -8413 19770 -8357 21017
rect -5457 21015 -5377 21017
rect -4791 21070 -4721 21072
rect -4371 21070 -4315 21800
rect -3479 21798 -3399 21800
rect -2749 21800 -1981 21856
rect -1925 21800 -1913 21856
rect -3847 21706 -3767 21720
rect -4060 21684 -4014 21695
rect -3847 21650 -3835 21706
rect -3779 21650 -3767 21706
rect -3663 21706 -3583 21720
rect -3663 21650 -3651 21706
rect -3595 21650 -3583 21706
rect -3479 21706 -3399 21720
rect -3479 21650 -3467 21706
rect -3411 21650 -3399 21706
rect -3232 21684 -3186 21695
rect -3845 21647 -3834 21650
rect -3780 21647 -3769 21650
rect -3661 21647 -3650 21650
rect -3596 21647 -3585 21650
rect -3477 21647 -3466 21650
rect -3412 21647 -3401 21650
rect -3922 21601 -3876 21612
rect -4014 21427 -3922 21601
rect -3922 21416 -3876 21427
rect -3738 21601 -3692 21612
rect -3738 21416 -3692 21427
rect -3554 21601 -3508 21612
rect -3370 21601 -3324 21612
rect -3387 21574 -3370 21576
rect -3324 21574 -3307 21576
rect -3387 21454 -3375 21574
rect -3319 21454 -3307 21574
rect -3387 21452 -3370 21454
rect -3554 21416 -3508 21427
rect -3324 21452 -3307 21454
rect -3370 21416 -3324 21427
rect -4060 21199 -4014 21344
rect -3845 21335 -3834 21381
rect -3780 21335 -3769 21381
rect -3845 21302 -3769 21335
rect -3661 21335 -3650 21381
rect -3596 21335 -3585 21381
rect -3661 21302 -3585 21335
rect -3477 21335 -3466 21381
rect -3412 21335 -3401 21381
rect -3477 21302 -3401 21335
rect -3232 21199 -3186 21344
rect -4072 21187 -3992 21199
rect -4072 21131 -4060 21187
rect -4004 21131 -3992 21187
rect -4072 21119 -3992 21131
rect -3254 21187 -3176 21199
rect -3254 21131 -3242 21187
rect -3186 21131 -3176 21187
rect -3254 21119 -3176 21131
rect -4791 21014 -4779 21070
rect -4723 21014 -4315 21070
rect -2749 21070 -2693 21800
rect -1993 21798 -1913 21800
rect -329 21800 575 21856
rect 631 21800 643 21856
rect -2361 21706 -2281 21720
rect -2574 21684 -2528 21695
rect -2361 21650 -2349 21706
rect -2293 21650 -2281 21706
rect -2177 21706 -2097 21720
rect -2177 21650 -2165 21706
rect -2109 21650 -2097 21706
rect -1993 21706 -1913 21720
rect -1993 21650 -1981 21706
rect -1925 21650 -1913 21706
rect -1746 21684 -1700 21695
rect -2359 21647 -2348 21650
rect -2294 21647 -2283 21650
rect -2175 21647 -2164 21650
rect -2110 21647 -2099 21650
rect -1991 21647 -1980 21650
rect -1926 21647 -1915 21650
rect -2436 21601 -2390 21612
rect -2528 21427 -2436 21601
rect -2436 21416 -2390 21427
rect -2252 21601 -2206 21612
rect -2252 21416 -2206 21427
rect -2068 21601 -2022 21612
rect -1884 21601 -1838 21612
rect -1901 21574 -1884 21576
rect -1838 21574 -1821 21576
rect -1901 21454 -1889 21574
rect -1833 21454 -1821 21574
rect -1901 21452 -1884 21454
rect -2068 21416 -2022 21427
rect -1838 21452 -1821 21454
rect -1884 21416 -1838 21427
rect -2574 21199 -2528 21344
rect -2359 21335 -2348 21381
rect -2294 21335 -2283 21381
rect -2359 21302 -2283 21335
rect -2175 21335 -2164 21381
rect -2110 21335 -2099 21381
rect -2175 21302 -2099 21335
rect -1991 21335 -1980 21381
rect -1926 21335 -1915 21381
rect -1991 21302 -1915 21335
rect -1746 21199 -1700 21344
rect -2586 21187 -2506 21199
rect -2586 21131 -2574 21187
rect -2518 21131 -2506 21187
rect -2586 21119 -2506 21131
rect -1768 21187 -1690 21199
rect -1768 21131 -1756 21187
rect -1700 21131 -1690 21187
rect -1768 21119 -1690 21131
rect -1415 21070 -1335 21080
rect -2749 21014 -1403 21070
rect -1347 21014 -1335 21070
rect -4791 21002 -4721 21014
rect -6933 20962 -6863 20964
rect -5633 20963 -5553 20965
rect -8277 20906 -6931 20962
rect -6875 20906 -6863 20962
rect -8277 19886 -8221 20906
rect -6933 20894 -6863 20906
rect -6791 20907 -5621 20963
rect -5565 20907 -5553 20963
rect -7613 20855 -7527 20859
rect -7613 20799 -7601 20855
rect -7545 20799 -7527 20855
rect -7613 20787 -7527 20799
rect -8102 20642 -8056 20653
rect -7887 20651 -7811 20684
rect -7887 20605 -7876 20651
rect -7822 20605 -7811 20651
rect -7703 20651 -7627 20684
rect -7703 20605 -7692 20651
rect -7638 20605 -7627 20651
rect -7519 20651 -7443 20684
rect -7519 20605 -7508 20651
rect -7454 20605 -7443 20651
rect -7274 20642 -7228 20653
rect -7964 20559 -7918 20570
rect -7981 20532 -7964 20534
rect -7780 20559 -7734 20570
rect -7918 20532 -7901 20534
rect -8056 20412 -7969 20532
rect -7913 20412 -7901 20532
rect -7981 20410 -7964 20412
rect -8056 20112 -7964 20232
rect -7918 20410 -7901 20412
rect -7797 20232 -7780 20234
rect -7596 20559 -7550 20570
rect -7613 20532 -7596 20534
rect -7412 20559 -7366 20570
rect -7550 20532 -7533 20534
rect -7613 20412 -7601 20532
rect -7545 20412 -7533 20532
rect -7613 20410 -7596 20412
rect -7734 20232 -7717 20234
rect -7797 20112 -7785 20232
rect -7729 20112 -7717 20232
rect -7797 20110 -7780 20112
rect -7964 20074 -7918 20085
rect -7734 20110 -7717 20112
rect -7780 20074 -7734 20085
rect -7550 20410 -7533 20412
rect -7429 20232 -7412 20234
rect -7291 20532 -7274 20534
rect -7228 20532 -7211 20534
rect -7291 20411 -7279 20532
rect -7223 20411 -7211 20532
rect -7291 20409 -7274 20411
rect -7366 20232 -7349 20234
rect -7429 20112 -7417 20232
rect -7361 20112 -7349 20232
rect -7429 20110 -7412 20112
rect -7596 20074 -7550 20085
rect -7366 20110 -7349 20112
rect -7412 20074 -7366 20085
rect -7887 20036 -7876 20039
rect -7822 20036 -7811 20039
rect -7703 20036 -7692 20039
rect -7638 20036 -7627 20039
rect -7519 20036 -7508 20039
rect -7454 20036 -7443 20039
rect -8102 19991 -8056 20002
rect -7889 19980 -7877 20036
rect -7821 19980 -7809 20036
rect -7889 19966 -7809 19980
rect -7705 19980 -7693 20036
rect -7637 19980 -7625 20036
rect -7705 19966 -7625 19980
rect -7521 19980 -7509 20036
rect -7453 19980 -7441 20036
rect -7228 20409 -7211 20411
rect -7274 19991 -7228 20002
rect -7521 19966 -7441 19980
rect -7889 19886 -7809 19888
rect -8277 19830 -7877 19886
rect -7821 19830 -7809 19886
rect -6791 19887 -6735 20907
rect -5633 20895 -5553 20907
rect -6127 20856 -6041 20860
rect -6127 20800 -6115 20856
rect -6059 20800 -6041 20856
rect -6127 20788 -6041 20800
rect -6616 20643 -6570 20654
rect -6401 20652 -6325 20685
rect -6401 20606 -6390 20652
rect -6336 20606 -6325 20652
rect -6217 20652 -6141 20685
rect -6217 20606 -6206 20652
rect -6152 20606 -6141 20652
rect -6033 20652 -5957 20685
rect -6033 20606 -6022 20652
rect -5968 20606 -5957 20652
rect -5788 20643 -5742 20654
rect -6478 20560 -6432 20571
rect -6495 20533 -6478 20535
rect -6294 20560 -6248 20571
rect -6432 20533 -6415 20535
rect -6570 20413 -6483 20533
rect -6427 20413 -6415 20533
rect -6495 20411 -6478 20413
rect -6570 20113 -6478 20233
rect -6432 20411 -6415 20413
rect -6311 20233 -6294 20235
rect -6110 20560 -6064 20571
rect -6127 20533 -6110 20535
rect -5926 20560 -5880 20571
rect -6064 20533 -6047 20535
rect -6127 20413 -6115 20533
rect -6059 20413 -6047 20533
rect -6127 20411 -6110 20413
rect -6248 20233 -6231 20235
rect -6311 20113 -6299 20233
rect -6243 20113 -6231 20233
rect -6311 20111 -6294 20113
rect -6478 20075 -6432 20086
rect -6248 20111 -6231 20113
rect -6294 20075 -6248 20086
rect -6064 20411 -6047 20413
rect -5943 20233 -5926 20235
rect -5805 20533 -5788 20535
rect -5742 20533 -5725 20535
rect -5805 20412 -5793 20533
rect -5737 20412 -5725 20533
rect -5805 20410 -5788 20412
rect -5880 20233 -5863 20235
rect -5943 20113 -5931 20233
rect -5875 20113 -5863 20233
rect -5943 20111 -5926 20113
rect -6110 20075 -6064 20086
rect -5880 20111 -5863 20113
rect -5926 20075 -5880 20086
rect -6401 20037 -6390 20040
rect -6336 20037 -6325 20040
rect -6217 20037 -6206 20040
rect -6152 20037 -6141 20040
rect -6033 20037 -6022 20040
rect -5968 20037 -5957 20040
rect -6616 19992 -6570 20003
rect -6403 19981 -6391 20037
rect -6335 19981 -6323 20037
rect -6403 19967 -6323 19981
rect -6219 19981 -6207 20037
rect -6151 19981 -6139 20037
rect -6219 19967 -6139 19981
rect -6035 19981 -6023 20037
rect -5967 19981 -5955 20037
rect -5742 20410 -5725 20412
rect -5788 19992 -5742 20003
rect -6035 19967 -5955 19981
rect -6403 19887 -6323 19889
rect -6791 19831 -6391 19887
rect -6335 19831 -6323 19887
rect -7889 19828 -7809 19830
rect -6403 19829 -6323 19831
rect -7705 19770 -7625 19772
rect -8413 19714 -7693 19770
rect -7637 19714 -7625 19770
rect -7705 19712 -7625 19714
rect -7376 19770 -7296 19772
rect -7109 19771 -7039 19782
rect -6219 19771 -6139 19773
rect -7109 19770 -6207 19771
rect -7376 19714 -7364 19770
rect -7308 19714 -7107 19770
rect -7051 19715 -6207 19770
rect -6151 19715 -6139 19771
rect -7051 19714 -6791 19715
rect -7376 19712 -7296 19714
rect -7109 19704 -7039 19714
rect -6219 19713 -6139 19715
rect -5890 19771 -5810 19773
rect -5447 19771 -5377 19781
rect -5890 19715 -5878 19771
rect -5822 19715 -5445 19771
rect -5389 19715 -5377 19771
rect -5890 19713 -5810 19715
rect -5447 19703 -5377 19715
rect -4371 19767 -4315 21014
rect -1415 21012 -1335 21014
rect -749 21070 -679 21072
rect -329 21070 -273 21800
rect 563 21798 643 21800
rect 1293 21800 2061 21856
rect 2117 21800 2129 21856
rect 195 21706 275 21720
rect -18 21684 28 21695
rect 195 21650 207 21706
rect 263 21650 275 21706
rect 379 21706 459 21720
rect 379 21650 391 21706
rect 447 21650 459 21706
rect 563 21706 643 21720
rect 563 21650 575 21706
rect 631 21650 643 21706
rect 810 21684 856 21695
rect 197 21647 208 21650
rect 262 21647 273 21650
rect 381 21647 392 21650
rect 446 21647 457 21650
rect 565 21647 576 21650
rect 630 21647 641 21650
rect 120 21601 166 21612
rect 28 21427 120 21601
rect 120 21416 166 21427
rect 304 21601 350 21612
rect 304 21416 350 21427
rect 488 21601 534 21612
rect 672 21601 718 21612
rect 655 21574 672 21576
rect 718 21574 735 21576
rect 655 21454 667 21574
rect 723 21454 735 21574
rect 655 21452 672 21454
rect 488 21416 534 21427
rect 718 21452 735 21454
rect 672 21416 718 21427
rect -18 21199 28 21344
rect 197 21335 208 21381
rect 262 21335 273 21381
rect 197 21302 273 21335
rect 381 21335 392 21381
rect 446 21335 457 21381
rect 381 21302 457 21335
rect 565 21335 576 21381
rect 630 21335 641 21381
rect 565 21302 641 21335
rect 810 21199 856 21344
rect -30 21187 50 21199
rect -30 21131 -18 21187
rect 38 21131 50 21187
rect -30 21119 50 21131
rect 788 21187 866 21199
rect 788 21131 800 21187
rect 856 21131 866 21187
rect 788 21119 866 21131
rect -749 21014 -737 21070
rect -681 21014 -273 21070
rect 1293 21070 1349 21800
rect 2049 21798 2129 21800
rect 3713 21800 4617 21856
rect 4673 21800 4685 21856
rect 1681 21706 1761 21720
rect 1468 21684 1514 21695
rect 1681 21650 1693 21706
rect 1749 21650 1761 21706
rect 1865 21706 1945 21720
rect 1865 21650 1877 21706
rect 1933 21650 1945 21706
rect 2049 21706 2129 21720
rect 2049 21650 2061 21706
rect 2117 21650 2129 21706
rect 2296 21684 2342 21695
rect 1683 21647 1694 21650
rect 1748 21647 1759 21650
rect 1867 21647 1878 21650
rect 1932 21647 1943 21650
rect 2051 21647 2062 21650
rect 2116 21647 2127 21650
rect 1606 21601 1652 21612
rect 1514 21427 1606 21601
rect 1606 21416 1652 21427
rect 1790 21601 1836 21612
rect 1790 21416 1836 21427
rect 1974 21601 2020 21612
rect 2158 21601 2204 21612
rect 2141 21574 2158 21576
rect 2204 21574 2221 21576
rect 2141 21454 2153 21574
rect 2209 21454 2221 21574
rect 2141 21452 2158 21454
rect 1974 21416 2020 21427
rect 2204 21452 2221 21454
rect 2158 21416 2204 21427
rect 1468 21199 1514 21344
rect 1683 21335 1694 21381
rect 1748 21335 1759 21381
rect 1683 21302 1759 21335
rect 1867 21335 1878 21381
rect 1932 21335 1943 21381
rect 1867 21302 1943 21335
rect 2051 21335 2062 21381
rect 2116 21335 2127 21381
rect 2051 21302 2127 21335
rect 2296 21199 2342 21344
rect 1456 21187 1536 21199
rect 1456 21131 1468 21187
rect 1524 21131 1536 21187
rect 1456 21119 1536 21131
rect 2274 21187 2352 21199
rect 2274 21131 2286 21187
rect 2342 21131 2352 21187
rect 2274 21119 2352 21131
rect 2627 21070 2707 21080
rect 1293 21014 2639 21070
rect 2695 21014 2707 21070
rect -749 21002 -679 21014
rect -2891 20959 -2821 20961
rect -1591 20960 -1511 20962
rect -4235 20903 -2889 20959
rect -2833 20903 -2821 20959
rect -4235 19883 -4179 20903
rect -2891 20891 -2821 20903
rect -2749 20904 -1579 20960
rect -1523 20904 -1511 20960
rect -3571 20852 -3485 20856
rect -3571 20796 -3559 20852
rect -3503 20796 -3485 20852
rect -3571 20784 -3485 20796
rect -4060 20639 -4014 20650
rect -3845 20648 -3769 20681
rect -3845 20602 -3834 20648
rect -3780 20602 -3769 20648
rect -3661 20648 -3585 20681
rect -3661 20602 -3650 20648
rect -3596 20602 -3585 20648
rect -3477 20648 -3401 20681
rect -3477 20602 -3466 20648
rect -3412 20602 -3401 20648
rect -3232 20639 -3186 20650
rect -3922 20556 -3876 20567
rect -3939 20529 -3922 20531
rect -3738 20556 -3692 20567
rect -3876 20529 -3859 20531
rect -4014 20409 -3927 20529
rect -3871 20409 -3859 20529
rect -3939 20407 -3922 20409
rect -4014 20109 -3922 20229
rect -3876 20407 -3859 20409
rect -3755 20229 -3738 20231
rect -3554 20556 -3508 20567
rect -3571 20529 -3554 20531
rect -3370 20556 -3324 20567
rect -3508 20529 -3491 20531
rect -3571 20409 -3559 20529
rect -3503 20409 -3491 20529
rect -3571 20407 -3554 20409
rect -3692 20229 -3675 20231
rect -3755 20109 -3743 20229
rect -3687 20109 -3675 20229
rect -3755 20107 -3738 20109
rect -3922 20071 -3876 20082
rect -3692 20107 -3675 20109
rect -3738 20071 -3692 20082
rect -3508 20407 -3491 20409
rect -3387 20229 -3370 20231
rect -3249 20529 -3232 20531
rect -3186 20529 -3169 20531
rect -3249 20408 -3237 20529
rect -3181 20408 -3169 20529
rect -3249 20406 -3232 20408
rect -3324 20229 -3307 20231
rect -3387 20109 -3375 20229
rect -3319 20109 -3307 20229
rect -3387 20107 -3370 20109
rect -3554 20071 -3508 20082
rect -3324 20107 -3307 20109
rect -3370 20071 -3324 20082
rect -3845 20033 -3834 20036
rect -3780 20033 -3769 20036
rect -3661 20033 -3650 20036
rect -3596 20033 -3585 20036
rect -3477 20033 -3466 20036
rect -3412 20033 -3401 20036
rect -4060 19988 -4014 19999
rect -3847 19977 -3835 20033
rect -3779 19977 -3767 20033
rect -3847 19963 -3767 19977
rect -3663 19977 -3651 20033
rect -3595 19977 -3583 20033
rect -3663 19963 -3583 19977
rect -3479 19977 -3467 20033
rect -3411 19977 -3399 20033
rect -3186 20406 -3169 20408
rect -3232 19988 -3186 19999
rect -3479 19963 -3399 19977
rect -3847 19883 -3767 19885
rect -4235 19827 -3835 19883
rect -3779 19827 -3767 19883
rect -2749 19884 -2693 20904
rect -1591 20892 -1511 20904
rect -2085 20853 -1999 20857
rect -2085 20797 -2073 20853
rect -2017 20797 -1999 20853
rect -2085 20785 -1999 20797
rect -2574 20640 -2528 20651
rect -2359 20649 -2283 20682
rect -2359 20603 -2348 20649
rect -2294 20603 -2283 20649
rect -2175 20649 -2099 20682
rect -2175 20603 -2164 20649
rect -2110 20603 -2099 20649
rect -1991 20649 -1915 20682
rect -1991 20603 -1980 20649
rect -1926 20603 -1915 20649
rect -1746 20640 -1700 20651
rect -2436 20557 -2390 20568
rect -2453 20530 -2436 20532
rect -2252 20557 -2206 20568
rect -2390 20530 -2373 20532
rect -2528 20410 -2441 20530
rect -2385 20410 -2373 20530
rect -2453 20408 -2436 20410
rect -2528 20110 -2436 20230
rect -2390 20408 -2373 20410
rect -2269 20230 -2252 20232
rect -2068 20557 -2022 20568
rect -2085 20530 -2068 20532
rect -1884 20557 -1838 20568
rect -2022 20530 -2005 20532
rect -2085 20410 -2073 20530
rect -2017 20410 -2005 20530
rect -2085 20408 -2068 20410
rect -2206 20230 -2189 20232
rect -2269 20110 -2257 20230
rect -2201 20110 -2189 20230
rect -2269 20108 -2252 20110
rect -2436 20072 -2390 20083
rect -2206 20108 -2189 20110
rect -2252 20072 -2206 20083
rect -2022 20408 -2005 20410
rect -1901 20230 -1884 20232
rect -1763 20530 -1746 20532
rect -1700 20530 -1683 20532
rect -1763 20409 -1751 20530
rect -1695 20409 -1683 20530
rect -1763 20407 -1746 20409
rect -1838 20230 -1821 20232
rect -1901 20110 -1889 20230
rect -1833 20110 -1821 20230
rect -1901 20108 -1884 20110
rect -2068 20072 -2022 20083
rect -1838 20108 -1821 20110
rect -1884 20072 -1838 20083
rect -2359 20034 -2348 20037
rect -2294 20034 -2283 20037
rect -2175 20034 -2164 20037
rect -2110 20034 -2099 20037
rect -1991 20034 -1980 20037
rect -1926 20034 -1915 20037
rect -2574 19989 -2528 20000
rect -2361 19978 -2349 20034
rect -2293 19978 -2281 20034
rect -2361 19964 -2281 19978
rect -2177 19978 -2165 20034
rect -2109 19978 -2097 20034
rect -2177 19964 -2097 19978
rect -1993 19978 -1981 20034
rect -1925 19978 -1913 20034
rect -1700 20407 -1683 20409
rect -1746 19989 -1700 20000
rect -1993 19964 -1913 19978
rect -2361 19884 -2281 19886
rect -2749 19828 -2349 19884
rect -2293 19828 -2281 19884
rect -3847 19825 -3767 19827
rect -2361 19826 -2281 19828
rect -3663 19767 -3583 19769
rect -4371 19711 -3651 19767
rect -3595 19711 -3583 19767
rect -3663 19709 -3583 19711
rect -3334 19767 -3254 19769
rect -3067 19768 -2997 19779
rect -2177 19768 -2097 19770
rect -3067 19767 -2165 19768
rect -3334 19711 -3322 19767
rect -3266 19711 -3065 19767
rect -3009 19712 -2165 19767
rect -2109 19712 -2097 19768
rect -3009 19711 -2749 19712
rect -3334 19709 -3254 19711
rect -3067 19701 -2997 19711
rect -2177 19710 -2097 19712
rect -1848 19768 -1768 19770
rect -1405 19768 -1335 19778
rect -1848 19712 -1836 19768
rect -1780 19712 -1403 19768
rect -1347 19712 -1335 19768
rect -1848 19710 -1768 19712
rect -1405 19700 -1335 19712
rect -329 19767 -273 21014
rect 2627 21012 2707 21014
rect 3293 21070 3363 21072
rect 3713 21070 3769 21800
rect 4605 21798 4685 21800
rect 5335 21800 6103 21856
rect 6159 21800 6171 21856
rect 4237 21706 4317 21720
rect 4024 21684 4070 21695
rect 4237 21650 4249 21706
rect 4305 21650 4317 21706
rect 4421 21706 4501 21720
rect 4421 21650 4433 21706
rect 4489 21650 4501 21706
rect 4605 21706 4685 21720
rect 4605 21650 4617 21706
rect 4673 21650 4685 21706
rect 4852 21684 4898 21695
rect 4239 21647 4250 21650
rect 4304 21647 4315 21650
rect 4423 21647 4434 21650
rect 4488 21647 4499 21650
rect 4607 21647 4618 21650
rect 4672 21647 4683 21650
rect 4162 21601 4208 21612
rect 4070 21427 4162 21601
rect 4162 21416 4208 21427
rect 4346 21601 4392 21612
rect 4346 21416 4392 21427
rect 4530 21601 4576 21612
rect 4714 21601 4760 21612
rect 4697 21574 4714 21576
rect 4760 21574 4777 21576
rect 4697 21454 4709 21574
rect 4765 21454 4777 21574
rect 4697 21452 4714 21454
rect 4530 21416 4576 21427
rect 4760 21452 4777 21454
rect 4714 21416 4760 21427
rect 4024 21199 4070 21344
rect 4239 21335 4250 21381
rect 4304 21335 4315 21381
rect 4239 21302 4315 21335
rect 4423 21335 4434 21381
rect 4488 21335 4499 21381
rect 4423 21302 4499 21335
rect 4607 21335 4618 21381
rect 4672 21335 4683 21381
rect 4607 21302 4683 21335
rect 4852 21199 4898 21344
rect 4012 21187 4092 21199
rect 4012 21131 4024 21187
rect 4080 21131 4092 21187
rect 4012 21119 4092 21131
rect 4830 21187 4908 21199
rect 4830 21131 4842 21187
rect 4898 21131 4908 21187
rect 4830 21119 4908 21131
rect 3293 21014 3305 21070
rect 3361 21014 3769 21070
rect 5335 21070 5391 21800
rect 6091 21798 6171 21800
rect 7755 21800 8659 21856
rect 8715 21800 8727 21856
rect 5723 21706 5803 21720
rect 5510 21684 5556 21695
rect 5723 21650 5735 21706
rect 5791 21650 5803 21706
rect 5907 21706 5987 21720
rect 5907 21650 5919 21706
rect 5975 21650 5987 21706
rect 6091 21706 6171 21720
rect 6091 21650 6103 21706
rect 6159 21650 6171 21706
rect 6338 21684 6384 21695
rect 5725 21647 5736 21650
rect 5790 21647 5801 21650
rect 5909 21647 5920 21650
rect 5974 21647 5985 21650
rect 6093 21647 6104 21650
rect 6158 21647 6169 21650
rect 5648 21601 5694 21612
rect 5556 21427 5648 21601
rect 5648 21416 5694 21427
rect 5832 21601 5878 21612
rect 5832 21416 5878 21427
rect 6016 21601 6062 21612
rect 6200 21601 6246 21612
rect 6183 21574 6200 21576
rect 6246 21574 6263 21576
rect 6183 21454 6195 21574
rect 6251 21454 6263 21574
rect 6183 21452 6200 21454
rect 6016 21416 6062 21427
rect 6246 21452 6263 21454
rect 6200 21416 6246 21427
rect 5510 21199 5556 21344
rect 5725 21335 5736 21381
rect 5790 21335 5801 21381
rect 5725 21302 5801 21335
rect 5909 21335 5920 21381
rect 5974 21335 5985 21381
rect 5909 21302 5985 21335
rect 6093 21335 6104 21381
rect 6158 21335 6169 21381
rect 6093 21302 6169 21335
rect 6338 21199 6384 21344
rect 5498 21187 5578 21199
rect 5498 21131 5510 21187
rect 5566 21131 5578 21187
rect 5498 21119 5578 21131
rect 6316 21187 6394 21199
rect 6316 21131 6328 21187
rect 6384 21131 6394 21187
rect 6316 21119 6394 21131
rect 6669 21070 6749 21080
rect 5335 21014 6681 21070
rect 6737 21014 6749 21070
rect 3293 21002 3363 21014
rect 1151 20959 1221 20961
rect 2451 20960 2531 20962
rect -193 20903 1153 20959
rect 1209 20903 1221 20959
rect -193 19883 -137 20903
rect 1151 20891 1221 20903
rect 1293 20904 2463 20960
rect 2519 20904 2531 20960
rect 471 20852 557 20856
rect 471 20796 483 20852
rect 539 20796 557 20852
rect 471 20784 557 20796
rect -18 20639 28 20650
rect 197 20648 273 20681
rect 197 20602 208 20648
rect 262 20602 273 20648
rect 381 20648 457 20681
rect 381 20602 392 20648
rect 446 20602 457 20648
rect 565 20648 641 20681
rect 565 20602 576 20648
rect 630 20602 641 20648
rect 810 20639 856 20650
rect 120 20556 166 20567
rect 103 20529 120 20531
rect 304 20556 350 20567
rect 166 20529 183 20531
rect 28 20409 115 20529
rect 171 20409 183 20529
rect 103 20407 120 20409
rect 28 20109 120 20229
rect 166 20407 183 20409
rect 287 20229 304 20231
rect 488 20556 534 20567
rect 471 20529 488 20531
rect 672 20556 718 20567
rect 534 20529 551 20531
rect 471 20409 483 20529
rect 539 20409 551 20529
rect 471 20407 488 20409
rect 350 20229 367 20231
rect 287 20109 299 20229
rect 355 20109 367 20229
rect 287 20107 304 20109
rect 120 20071 166 20082
rect 350 20107 367 20109
rect 304 20071 350 20082
rect 534 20407 551 20409
rect 655 20229 672 20231
rect 793 20529 810 20531
rect 856 20529 873 20531
rect 793 20408 805 20529
rect 861 20408 873 20529
rect 793 20406 810 20408
rect 718 20229 735 20231
rect 655 20109 667 20229
rect 723 20109 735 20229
rect 655 20107 672 20109
rect 488 20071 534 20082
rect 718 20107 735 20109
rect 672 20071 718 20082
rect 197 20033 208 20036
rect 262 20033 273 20036
rect 381 20033 392 20036
rect 446 20033 457 20036
rect 565 20033 576 20036
rect 630 20033 641 20036
rect -18 19988 28 19999
rect 195 19977 207 20033
rect 263 19977 275 20033
rect 195 19963 275 19977
rect 379 19977 391 20033
rect 447 19977 459 20033
rect 379 19963 459 19977
rect 563 19977 575 20033
rect 631 19977 643 20033
rect 856 20406 873 20408
rect 810 19988 856 19999
rect 563 19963 643 19977
rect 195 19883 275 19885
rect -193 19827 207 19883
rect 263 19827 275 19883
rect 1293 19884 1349 20904
rect 2451 20892 2531 20904
rect 1957 20853 2043 20857
rect 1957 20797 1969 20853
rect 2025 20797 2043 20853
rect 1957 20785 2043 20797
rect 1468 20640 1514 20651
rect 1683 20649 1759 20682
rect 1683 20603 1694 20649
rect 1748 20603 1759 20649
rect 1867 20649 1943 20682
rect 1867 20603 1878 20649
rect 1932 20603 1943 20649
rect 2051 20649 2127 20682
rect 2051 20603 2062 20649
rect 2116 20603 2127 20649
rect 2296 20640 2342 20651
rect 1606 20557 1652 20568
rect 1589 20530 1606 20532
rect 1790 20557 1836 20568
rect 1652 20530 1669 20532
rect 1514 20410 1601 20530
rect 1657 20410 1669 20530
rect 1589 20408 1606 20410
rect 1514 20110 1606 20230
rect 1652 20408 1669 20410
rect 1773 20230 1790 20232
rect 1974 20557 2020 20568
rect 1957 20530 1974 20532
rect 2158 20557 2204 20568
rect 2020 20530 2037 20532
rect 1957 20410 1969 20530
rect 2025 20410 2037 20530
rect 1957 20408 1974 20410
rect 1836 20230 1853 20232
rect 1773 20110 1785 20230
rect 1841 20110 1853 20230
rect 1773 20108 1790 20110
rect 1606 20072 1652 20083
rect 1836 20108 1853 20110
rect 1790 20072 1836 20083
rect 2020 20408 2037 20410
rect 2141 20230 2158 20232
rect 2279 20530 2296 20532
rect 2342 20530 2359 20532
rect 2279 20409 2291 20530
rect 2347 20409 2359 20530
rect 2279 20407 2296 20409
rect 2204 20230 2221 20232
rect 2141 20110 2153 20230
rect 2209 20110 2221 20230
rect 2141 20108 2158 20110
rect 1974 20072 2020 20083
rect 2204 20108 2221 20110
rect 2158 20072 2204 20083
rect 1683 20034 1694 20037
rect 1748 20034 1759 20037
rect 1867 20034 1878 20037
rect 1932 20034 1943 20037
rect 2051 20034 2062 20037
rect 2116 20034 2127 20037
rect 1468 19989 1514 20000
rect 1681 19978 1693 20034
rect 1749 19978 1761 20034
rect 1681 19964 1761 19978
rect 1865 19978 1877 20034
rect 1933 19978 1945 20034
rect 1865 19964 1945 19978
rect 2049 19978 2061 20034
rect 2117 19978 2129 20034
rect 2342 20407 2359 20409
rect 2296 19989 2342 20000
rect 2049 19964 2129 19978
rect 1681 19884 1761 19886
rect 1293 19828 1693 19884
rect 1749 19828 1761 19884
rect 195 19825 275 19827
rect 1681 19826 1761 19828
rect 379 19767 459 19769
rect -329 19711 391 19767
rect 447 19711 459 19767
rect 379 19709 459 19711
rect 708 19767 788 19769
rect 975 19768 1045 19779
rect 1865 19768 1945 19770
rect 975 19767 1877 19768
rect 708 19711 720 19767
rect 776 19711 977 19767
rect 1033 19712 1877 19767
rect 1933 19712 1945 19768
rect 1033 19711 1293 19712
rect 708 19709 788 19711
rect 975 19701 1045 19711
rect 1865 19710 1945 19712
rect 2194 19768 2274 19770
rect 2637 19768 2707 19778
rect 2194 19712 2206 19768
rect 2262 19712 2639 19768
rect 2695 19712 2707 19768
rect 2194 19710 2274 19712
rect 2637 19700 2707 19712
rect 3713 19767 3769 21014
rect 6669 21012 6749 21014
rect 7335 21070 7405 21072
rect 7755 21070 7811 21800
rect 8647 21798 8727 21800
rect 9377 21800 10145 21856
rect 10201 21800 10213 21856
rect 8279 21706 8359 21720
rect 8066 21684 8112 21695
rect 8279 21650 8291 21706
rect 8347 21650 8359 21706
rect 8463 21706 8543 21720
rect 8463 21650 8475 21706
rect 8531 21650 8543 21706
rect 8647 21706 8727 21720
rect 8647 21650 8659 21706
rect 8715 21650 8727 21706
rect 8894 21684 8940 21695
rect 8281 21647 8292 21650
rect 8346 21647 8357 21650
rect 8465 21647 8476 21650
rect 8530 21647 8541 21650
rect 8649 21647 8660 21650
rect 8714 21647 8725 21650
rect 8204 21601 8250 21612
rect 8112 21427 8204 21601
rect 8204 21416 8250 21427
rect 8388 21601 8434 21612
rect 8388 21416 8434 21427
rect 8572 21601 8618 21612
rect 8756 21601 8802 21612
rect 8739 21574 8756 21576
rect 8802 21574 8819 21576
rect 8739 21454 8751 21574
rect 8807 21454 8819 21574
rect 8739 21452 8756 21454
rect 8572 21416 8618 21427
rect 8802 21452 8819 21454
rect 8756 21416 8802 21427
rect 8066 21199 8112 21344
rect 8281 21335 8292 21381
rect 8346 21335 8357 21381
rect 8281 21302 8357 21335
rect 8465 21335 8476 21381
rect 8530 21335 8541 21381
rect 8465 21302 8541 21335
rect 8649 21335 8660 21381
rect 8714 21335 8725 21381
rect 8649 21302 8725 21335
rect 8894 21199 8940 21344
rect 8054 21187 8134 21199
rect 8054 21131 8066 21187
rect 8122 21131 8134 21187
rect 8054 21119 8134 21131
rect 8872 21187 8950 21199
rect 8872 21131 8884 21187
rect 8940 21131 8950 21187
rect 8872 21119 8950 21131
rect 7335 21014 7347 21070
rect 7403 21014 7811 21070
rect 9377 21070 9433 21800
rect 10133 21798 10213 21800
rect 11797 21800 12701 21856
rect 12757 21800 12769 21856
rect 9765 21706 9845 21720
rect 9552 21684 9598 21695
rect 9765 21650 9777 21706
rect 9833 21650 9845 21706
rect 9949 21706 10029 21720
rect 9949 21650 9961 21706
rect 10017 21650 10029 21706
rect 10133 21706 10213 21720
rect 10133 21650 10145 21706
rect 10201 21650 10213 21706
rect 10380 21684 10426 21695
rect 9767 21647 9778 21650
rect 9832 21647 9843 21650
rect 9951 21647 9962 21650
rect 10016 21647 10027 21650
rect 10135 21647 10146 21650
rect 10200 21647 10211 21650
rect 9690 21601 9736 21612
rect 9598 21427 9690 21601
rect 9690 21416 9736 21427
rect 9874 21601 9920 21612
rect 9874 21416 9920 21427
rect 10058 21601 10104 21612
rect 10242 21601 10288 21612
rect 10225 21574 10242 21576
rect 10288 21574 10305 21576
rect 10225 21454 10237 21574
rect 10293 21454 10305 21574
rect 10225 21452 10242 21454
rect 10058 21416 10104 21427
rect 10288 21452 10305 21454
rect 10242 21416 10288 21427
rect 9552 21199 9598 21344
rect 9767 21335 9778 21381
rect 9832 21335 9843 21381
rect 9767 21302 9843 21335
rect 9951 21335 9962 21381
rect 10016 21335 10027 21381
rect 9951 21302 10027 21335
rect 10135 21335 10146 21381
rect 10200 21335 10211 21381
rect 10135 21302 10211 21335
rect 10380 21199 10426 21344
rect 9540 21187 9620 21199
rect 9540 21131 9552 21187
rect 9608 21131 9620 21187
rect 9540 21119 9620 21131
rect 10358 21187 10436 21199
rect 10358 21131 10370 21187
rect 10426 21131 10436 21187
rect 10358 21119 10436 21131
rect 10711 21070 10791 21080
rect 9377 21014 10723 21070
rect 10779 21014 10791 21070
rect 7335 21002 7405 21014
rect 5193 20959 5263 20961
rect 6493 20960 6573 20962
rect 3849 20903 5195 20959
rect 5251 20903 5263 20959
rect 3849 19883 3905 20903
rect 5193 20891 5263 20903
rect 5335 20904 6505 20960
rect 6561 20904 6573 20960
rect 4513 20852 4599 20856
rect 4513 20796 4525 20852
rect 4581 20796 4599 20852
rect 4513 20784 4599 20796
rect 4024 20639 4070 20650
rect 4239 20648 4315 20681
rect 4239 20602 4250 20648
rect 4304 20602 4315 20648
rect 4423 20648 4499 20681
rect 4423 20602 4434 20648
rect 4488 20602 4499 20648
rect 4607 20648 4683 20681
rect 4607 20602 4618 20648
rect 4672 20602 4683 20648
rect 4852 20639 4898 20650
rect 4162 20556 4208 20567
rect 4145 20529 4162 20531
rect 4346 20556 4392 20567
rect 4208 20529 4225 20531
rect 4070 20409 4157 20529
rect 4213 20409 4225 20529
rect 4145 20407 4162 20409
rect 4070 20109 4162 20229
rect 4208 20407 4225 20409
rect 4329 20229 4346 20231
rect 4530 20556 4576 20567
rect 4513 20529 4530 20531
rect 4714 20556 4760 20567
rect 4576 20529 4593 20531
rect 4513 20409 4525 20529
rect 4581 20409 4593 20529
rect 4513 20407 4530 20409
rect 4392 20229 4409 20231
rect 4329 20109 4341 20229
rect 4397 20109 4409 20229
rect 4329 20107 4346 20109
rect 4162 20071 4208 20082
rect 4392 20107 4409 20109
rect 4346 20071 4392 20082
rect 4576 20407 4593 20409
rect 4697 20229 4714 20231
rect 4835 20529 4852 20531
rect 4898 20529 4915 20531
rect 4835 20408 4847 20529
rect 4903 20408 4915 20529
rect 4835 20406 4852 20408
rect 4760 20229 4777 20231
rect 4697 20109 4709 20229
rect 4765 20109 4777 20229
rect 4697 20107 4714 20109
rect 4530 20071 4576 20082
rect 4760 20107 4777 20109
rect 4714 20071 4760 20082
rect 4239 20033 4250 20036
rect 4304 20033 4315 20036
rect 4423 20033 4434 20036
rect 4488 20033 4499 20036
rect 4607 20033 4618 20036
rect 4672 20033 4683 20036
rect 4024 19988 4070 19999
rect 4237 19977 4249 20033
rect 4305 19977 4317 20033
rect 4237 19963 4317 19977
rect 4421 19977 4433 20033
rect 4489 19977 4501 20033
rect 4421 19963 4501 19977
rect 4605 19977 4617 20033
rect 4673 19977 4685 20033
rect 4898 20406 4915 20408
rect 4852 19988 4898 19999
rect 4605 19963 4685 19977
rect 4237 19883 4317 19885
rect 3849 19827 4249 19883
rect 4305 19827 4317 19883
rect 5335 19884 5391 20904
rect 6493 20892 6573 20904
rect 5999 20853 6085 20857
rect 5999 20797 6011 20853
rect 6067 20797 6085 20853
rect 5999 20785 6085 20797
rect 5510 20640 5556 20651
rect 5725 20649 5801 20682
rect 5725 20603 5736 20649
rect 5790 20603 5801 20649
rect 5909 20649 5985 20682
rect 5909 20603 5920 20649
rect 5974 20603 5985 20649
rect 6093 20649 6169 20682
rect 6093 20603 6104 20649
rect 6158 20603 6169 20649
rect 6338 20640 6384 20651
rect 5648 20557 5694 20568
rect 5631 20530 5648 20532
rect 5832 20557 5878 20568
rect 5694 20530 5711 20532
rect 5556 20410 5643 20530
rect 5699 20410 5711 20530
rect 5631 20408 5648 20410
rect 5556 20110 5648 20230
rect 5694 20408 5711 20410
rect 5815 20230 5832 20232
rect 6016 20557 6062 20568
rect 5999 20530 6016 20532
rect 6200 20557 6246 20568
rect 6062 20530 6079 20532
rect 5999 20410 6011 20530
rect 6067 20410 6079 20530
rect 5999 20408 6016 20410
rect 5878 20230 5895 20232
rect 5815 20110 5827 20230
rect 5883 20110 5895 20230
rect 5815 20108 5832 20110
rect 5648 20072 5694 20083
rect 5878 20108 5895 20110
rect 5832 20072 5878 20083
rect 6062 20408 6079 20410
rect 6183 20230 6200 20232
rect 6321 20530 6338 20532
rect 6384 20530 6401 20532
rect 6321 20409 6333 20530
rect 6389 20409 6401 20530
rect 6321 20407 6338 20409
rect 6246 20230 6263 20232
rect 6183 20110 6195 20230
rect 6251 20110 6263 20230
rect 6183 20108 6200 20110
rect 6016 20072 6062 20083
rect 6246 20108 6263 20110
rect 6200 20072 6246 20083
rect 5725 20034 5736 20037
rect 5790 20034 5801 20037
rect 5909 20034 5920 20037
rect 5974 20034 5985 20037
rect 6093 20034 6104 20037
rect 6158 20034 6169 20037
rect 5510 19989 5556 20000
rect 5723 19978 5735 20034
rect 5791 19978 5803 20034
rect 5723 19964 5803 19978
rect 5907 19978 5919 20034
rect 5975 19978 5987 20034
rect 5907 19964 5987 19978
rect 6091 19978 6103 20034
rect 6159 19978 6171 20034
rect 6384 20407 6401 20409
rect 6338 19989 6384 20000
rect 6091 19964 6171 19978
rect 5723 19884 5803 19886
rect 5335 19828 5735 19884
rect 5791 19828 5803 19884
rect 4237 19825 4317 19827
rect 5723 19826 5803 19828
rect 4421 19767 4501 19769
rect 3713 19711 4433 19767
rect 4489 19711 4501 19767
rect 4421 19709 4501 19711
rect 4750 19767 4830 19769
rect 5017 19768 5087 19779
rect 5907 19768 5987 19770
rect 5017 19767 5919 19768
rect 4750 19711 4762 19767
rect 4818 19711 5019 19767
rect 5075 19712 5919 19767
rect 5975 19712 5987 19768
rect 5075 19711 5335 19712
rect 4750 19709 4830 19711
rect 5017 19701 5087 19711
rect 5907 19710 5987 19712
rect 6236 19768 6316 19770
rect 6679 19768 6749 19778
rect 6236 19712 6248 19768
rect 6304 19712 6681 19768
rect 6737 19712 6749 19768
rect 6236 19710 6316 19712
rect 6679 19700 6749 19712
rect 7755 19767 7811 21014
rect 10711 21012 10791 21014
rect 11377 21070 11447 21072
rect 11797 21070 11853 21800
rect 12689 21798 12769 21800
rect 13419 21800 14187 21856
rect 14243 21800 14255 21856
rect 12321 21706 12401 21720
rect 12108 21684 12154 21695
rect 12321 21650 12333 21706
rect 12389 21650 12401 21706
rect 12505 21706 12585 21720
rect 12505 21650 12517 21706
rect 12573 21650 12585 21706
rect 12689 21706 12769 21720
rect 12689 21650 12701 21706
rect 12757 21650 12769 21706
rect 12936 21684 12982 21695
rect 12323 21647 12334 21650
rect 12388 21647 12399 21650
rect 12507 21647 12518 21650
rect 12572 21647 12583 21650
rect 12691 21647 12702 21650
rect 12756 21647 12767 21650
rect 12246 21601 12292 21612
rect 12154 21427 12246 21601
rect 12246 21416 12292 21427
rect 12430 21601 12476 21612
rect 12430 21416 12476 21427
rect 12614 21601 12660 21612
rect 12798 21601 12844 21612
rect 12781 21574 12798 21576
rect 12844 21574 12861 21576
rect 12781 21454 12793 21574
rect 12849 21454 12861 21574
rect 12781 21452 12798 21454
rect 12614 21416 12660 21427
rect 12844 21452 12861 21454
rect 12798 21416 12844 21427
rect 12108 21199 12154 21344
rect 12323 21335 12334 21381
rect 12388 21335 12399 21381
rect 12323 21302 12399 21335
rect 12507 21335 12518 21381
rect 12572 21335 12583 21381
rect 12507 21302 12583 21335
rect 12691 21335 12702 21381
rect 12756 21335 12767 21381
rect 12691 21302 12767 21335
rect 12936 21199 12982 21344
rect 12096 21187 12176 21199
rect 12096 21131 12108 21187
rect 12164 21131 12176 21187
rect 12096 21119 12176 21131
rect 12914 21187 12992 21199
rect 12914 21131 12926 21187
rect 12982 21131 12992 21187
rect 12914 21119 12992 21131
rect 11377 21014 11389 21070
rect 11445 21014 11853 21070
rect 13419 21070 13475 21800
rect 14175 21798 14255 21800
rect 15839 21800 16743 21856
rect 16799 21800 16811 21856
rect 13807 21706 13887 21720
rect 13594 21684 13640 21695
rect 13807 21650 13819 21706
rect 13875 21650 13887 21706
rect 13991 21706 14071 21720
rect 13991 21650 14003 21706
rect 14059 21650 14071 21706
rect 14175 21706 14255 21720
rect 14175 21650 14187 21706
rect 14243 21650 14255 21706
rect 14422 21684 14468 21695
rect 13809 21647 13820 21650
rect 13874 21647 13885 21650
rect 13993 21647 14004 21650
rect 14058 21647 14069 21650
rect 14177 21647 14188 21650
rect 14242 21647 14253 21650
rect 13732 21601 13778 21612
rect 13640 21427 13732 21601
rect 13732 21416 13778 21427
rect 13916 21601 13962 21612
rect 13916 21416 13962 21427
rect 14100 21601 14146 21612
rect 14284 21601 14330 21612
rect 14267 21574 14284 21576
rect 14330 21574 14347 21576
rect 14267 21454 14279 21574
rect 14335 21454 14347 21574
rect 14267 21452 14284 21454
rect 14100 21416 14146 21427
rect 14330 21452 14347 21454
rect 14284 21416 14330 21427
rect 13594 21199 13640 21344
rect 13809 21335 13820 21381
rect 13874 21335 13885 21381
rect 13809 21302 13885 21335
rect 13993 21335 14004 21381
rect 14058 21335 14069 21381
rect 13993 21302 14069 21335
rect 14177 21335 14188 21381
rect 14242 21335 14253 21381
rect 14177 21302 14253 21335
rect 14422 21199 14468 21344
rect 13582 21187 13662 21199
rect 13582 21131 13594 21187
rect 13650 21131 13662 21187
rect 13582 21119 13662 21131
rect 14400 21187 14478 21199
rect 14400 21131 14412 21187
rect 14468 21131 14478 21187
rect 14400 21119 14478 21131
rect 14753 21070 14833 21080
rect 13419 21014 14765 21070
rect 14821 21014 14833 21070
rect 11377 21002 11447 21014
rect 9235 20959 9305 20961
rect 10535 20960 10615 20962
rect 7891 20903 9237 20959
rect 9293 20903 9305 20959
rect 7891 19883 7947 20903
rect 9235 20891 9305 20903
rect 9377 20904 10547 20960
rect 10603 20904 10615 20960
rect 8555 20852 8641 20856
rect 8555 20796 8567 20852
rect 8623 20796 8641 20852
rect 8555 20784 8641 20796
rect 8066 20639 8112 20650
rect 8281 20648 8357 20681
rect 8281 20602 8292 20648
rect 8346 20602 8357 20648
rect 8465 20648 8541 20681
rect 8465 20602 8476 20648
rect 8530 20602 8541 20648
rect 8649 20648 8725 20681
rect 8649 20602 8660 20648
rect 8714 20602 8725 20648
rect 8894 20639 8940 20650
rect 8204 20556 8250 20567
rect 8187 20529 8204 20531
rect 8388 20556 8434 20567
rect 8250 20529 8267 20531
rect 8112 20409 8199 20529
rect 8255 20409 8267 20529
rect 8187 20407 8204 20409
rect 8112 20109 8204 20229
rect 8250 20407 8267 20409
rect 8371 20229 8388 20231
rect 8572 20556 8618 20567
rect 8555 20529 8572 20531
rect 8756 20556 8802 20567
rect 8618 20529 8635 20531
rect 8555 20409 8567 20529
rect 8623 20409 8635 20529
rect 8555 20407 8572 20409
rect 8434 20229 8451 20231
rect 8371 20109 8383 20229
rect 8439 20109 8451 20229
rect 8371 20107 8388 20109
rect 8204 20071 8250 20082
rect 8434 20107 8451 20109
rect 8388 20071 8434 20082
rect 8618 20407 8635 20409
rect 8739 20229 8756 20231
rect 8877 20529 8894 20531
rect 8940 20529 8957 20531
rect 8877 20408 8889 20529
rect 8945 20408 8957 20529
rect 8877 20406 8894 20408
rect 8802 20229 8819 20231
rect 8739 20109 8751 20229
rect 8807 20109 8819 20229
rect 8739 20107 8756 20109
rect 8572 20071 8618 20082
rect 8802 20107 8819 20109
rect 8756 20071 8802 20082
rect 8281 20033 8292 20036
rect 8346 20033 8357 20036
rect 8465 20033 8476 20036
rect 8530 20033 8541 20036
rect 8649 20033 8660 20036
rect 8714 20033 8725 20036
rect 8066 19988 8112 19999
rect 8279 19977 8291 20033
rect 8347 19977 8359 20033
rect 8279 19963 8359 19977
rect 8463 19977 8475 20033
rect 8531 19977 8543 20033
rect 8463 19963 8543 19977
rect 8647 19977 8659 20033
rect 8715 19977 8727 20033
rect 8940 20406 8957 20408
rect 8894 19988 8940 19999
rect 8647 19963 8727 19977
rect 8279 19883 8359 19885
rect 7891 19827 8291 19883
rect 8347 19827 8359 19883
rect 9377 19884 9433 20904
rect 10535 20892 10615 20904
rect 10041 20853 10127 20857
rect 10041 20797 10053 20853
rect 10109 20797 10127 20853
rect 10041 20785 10127 20797
rect 9552 20640 9598 20651
rect 9767 20649 9843 20682
rect 9767 20603 9778 20649
rect 9832 20603 9843 20649
rect 9951 20649 10027 20682
rect 9951 20603 9962 20649
rect 10016 20603 10027 20649
rect 10135 20649 10211 20682
rect 10135 20603 10146 20649
rect 10200 20603 10211 20649
rect 10380 20640 10426 20651
rect 9690 20557 9736 20568
rect 9673 20530 9690 20532
rect 9874 20557 9920 20568
rect 9736 20530 9753 20532
rect 9598 20410 9685 20530
rect 9741 20410 9753 20530
rect 9673 20408 9690 20410
rect 9598 20110 9690 20230
rect 9736 20408 9753 20410
rect 9857 20230 9874 20232
rect 10058 20557 10104 20568
rect 10041 20530 10058 20532
rect 10242 20557 10288 20568
rect 10104 20530 10121 20532
rect 10041 20410 10053 20530
rect 10109 20410 10121 20530
rect 10041 20408 10058 20410
rect 9920 20230 9937 20232
rect 9857 20110 9869 20230
rect 9925 20110 9937 20230
rect 9857 20108 9874 20110
rect 9690 20072 9736 20083
rect 9920 20108 9937 20110
rect 9874 20072 9920 20083
rect 10104 20408 10121 20410
rect 10225 20230 10242 20232
rect 10363 20530 10380 20532
rect 10426 20530 10443 20532
rect 10363 20409 10375 20530
rect 10431 20409 10443 20530
rect 10363 20407 10380 20409
rect 10288 20230 10305 20232
rect 10225 20110 10237 20230
rect 10293 20110 10305 20230
rect 10225 20108 10242 20110
rect 10058 20072 10104 20083
rect 10288 20108 10305 20110
rect 10242 20072 10288 20083
rect 9767 20034 9778 20037
rect 9832 20034 9843 20037
rect 9951 20034 9962 20037
rect 10016 20034 10027 20037
rect 10135 20034 10146 20037
rect 10200 20034 10211 20037
rect 9552 19989 9598 20000
rect 9765 19978 9777 20034
rect 9833 19978 9845 20034
rect 9765 19964 9845 19978
rect 9949 19978 9961 20034
rect 10017 19978 10029 20034
rect 9949 19964 10029 19978
rect 10133 19978 10145 20034
rect 10201 19978 10213 20034
rect 10426 20407 10443 20409
rect 10380 19989 10426 20000
rect 10133 19964 10213 19978
rect 9765 19884 9845 19886
rect 9377 19828 9777 19884
rect 9833 19828 9845 19884
rect 8279 19825 8359 19827
rect 9765 19826 9845 19828
rect 8463 19767 8543 19769
rect 7755 19711 8475 19767
rect 8531 19711 8543 19767
rect 8463 19709 8543 19711
rect 8792 19767 8872 19769
rect 9059 19768 9129 19779
rect 9949 19768 10029 19770
rect 9059 19767 9961 19768
rect 8792 19711 8804 19767
rect 8860 19711 9061 19767
rect 9117 19712 9961 19767
rect 10017 19712 10029 19768
rect 9117 19711 9377 19712
rect 8792 19709 8872 19711
rect 9059 19701 9129 19711
rect 9949 19710 10029 19712
rect 10278 19768 10358 19770
rect 10721 19768 10791 19778
rect 10278 19712 10290 19768
rect 10346 19712 10723 19768
rect 10779 19712 10791 19768
rect 10278 19710 10358 19712
rect 10721 19700 10791 19712
rect 11797 19767 11853 21014
rect 14753 21012 14833 21014
rect 15375 21070 15453 21082
rect 15839 21070 15895 21800
rect 16731 21798 16811 21800
rect 17461 21800 18229 21856
rect 18285 21800 18297 21856
rect 16363 21706 16443 21720
rect 16150 21684 16196 21695
rect 16363 21650 16375 21706
rect 16431 21650 16443 21706
rect 16547 21706 16627 21720
rect 16547 21650 16559 21706
rect 16615 21650 16627 21706
rect 16731 21706 16811 21720
rect 16731 21650 16743 21706
rect 16799 21650 16811 21706
rect 16978 21684 17024 21695
rect 16365 21647 16376 21650
rect 16430 21647 16441 21650
rect 16549 21647 16560 21650
rect 16614 21647 16625 21650
rect 16733 21647 16744 21650
rect 16798 21647 16809 21650
rect 16288 21601 16334 21612
rect 16196 21427 16288 21601
rect 16288 21416 16334 21427
rect 16472 21601 16518 21612
rect 16472 21416 16518 21427
rect 16656 21601 16702 21612
rect 16840 21601 16886 21612
rect 16823 21574 16840 21576
rect 16886 21574 16903 21576
rect 16823 21454 16835 21574
rect 16891 21454 16903 21574
rect 16823 21452 16840 21454
rect 16656 21416 16702 21427
rect 16886 21452 16903 21454
rect 16840 21416 16886 21427
rect 16150 21199 16196 21344
rect 16365 21335 16376 21381
rect 16430 21335 16441 21381
rect 16365 21302 16441 21335
rect 16549 21335 16560 21381
rect 16614 21335 16625 21381
rect 16549 21302 16625 21335
rect 16733 21335 16744 21381
rect 16798 21335 16809 21381
rect 16733 21302 16809 21335
rect 16978 21199 17024 21344
rect 16138 21187 16218 21199
rect 16138 21131 16150 21187
rect 16206 21131 16218 21187
rect 16138 21119 16218 21131
rect 16956 21187 17034 21199
rect 16956 21131 16968 21187
rect 17024 21131 17034 21187
rect 16956 21119 17034 21131
rect 15375 21014 15386 21070
rect 15442 21014 15895 21070
rect 17461 21070 17517 21800
rect 18217 21798 18297 21800
rect 17849 21706 17929 21720
rect 17636 21684 17682 21695
rect 17849 21650 17861 21706
rect 17917 21650 17929 21706
rect 18033 21706 18113 21720
rect 18033 21650 18045 21706
rect 18101 21650 18113 21706
rect 18217 21706 18297 21720
rect 18217 21650 18229 21706
rect 18285 21650 18297 21706
rect 18464 21684 18510 21695
rect 17851 21647 17862 21650
rect 17916 21647 17927 21650
rect 18035 21647 18046 21650
rect 18100 21647 18111 21650
rect 18219 21647 18230 21650
rect 18284 21647 18295 21650
rect 17774 21601 17820 21612
rect 17682 21427 17774 21601
rect 17774 21416 17820 21427
rect 17958 21601 18004 21612
rect 17958 21416 18004 21427
rect 18142 21601 18188 21612
rect 18326 21601 18372 21612
rect 18309 21574 18326 21576
rect 18372 21574 18389 21576
rect 18309 21454 18321 21574
rect 18377 21454 18389 21574
rect 18309 21452 18326 21454
rect 18142 21416 18188 21427
rect 18372 21452 18389 21454
rect 18326 21416 18372 21427
rect 17636 21199 17682 21344
rect 17851 21335 17862 21381
rect 17916 21335 17927 21381
rect 17851 21302 17927 21335
rect 18035 21335 18046 21381
rect 18100 21335 18111 21381
rect 18035 21302 18111 21335
rect 18219 21335 18230 21381
rect 18284 21335 18295 21381
rect 18219 21302 18295 21335
rect 18464 21199 18510 21344
rect 17624 21187 17704 21199
rect 17624 21131 17636 21187
rect 17692 21131 17704 21187
rect 17624 21119 17704 21131
rect 18442 21187 18520 21199
rect 18442 21131 18454 21187
rect 18510 21131 18520 21187
rect 18442 21119 18520 21131
rect 18795 21070 18875 21080
rect 17461 21014 18807 21070
rect 18863 21014 18875 21070
rect 15375 21002 15453 21014
rect 13277 20959 13347 20961
rect 14577 20960 14657 20962
rect 11933 20903 13279 20959
rect 13335 20903 13347 20959
rect 11933 19883 11989 20903
rect 13277 20891 13347 20903
rect 13419 20904 14589 20960
rect 14645 20904 14657 20960
rect 12597 20852 12683 20856
rect 12597 20796 12609 20852
rect 12665 20796 12683 20852
rect 12597 20784 12683 20796
rect 12108 20639 12154 20650
rect 12323 20648 12399 20681
rect 12323 20602 12334 20648
rect 12388 20602 12399 20648
rect 12507 20648 12583 20681
rect 12507 20602 12518 20648
rect 12572 20602 12583 20648
rect 12691 20648 12767 20681
rect 12691 20602 12702 20648
rect 12756 20602 12767 20648
rect 12936 20639 12982 20650
rect 12246 20556 12292 20567
rect 12229 20529 12246 20531
rect 12430 20556 12476 20567
rect 12292 20529 12309 20531
rect 12154 20409 12241 20529
rect 12297 20409 12309 20529
rect 12229 20407 12246 20409
rect 12154 20109 12246 20229
rect 12292 20407 12309 20409
rect 12413 20229 12430 20231
rect 12614 20556 12660 20567
rect 12597 20529 12614 20531
rect 12798 20556 12844 20567
rect 12660 20529 12677 20531
rect 12597 20409 12609 20529
rect 12665 20409 12677 20529
rect 12597 20407 12614 20409
rect 12476 20229 12493 20231
rect 12413 20109 12425 20229
rect 12481 20109 12493 20229
rect 12413 20107 12430 20109
rect 12246 20071 12292 20082
rect 12476 20107 12493 20109
rect 12430 20071 12476 20082
rect 12660 20407 12677 20409
rect 12781 20229 12798 20231
rect 12919 20529 12936 20531
rect 12982 20529 12999 20531
rect 12919 20408 12931 20529
rect 12987 20408 12999 20529
rect 12919 20406 12936 20408
rect 12844 20229 12861 20231
rect 12781 20109 12793 20229
rect 12849 20109 12861 20229
rect 12781 20107 12798 20109
rect 12614 20071 12660 20082
rect 12844 20107 12861 20109
rect 12798 20071 12844 20082
rect 12323 20033 12334 20036
rect 12388 20033 12399 20036
rect 12507 20033 12518 20036
rect 12572 20033 12583 20036
rect 12691 20033 12702 20036
rect 12756 20033 12767 20036
rect 12108 19988 12154 19999
rect 12321 19977 12333 20033
rect 12389 19977 12401 20033
rect 12321 19963 12401 19977
rect 12505 19977 12517 20033
rect 12573 19977 12585 20033
rect 12505 19963 12585 19977
rect 12689 19977 12701 20033
rect 12757 19977 12769 20033
rect 12982 20406 12999 20408
rect 12936 19988 12982 19999
rect 12689 19963 12769 19977
rect 12321 19883 12401 19885
rect 11933 19827 12333 19883
rect 12389 19827 12401 19883
rect 13419 19884 13475 20904
rect 14577 20892 14657 20904
rect 14083 20853 14169 20857
rect 14083 20797 14095 20853
rect 14151 20797 14169 20853
rect 14083 20785 14169 20797
rect 13594 20640 13640 20651
rect 13809 20649 13885 20682
rect 13809 20603 13820 20649
rect 13874 20603 13885 20649
rect 13993 20649 14069 20682
rect 13993 20603 14004 20649
rect 14058 20603 14069 20649
rect 14177 20649 14253 20682
rect 14177 20603 14188 20649
rect 14242 20603 14253 20649
rect 14422 20640 14468 20651
rect 13732 20557 13778 20568
rect 13715 20530 13732 20532
rect 13916 20557 13962 20568
rect 13778 20530 13795 20532
rect 13640 20410 13727 20530
rect 13783 20410 13795 20530
rect 13715 20408 13732 20410
rect 13640 20110 13732 20230
rect 13778 20408 13795 20410
rect 13899 20230 13916 20232
rect 14100 20557 14146 20568
rect 14083 20530 14100 20532
rect 14284 20557 14330 20568
rect 14146 20530 14163 20532
rect 14083 20410 14095 20530
rect 14151 20410 14163 20530
rect 14083 20408 14100 20410
rect 13962 20230 13979 20232
rect 13899 20110 13911 20230
rect 13967 20110 13979 20230
rect 13899 20108 13916 20110
rect 13732 20072 13778 20083
rect 13962 20108 13979 20110
rect 13916 20072 13962 20083
rect 14146 20408 14163 20410
rect 14267 20230 14284 20232
rect 14405 20530 14422 20532
rect 14468 20530 14485 20532
rect 14405 20409 14417 20530
rect 14473 20409 14485 20530
rect 14405 20407 14422 20409
rect 14330 20230 14347 20232
rect 14267 20110 14279 20230
rect 14335 20110 14347 20230
rect 14267 20108 14284 20110
rect 14100 20072 14146 20083
rect 14330 20108 14347 20110
rect 14284 20072 14330 20083
rect 13809 20034 13820 20037
rect 13874 20034 13885 20037
rect 13993 20034 14004 20037
rect 14058 20034 14069 20037
rect 14177 20034 14188 20037
rect 14242 20034 14253 20037
rect 13594 19989 13640 20000
rect 13807 19978 13819 20034
rect 13875 19978 13887 20034
rect 13807 19964 13887 19978
rect 13991 19978 14003 20034
rect 14059 19978 14071 20034
rect 13991 19964 14071 19978
rect 14175 19978 14187 20034
rect 14243 19978 14255 20034
rect 14468 20407 14485 20409
rect 14422 19989 14468 20000
rect 14175 19964 14255 19978
rect 13807 19884 13887 19886
rect 13419 19828 13819 19884
rect 13875 19828 13887 19884
rect 12321 19825 12401 19827
rect 13807 19826 13887 19828
rect 12505 19767 12585 19769
rect 11797 19711 12517 19767
rect 12573 19711 12585 19767
rect 12505 19709 12585 19711
rect 12834 19767 12914 19769
rect 13101 19768 13171 19779
rect 13991 19768 14071 19770
rect 13101 19767 14003 19768
rect 12834 19711 12846 19767
rect 12902 19711 13103 19767
rect 13159 19712 14003 19767
rect 14059 19712 14071 19768
rect 13159 19711 13419 19712
rect 12834 19709 12914 19711
rect 13101 19701 13171 19711
rect 13991 19710 14071 19712
rect 14320 19768 14400 19770
rect 14763 19768 14833 19778
rect 14320 19712 14332 19768
rect 14388 19712 14765 19768
rect 14821 19712 14833 19768
rect 14320 19710 14400 19712
rect 14763 19700 14833 19712
rect 15839 19767 15895 21014
rect 18795 21012 18875 21014
rect 17319 20959 17389 20961
rect 18619 20960 18699 20962
rect 15975 20903 17321 20959
rect 17377 20903 17389 20959
rect 15975 19883 16031 20903
rect 17319 20891 17389 20903
rect 17461 20904 18631 20960
rect 18687 20904 18699 20960
rect 16639 20852 16725 20856
rect 16639 20796 16651 20852
rect 16707 20796 16725 20852
rect 16639 20784 16725 20796
rect 16150 20639 16196 20650
rect 16365 20648 16441 20681
rect 16365 20602 16376 20648
rect 16430 20602 16441 20648
rect 16549 20648 16625 20681
rect 16549 20602 16560 20648
rect 16614 20602 16625 20648
rect 16733 20648 16809 20681
rect 16733 20602 16744 20648
rect 16798 20602 16809 20648
rect 16978 20639 17024 20650
rect 16288 20556 16334 20567
rect 16271 20529 16288 20531
rect 16472 20556 16518 20567
rect 16334 20529 16351 20531
rect 16196 20409 16283 20529
rect 16339 20409 16351 20529
rect 16271 20407 16288 20409
rect 16196 20109 16288 20229
rect 16334 20407 16351 20409
rect 16455 20229 16472 20231
rect 16656 20556 16702 20567
rect 16639 20529 16656 20531
rect 16840 20556 16886 20567
rect 16702 20529 16719 20531
rect 16639 20409 16651 20529
rect 16707 20409 16719 20529
rect 16639 20407 16656 20409
rect 16518 20229 16535 20231
rect 16455 20109 16467 20229
rect 16523 20109 16535 20229
rect 16455 20107 16472 20109
rect 16288 20071 16334 20082
rect 16518 20107 16535 20109
rect 16472 20071 16518 20082
rect 16702 20407 16719 20409
rect 16823 20229 16840 20231
rect 16961 20529 16978 20531
rect 17024 20529 17041 20531
rect 16961 20408 16973 20529
rect 17029 20408 17041 20529
rect 16961 20406 16978 20408
rect 16886 20229 16903 20231
rect 16823 20109 16835 20229
rect 16891 20109 16903 20229
rect 16823 20107 16840 20109
rect 16656 20071 16702 20082
rect 16886 20107 16903 20109
rect 16840 20071 16886 20082
rect 16365 20033 16376 20036
rect 16430 20033 16441 20036
rect 16549 20033 16560 20036
rect 16614 20033 16625 20036
rect 16733 20033 16744 20036
rect 16798 20033 16809 20036
rect 16150 19988 16196 19999
rect 16363 19977 16375 20033
rect 16431 19977 16443 20033
rect 16363 19963 16443 19977
rect 16547 19977 16559 20033
rect 16615 19977 16627 20033
rect 16547 19963 16627 19977
rect 16731 19977 16743 20033
rect 16799 19977 16811 20033
rect 17024 20406 17041 20408
rect 16978 19988 17024 19999
rect 16731 19963 16811 19977
rect 16363 19883 16443 19885
rect 15975 19827 16375 19883
rect 16431 19827 16443 19883
rect 17461 19884 17517 20904
rect 18619 20892 18699 20904
rect 18125 20853 18211 20857
rect 18125 20797 18137 20853
rect 18193 20797 18211 20853
rect 18125 20785 18211 20797
rect 17636 20640 17682 20651
rect 17851 20649 17927 20682
rect 17851 20603 17862 20649
rect 17916 20603 17927 20649
rect 18035 20649 18111 20682
rect 18035 20603 18046 20649
rect 18100 20603 18111 20649
rect 18219 20649 18295 20682
rect 18219 20603 18230 20649
rect 18284 20603 18295 20649
rect 18464 20640 18510 20651
rect 17774 20557 17820 20568
rect 17757 20530 17774 20532
rect 17958 20557 18004 20568
rect 17820 20530 17837 20532
rect 17682 20410 17769 20530
rect 17825 20410 17837 20530
rect 17757 20408 17774 20410
rect 17682 20110 17774 20230
rect 17820 20408 17837 20410
rect 17941 20230 17958 20232
rect 18142 20557 18188 20568
rect 18125 20530 18142 20532
rect 18326 20557 18372 20568
rect 18188 20530 18205 20532
rect 18125 20410 18137 20530
rect 18193 20410 18205 20530
rect 18125 20408 18142 20410
rect 18004 20230 18021 20232
rect 17941 20110 17953 20230
rect 18009 20110 18021 20230
rect 17941 20108 17958 20110
rect 17774 20072 17820 20083
rect 18004 20108 18021 20110
rect 17958 20072 18004 20083
rect 18188 20408 18205 20410
rect 18309 20230 18326 20232
rect 18447 20530 18464 20532
rect 18510 20530 18527 20532
rect 18447 20409 18459 20530
rect 18515 20409 18527 20530
rect 18447 20407 18464 20409
rect 18372 20230 18389 20232
rect 18309 20110 18321 20230
rect 18377 20110 18389 20230
rect 18309 20108 18326 20110
rect 18142 20072 18188 20083
rect 18372 20108 18389 20110
rect 18326 20072 18372 20083
rect 17851 20034 17862 20037
rect 17916 20034 17927 20037
rect 18035 20034 18046 20037
rect 18100 20034 18111 20037
rect 18219 20034 18230 20037
rect 18284 20034 18295 20037
rect 17636 19989 17682 20000
rect 17849 19978 17861 20034
rect 17917 19978 17929 20034
rect 17849 19964 17929 19978
rect 18033 19978 18045 20034
rect 18101 19978 18113 20034
rect 18033 19964 18113 19978
rect 18217 19978 18229 20034
rect 18285 19978 18297 20034
rect 18510 20407 18527 20409
rect 18464 19989 18510 20000
rect 18217 19964 18297 19978
rect 17849 19884 17929 19886
rect 17461 19828 17861 19884
rect 17917 19828 17929 19884
rect 16363 19825 16443 19827
rect 17849 19826 17929 19828
rect 16547 19767 16627 19769
rect 15839 19711 16559 19767
rect 16615 19711 16627 19767
rect 16547 19709 16627 19711
rect 16876 19767 16956 19769
rect 17143 19768 17213 19779
rect 18033 19768 18113 19770
rect 17143 19767 18045 19768
rect 16876 19711 16888 19767
rect 16944 19711 17145 19767
rect 17201 19712 18045 19767
rect 18101 19712 18113 19768
rect 17201 19711 17461 19712
rect 16876 19709 16956 19711
rect 17143 19701 17213 19711
rect 18033 19710 18113 19712
rect 18362 19768 18442 19770
rect 18805 19768 18875 19778
rect 18362 19712 18374 19768
rect 18430 19712 18807 19768
rect 18863 19712 18875 19768
rect 18362 19710 18442 19712
rect 18805 19700 18875 19712
rect -8561 19654 -8491 19666
rect -7521 19654 -7441 19656
rect -6035 19655 -5955 19657
rect -8561 19598 -8549 19654
rect -8493 19598 -7509 19654
rect -7453 19598 -7441 19654
rect -8561 19586 -8491 19598
rect -8277 18867 -8221 19598
rect -7521 19596 -7441 19598
rect -6791 19599 -6023 19655
rect -5967 19599 -5955 19655
rect -7889 19504 -7809 19518
rect -8102 19482 -8056 19493
rect -7889 19448 -7877 19504
rect -7821 19448 -7809 19504
rect -7705 19504 -7625 19518
rect -7705 19448 -7693 19504
rect -7637 19448 -7625 19504
rect -7521 19504 -7441 19518
rect -7521 19448 -7509 19504
rect -7453 19448 -7441 19504
rect -7274 19482 -7228 19493
rect -7887 19445 -7876 19448
rect -7822 19445 -7811 19448
rect -7703 19445 -7692 19448
rect -7638 19445 -7627 19448
rect -7519 19445 -7508 19448
rect -7454 19445 -7443 19448
rect -7964 19399 -7918 19410
rect -8056 19225 -7964 19399
rect -7964 19214 -7918 19225
rect -7780 19399 -7734 19410
rect -7780 19214 -7734 19225
rect -7596 19399 -7550 19410
rect -7412 19399 -7366 19410
rect -7429 19372 -7412 19374
rect -7366 19372 -7349 19374
rect -7429 19252 -7417 19372
rect -7361 19252 -7349 19372
rect -7429 19250 -7412 19252
rect -7596 19214 -7550 19225
rect -7366 19250 -7349 19252
rect -7412 19214 -7366 19225
rect -8102 18997 -8056 19142
rect -7887 19133 -7876 19179
rect -7822 19133 -7811 19179
rect -7887 19100 -7811 19133
rect -7703 19133 -7692 19179
rect -7638 19133 -7627 19179
rect -7703 19100 -7627 19133
rect -7519 19133 -7508 19179
rect -7454 19133 -7443 19179
rect -7519 19100 -7443 19133
rect -7274 18997 -7228 19142
rect -8114 18985 -8034 18997
rect -8114 18929 -8102 18985
rect -8046 18929 -8034 18985
rect -8114 18917 -8034 18929
rect -7296 18985 -7218 18997
rect -7296 18929 -7284 18985
rect -7228 18929 -7218 18985
rect -7296 18917 -7218 18929
rect -6943 18867 -6863 18877
rect -8277 18811 -6931 18867
rect -6875 18811 -6863 18867
rect -6943 18809 -6863 18811
rect -7109 18758 -7039 18760
rect -8277 18757 -7039 18758
rect -8277 18703 -7107 18757
rect -7051 18703 -7039 18757
rect -8277 18702 -7039 18703
rect -8277 17681 -8221 18702
rect -7109 18694 -7039 18702
rect -7613 18650 -7527 18654
rect -7613 18594 -7601 18650
rect -7545 18594 -7527 18650
rect -7613 18582 -7527 18594
rect -8102 18437 -8056 18448
rect -7887 18446 -7811 18479
rect -7887 18400 -7876 18446
rect -7822 18400 -7811 18446
rect -7703 18446 -7627 18479
rect -7703 18400 -7692 18446
rect -7638 18400 -7627 18446
rect -7519 18446 -7443 18479
rect -7519 18400 -7508 18446
rect -7454 18400 -7443 18446
rect -7274 18437 -7228 18448
rect -7964 18354 -7918 18365
rect -7981 18327 -7964 18329
rect -7780 18354 -7734 18365
rect -7918 18327 -7901 18329
rect -8056 18207 -7969 18327
rect -7913 18207 -7901 18327
rect -7981 18205 -7964 18207
rect -8056 17907 -7964 18027
rect -7918 18205 -7901 18207
rect -7797 18027 -7780 18029
rect -7596 18354 -7550 18365
rect -7613 18327 -7596 18329
rect -7412 18354 -7366 18365
rect -7550 18327 -7533 18329
rect -7613 18207 -7601 18327
rect -7545 18207 -7533 18327
rect -7613 18205 -7596 18207
rect -7734 18027 -7717 18029
rect -7797 17907 -7785 18027
rect -7729 17907 -7717 18027
rect -7797 17905 -7780 17907
rect -7964 17869 -7918 17880
rect -7734 17905 -7717 17907
rect -7780 17869 -7734 17880
rect -7550 18205 -7533 18207
rect -7429 18027 -7412 18029
rect -7291 18327 -7274 18329
rect -7228 18327 -7211 18329
rect -7291 18206 -7279 18327
rect -7223 18206 -7211 18327
rect -7291 18204 -7274 18206
rect -7366 18027 -7349 18029
rect -7429 17907 -7417 18027
rect -7361 17907 -7349 18027
rect -7429 17905 -7412 17907
rect -7596 17869 -7550 17880
rect -7366 17905 -7349 17907
rect -7412 17869 -7366 17880
rect -7887 17831 -7876 17834
rect -7822 17831 -7811 17834
rect -7703 17831 -7692 17834
rect -7638 17831 -7627 17834
rect -7519 17831 -7508 17834
rect -7454 17831 -7443 17834
rect -8102 17786 -8056 17797
rect -7889 17775 -7877 17831
rect -7821 17775 -7809 17831
rect -7889 17761 -7809 17775
rect -7705 17775 -7693 17831
rect -7637 17775 -7625 17831
rect -7705 17761 -7625 17775
rect -7521 17775 -7509 17831
rect -7453 17775 -7441 17831
rect -7228 18204 -7211 18206
rect -7274 17786 -7228 17797
rect -7521 17761 -7441 17775
rect -7889 17681 -7809 17683
rect -8277 17625 -7877 17681
rect -7821 17625 -7809 17681
rect -7889 17623 -7809 17625
rect -8697 17565 -8627 17579
rect -7705 17565 -7625 17567
rect -8697 17509 -8685 17565
rect -8629 17509 -7693 17565
rect -7637 17509 -7625 17565
rect -8697 17497 -8627 17509
rect -7705 17507 -7625 17509
rect -7376 17565 -7296 17567
rect -6933 17565 -6873 17577
rect -7376 17509 -7364 17565
rect -7308 17509 -6931 17565
rect -6875 17509 -6873 17565
rect -7376 17507 -7296 17509
rect -6933 17497 -6873 17509
rect -9513 17449 -9443 17461
rect -7521 17449 -7441 17451
rect -9513 17393 -9501 17449
rect -9445 17393 -7509 17449
rect -7453 17393 -7441 17449
rect -9513 17381 -9443 17393
rect -7521 17391 -7441 17393
rect -7889 17299 -7809 17313
rect -8102 17277 -8056 17288
rect -7889 17243 -7877 17299
rect -7821 17243 -7809 17299
rect -7705 17299 -7625 17313
rect -7705 17243 -7693 17299
rect -7637 17243 -7625 17299
rect -7521 17299 -7441 17313
rect -7521 17243 -7509 17299
rect -7453 17243 -7441 17299
rect -7274 17277 -7228 17288
rect -7887 17240 -7876 17243
rect -7822 17240 -7811 17243
rect -7703 17240 -7692 17243
rect -7638 17240 -7627 17243
rect -7519 17240 -7508 17243
rect -7454 17240 -7443 17243
rect -7964 17194 -7918 17205
rect -8056 17020 -7964 17194
rect -7964 17009 -7918 17020
rect -7780 17194 -7734 17205
rect -7780 17009 -7734 17020
rect -7596 17194 -7550 17205
rect -7412 17194 -7366 17205
rect -7429 17167 -7412 17169
rect -7366 17167 -7349 17169
rect -7429 17047 -7417 17167
rect -7361 17047 -7349 17167
rect -7429 17045 -7412 17047
rect -7596 17009 -7550 17020
rect -7366 17045 -7349 17047
rect -7412 17009 -7366 17020
rect -8102 16792 -8056 16937
rect -7887 16928 -7876 16974
rect -7822 16928 -7811 16974
rect -7887 16895 -7811 16928
rect -7703 16928 -7692 16974
rect -7638 16928 -7627 16974
rect -7703 16895 -7627 16928
rect -7519 16928 -7508 16974
rect -7454 16928 -7443 16974
rect -7519 16895 -7443 16928
rect -7274 16792 -7228 16937
rect -8114 16780 -8034 16792
rect -8114 16724 -8102 16780
rect -8046 16724 -8034 16780
rect -8114 16712 -8034 16724
rect -7296 16780 -7216 16792
rect -7296 16724 -7284 16780
rect -7228 16724 -7216 16780
rect -7296 16712 -7216 16724
rect -8969 16662 -8899 16674
rect -8687 16662 -8627 16666
rect -6791 16662 -6735 19599
rect -6035 19597 -5955 19599
rect -4519 19651 -4449 19663
rect -3479 19651 -3399 19653
rect -1993 19652 -1913 19654
rect -4519 19595 -4507 19651
rect -4451 19595 -3467 19651
rect -3411 19595 -3399 19651
rect -4519 19583 -4449 19595
rect -6403 19505 -6323 19519
rect -6616 19483 -6570 19494
rect -6403 19449 -6391 19505
rect -6335 19449 -6323 19505
rect -6219 19505 -6139 19519
rect -6219 19449 -6207 19505
rect -6151 19449 -6139 19505
rect -6035 19505 -5955 19519
rect -6035 19449 -6023 19505
rect -5967 19449 -5955 19505
rect -5788 19483 -5742 19494
rect -6401 19446 -6390 19449
rect -6336 19446 -6325 19449
rect -6217 19446 -6206 19449
rect -6152 19446 -6141 19449
rect -6033 19446 -6022 19449
rect -5968 19446 -5957 19449
rect -6478 19400 -6432 19411
rect -6570 19226 -6478 19400
rect -6478 19215 -6432 19226
rect -6294 19400 -6248 19411
rect -6294 19215 -6248 19226
rect -6110 19400 -6064 19411
rect -5926 19400 -5880 19411
rect -5943 19373 -5926 19375
rect -5880 19373 -5863 19375
rect -5943 19253 -5931 19373
rect -5875 19253 -5863 19373
rect -5943 19251 -5926 19253
rect -6110 19215 -6064 19226
rect -5880 19251 -5863 19253
rect -5926 19215 -5880 19226
rect -6616 18998 -6570 19143
rect -6401 19134 -6390 19180
rect -6336 19134 -6325 19180
rect -6401 19101 -6325 19134
rect -6217 19134 -6206 19180
rect -6152 19134 -6141 19180
rect -6217 19101 -6141 19134
rect -6033 19134 -6022 19180
rect -5968 19134 -5957 19180
rect -6033 19101 -5957 19134
rect -5788 18998 -5742 19143
rect -6628 18986 -6548 18998
rect -6628 18930 -6616 18986
rect -6560 18930 -6548 18986
rect -6628 18918 -6548 18930
rect -5810 18986 -5732 18998
rect -5810 18930 -5798 18986
rect -5742 18930 -5732 18986
rect -5810 18918 -5732 18930
rect -4235 18864 -4179 19595
rect -3479 19593 -3399 19595
rect -2749 19596 -1981 19652
rect -1925 19596 -1913 19652
rect -3847 19501 -3767 19515
rect -4060 19479 -4014 19490
rect -3847 19445 -3835 19501
rect -3779 19445 -3767 19501
rect -3663 19501 -3583 19515
rect -3663 19445 -3651 19501
rect -3595 19445 -3583 19501
rect -3479 19501 -3399 19515
rect -3479 19445 -3467 19501
rect -3411 19445 -3399 19501
rect -3232 19479 -3186 19490
rect -3845 19442 -3834 19445
rect -3780 19442 -3769 19445
rect -3661 19442 -3650 19445
rect -3596 19442 -3585 19445
rect -3477 19442 -3466 19445
rect -3412 19442 -3401 19445
rect -3922 19396 -3876 19407
rect -4014 19222 -3922 19396
rect -3922 19211 -3876 19222
rect -3738 19396 -3692 19407
rect -3738 19211 -3692 19222
rect -3554 19396 -3508 19407
rect -3370 19396 -3324 19407
rect -3387 19369 -3370 19371
rect -3324 19369 -3307 19371
rect -3387 19249 -3375 19369
rect -3319 19249 -3307 19369
rect -3387 19247 -3370 19249
rect -3554 19211 -3508 19222
rect -3324 19247 -3307 19249
rect -3370 19211 -3324 19222
rect -4060 18994 -4014 19139
rect -3845 19130 -3834 19176
rect -3780 19130 -3769 19176
rect -3845 19097 -3769 19130
rect -3661 19130 -3650 19176
rect -3596 19130 -3585 19176
rect -3661 19097 -3585 19130
rect -3477 19130 -3466 19176
rect -3412 19130 -3401 19176
rect -3477 19097 -3401 19130
rect -3232 18994 -3186 19139
rect -4072 18982 -3992 18994
rect -4072 18926 -4060 18982
rect -4004 18926 -3992 18982
rect -4072 18914 -3992 18926
rect -3254 18982 -3176 18994
rect -3254 18926 -3242 18982
rect -3186 18926 -3176 18982
rect -3254 18914 -3176 18926
rect -2901 18864 -2821 18874
rect -4235 18808 -2889 18864
rect -2833 18808 -2821 18864
rect -2901 18806 -2821 18808
rect -3067 18755 -2997 18757
rect -4235 18754 -2997 18755
rect -4235 18700 -3065 18754
rect -3009 18700 -2997 18754
rect -4235 18699 -2997 18700
rect -4235 17678 -4179 18699
rect -3067 18691 -2997 18699
rect -3571 18647 -3485 18651
rect -3571 18591 -3559 18647
rect -3503 18591 -3485 18647
rect -3571 18579 -3485 18591
rect -4060 18434 -4014 18445
rect -3845 18443 -3769 18476
rect -3845 18397 -3834 18443
rect -3780 18397 -3769 18443
rect -3661 18443 -3585 18476
rect -3661 18397 -3650 18443
rect -3596 18397 -3585 18443
rect -3477 18443 -3401 18476
rect -3477 18397 -3466 18443
rect -3412 18397 -3401 18443
rect -3232 18434 -3186 18445
rect -3922 18351 -3876 18362
rect -3939 18324 -3922 18326
rect -3738 18351 -3692 18362
rect -3876 18324 -3859 18326
rect -4014 18204 -3927 18324
rect -3871 18204 -3859 18324
rect -3939 18202 -3922 18204
rect -4014 17904 -3922 18024
rect -3876 18202 -3859 18204
rect -3755 18024 -3738 18026
rect -3554 18351 -3508 18362
rect -3571 18324 -3554 18326
rect -3370 18351 -3324 18362
rect -3508 18324 -3491 18326
rect -3571 18204 -3559 18324
rect -3503 18204 -3491 18324
rect -3571 18202 -3554 18204
rect -3692 18024 -3675 18026
rect -3755 17904 -3743 18024
rect -3687 17904 -3675 18024
rect -3755 17902 -3738 17904
rect -3922 17866 -3876 17877
rect -3692 17902 -3675 17904
rect -3738 17866 -3692 17877
rect -3508 18202 -3491 18204
rect -3387 18024 -3370 18026
rect -3249 18324 -3232 18326
rect -3186 18324 -3169 18326
rect -3249 18203 -3237 18324
rect -3181 18203 -3169 18324
rect -3249 18201 -3232 18203
rect -3324 18024 -3307 18026
rect -3387 17904 -3375 18024
rect -3319 17904 -3307 18024
rect -3387 17902 -3370 17904
rect -3554 17866 -3508 17877
rect -3324 17902 -3307 17904
rect -3370 17866 -3324 17877
rect -3845 17828 -3834 17831
rect -3780 17828 -3769 17831
rect -3661 17828 -3650 17831
rect -3596 17828 -3585 17831
rect -3477 17828 -3466 17831
rect -3412 17828 -3401 17831
rect -4060 17783 -4014 17794
rect -3847 17772 -3835 17828
rect -3779 17772 -3767 17828
rect -3847 17758 -3767 17772
rect -3663 17772 -3651 17828
rect -3595 17772 -3583 17828
rect -3663 17758 -3583 17772
rect -3479 17772 -3467 17828
rect -3411 17772 -3399 17828
rect -3186 18201 -3169 18203
rect -3232 17783 -3186 17794
rect -3479 17758 -3399 17772
rect -3847 17678 -3767 17680
rect -4235 17622 -3835 17678
rect -3779 17622 -3767 17678
rect -3847 17620 -3767 17622
rect -4655 17562 -4585 17576
rect -3663 17562 -3583 17564
rect -4655 17506 -4643 17562
rect -4587 17506 -3651 17562
rect -3595 17506 -3583 17562
rect -4655 17494 -4585 17506
rect -3663 17504 -3583 17506
rect -3334 17562 -3254 17564
rect -2891 17562 -2831 17574
rect -3334 17506 -3322 17562
rect -3266 17506 -2889 17562
rect -2833 17506 -2831 17562
rect -3334 17504 -3254 17506
rect -2891 17494 -2831 17506
rect -5501 17446 -5431 17458
rect -3479 17446 -3399 17448
rect -5501 17390 -5489 17446
rect -5433 17390 -3467 17446
rect -3411 17390 -3399 17446
rect -5501 17378 -5431 17390
rect -3479 17388 -3399 17390
rect -3847 17296 -3767 17310
rect -4060 17274 -4014 17285
rect -3847 17240 -3835 17296
rect -3779 17240 -3767 17296
rect -3663 17296 -3583 17310
rect -3663 17240 -3651 17296
rect -3595 17240 -3583 17296
rect -3479 17296 -3399 17310
rect -3479 17240 -3467 17296
rect -3411 17240 -3399 17296
rect -3232 17274 -3186 17285
rect -3845 17237 -3834 17240
rect -3780 17237 -3769 17240
rect -3661 17237 -3650 17240
rect -3596 17237 -3585 17240
rect -3477 17237 -3466 17240
rect -3412 17237 -3401 17240
rect -3922 17191 -3876 17202
rect -4014 17017 -3922 17191
rect -3922 17006 -3876 17017
rect -3738 17191 -3692 17202
rect -3738 17006 -3692 17017
rect -3554 17191 -3508 17202
rect -3370 17191 -3324 17202
rect -3387 17164 -3370 17166
rect -3324 17164 -3307 17166
rect -3387 17044 -3375 17164
rect -3319 17044 -3307 17164
rect -3387 17042 -3370 17044
rect -3554 17006 -3508 17017
rect -3324 17042 -3307 17044
rect -3370 17006 -3324 17017
rect -4060 16789 -4014 16934
rect -3845 16925 -3834 16971
rect -3780 16925 -3769 16971
rect -3845 16892 -3769 16925
rect -3661 16925 -3650 16971
rect -3596 16925 -3585 16971
rect -3661 16892 -3585 16925
rect -3477 16925 -3466 16971
rect -3412 16925 -3401 16971
rect -3477 16892 -3401 16925
rect -3232 16789 -3186 16934
rect -4072 16777 -3992 16789
rect -4072 16721 -4060 16777
rect -4004 16721 -3992 16777
rect -4072 16709 -3992 16721
rect -3254 16777 -3174 16789
rect -3254 16721 -3242 16777
rect -3186 16721 -3174 16777
rect -3254 16709 -3174 16721
rect -8969 16606 -8957 16662
rect -8901 16606 -8685 16662
rect -8629 16606 -6735 16662
rect -4957 16659 -4887 16671
rect -4645 16659 -4585 16663
rect -2749 16659 -2693 19596
rect -1993 19594 -1913 19596
rect -477 19651 -407 19663
rect 563 19651 643 19653
rect 2049 19652 2129 19654
rect -477 19595 -465 19651
rect -409 19595 575 19651
rect 631 19595 643 19651
rect -477 19583 -407 19595
rect -2361 19502 -2281 19516
rect -2574 19480 -2528 19491
rect -2361 19446 -2349 19502
rect -2293 19446 -2281 19502
rect -2177 19502 -2097 19516
rect -2177 19446 -2165 19502
rect -2109 19446 -2097 19502
rect -1993 19502 -1913 19516
rect -1993 19446 -1981 19502
rect -1925 19446 -1913 19502
rect -1746 19480 -1700 19491
rect -2359 19443 -2348 19446
rect -2294 19443 -2283 19446
rect -2175 19443 -2164 19446
rect -2110 19443 -2099 19446
rect -1991 19443 -1980 19446
rect -1926 19443 -1915 19446
rect -2436 19397 -2390 19408
rect -2528 19223 -2436 19397
rect -2436 19212 -2390 19223
rect -2252 19397 -2206 19408
rect -2252 19212 -2206 19223
rect -2068 19397 -2022 19408
rect -1884 19397 -1838 19408
rect -1901 19370 -1884 19372
rect -1838 19370 -1821 19372
rect -1901 19250 -1889 19370
rect -1833 19250 -1821 19370
rect -1901 19248 -1884 19250
rect -2068 19212 -2022 19223
rect -1838 19248 -1821 19250
rect -1884 19212 -1838 19223
rect -2574 18995 -2528 19140
rect -2359 19131 -2348 19177
rect -2294 19131 -2283 19177
rect -2359 19098 -2283 19131
rect -2175 19131 -2164 19177
rect -2110 19131 -2099 19177
rect -2175 19098 -2099 19131
rect -1991 19131 -1980 19177
rect -1926 19131 -1915 19177
rect -1991 19098 -1915 19131
rect -1746 18995 -1700 19140
rect -2586 18983 -2506 18995
rect -2586 18927 -2574 18983
rect -2518 18927 -2506 18983
rect -2586 18915 -2506 18927
rect -1768 18983 -1690 18995
rect -1768 18927 -1756 18983
rect -1700 18927 -1690 18983
rect -1768 18915 -1690 18927
rect -193 18864 -137 19595
rect 563 19593 643 19595
rect 1293 19596 2061 19652
rect 2117 19596 2129 19652
rect 195 19501 275 19515
rect -18 19479 28 19490
rect 195 19445 207 19501
rect 263 19445 275 19501
rect 379 19501 459 19515
rect 379 19445 391 19501
rect 447 19445 459 19501
rect 563 19501 643 19515
rect 563 19445 575 19501
rect 631 19445 643 19501
rect 810 19479 856 19490
rect 197 19442 208 19445
rect 262 19442 273 19445
rect 381 19442 392 19445
rect 446 19442 457 19445
rect 565 19442 576 19445
rect 630 19442 641 19445
rect 120 19396 166 19407
rect 28 19222 120 19396
rect 120 19211 166 19222
rect 304 19396 350 19407
rect 304 19211 350 19222
rect 488 19396 534 19407
rect 672 19396 718 19407
rect 655 19369 672 19371
rect 718 19369 735 19371
rect 655 19249 667 19369
rect 723 19249 735 19369
rect 655 19247 672 19249
rect 488 19211 534 19222
rect 718 19247 735 19249
rect 672 19211 718 19222
rect -18 18994 28 19139
rect 197 19130 208 19176
rect 262 19130 273 19176
rect 197 19097 273 19130
rect 381 19130 392 19176
rect 446 19130 457 19176
rect 381 19097 457 19130
rect 565 19130 576 19176
rect 630 19130 641 19176
rect 565 19097 641 19130
rect 810 18994 856 19139
rect -30 18982 50 18994
rect -30 18926 -18 18982
rect 38 18926 50 18982
rect -30 18914 50 18926
rect 788 18982 866 18994
rect 788 18926 800 18982
rect 856 18926 866 18982
rect 788 18914 866 18926
rect 1141 18864 1221 18874
rect -193 18808 1153 18864
rect 1209 18808 1221 18864
rect 1141 18806 1221 18808
rect 975 18755 1045 18757
rect -193 18754 1045 18755
rect -193 18700 977 18754
rect 1033 18700 1045 18754
rect -193 18699 1045 18700
rect -193 17678 -137 18699
rect 975 18691 1045 18699
rect 471 18647 557 18651
rect 471 18591 483 18647
rect 539 18591 557 18647
rect 471 18579 557 18591
rect -18 18434 28 18445
rect 197 18443 273 18476
rect 197 18397 208 18443
rect 262 18397 273 18443
rect 381 18443 457 18476
rect 381 18397 392 18443
rect 446 18397 457 18443
rect 565 18443 641 18476
rect 565 18397 576 18443
rect 630 18397 641 18443
rect 810 18434 856 18445
rect 120 18351 166 18362
rect 103 18324 120 18326
rect 304 18351 350 18362
rect 166 18324 183 18326
rect 28 18204 115 18324
rect 171 18204 183 18324
rect 103 18202 120 18204
rect 28 17904 120 18024
rect 166 18202 183 18204
rect 287 18024 304 18026
rect 488 18351 534 18362
rect 471 18324 488 18326
rect 672 18351 718 18362
rect 534 18324 551 18326
rect 471 18204 483 18324
rect 539 18204 551 18324
rect 471 18202 488 18204
rect 350 18024 367 18026
rect 287 17904 299 18024
rect 355 17904 367 18024
rect 287 17902 304 17904
rect 120 17866 166 17877
rect 350 17902 367 17904
rect 304 17866 350 17877
rect 534 18202 551 18204
rect 655 18024 672 18026
rect 793 18324 810 18326
rect 856 18324 873 18326
rect 793 18203 805 18324
rect 861 18203 873 18324
rect 793 18201 810 18203
rect 718 18024 735 18026
rect 655 17904 667 18024
rect 723 17904 735 18024
rect 655 17902 672 17904
rect 488 17866 534 17877
rect 718 17902 735 17904
rect 672 17866 718 17877
rect 197 17828 208 17831
rect 262 17828 273 17831
rect 381 17828 392 17831
rect 446 17828 457 17831
rect 565 17828 576 17831
rect 630 17828 641 17831
rect -18 17783 28 17794
rect 195 17772 207 17828
rect 263 17772 275 17828
rect 195 17758 275 17772
rect 379 17772 391 17828
rect 447 17772 459 17828
rect 379 17758 459 17772
rect 563 17772 575 17828
rect 631 17772 643 17828
rect 856 18201 873 18203
rect 810 17783 856 17794
rect 563 17758 643 17772
rect 195 17678 275 17680
rect -193 17622 207 17678
rect 263 17622 275 17678
rect 195 17620 275 17622
rect -613 17562 -543 17576
rect 379 17562 459 17564
rect -613 17506 -601 17562
rect -545 17506 391 17562
rect 447 17506 459 17562
rect -613 17494 -543 17506
rect 379 17504 459 17506
rect 708 17562 788 17564
rect 1151 17562 1211 17574
rect 708 17506 720 17562
rect 776 17506 1153 17562
rect 1209 17506 1211 17562
rect 708 17504 788 17506
rect 1151 17494 1211 17506
rect -1459 17446 -1389 17458
rect 563 17446 643 17448
rect -1459 17390 -1447 17446
rect -1391 17390 575 17446
rect 631 17390 643 17446
rect -1459 17378 -1389 17390
rect 563 17388 643 17390
rect 195 17296 275 17310
rect -18 17274 28 17285
rect 195 17240 207 17296
rect 263 17240 275 17296
rect 379 17296 459 17310
rect 379 17240 391 17296
rect 447 17240 459 17296
rect 563 17296 643 17310
rect 563 17240 575 17296
rect 631 17240 643 17296
rect 810 17274 856 17285
rect 197 17237 208 17240
rect 262 17237 273 17240
rect 381 17237 392 17240
rect 446 17237 457 17240
rect 565 17237 576 17240
rect 630 17237 641 17240
rect 120 17191 166 17202
rect 28 17017 120 17191
rect 120 17006 166 17017
rect 304 17191 350 17202
rect 304 17006 350 17017
rect 488 17191 534 17202
rect 672 17191 718 17202
rect 655 17164 672 17166
rect 718 17164 735 17166
rect 655 17044 667 17164
rect 723 17044 735 17164
rect 655 17042 672 17044
rect 488 17006 534 17017
rect 718 17042 735 17044
rect 672 17006 718 17017
rect -18 16789 28 16934
rect 197 16925 208 16971
rect 262 16925 273 16971
rect 197 16892 273 16925
rect 381 16925 392 16971
rect 446 16925 457 16971
rect 381 16892 457 16925
rect 565 16925 576 16971
rect 630 16925 641 16971
rect 565 16892 641 16925
rect 810 16789 856 16934
rect -30 16777 50 16789
rect -30 16721 -18 16777
rect 38 16721 50 16777
rect -30 16709 50 16721
rect 788 16777 868 16789
rect 788 16721 800 16777
rect 856 16721 868 16777
rect 788 16709 868 16721
rect -8969 16604 -8899 16606
rect -8687 16594 -8627 16606
rect -4957 16603 -4945 16659
rect -4889 16603 -4643 16659
rect -4587 16603 -2693 16659
rect -915 16659 -845 16671
rect -603 16659 -543 16663
rect 1293 16659 1349 19596
rect 2049 19594 2129 19596
rect 3565 19651 3635 19663
rect 4605 19651 4685 19653
rect 6091 19652 6171 19654
rect 3565 19595 3577 19651
rect 3633 19595 4617 19651
rect 4673 19595 4685 19651
rect 3565 19583 3635 19595
rect 1681 19502 1761 19516
rect 1468 19480 1514 19491
rect 1681 19446 1693 19502
rect 1749 19446 1761 19502
rect 1865 19502 1945 19516
rect 1865 19446 1877 19502
rect 1933 19446 1945 19502
rect 2049 19502 2129 19516
rect 2049 19446 2061 19502
rect 2117 19446 2129 19502
rect 2296 19480 2342 19491
rect 1683 19443 1694 19446
rect 1748 19443 1759 19446
rect 1867 19443 1878 19446
rect 1932 19443 1943 19446
rect 2051 19443 2062 19446
rect 2116 19443 2127 19446
rect 1606 19397 1652 19408
rect 1514 19223 1606 19397
rect 1606 19212 1652 19223
rect 1790 19397 1836 19408
rect 1790 19212 1836 19223
rect 1974 19397 2020 19408
rect 2158 19397 2204 19408
rect 2141 19370 2158 19372
rect 2204 19370 2221 19372
rect 2141 19250 2153 19370
rect 2209 19250 2221 19370
rect 2141 19248 2158 19250
rect 1974 19212 2020 19223
rect 2204 19248 2221 19250
rect 2158 19212 2204 19223
rect 1468 18995 1514 19140
rect 1683 19131 1694 19177
rect 1748 19131 1759 19177
rect 1683 19098 1759 19131
rect 1867 19131 1878 19177
rect 1932 19131 1943 19177
rect 1867 19098 1943 19131
rect 2051 19131 2062 19177
rect 2116 19131 2127 19177
rect 2051 19098 2127 19131
rect 2296 18995 2342 19140
rect 1456 18983 1536 18995
rect 1456 18927 1468 18983
rect 1524 18927 1536 18983
rect 1456 18915 1536 18927
rect 2274 18983 2352 18995
rect 2274 18927 2286 18983
rect 2342 18927 2352 18983
rect 2274 18915 2352 18927
rect 3849 18864 3905 19595
rect 4605 19593 4685 19595
rect 5335 19596 6103 19652
rect 6159 19596 6171 19652
rect 4237 19501 4317 19515
rect 4024 19479 4070 19490
rect 4237 19445 4249 19501
rect 4305 19445 4317 19501
rect 4421 19501 4501 19515
rect 4421 19445 4433 19501
rect 4489 19445 4501 19501
rect 4605 19501 4685 19515
rect 4605 19445 4617 19501
rect 4673 19445 4685 19501
rect 4852 19479 4898 19490
rect 4239 19442 4250 19445
rect 4304 19442 4315 19445
rect 4423 19442 4434 19445
rect 4488 19442 4499 19445
rect 4607 19442 4618 19445
rect 4672 19442 4683 19445
rect 4162 19396 4208 19407
rect 4070 19222 4162 19396
rect 4162 19211 4208 19222
rect 4346 19396 4392 19407
rect 4346 19211 4392 19222
rect 4530 19396 4576 19407
rect 4714 19396 4760 19407
rect 4697 19369 4714 19371
rect 4760 19369 4777 19371
rect 4697 19249 4709 19369
rect 4765 19249 4777 19369
rect 4697 19247 4714 19249
rect 4530 19211 4576 19222
rect 4760 19247 4777 19249
rect 4714 19211 4760 19222
rect 4024 18994 4070 19139
rect 4239 19130 4250 19176
rect 4304 19130 4315 19176
rect 4239 19097 4315 19130
rect 4423 19130 4434 19176
rect 4488 19130 4499 19176
rect 4423 19097 4499 19130
rect 4607 19130 4618 19176
rect 4672 19130 4683 19176
rect 4607 19097 4683 19130
rect 4852 18994 4898 19139
rect 4012 18982 4092 18994
rect 4012 18926 4024 18982
rect 4080 18926 4092 18982
rect 4012 18914 4092 18926
rect 4830 18982 4908 18994
rect 4830 18926 4842 18982
rect 4898 18926 4908 18982
rect 4830 18914 4908 18926
rect 5183 18864 5263 18874
rect 3849 18808 5195 18864
rect 5251 18808 5263 18864
rect 5183 18806 5263 18808
rect 5017 18755 5087 18757
rect 3849 18754 5087 18755
rect 3849 18700 5019 18754
rect 5075 18700 5087 18754
rect 3849 18699 5087 18700
rect 3849 17678 3905 18699
rect 5017 18691 5087 18699
rect 4513 18647 4599 18651
rect 4513 18591 4525 18647
rect 4581 18591 4599 18647
rect 4513 18579 4599 18591
rect 4024 18434 4070 18445
rect 4239 18443 4315 18476
rect 4239 18397 4250 18443
rect 4304 18397 4315 18443
rect 4423 18443 4499 18476
rect 4423 18397 4434 18443
rect 4488 18397 4499 18443
rect 4607 18443 4683 18476
rect 4607 18397 4618 18443
rect 4672 18397 4683 18443
rect 4852 18434 4898 18445
rect 4162 18351 4208 18362
rect 4145 18324 4162 18326
rect 4346 18351 4392 18362
rect 4208 18324 4225 18326
rect 4070 18204 4157 18324
rect 4213 18204 4225 18324
rect 4145 18202 4162 18204
rect 4070 17904 4162 18024
rect 4208 18202 4225 18204
rect 4329 18024 4346 18026
rect 4530 18351 4576 18362
rect 4513 18324 4530 18326
rect 4714 18351 4760 18362
rect 4576 18324 4593 18326
rect 4513 18204 4525 18324
rect 4581 18204 4593 18324
rect 4513 18202 4530 18204
rect 4392 18024 4409 18026
rect 4329 17904 4341 18024
rect 4397 17904 4409 18024
rect 4329 17902 4346 17904
rect 4162 17866 4208 17877
rect 4392 17902 4409 17904
rect 4346 17866 4392 17877
rect 4576 18202 4593 18204
rect 4697 18024 4714 18026
rect 4835 18324 4852 18326
rect 4898 18324 4915 18326
rect 4835 18203 4847 18324
rect 4903 18203 4915 18324
rect 4835 18201 4852 18203
rect 4760 18024 4777 18026
rect 4697 17904 4709 18024
rect 4765 17904 4777 18024
rect 4697 17902 4714 17904
rect 4530 17866 4576 17877
rect 4760 17902 4777 17904
rect 4714 17866 4760 17877
rect 4239 17828 4250 17831
rect 4304 17828 4315 17831
rect 4423 17828 4434 17831
rect 4488 17828 4499 17831
rect 4607 17828 4618 17831
rect 4672 17828 4683 17831
rect 4024 17783 4070 17794
rect 4237 17772 4249 17828
rect 4305 17772 4317 17828
rect 4237 17758 4317 17772
rect 4421 17772 4433 17828
rect 4489 17772 4501 17828
rect 4421 17758 4501 17772
rect 4605 17772 4617 17828
rect 4673 17772 4685 17828
rect 4898 18201 4915 18203
rect 4852 17783 4898 17794
rect 4605 17758 4685 17772
rect 4237 17678 4317 17680
rect 3849 17622 4249 17678
rect 4305 17622 4317 17678
rect 4237 17620 4317 17622
rect 3429 17562 3499 17576
rect 4421 17562 4501 17564
rect 3429 17506 3441 17562
rect 3497 17506 4433 17562
rect 4489 17506 4501 17562
rect 3429 17494 3499 17506
rect 4421 17504 4501 17506
rect 4750 17562 4830 17564
rect 5193 17562 5253 17574
rect 4750 17506 4762 17562
rect 4818 17506 5195 17562
rect 5251 17506 5253 17562
rect 4750 17504 4830 17506
rect 5193 17494 5253 17506
rect 2583 17446 2653 17458
rect 4605 17446 4685 17448
rect 2583 17390 2595 17446
rect 2651 17390 4617 17446
rect 4673 17390 4685 17446
rect 2583 17378 2653 17390
rect 4605 17388 4685 17390
rect 4237 17296 4317 17310
rect 4024 17274 4070 17285
rect 4237 17240 4249 17296
rect 4305 17240 4317 17296
rect 4421 17296 4501 17310
rect 4421 17240 4433 17296
rect 4489 17240 4501 17296
rect 4605 17296 4685 17310
rect 4605 17240 4617 17296
rect 4673 17240 4685 17296
rect 4852 17274 4898 17285
rect 4239 17237 4250 17240
rect 4304 17237 4315 17240
rect 4423 17237 4434 17240
rect 4488 17237 4499 17240
rect 4607 17237 4618 17240
rect 4672 17237 4683 17240
rect 4162 17191 4208 17202
rect 4070 17017 4162 17191
rect 4162 17006 4208 17017
rect 4346 17191 4392 17202
rect 4346 17006 4392 17017
rect 4530 17191 4576 17202
rect 4714 17191 4760 17202
rect 4697 17164 4714 17166
rect 4760 17164 4777 17166
rect 4697 17044 4709 17164
rect 4765 17044 4777 17164
rect 4697 17042 4714 17044
rect 4530 17006 4576 17017
rect 4760 17042 4777 17044
rect 4714 17006 4760 17017
rect 4024 16789 4070 16934
rect 4239 16925 4250 16971
rect 4304 16925 4315 16971
rect 4239 16892 4315 16925
rect 4423 16925 4434 16971
rect 4488 16925 4499 16971
rect 4423 16892 4499 16925
rect 4607 16925 4618 16971
rect 4672 16925 4683 16971
rect 4607 16892 4683 16925
rect 4852 16789 4898 16934
rect 4012 16777 4092 16789
rect 4012 16721 4024 16777
rect 4080 16721 4092 16777
rect 4012 16709 4092 16721
rect 4830 16777 4910 16789
rect 4830 16721 4842 16777
rect 4898 16721 4910 16777
rect 4830 16709 4910 16721
rect -915 16603 -903 16659
rect -847 16603 -601 16659
rect -545 16603 1349 16659
rect 3127 16659 3197 16671
rect 3439 16659 3499 16663
rect 5335 16659 5391 19596
rect 6091 19594 6171 19596
rect 7607 19651 7677 19663
rect 8647 19651 8727 19653
rect 10133 19652 10213 19654
rect 7607 19595 7619 19651
rect 7675 19595 8659 19651
rect 8715 19595 8727 19651
rect 7607 19583 7677 19595
rect 5723 19502 5803 19516
rect 5510 19480 5556 19491
rect 5723 19446 5735 19502
rect 5791 19446 5803 19502
rect 5907 19502 5987 19516
rect 5907 19446 5919 19502
rect 5975 19446 5987 19502
rect 6091 19502 6171 19516
rect 6091 19446 6103 19502
rect 6159 19446 6171 19502
rect 6338 19480 6384 19491
rect 5725 19443 5736 19446
rect 5790 19443 5801 19446
rect 5909 19443 5920 19446
rect 5974 19443 5985 19446
rect 6093 19443 6104 19446
rect 6158 19443 6169 19446
rect 5648 19397 5694 19408
rect 5556 19223 5648 19397
rect 5648 19212 5694 19223
rect 5832 19397 5878 19408
rect 5832 19212 5878 19223
rect 6016 19397 6062 19408
rect 6200 19397 6246 19408
rect 6183 19370 6200 19372
rect 6246 19370 6263 19372
rect 6183 19250 6195 19370
rect 6251 19250 6263 19370
rect 6183 19248 6200 19250
rect 6016 19212 6062 19223
rect 6246 19248 6263 19250
rect 6200 19212 6246 19223
rect 5510 18995 5556 19140
rect 5725 19131 5736 19177
rect 5790 19131 5801 19177
rect 5725 19098 5801 19131
rect 5909 19131 5920 19177
rect 5974 19131 5985 19177
rect 5909 19098 5985 19131
rect 6093 19131 6104 19177
rect 6158 19131 6169 19177
rect 6093 19098 6169 19131
rect 6338 18995 6384 19140
rect 5498 18983 5578 18995
rect 5498 18927 5510 18983
rect 5566 18927 5578 18983
rect 5498 18915 5578 18927
rect 6316 18983 6394 18995
rect 6316 18927 6328 18983
rect 6384 18927 6394 18983
rect 6316 18915 6394 18927
rect 7891 18864 7947 19595
rect 8647 19593 8727 19595
rect 9377 19596 10145 19652
rect 10201 19596 10213 19652
rect 8279 19501 8359 19515
rect 8066 19479 8112 19490
rect 8279 19445 8291 19501
rect 8347 19445 8359 19501
rect 8463 19501 8543 19515
rect 8463 19445 8475 19501
rect 8531 19445 8543 19501
rect 8647 19501 8727 19515
rect 8647 19445 8659 19501
rect 8715 19445 8727 19501
rect 8894 19479 8940 19490
rect 8281 19442 8292 19445
rect 8346 19442 8357 19445
rect 8465 19442 8476 19445
rect 8530 19442 8541 19445
rect 8649 19442 8660 19445
rect 8714 19442 8725 19445
rect 8204 19396 8250 19407
rect 8112 19222 8204 19396
rect 8204 19211 8250 19222
rect 8388 19396 8434 19407
rect 8388 19211 8434 19222
rect 8572 19396 8618 19407
rect 8756 19396 8802 19407
rect 8739 19369 8756 19371
rect 8802 19369 8819 19371
rect 8739 19249 8751 19369
rect 8807 19249 8819 19369
rect 8739 19247 8756 19249
rect 8572 19211 8618 19222
rect 8802 19247 8819 19249
rect 8756 19211 8802 19222
rect 8066 18994 8112 19139
rect 8281 19130 8292 19176
rect 8346 19130 8357 19176
rect 8281 19097 8357 19130
rect 8465 19130 8476 19176
rect 8530 19130 8541 19176
rect 8465 19097 8541 19130
rect 8649 19130 8660 19176
rect 8714 19130 8725 19176
rect 8649 19097 8725 19130
rect 8894 18994 8940 19139
rect 8054 18982 8134 18994
rect 8054 18926 8066 18982
rect 8122 18926 8134 18982
rect 8054 18914 8134 18926
rect 8872 18982 8950 18994
rect 8872 18926 8884 18982
rect 8940 18926 8950 18982
rect 8872 18914 8950 18926
rect 9225 18864 9305 18874
rect 7891 18808 9237 18864
rect 9293 18808 9305 18864
rect 9225 18806 9305 18808
rect 9059 18755 9129 18757
rect 7891 18754 9129 18755
rect 7891 18700 9061 18754
rect 9117 18700 9129 18754
rect 7891 18699 9129 18700
rect 7891 17678 7947 18699
rect 9059 18691 9129 18699
rect 8555 18647 8641 18651
rect 8555 18591 8567 18647
rect 8623 18591 8641 18647
rect 8555 18579 8641 18591
rect 8066 18434 8112 18445
rect 8281 18443 8357 18476
rect 8281 18397 8292 18443
rect 8346 18397 8357 18443
rect 8465 18443 8541 18476
rect 8465 18397 8476 18443
rect 8530 18397 8541 18443
rect 8649 18443 8725 18476
rect 8649 18397 8660 18443
rect 8714 18397 8725 18443
rect 8894 18434 8940 18445
rect 8204 18351 8250 18362
rect 8187 18324 8204 18326
rect 8388 18351 8434 18362
rect 8250 18324 8267 18326
rect 8112 18204 8199 18324
rect 8255 18204 8267 18324
rect 8187 18202 8204 18204
rect 8112 17904 8204 18024
rect 8250 18202 8267 18204
rect 8371 18024 8388 18026
rect 8572 18351 8618 18362
rect 8555 18324 8572 18326
rect 8756 18351 8802 18362
rect 8618 18324 8635 18326
rect 8555 18204 8567 18324
rect 8623 18204 8635 18324
rect 8555 18202 8572 18204
rect 8434 18024 8451 18026
rect 8371 17904 8383 18024
rect 8439 17904 8451 18024
rect 8371 17902 8388 17904
rect 8204 17866 8250 17877
rect 8434 17902 8451 17904
rect 8388 17866 8434 17877
rect 8618 18202 8635 18204
rect 8739 18024 8756 18026
rect 8877 18324 8894 18326
rect 8940 18324 8957 18326
rect 8877 18203 8889 18324
rect 8945 18203 8957 18324
rect 8877 18201 8894 18203
rect 8802 18024 8819 18026
rect 8739 17904 8751 18024
rect 8807 17904 8819 18024
rect 8739 17902 8756 17904
rect 8572 17866 8618 17877
rect 8802 17902 8819 17904
rect 8756 17866 8802 17877
rect 8281 17828 8292 17831
rect 8346 17828 8357 17831
rect 8465 17828 8476 17831
rect 8530 17828 8541 17831
rect 8649 17828 8660 17831
rect 8714 17828 8725 17831
rect 8066 17783 8112 17794
rect 8279 17772 8291 17828
rect 8347 17772 8359 17828
rect 8279 17758 8359 17772
rect 8463 17772 8475 17828
rect 8531 17772 8543 17828
rect 8463 17758 8543 17772
rect 8647 17772 8659 17828
rect 8715 17772 8727 17828
rect 8940 18201 8957 18203
rect 8894 17783 8940 17794
rect 8647 17758 8727 17772
rect 8279 17678 8359 17680
rect 7891 17622 8291 17678
rect 8347 17622 8359 17678
rect 8279 17620 8359 17622
rect 7471 17562 7541 17576
rect 8463 17562 8543 17564
rect 7471 17506 7483 17562
rect 7539 17506 8475 17562
rect 8531 17506 8543 17562
rect 7471 17494 7541 17506
rect 8463 17504 8543 17506
rect 8792 17562 8872 17564
rect 9235 17562 9295 17574
rect 8792 17506 8804 17562
rect 8860 17506 9237 17562
rect 9293 17506 9295 17562
rect 8792 17504 8872 17506
rect 9235 17494 9295 17506
rect 6625 17446 6695 17458
rect 8647 17446 8727 17448
rect 6625 17390 6637 17446
rect 6693 17390 8659 17446
rect 8715 17390 8727 17446
rect 6625 17378 6695 17390
rect 8647 17388 8727 17390
rect 8279 17296 8359 17310
rect 8066 17274 8112 17285
rect 8279 17240 8291 17296
rect 8347 17240 8359 17296
rect 8463 17296 8543 17310
rect 8463 17240 8475 17296
rect 8531 17240 8543 17296
rect 8647 17296 8727 17310
rect 8647 17240 8659 17296
rect 8715 17240 8727 17296
rect 8894 17274 8940 17285
rect 8281 17237 8292 17240
rect 8346 17237 8357 17240
rect 8465 17237 8476 17240
rect 8530 17237 8541 17240
rect 8649 17237 8660 17240
rect 8714 17237 8725 17240
rect 8204 17191 8250 17202
rect 8112 17017 8204 17191
rect 8204 17006 8250 17017
rect 8388 17191 8434 17202
rect 8388 17006 8434 17017
rect 8572 17191 8618 17202
rect 8756 17191 8802 17202
rect 8739 17164 8756 17166
rect 8802 17164 8819 17166
rect 8739 17044 8751 17164
rect 8807 17044 8819 17164
rect 8739 17042 8756 17044
rect 8572 17006 8618 17017
rect 8802 17042 8819 17044
rect 8756 17006 8802 17017
rect 8066 16789 8112 16934
rect 8281 16925 8292 16971
rect 8346 16925 8357 16971
rect 8281 16892 8357 16925
rect 8465 16925 8476 16971
rect 8530 16925 8541 16971
rect 8465 16892 8541 16925
rect 8649 16925 8660 16971
rect 8714 16925 8725 16971
rect 8649 16892 8725 16925
rect 8894 16789 8940 16934
rect 8054 16777 8134 16789
rect 8054 16721 8066 16777
rect 8122 16721 8134 16777
rect 8054 16709 8134 16721
rect 8872 16777 8952 16789
rect 8872 16721 8884 16777
rect 8940 16721 8952 16777
rect 8872 16709 8952 16721
rect 3127 16603 3139 16659
rect 3195 16603 3441 16659
rect 3497 16603 5391 16659
rect 7169 16659 7239 16671
rect 7481 16659 7541 16663
rect 9377 16659 9433 19596
rect 10133 19594 10213 19596
rect 11649 19651 11719 19663
rect 12689 19651 12769 19653
rect 14175 19652 14255 19654
rect 11649 19595 11661 19651
rect 11717 19595 12701 19651
rect 12757 19595 12769 19651
rect 11649 19583 11719 19595
rect 9765 19502 9845 19516
rect 9552 19480 9598 19491
rect 9765 19446 9777 19502
rect 9833 19446 9845 19502
rect 9949 19502 10029 19516
rect 9949 19446 9961 19502
rect 10017 19446 10029 19502
rect 10133 19502 10213 19516
rect 10133 19446 10145 19502
rect 10201 19446 10213 19502
rect 10380 19480 10426 19491
rect 9767 19443 9778 19446
rect 9832 19443 9843 19446
rect 9951 19443 9962 19446
rect 10016 19443 10027 19446
rect 10135 19443 10146 19446
rect 10200 19443 10211 19446
rect 9690 19397 9736 19408
rect 9598 19223 9690 19397
rect 9690 19212 9736 19223
rect 9874 19397 9920 19408
rect 9874 19212 9920 19223
rect 10058 19397 10104 19408
rect 10242 19397 10288 19408
rect 10225 19370 10242 19372
rect 10288 19370 10305 19372
rect 10225 19250 10237 19370
rect 10293 19250 10305 19370
rect 10225 19248 10242 19250
rect 10058 19212 10104 19223
rect 10288 19248 10305 19250
rect 10242 19212 10288 19223
rect 9552 18995 9598 19140
rect 9767 19131 9778 19177
rect 9832 19131 9843 19177
rect 9767 19098 9843 19131
rect 9951 19131 9962 19177
rect 10016 19131 10027 19177
rect 9951 19098 10027 19131
rect 10135 19131 10146 19177
rect 10200 19131 10211 19177
rect 10135 19098 10211 19131
rect 10380 18995 10426 19140
rect 9540 18983 9620 18995
rect 9540 18927 9552 18983
rect 9608 18927 9620 18983
rect 9540 18915 9620 18927
rect 10358 18983 10436 18995
rect 10358 18927 10370 18983
rect 10426 18927 10436 18983
rect 10358 18915 10436 18927
rect 11933 18864 11989 19595
rect 12689 19593 12769 19595
rect 13419 19596 14187 19652
rect 14243 19596 14255 19652
rect 12321 19501 12401 19515
rect 12108 19479 12154 19490
rect 12321 19445 12333 19501
rect 12389 19445 12401 19501
rect 12505 19501 12585 19515
rect 12505 19445 12517 19501
rect 12573 19445 12585 19501
rect 12689 19501 12769 19515
rect 12689 19445 12701 19501
rect 12757 19445 12769 19501
rect 12936 19479 12982 19490
rect 12323 19442 12334 19445
rect 12388 19442 12399 19445
rect 12507 19442 12518 19445
rect 12572 19442 12583 19445
rect 12691 19442 12702 19445
rect 12756 19442 12767 19445
rect 12246 19396 12292 19407
rect 12154 19222 12246 19396
rect 12246 19211 12292 19222
rect 12430 19396 12476 19407
rect 12430 19211 12476 19222
rect 12614 19396 12660 19407
rect 12798 19396 12844 19407
rect 12781 19369 12798 19371
rect 12844 19369 12861 19371
rect 12781 19249 12793 19369
rect 12849 19249 12861 19369
rect 12781 19247 12798 19249
rect 12614 19211 12660 19222
rect 12844 19247 12861 19249
rect 12798 19211 12844 19222
rect 12108 18994 12154 19139
rect 12323 19130 12334 19176
rect 12388 19130 12399 19176
rect 12323 19097 12399 19130
rect 12507 19130 12518 19176
rect 12572 19130 12583 19176
rect 12507 19097 12583 19130
rect 12691 19130 12702 19176
rect 12756 19130 12767 19176
rect 12691 19097 12767 19130
rect 12936 18994 12982 19139
rect 12096 18982 12176 18994
rect 12096 18926 12108 18982
rect 12164 18926 12176 18982
rect 12096 18914 12176 18926
rect 12914 18982 12992 18994
rect 12914 18926 12926 18982
rect 12982 18926 12992 18982
rect 12914 18914 12992 18926
rect 13267 18864 13347 18874
rect 11933 18808 13279 18864
rect 13335 18808 13347 18864
rect 13267 18806 13347 18808
rect 13101 18755 13171 18757
rect 11933 18754 13171 18755
rect 11933 18700 13103 18754
rect 13159 18700 13171 18754
rect 11933 18699 13171 18700
rect 11933 17678 11989 18699
rect 13101 18691 13171 18699
rect 12597 18647 12683 18651
rect 12597 18591 12609 18647
rect 12665 18591 12683 18647
rect 12597 18579 12683 18591
rect 12108 18434 12154 18445
rect 12323 18443 12399 18476
rect 12323 18397 12334 18443
rect 12388 18397 12399 18443
rect 12507 18443 12583 18476
rect 12507 18397 12518 18443
rect 12572 18397 12583 18443
rect 12691 18443 12767 18476
rect 12691 18397 12702 18443
rect 12756 18397 12767 18443
rect 12936 18434 12982 18445
rect 12246 18351 12292 18362
rect 12229 18324 12246 18326
rect 12430 18351 12476 18362
rect 12292 18324 12309 18326
rect 12154 18204 12241 18324
rect 12297 18204 12309 18324
rect 12229 18202 12246 18204
rect 12154 17904 12246 18024
rect 12292 18202 12309 18204
rect 12413 18024 12430 18026
rect 12614 18351 12660 18362
rect 12597 18324 12614 18326
rect 12798 18351 12844 18362
rect 12660 18324 12677 18326
rect 12597 18204 12609 18324
rect 12665 18204 12677 18324
rect 12597 18202 12614 18204
rect 12476 18024 12493 18026
rect 12413 17904 12425 18024
rect 12481 17904 12493 18024
rect 12413 17902 12430 17904
rect 12246 17866 12292 17877
rect 12476 17902 12493 17904
rect 12430 17866 12476 17877
rect 12660 18202 12677 18204
rect 12781 18024 12798 18026
rect 12919 18324 12936 18326
rect 12982 18324 12999 18326
rect 12919 18203 12931 18324
rect 12987 18203 12999 18324
rect 12919 18201 12936 18203
rect 12844 18024 12861 18026
rect 12781 17904 12793 18024
rect 12849 17904 12861 18024
rect 12781 17902 12798 17904
rect 12614 17866 12660 17877
rect 12844 17902 12861 17904
rect 12798 17866 12844 17877
rect 12323 17828 12334 17831
rect 12388 17828 12399 17831
rect 12507 17828 12518 17831
rect 12572 17828 12583 17831
rect 12691 17828 12702 17831
rect 12756 17828 12767 17831
rect 12108 17783 12154 17794
rect 12321 17772 12333 17828
rect 12389 17772 12401 17828
rect 12321 17758 12401 17772
rect 12505 17772 12517 17828
rect 12573 17772 12585 17828
rect 12505 17758 12585 17772
rect 12689 17772 12701 17828
rect 12757 17772 12769 17828
rect 12982 18201 12999 18203
rect 12936 17783 12982 17794
rect 12689 17758 12769 17772
rect 12321 17678 12401 17680
rect 11933 17622 12333 17678
rect 12389 17622 12401 17678
rect 12321 17620 12401 17622
rect 11513 17562 11583 17576
rect 12505 17562 12585 17564
rect 11513 17506 11525 17562
rect 11581 17506 12517 17562
rect 12573 17506 12585 17562
rect 11513 17494 11583 17506
rect 12505 17504 12585 17506
rect 12834 17562 12914 17564
rect 13277 17562 13337 17574
rect 12834 17506 12846 17562
rect 12902 17506 13279 17562
rect 13335 17506 13337 17562
rect 12834 17504 12914 17506
rect 13277 17494 13337 17506
rect 10667 17446 10737 17458
rect 12689 17446 12769 17448
rect 10667 17390 10679 17446
rect 10735 17390 12701 17446
rect 12757 17390 12769 17446
rect 10667 17378 10737 17390
rect 12689 17388 12769 17390
rect 12321 17296 12401 17310
rect 12108 17274 12154 17285
rect 12321 17240 12333 17296
rect 12389 17240 12401 17296
rect 12505 17296 12585 17310
rect 12505 17240 12517 17296
rect 12573 17240 12585 17296
rect 12689 17296 12769 17310
rect 12689 17240 12701 17296
rect 12757 17240 12769 17296
rect 12936 17274 12982 17285
rect 12323 17237 12334 17240
rect 12388 17237 12399 17240
rect 12507 17237 12518 17240
rect 12572 17237 12583 17240
rect 12691 17237 12702 17240
rect 12756 17237 12767 17240
rect 12246 17191 12292 17202
rect 12154 17017 12246 17191
rect 12246 17006 12292 17017
rect 12430 17191 12476 17202
rect 12430 17006 12476 17017
rect 12614 17191 12660 17202
rect 12798 17191 12844 17202
rect 12781 17164 12798 17166
rect 12844 17164 12861 17166
rect 12781 17044 12793 17164
rect 12849 17044 12861 17164
rect 12781 17042 12798 17044
rect 12614 17006 12660 17017
rect 12844 17042 12861 17044
rect 12798 17006 12844 17017
rect 12108 16789 12154 16934
rect 12323 16925 12334 16971
rect 12388 16925 12399 16971
rect 12323 16892 12399 16925
rect 12507 16925 12518 16971
rect 12572 16925 12583 16971
rect 12507 16892 12583 16925
rect 12691 16925 12702 16971
rect 12756 16925 12767 16971
rect 12691 16892 12767 16925
rect 12936 16789 12982 16934
rect 12096 16777 12176 16789
rect 12096 16721 12108 16777
rect 12164 16721 12176 16777
rect 12096 16709 12176 16721
rect 12914 16777 12994 16789
rect 12914 16721 12926 16777
rect 12982 16721 12994 16777
rect 12914 16709 12994 16721
rect 7169 16603 7181 16659
rect 7237 16603 7483 16659
rect 7539 16603 9433 16659
rect 11211 16659 11281 16671
rect 11523 16659 11583 16663
rect 13419 16659 13475 19596
rect 14175 19594 14255 19596
rect 15691 19651 15761 19663
rect 16731 19651 16811 19653
rect 18217 19652 18297 19654
rect 15691 19595 15703 19651
rect 15759 19595 16743 19651
rect 16799 19595 16811 19651
rect 15691 19583 15761 19595
rect 13807 19502 13887 19516
rect 13594 19480 13640 19491
rect 13807 19446 13819 19502
rect 13875 19446 13887 19502
rect 13991 19502 14071 19516
rect 13991 19446 14003 19502
rect 14059 19446 14071 19502
rect 14175 19502 14255 19516
rect 14175 19446 14187 19502
rect 14243 19446 14255 19502
rect 14422 19480 14468 19491
rect 13809 19443 13820 19446
rect 13874 19443 13885 19446
rect 13993 19443 14004 19446
rect 14058 19443 14069 19446
rect 14177 19443 14188 19446
rect 14242 19443 14253 19446
rect 13732 19397 13778 19408
rect 13640 19223 13732 19397
rect 13732 19212 13778 19223
rect 13916 19397 13962 19408
rect 13916 19212 13962 19223
rect 14100 19397 14146 19408
rect 14284 19397 14330 19408
rect 14267 19370 14284 19372
rect 14330 19370 14347 19372
rect 14267 19250 14279 19370
rect 14335 19250 14347 19370
rect 14267 19248 14284 19250
rect 14100 19212 14146 19223
rect 14330 19248 14347 19250
rect 14284 19212 14330 19223
rect 13594 18995 13640 19140
rect 13809 19131 13820 19177
rect 13874 19131 13885 19177
rect 13809 19098 13885 19131
rect 13993 19131 14004 19177
rect 14058 19131 14069 19177
rect 13993 19098 14069 19131
rect 14177 19131 14188 19177
rect 14242 19131 14253 19177
rect 14177 19098 14253 19131
rect 14422 18995 14468 19140
rect 13582 18983 13662 18995
rect 13582 18927 13594 18983
rect 13650 18927 13662 18983
rect 13582 18915 13662 18927
rect 14400 18983 14478 18995
rect 14400 18927 14412 18983
rect 14468 18927 14478 18983
rect 14400 18915 14478 18927
rect 15975 18864 16031 19595
rect 16731 19593 16811 19595
rect 17461 19596 18229 19652
rect 18285 19596 18297 19652
rect 16363 19501 16443 19515
rect 16150 19479 16196 19490
rect 16363 19445 16375 19501
rect 16431 19445 16443 19501
rect 16547 19501 16627 19515
rect 16547 19445 16559 19501
rect 16615 19445 16627 19501
rect 16731 19501 16811 19515
rect 16731 19445 16743 19501
rect 16799 19445 16811 19501
rect 16978 19479 17024 19490
rect 16365 19442 16376 19445
rect 16430 19442 16441 19445
rect 16549 19442 16560 19445
rect 16614 19442 16625 19445
rect 16733 19442 16744 19445
rect 16798 19442 16809 19445
rect 16288 19396 16334 19407
rect 16196 19222 16288 19396
rect 16288 19211 16334 19222
rect 16472 19396 16518 19407
rect 16472 19211 16518 19222
rect 16656 19396 16702 19407
rect 16840 19396 16886 19407
rect 16823 19369 16840 19371
rect 16886 19369 16903 19371
rect 16823 19249 16835 19369
rect 16891 19249 16903 19369
rect 16823 19247 16840 19249
rect 16656 19211 16702 19222
rect 16886 19247 16903 19249
rect 16840 19211 16886 19222
rect 16150 18994 16196 19139
rect 16365 19130 16376 19176
rect 16430 19130 16441 19176
rect 16365 19097 16441 19130
rect 16549 19130 16560 19176
rect 16614 19130 16625 19176
rect 16549 19097 16625 19130
rect 16733 19130 16744 19176
rect 16798 19130 16809 19176
rect 16733 19097 16809 19130
rect 16978 18994 17024 19139
rect 16138 18982 16218 18994
rect 16138 18926 16150 18982
rect 16206 18926 16218 18982
rect 16138 18914 16218 18926
rect 16956 18982 17034 18994
rect 16956 18926 16968 18982
rect 17024 18926 17034 18982
rect 16956 18914 17034 18926
rect 17309 18864 17389 18874
rect 15975 18808 17321 18864
rect 17377 18808 17389 18864
rect 17309 18806 17389 18808
rect 17143 18755 17213 18757
rect 15975 18754 17213 18755
rect 15975 18700 17145 18754
rect 17201 18700 17213 18754
rect 15975 18699 17213 18700
rect 15975 17678 16031 18699
rect 17143 18691 17213 18699
rect 16639 18647 16725 18651
rect 16639 18591 16651 18647
rect 16707 18591 16725 18647
rect 16639 18579 16725 18591
rect 16150 18434 16196 18445
rect 16365 18443 16441 18476
rect 16365 18397 16376 18443
rect 16430 18397 16441 18443
rect 16549 18443 16625 18476
rect 16549 18397 16560 18443
rect 16614 18397 16625 18443
rect 16733 18443 16809 18476
rect 16733 18397 16744 18443
rect 16798 18397 16809 18443
rect 16978 18434 17024 18445
rect 16288 18351 16334 18362
rect 16271 18324 16288 18326
rect 16472 18351 16518 18362
rect 16334 18324 16351 18326
rect 16196 18204 16283 18324
rect 16339 18204 16351 18324
rect 16271 18202 16288 18204
rect 16196 17904 16288 18024
rect 16334 18202 16351 18204
rect 16455 18024 16472 18026
rect 16656 18351 16702 18362
rect 16639 18324 16656 18326
rect 16840 18351 16886 18362
rect 16702 18324 16719 18326
rect 16639 18204 16651 18324
rect 16707 18204 16719 18324
rect 16639 18202 16656 18204
rect 16518 18024 16535 18026
rect 16455 17904 16467 18024
rect 16523 17904 16535 18024
rect 16455 17902 16472 17904
rect 16288 17866 16334 17877
rect 16518 17902 16535 17904
rect 16472 17866 16518 17877
rect 16702 18202 16719 18204
rect 16823 18024 16840 18026
rect 16961 18324 16978 18326
rect 17024 18324 17041 18326
rect 16961 18203 16973 18324
rect 17029 18203 17041 18324
rect 16961 18201 16978 18203
rect 16886 18024 16903 18026
rect 16823 17904 16835 18024
rect 16891 17904 16903 18024
rect 16823 17902 16840 17904
rect 16656 17866 16702 17877
rect 16886 17902 16903 17904
rect 16840 17866 16886 17877
rect 16365 17828 16376 17831
rect 16430 17828 16441 17831
rect 16549 17828 16560 17831
rect 16614 17828 16625 17831
rect 16733 17828 16744 17831
rect 16798 17828 16809 17831
rect 16150 17783 16196 17794
rect 16363 17772 16375 17828
rect 16431 17772 16443 17828
rect 16363 17758 16443 17772
rect 16547 17772 16559 17828
rect 16615 17772 16627 17828
rect 16547 17758 16627 17772
rect 16731 17772 16743 17828
rect 16799 17772 16811 17828
rect 17024 18201 17041 18203
rect 16978 17783 17024 17794
rect 16731 17758 16811 17772
rect 16363 17678 16443 17680
rect 15975 17622 16375 17678
rect 16431 17622 16443 17678
rect 16363 17620 16443 17622
rect 15555 17562 15625 17576
rect 16547 17562 16627 17564
rect 15555 17506 15567 17562
rect 15623 17506 16559 17562
rect 16615 17506 16627 17562
rect 15555 17494 15625 17506
rect 16547 17504 16627 17506
rect 16876 17562 16956 17564
rect 17319 17562 17379 17574
rect 16876 17506 16888 17562
rect 16944 17506 17321 17562
rect 17377 17506 17379 17562
rect 16876 17504 16956 17506
rect 17319 17494 17379 17506
rect 15375 17446 15453 17458
rect 16731 17446 16811 17448
rect 15375 17390 15386 17446
rect 15442 17390 16743 17446
rect 16799 17390 16811 17446
rect 15375 17378 15453 17390
rect 16731 17388 16811 17390
rect 16363 17296 16443 17310
rect 16150 17274 16196 17285
rect 16363 17240 16375 17296
rect 16431 17240 16443 17296
rect 16547 17296 16627 17310
rect 16547 17240 16559 17296
rect 16615 17240 16627 17296
rect 16731 17296 16811 17310
rect 16731 17240 16743 17296
rect 16799 17240 16811 17296
rect 16978 17274 17024 17285
rect 16365 17237 16376 17240
rect 16430 17237 16441 17240
rect 16549 17237 16560 17240
rect 16614 17237 16625 17240
rect 16733 17237 16744 17240
rect 16798 17237 16809 17240
rect 16288 17191 16334 17202
rect 16196 17017 16288 17191
rect 16288 17006 16334 17017
rect 16472 17191 16518 17202
rect 16472 17006 16518 17017
rect 16656 17191 16702 17202
rect 16840 17191 16886 17202
rect 16823 17164 16840 17166
rect 16886 17164 16903 17166
rect 16823 17044 16835 17164
rect 16891 17044 16903 17164
rect 16823 17042 16840 17044
rect 16656 17006 16702 17017
rect 16886 17042 16903 17044
rect 16840 17006 16886 17017
rect 16150 16789 16196 16934
rect 16365 16925 16376 16971
rect 16430 16925 16441 16971
rect 16365 16892 16441 16925
rect 16549 16925 16560 16971
rect 16614 16925 16625 16971
rect 16549 16892 16625 16925
rect 16733 16925 16744 16971
rect 16798 16925 16809 16971
rect 16733 16892 16809 16925
rect 16978 16789 17024 16934
rect 16138 16777 16218 16789
rect 16138 16721 16150 16777
rect 16206 16721 16218 16777
rect 16138 16709 16218 16721
rect 16956 16777 17036 16789
rect 16956 16721 16968 16777
rect 17024 16721 17036 16777
rect 16956 16709 17036 16721
rect 11211 16603 11223 16659
rect 11279 16603 11525 16659
rect 11581 16603 13475 16659
rect 15253 16659 15323 16671
rect 15565 16659 15625 16663
rect 17461 16659 17517 19596
rect 18217 19594 18297 19596
rect 17849 19502 17929 19516
rect 17636 19480 17682 19491
rect 17849 19446 17861 19502
rect 17917 19446 17929 19502
rect 18033 19502 18113 19516
rect 18033 19446 18045 19502
rect 18101 19446 18113 19502
rect 18217 19502 18297 19516
rect 18217 19446 18229 19502
rect 18285 19446 18297 19502
rect 18464 19480 18510 19491
rect 17851 19443 17862 19446
rect 17916 19443 17927 19446
rect 18035 19443 18046 19446
rect 18100 19443 18111 19446
rect 18219 19443 18230 19446
rect 18284 19443 18295 19446
rect 17774 19397 17820 19408
rect 17682 19223 17774 19397
rect 17774 19212 17820 19223
rect 17958 19397 18004 19408
rect 17958 19212 18004 19223
rect 18142 19397 18188 19408
rect 18326 19397 18372 19408
rect 18309 19370 18326 19372
rect 18372 19370 18389 19372
rect 18309 19250 18321 19370
rect 18377 19250 18389 19370
rect 18309 19248 18326 19250
rect 18142 19212 18188 19223
rect 18372 19248 18389 19250
rect 18326 19212 18372 19223
rect 17636 18995 17682 19140
rect 17851 19131 17862 19177
rect 17916 19131 17927 19177
rect 17851 19098 17927 19131
rect 18035 19131 18046 19177
rect 18100 19131 18111 19177
rect 18035 19098 18111 19131
rect 18219 19131 18230 19177
rect 18284 19131 18295 19177
rect 18219 19098 18295 19131
rect 18464 18995 18510 19140
rect 17624 18983 17704 18995
rect 17624 18927 17636 18983
rect 17692 18927 17704 18983
rect 17624 18915 17704 18927
rect 18442 18983 18520 18995
rect 18442 18927 18454 18983
rect 18510 18927 18520 18983
rect 18442 18915 18520 18927
rect 15253 16603 15265 16659
rect 15321 16603 15567 16659
rect 15623 16603 17517 16659
rect -4957 16601 -4887 16603
rect -4645 16591 -4585 16603
rect -915 16601 -845 16603
rect -603 16591 -543 16603
rect 3127 16601 3197 16603
rect 3439 16591 3499 16603
rect 7169 16601 7239 16603
rect 7481 16591 7541 16603
rect 11211 16601 11281 16603
rect 11523 16591 11583 16603
rect 15253 16591 15323 16603
rect 15565 16591 15625 16603
rect -12294 15738 -10747 15794
rect -12845 14717 -12775 14729
rect -12294 14717 -12238 15738
rect -11625 15686 -11539 15690
rect -11625 15630 -11613 15686
rect -11557 15630 -11539 15686
rect -11625 15618 -11539 15630
rect -12114 15473 -12068 15484
rect -11899 15482 -11823 15515
rect -11899 15436 -11888 15482
rect -11834 15436 -11823 15482
rect -11715 15482 -11639 15515
rect -11715 15436 -11704 15482
rect -11650 15436 -11639 15482
rect -11531 15482 -11455 15515
rect -11531 15436 -11520 15482
rect -11466 15436 -11455 15482
rect -11286 15473 -11240 15484
rect -11976 15390 -11930 15401
rect -11993 15363 -11976 15365
rect -11792 15390 -11746 15401
rect -11930 15363 -11913 15365
rect -12068 15243 -11981 15363
rect -11925 15243 -11913 15363
rect -11993 15241 -11976 15243
rect -12068 14943 -11976 15063
rect -11930 15241 -11913 15243
rect -11809 15063 -11792 15065
rect -11608 15390 -11562 15401
rect -11625 15363 -11608 15365
rect -11424 15390 -11378 15401
rect -11562 15363 -11545 15365
rect -11625 15243 -11613 15363
rect -11557 15243 -11545 15363
rect -11625 15241 -11608 15243
rect -11746 15063 -11729 15065
rect -11809 14943 -11797 15063
rect -11741 14943 -11729 15063
rect -11809 14941 -11792 14943
rect -11976 14905 -11930 14916
rect -11746 14941 -11729 14943
rect -11792 14905 -11746 14916
rect -11562 15241 -11545 15243
rect -11441 15063 -11424 15065
rect -11303 15363 -11286 15365
rect -11240 15363 -11223 15365
rect -11303 15242 -11291 15363
rect -11235 15242 -11223 15363
rect -11303 15240 -11286 15242
rect -11378 15063 -11361 15065
rect -11441 14943 -11429 15063
rect -11373 14943 -11361 15063
rect -11441 14941 -11424 14943
rect -11608 14905 -11562 14916
rect -11378 14941 -11361 14943
rect -11424 14905 -11378 14916
rect -11899 14867 -11888 14870
rect -11834 14867 -11823 14870
rect -11715 14867 -11704 14870
rect -11650 14867 -11639 14870
rect -11531 14867 -11520 14870
rect -11466 14867 -11455 14870
rect -12114 14822 -12068 14833
rect -11901 14811 -11889 14867
rect -11833 14811 -11821 14867
rect -11901 14797 -11821 14811
rect -11717 14811 -11705 14867
rect -11649 14811 -11637 14867
rect -11717 14797 -11637 14811
rect -11533 14811 -11521 14867
rect -11465 14811 -11453 14867
rect -11240 15240 -11223 15242
rect -11286 14822 -11240 14833
rect -11533 14797 -11453 14811
rect -11901 14717 -11821 14719
rect -12845 14661 -12833 14717
rect -12777 14661 -11889 14717
rect -11833 14661 -11821 14717
rect -12845 14649 -12775 14661
rect -11901 14659 -11821 14661
rect -12573 14601 -12503 14613
rect -11717 14601 -11637 14603
rect -12573 14545 -12561 14601
rect -12505 14545 -11705 14601
rect -11649 14545 -11637 14601
rect -12573 14533 -12503 14545
rect -11717 14543 -11637 14545
rect -11388 14601 -11308 14603
rect -11121 14601 -11051 14613
rect -11388 14545 -11376 14601
rect -11320 14545 -11119 14601
rect -11063 14545 -11051 14601
rect -11388 14543 -11308 14545
rect -11121 14535 -11051 14545
rect -11533 14485 -11453 14487
rect -12289 14429 -11521 14485
rect -11465 14429 -11453 14485
rect -12289 13698 -12233 14429
rect -11533 14427 -11453 14429
rect -11901 14335 -11821 14349
rect -12114 14313 -12068 14324
rect -11901 14279 -11889 14335
rect -11833 14279 -11821 14335
rect -11717 14335 -11637 14349
rect -11717 14279 -11705 14335
rect -11649 14279 -11637 14335
rect -11533 14335 -11453 14349
rect -11533 14279 -11521 14335
rect -11465 14279 -11453 14335
rect -11286 14313 -11240 14324
rect -11899 14276 -11888 14279
rect -11834 14276 -11823 14279
rect -11715 14276 -11704 14279
rect -11650 14276 -11639 14279
rect -11531 14276 -11520 14279
rect -11466 14276 -11455 14279
rect -11976 14230 -11930 14241
rect -12068 14056 -11976 14230
rect -11976 14045 -11930 14056
rect -11792 14230 -11746 14241
rect -11792 14045 -11746 14056
rect -11608 14230 -11562 14241
rect -11424 14230 -11378 14241
rect -11441 14203 -11424 14205
rect -11378 14203 -11361 14205
rect -11441 14083 -11429 14203
rect -11373 14083 -11361 14203
rect -11441 14081 -11424 14083
rect -11608 14045 -11562 14056
rect -11378 14081 -11361 14083
rect -11424 14045 -11378 14056
rect -12114 13828 -12068 13973
rect -11899 13964 -11888 14010
rect -11834 13964 -11823 14010
rect -11899 13931 -11823 13964
rect -11715 13964 -11704 14010
rect -11650 13964 -11639 14010
rect -11715 13931 -11639 13964
rect -11531 13964 -11520 14010
rect -11466 13964 -11455 14010
rect -11531 13931 -11455 13964
rect -11286 13828 -11240 13973
rect -12126 13816 -12046 13828
rect -12126 13760 -12114 13816
rect -12058 13760 -12046 13816
rect -12126 13748 -12046 13760
rect -11308 13816 -11228 13828
rect -11308 13760 -11296 13816
rect -11240 13760 -11228 13816
rect -11308 13748 -11228 13760
rect -10955 13698 -10875 13708
rect -12289 13642 -10943 13698
rect -10887 13642 -10875 13698
rect -10955 13640 -10875 13642
rect -11121 13589 -11051 13591
rect -12289 13588 -11051 13589
rect -12289 13534 -11119 13588
rect -11063 13534 -11051 13588
rect -12289 13533 -11051 13534
rect -12289 12512 -12233 13533
rect -11121 13525 -11051 13533
rect -11625 13481 -11539 13485
rect -11625 13425 -11613 13481
rect -11557 13425 -11539 13481
rect -11625 13413 -11539 13425
rect -12114 13268 -12068 13279
rect -11899 13277 -11823 13310
rect -11899 13231 -11888 13277
rect -11834 13231 -11823 13277
rect -11715 13277 -11639 13310
rect -11715 13231 -11704 13277
rect -11650 13231 -11639 13277
rect -11531 13277 -11455 13310
rect -11531 13231 -11520 13277
rect -11466 13231 -11455 13277
rect -11286 13268 -11240 13279
rect -11976 13185 -11930 13196
rect -11993 13158 -11976 13160
rect -11792 13185 -11746 13196
rect -11930 13158 -11913 13160
rect -12068 13038 -11981 13158
rect -11925 13038 -11913 13158
rect -11993 13036 -11976 13038
rect -12068 12738 -11976 12858
rect -11930 13036 -11913 13038
rect -11809 12858 -11792 12860
rect -11608 13185 -11562 13196
rect -11625 13158 -11608 13160
rect -11424 13185 -11378 13196
rect -11562 13158 -11545 13160
rect -11625 13038 -11613 13158
rect -11557 13038 -11545 13158
rect -11625 13036 -11608 13038
rect -11746 12858 -11729 12860
rect -11809 12738 -11797 12858
rect -11741 12738 -11729 12858
rect -11809 12736 -11792 12738
rect -11976 12700 -11930 12711
rect -11746 12736 -11729 12738
rect -11792 12700 -11746 12711
rect -11562 13036 -11545 13038
rect -11441 12858 -11424 12860
rect -11303 13158 -11286 13160
rect -11240 13158 -11223 13160
rect -11303 13037 -11291 13158
rect -11235 13037 -11223 13158
rect -11303 13035 -11286 13037
rect -11378 12858 -11361 12860
rect -11441 12738 -11429 12858
rect -11373 12738 -11361 12858
rect -11441 12736 -11424 12738
rect -11608 12700 -11562 12711
rect -11378 12736 -11361 12738
rect -11424 12700 -11378 12711
rect -11899 12662 -11888 12665
rect -11834 12662 -11823 12665
rect -11715 12662 -11704 12665
rect -11650 12662 -11639 12665
rect -11531 12662 -11520 12665
rect -11466 12662 -11455 12665
rect -12114 12617 -12068 12628
rect -11901 12606 -11889 12662
rect -11833 12606 -11821 12662
rect -11901 12592 -11821 12606
rect -11717 12606 -11705 12662
rect -11649 12606 -11637 12662
rect -11717 12592 -11637 12606
rect -11533 12606 -11521 12662
rect -11465 12606 -11453 12662
rect -11240 13035 -11223 13037
rect -11286 12617 -11240 12628
rect -11533 12592 -11453 12606
rect -11901 12512 -11821 12514
rect -12289 12456 -11889 12512
rect -11833 12456 -11821 12512
rect -10803 12512 -10747 15738
rect -8282 15738 -6735 15794
rect -8777 14717 -8691 14729
rect -8282 14717 -8226 15738
rect -7613 15686 -7527 15690
rect -7613 15630 -7601 15686
rect -7545 15630 -7527 15686
rect -7613 15618 -7527 15630
rect -8102 15473 -8056 15484
rect -7887 15482 -7811 15515
rect -7887 15436 -7876 15482
rect -7822 15436 -7811 15482
rect -7703 15482 -7627 15515
rect -7703 15436 -7692 15482
rect -7638 15436 -7627 15482
rect -7519 15482 -7443 15515
rect -7519 15436 -7508 15482
rect -7454 15436 -7443 15482
rect -7274 15473 -7228 15484
rect -7964 15390 -7918 15401
rect -7981 15363 -7964 15365
rect -7780 15390 -7734 15401
rect -7918 15363 -7901 15365
rect -8056 15243 -7969 15363
rect -7913 15243 -7901 15363
rect -7981 15241 -7964 15243
rect -8056 14943 -7964 15063
rect -7918 15241 -7901 15243
rect -7797 15063 -7780 15065
rect -7596 15390 -7550 15401
rect -7613 15363 -7596 15365
rect -7412 15390 -7366 15401
rect -7550 15363 -7533 15365
rect -7613 15243 -7601 15363
rect -7545 15243 -7533 15363
rect -7613 15241 -7596 15243
rect -7734 15063 -7717 15065
rect -7797 14943 -7785 15063
rect -7729 14943 -7717 15063
rect -7797 14941 -7780 14943
rect -7964 14905 -7918 14916
rect -7734 14941 -7717 14943
rect -7780 14905 -7734 14916
rect -7550 15241 -7533 15243
rect -7429 15063 -7412 15065
rect -7291 15363 -7274 15365
rect -7228 15363 -7211 15365
rect -7291 15242 -7279 15363
rect -7223 15242 -7211 15363
rect -7291 15240 -7274 15242
rect -7366 15063 -7349 15065
rect -7429 14943 -7417 15063
rect -7361 14943 -7349 15063
rect -7429 14941 -7412 14943
rect -7596 14905 -7550 14916
rect -7366 14941 -7349 14943
rect -7412 14905 -7366 14916
rect -7887 14867 -7876 14870
rect -7822 14867 -7811 14870
rect -7703 14867 -7692 14870
rect -7638 14867 -7627 14870
rect -7519 14867 -7508 14870
rect -7454 14867 -7443 14870
rect -8102 14822 -8056 14833
rect -7889 14811 -7877 14867
rect -7821 14811 -7809 14867
rect -7889 14797 -7809 14811
rect -7705 14811 -7693 14867
rect -7637 14811 -7625 14867
rect -7705 14797 -7625 14811
rect -7521 14811 -7509 14867
rect -7453 14811 -7441 14867
rect -7228 15240 -7211 15242
rect -7274 14822 -7228 14833
rect -7521 14797 -7441 14811
rect -7889 14717 -7809 14719
rect -8777 14661 -8765 14717
rect -8709 14661 -7877 14717
rect -7821 14661 -7809 14717
rect -8777 14649 -8691 14661
rect -7889 14659 -7809 14661
rect -8561 14601 -8491 14613
rect -7705 14601 -7625 14603
rect -8561 14545 -8549 14601
rect -8493 14545 -7693 14601
rect -7637 14545 -7625 14601
rect -8561 14533 -8491 14545
rect -7705 14543 -7625 14545
rect -7376 14601 -7296 14603
rect -7109 14601 -7039 14613
rect -7376 14545 -7364 14601
rect -7308 14545 -7107 14601
rect -7051 14545 -7039 14601
rect -7376 14543 -7296 14545
rect -7109 14535 -7039 14545
rect -7521 14485 -7441 14487
rect -8277 14429 -7509 14485
rect -7453 14429 -7441 14485
rect -8277 13698 -8221 14429
rect -7521 14427 -7441 14429
rect -7889 14335 -7809 14349
rect -8102 14313 -8056 14324
rect -7889 14279 -7877 14335
rect -7821 14279 -7809 14335
rect -7705 14335 -7625 14349
rect -7705 14279 -7693 14335
rect -7637 14279 -7625 14335
rect -7521 14335 -7441 14349
rect -7521 14279 -7509 14335
rect -7453 14279 -7441 14335
rect -7274 14313 -7228 14324
rect -7887 14276 -7876 14279
rect -7822 14276 -7811 14279
rect -7703 14276 -7692 14279
rect -7638 14276 -7627 14279
rect -7519 14276 -7508 14279
rect -7454 14276 -7443 14279
rect -7964 14230 -7918 14241
rect -8056 14056 -7964 14230
rect -7964 14045 -7918 14056
rect -7780 14230 -7734 14241
rect -7780 14045 -7734 14056
rect -7596 14230 -7550 14241
rect -7412 14230 -7366 14241
rect -7429 14203 -7412 14205
rect -7366 14203 -7349 14205
rect -7429 14083 -7417 14203
rect -7361 14083 -7349 14203
rect -7429 14081 -7412 14083
rect -7596 14045 -7550 14056
rect -7366 14081 -7349 14083
rect -7412 14045 -7366 14056
rect -8102 13828 -8056 13973
rect -7887 13964 -7876 14010
rect -7822 13964 -7811 14010
rect -7887 13931 -7811 13964
rect -7703 13964 -7692 14010
rect -7638 13964 -7627 14010
rect -7703 13931 -7627 13964
rect -7519 13964 -7508 14010
rect -7454 13964 -7443 14010
rect -7519 13931 -7443 13964
rect -7274 13828 -7228 13973
rect -8114 13816 -8034 13828
rect -8114 13760 -8102 13816
rect -8046 13760 -8034 13816
rect -8114 13748 -8034 13760
rect -7296 13816 -7216 13828
rect -7296 13760 -7284 13816
rect -7228 13760 -7216 13816
rect -7296 13748 -7216 13760
rect -6943 13698 -6863 13708
rect -8277 13642 -6931 13698
rect -6875 13642 -6863 13698
rect -6943 13640 -6863 13642
rect -7109 13589 -7039 13591
rect -8277 13588 -7039 13589
rect -8277 13534 -7107 13588
rect -7051 13534 -7039 13588
rect -8277 13533 -7039 13534
rect -10139 13481 -10053 13485
rect -10139 13425 -10127 13481
rect -10071 13425 -10053 13481
rect -10139 13413 -10053 13425
rect -10628 13268 -10582 13279
rect -10413 13277 -10337 13310
rect -10413 13231 -10402 13277
rect -10348 13231 -10337 13277
rect -10229 13277 -10153 13310
rect -10229 13231 -10218 13277
rect -10164 13231 -10153 13277
rect -10045 13277 -9969 13310
rect -10045 13231 -10034 13277
rect -9980 13231 -9969 13277
rect -9800 13268 -9754 13279
rect -10490 13185 -10444 13196
rect -10507 13158 -10490 13160
rect -10306 13185 -10260 13196
rect -10444 13158 -10427 13160
rect -10582 13038 -10495 13158
rect -10439 13038 -10427 13158
rect -10507 13036 -10490 13038
rect -10582 12738 -10490 12858
rect -10444 13036 -10427 13038
rect -10323 12858 -10306 12860
rect -10122 13185 -10076 13196
rect -10139 13158 -10122 13160
rect -9938 13185 -9892 13196
rect -10076 13158 -10059 13160
rect -10139 13038 -10127 13158
rect -10071 13038 -10059 13158
rect -10139 13036 -10122 13038
rect -10260 12858 -10243 12860
rect -10323 12738 -10311 12858
rect -10255 12738 -10243 12858
rect -10323 12736 -10306 12738
rect -10490 12700 -10444 12711
rect -10260 12736 -10243 12738
rect -10306 12700 -10260 12711
rect -10076 13036 -10059 13038
rect -9955 12858 -9938 12860
rect -9817 13158 -9800 13160
rect -9754 13158 -9737 13160
rect -9817 13037 -9805 13158
rect -9749 13037 -9737 13158
rect -9817 13035 -9800 13037
rect -9892 12858 -9875 12860
rect -9955 12738 -9943 12858
rect -9887 12738 -9875 12858
rect -9955 12736 -9938 12738
rect -10122 12700 -10076 12711
rect -9892 12736 -9875 12738
rect -9938 12700 -9892 12711
rect -10413 12662 -10402 12665
rect -10348 12662 -10337 12665
rect -10229 12662 -10218 12665
rect -10164 12662 -10153 12665
rect -10045 12662 -10034 12665
rect -9980 12662 -9969 12665
rect -10628 12617 -10582 12628
rect -10415 12606 -10403 12662
rect -10347 12606 -10335 12662
rect -10415 12592 -10335 12606
rect -10231 12606 -10219 12662
rect -10163 12606 -10151 12662
rect -10231 12592 -10151 12606
rect -10047 12606 -10035 12662
rect -9979 12606 -9967 12662
rect -9754 13035 -9737 13037
rect -9800 12617 -9754 12628
rect -10047 12592 -9967 12606
rect -10415 12512 -10335 12514
rect -10803 12456 -10403 12512
rect -10347 12456 -10335 12512
rect -8277 12512 -8221 13533
rect -7109 13525 -7039 13533
rect -7613 13481 -7527 13485
rect -7613 13425 -7601 13481
rect -7545 13425 -7527 13481
rect -7613 13413 -7527 13425
rect -8102 13268 -8056 13279
rect -7887 13277 -7811 13310
rect -7887 13231 -7876 13277
rect -7822 13231 -7811 13277
rect -7703 13277 -7627 13310
rect -7703 13231 -7692 13277
rect -7638 13231 -7627 13277
rect -7519 13277 -7443 13310
rect -7519 13231 -7508 13277
rect -7454 13231 -7443 13277
rect -7274 13268 -7228 13279
rect -7964 13185 -7918 13196
rect -7981 13158 -7964 13160
rect -7780 13185 -7734 13196
rect -7918 13158 -7901 13160
rect -8056 13038 -7969 13158
rect -7913 13038 -7901 13158
rect -7981 13036 -7964 13038
rect -8056 12738 -7964 12858
rect -7918 13036 -7901 13038
rect -7797 12858 -7780 12860
rect -7596 13185 -7550 13196
rect -7613 13158 -7596 13160
rect -7412 13185 -7366 13196
rect -7550 13158 -7533 13160
rect -7613 13038 -7601 13158
rect -7545 13038 -7533 13158
rect -7613 13036 -7596 13038
rect -7734 12858 -7717 12860
rect -7797 12738 -7785 12858
rect -7729 12738 -7717 12858
rect -7797 12736 -7780 12738
rect -7964 12700 -7918 12711
rect -7734 12736 -7717 12738
rect -7780 12700 -7734 12711
rect -7550 13036 -7533 13038
rect -7429 12858 -7412 12860
rect -7291 13158 -7274 13160
rect -7228 13158 -7211 13160
rect -7291 13037 -7279 13158
rect -7223 13037 -7211 13158
rect -7291 13035 -7274 13037
rect -7366 12858 -7349 12860
rect -7429 12738 -7417 12858
rect -7361 12738 -7349 12858
rect -7429 12736 -7412 12738
rect -7596 12700 -7550 12711
rect -7366 12736 -7349 12738
rect -7412 12700 -7366 12711
rect -7887 12662 -7876 12665
rect -7822 12662 -7811 12665
rect -7703 12662 -7692 12665
rect -7638 12662 -7627 12665
rect -7519 12662 -7508 12665
rect -7454 12662 -7443 12665
rect -8102 12617 -8056 12628
rect -7889 12606 -7877 12662
rect -7821 12606 -7809 12662
rect -7889 12592 -7809 12606
rect -7705 12606 -7693 12662
rect -7637 12606 -7625 12662
rect -7705 12592 -7625 12606
rect -7521 12606 -7509 12662
rect -7453 12606 -7441 12662
rect -7228 13035 -7211 13037
rect -7274 12617 -7228 12628
rect -7521 12592 -7441 12606
rect -7889 12512 -7809 12514
rect -8277 12456 -7877 12512
rect -7821 12456 -7809 12512
rect -6791 12512 -6735 15738
rect -4240 15738 -2693 15794
rect -4735 14717 -4649 14729
rect -4240 14717 -4184 15738
rect -3571 15686 -3485 15690
rect -3571 15630 -3559 15686
rect -3503 15630 -3485 15686
rect -3571 15618 -3485 15630
rect -4060 15473 -4014 15484
rect -3845 15482 -3769 15515
rect -3845 15436 -3834 15482
rect -3780 15436 -3769 15482
rect -3661 15482 -3585 15515
rect -3661 15436 -3650 15482
rect -3596 15436 -3585 15482
rect -3477 15482 -3401 15515
rect -3477 15436 -3466 15482
rect -3412 15436 -3401 15482
rect -3232 15473 -3186 15484
rect -3922 15390 -3876 15401
rect -3939 15363 -3922 15365
rect -3738 15390 -3692 15401
rect -3876 15363 -3859 15365
rect -4014 15243 -3927 15363
rect -3871 15243 -3859 15363
rect -3939 15241 -3922 15243
rect -4014 14943 -3922 15063
rect -3876 15241 -3859 15243
rect -3755 15063 -3738 15065
rect -3554 15390 -3508 15401
rect -3571 15363 -3554 15365
rect -3370 15390 -3324 15401
rect -3508 15363 -3491 15365
rect -3571 15243 -3559 15363
rect -3503 15243 -3491 15363
rect -3571 15241 -3554 15243
rect -3692 15063 -3675 15065
rect -3755 14943 -3743 15063
rect -3687 14943 -3675 15063
rect -3755 14941 -3738 14943
rect -3922 14905 -3876 14916
rect -3692 14941 -3675 14943
rect -3738 14905 -3692 14916
rect -3508 15241 -3491 15243
rect -3387 15063 -3370 15065
rect -3249 15363 -3232 15365
rect -3186 15363 -3169 15365
rect -3249 15242 -3237 15363
rect -3181 15242 -3169 15363
rect -3249 15240 -3232 15242
rect -3324 15063 -3307 15065
rect -3387 14943 -3375 15063
rect -3319 14943 -3307 15063
rect -3387 14941 -3370 14943
rect -3554 14905 -3508 14916
rect -3324 14941 -3307 14943
rect -3370 14905 -3324 14916
rect -3845 14867 -3834 14870
rect -3780 14867 -3769 14870
rect -3661 14867 -3650 14870
rect -3596 14867 -3585 14870
rect -3477 14867 -3466 14870
rect -3412 14867 -3401 14870
rect -4060 14822 -4014 14833
rect -3847 14811 -3835 14867
rect -3779 14811 -3767 14867
rect -3847 14797 -3767 14811
rect -3663 14811 -3651 14867
rect -3595 14811 -3583 14867
rect -3663 14797 -3583 14811
rect -3479 14811 -3467 14867
rect -3411 14811 -3399 14867
rect -3186 15240 -3169 15242
rect -3232 14822 -3186 14833
rect -3479 14797 -3399 14811
rect -3847 14717 -3767 14719
rect -4735 14661 -4723 14717
rect -4667 14661 -3835 14717
rect -3779 14661 -3767 14717
rect -4735 14649 -4649 14661
rect -3847 14659 -3767 14661
rect -4519 14601 -4449 14613
rect -3663 14601 -3583 14603
rect -4519 14545 -4507 14601
rect -4451 14545 -3651 14601
rect -3595 14545 -3583 14601
rect -4519 14533 -4449 14545
rect -3663 14543 -3583 14545
rect -3334 14601 -3254 14603
rect -3067 14601 -2997 14613
rect -3334 14545 -3322 14601
rect -3266 14545 -3065 14601
rect -3009 14545 -2997 14601
rect -3334 14543 -3254 14545
rect -3067 14535 -2997 14545
rect -3479 14485 -3399 14487
rect -4235 14429 -3467 14485
rect -3411 14429 -3399 14485
rect -4235 13698 -4179 14429
rect -3479 14427 -3399 14429
rect -3847 14335 -3767 14349
rect -4060 14313 -4014 14324
rect -3847 14279 -3835 14335
rect -3779 14279 -3767 14335
rect -3663 14335 -3583 14349
rect -3663 14279 -3651 14335
rect -3595 14279 -3583 14335
rect -3479 14335 -3399 14349
rect -3479 14279 -3467 14335
rect -3411 14279 -3399 14335
rect -3232 14313 -3186 14324
rect -3845 14276 -3834 14279
rect -3780 14276 -3769 14279
rect -3661 14276 -3650 14279
rect -3596 14276 -3585 14279
rect -3477 14276 -3466 14279
rect -3412 14276 -3401 14279
rect -3922 14230 -3876 14241
rect -4014 14056 -3922 14230
rect -3922 14045 -3876 14056
rect -3738 14230 -3692 14241
rect -3738 14045 -3692 14056
rect -3554 14230 -3508 14241
rect -3370 14230 -3324 14241
rect -3387 14203 -3370 14205
rect -3324 14203 -3307 14205
rect -3387 14083 -3375 14203
rect -3319 14083 -3307 14203
rect -3387 14081 -3370 14083
rect -3554 14045 -3508 14056
rect -3324 14081 -3307 14083
rect -3370 14045 -3324 14056
rect -4060 13828 -4014 13973
rect -3845 13964 -3834 14010
rect -3780 13964 -3769 14010
rect -3845 13931 -3769 13964
rect -3661 13964 -3650 14010
rect -3596 13964 -3585 14010
rect -3661 13931 -3585 13964
rect -3477 13964 -3466 14010
rect -3412 13964 -3401 14010
rect -3477 13931 -3401 13964
rect -3232 13828 -3186 13973
rect -4072 13816 -3992 13828
rect -4072 13760 -4060 13816
rect -4004 13760 -3992 13816
rect -4072 13748 -3992 13760
rect -3254 13816 -3174 13828
rect -3254 13760 -3242 13816
rect -3186 13760 -3174 13816
rect -3254 13748 -3174 13760
rect -2901 13698 -2821 13708
rect -4235 13642 -2889 13698
rect -2833 13642 -2821 13698
rect -2901 13640 -2821 13642
rect -3067 13589 -2997 13591
rect -4235 13588 -2997 13589
rect -4235 13534 -3065 13588
rect -3009 13534 -2997 13588
rect -4235 13533 -2997 13534
rect -6127 13481 -6041 13485
rect -6127 13425 -6115 13481
rect -6059 13425 -6041 13481
rect -6127 13413 -6041 13425
rect -6616 13268 -6570 13279
rect -6401 13277 -6325 13310
rect -6401 13231 -6390 13277
rect -6336 13231 -6325 13277
rect -6217 13277 -6141 13310
rect -6217 13231 -6206 13277
rect -6152 13231 -6141 13277
rect -6033 13277 -5957 13310
rect -6033 13231 -6022 13277
rect -5968 13231 -5957 13277
rect -5788 13268 -5742 13279
rect -6478 13185 -6432 13196
rect -6495 13158 -6478 13160
rect -6294 13185 -6248 13196
rect -6432 13158 -6415 13160
rect -6570 13038 -6483 13158
rect -6427 13038 -6415 13158
rect -6495 13036 -6478 13038
rect -6570 12738 -6478 12858
rect -6432 13036 -6415 13038
rect -6311 12858 -6294 12860
rect -6110 13185 -6064 13196
rect -6127 13158 -6110 13160
rect -5926 13185 -5880 13196
rect -6064 13158 -6047 13160
rect -6127 13038 -6115 13158
rect -6059 13038 -6047 13158
rect -6127 13036 -6110 13038
rect -6248 12858 -6231 12860
rect -6311 12738 -6299 12858
rect -6243 12738 -6231 12858
rect -6311 12736 -6294 12738
rect -6478 12700 -6432 12711
rect -6248 12736 -6231 12738
rect -6294 12700 -6248 12711
rect -6064 13036 -6047 13038
rect -5943 12858 -5926 12860
rect -5805 13158 -5788 13160
rect -5742 13158 -5725 13160
rect -5805 13037 -5793 13158
rect -5737 13037 -5725 13158
rect -5805 13035 -5788 13037
rect -5880 12858 -5863 12860
rect -5943 12738 -5931 12858
rect -5875 12738 -5863 12858
rect -5943 12736 -5926 12738
rect -6110 12700 -6064 12711
rect -5880 12736 -5863 12738
rect -5926 12700 -5880 12711
rect -6401 12662 -6390 12665
rect -6336 12662 -6325 12665
rect -6217 12662 -6206 12665
rect -6152 12662 -6141 12665
rect -6033 12662 -6022 12665
rect -5968 12662 -5957 12665
rect -6616 12617 -6570 12628
rect -6403 12606 -6391 12662
rect -6335 12606 -6323 12662
rect -6403 12592 -6323 12606
rect -6219 12606 -6207 12662
rect -6151 12606 -6139 12662
rect -6219 12592 -6139 12606
rect -6035 12606 -6023 12662
rect -5967 12606 -5955 12662
rect -5742 13035 -5725 13037
rect -5788 12617 -5742 12628
rect -6035 12592 -5955 12606
rect -6403 12512 -6323 12514
rect -6791 12456 -6391 12512
rect -6335 12456 -6323 12512
rect -4235 12512 -4179 13533
rect -3067 13525 -2997 13533
rect -3571 13481 -3485 13485
rect -3571 13425 -3559 13481
rect -3503 13425 -3485 13481
rect -3571 13413 -3485 13425
rect -4060 13268 -4014 13279
rect -3845 13277 -3769 13310
rect -3845 13231 -3834 13277
rect -3780 13231 -3769 13277
rect -3661 13277 -3585 13310
rect -3661 13231 -3650 13277
rect -3596 13231 -3585 13277
rect -3477 13277 -3401 13310
rect -3477 13231 -3466 13277
rect -3412 13231 -3401 13277
rect -3232 13268 -3186 13279
rect -3922 13185 -3876 13196
rect -3939 13158 -3922 13160
rect -3738 13185 -3692 13196
rect -3876 13158 -3859 13160
rect -4014 13038 -3927 13158
rect -3871 13038 -3859 13158
rect -3939 13036 -3922 13038
rect -4014 12738 -3922 12858
rect -3876 13036 -3859 13038
rect -3755 12858 -3738 12860
rect -3554 13185 -3508 13196
rect -3571 13158 -3554 13160
rect -3370 13185 -3324 13196
rect -3508 13158 -3491 13160
rect -3571 13038 -3559 13158
rect -3503 13038 -3491 13158
rect -3571 13036 -3554 13038
rect -3692 12858 -3675 12860
rect -3755 12738 -3743 12858
rect -3687 12738 -3675 12858
rect -3755 12736 -3738 12738
rect -3922 12700 -3876 12711
rect -3692 12736 -3675 12738
rect -3738 12700 -3692 12711
rect -3508 13036 -3491 13038
rect -3387 12858 -3370 12860
rect -3249 13158 -3232 13160
rect -3186 13158 -3169 13160
rect -3249 13037 -3237 13158
rect -3181 13037 -3169 13158
rect -3249 13035 -3232 13037
rect -3324 12858 -3307 12860
rect -3387 12738 -3375 12858
rect -3319 12738 -3307 12858
rect -3387 12736 -3370 12738
rect -3554 12700 -3508 12711
rect -3324 12736 -3307 12738
rect -3370 12700 -3324 12711
rect -3845 12662 -3834 12665
rect -3780 12662 -3769 12665
rect -3661 12662 -3650 12665
rect -3596 12662 -3585 12665
rect -3477 12662 -3466 12665
rect -3412 12662 -3401 12665
rect -4060 12617 -4014 12628
rect -3847 12606 -3835 12662
rect -3779 12606 -3767 12662
rect -3847 12592 -3767 12606
rect -3663 12606 -3651 12662
rect -3595 12606 -3583 12662
rect -3663 12592 -3583 12606
rect -3479 12606 -3467 12662
rect -3411 12606 -3399 12662
rect -3186 13035 -3169 13037
rect -3232 12617 -3186 12628
rect -3479 12592 -3399 12606
rect -3847 12512 -3767 12514
rect -4235 12456 -3835 12512
rect -3779 12456 -3767 12512
rect -2749 12512 -2693 15738
rect -198 15738 1349 15794
rect -693 14717 -607 14729
rect -198 14717 -142 15738
rect 471 15686 557 15690
rect 471 15630 483 15686
rect 539 15630 557 15686
rect 471 15618 557 15630
rect -18 15473 28 15484
rect 197 15482 273 15515
rect 197 15436 208 15482
rect 262 15436 273 15482
rect 381 15482 457 15515
rect 381 15436 392 15482
rect 446 15436 457 15482
rect 565 15482 641 15515
rect 565 15436 576 15482
rect 630 15436 641 15482
rect 810 15473 856 15484
rect 120 15390 166 15401
rect 103 15363 120 15365
rect 304 15390 350 15401
rect 166 15363 183 15365
rect 28 15243 115 15363
rect 171 15243 183 15363
rect 103 15241 120 15243
rect 28 14943 120 15063
rect 166 15241 183 15243
rect 287 15063 304 15065
rect 488 15390 534 15401
rect 471 15363 488 15365
rect 672 15390 718 15401
rect 534 15363 551 15365
rect 471 15243 483 15363
rect 539 15243 551 15363
rect 471 15241 488 15243
rect 350 15063 367 15065
rect 287 14943 299 15063
rect 355 14943 367 15063
rect 287 14941 304 14943
rect 120 14905 166 14916
rect 350 14941 367 14943
rect 304 14905 350 14916
rect 534 15241 551 15243
rect 655 15063 672 15065
rect 793 15363 810 15365
rect 856 15363 873 15365
rect 793 15242 805 15363
rect 861 15242 873 15363
rect 793 15240 810 15242
rect 718 15063 735 15065
rect 655 14943 667 15063
rect 723 14943 735 15063
rect 655 14941 672 14943
rect 488 14905 534 14916
rect 718 14941 735 14943
rect 672 14905 718 14916
rect 197 14867 208 14870
rect 262 14867 273 14870
rect 381 14867 392 14870
rect 446 14867 457 14870
rect 565 14867 576 14870
rect 630 14867 641 14870
rect -18 14822 28 14833
rect 195 14811 207 14867
rect 263 14811 275 14867
rect 195 14797 275 14811
rect 379 14811 391 14867
rect 447 14811 459 14867
rect 379 14797 459 14811
rect 563 14811 575 14867
rect 631 14811 643 14867
rect 856 15240 873 15242
rect 810 14822 856 14833
rect 563 14797 643 14811
rect 195 14717 275 14719
rect -693 14661 -681 14717
rect -625 14661 207 14717
rect 263 14661 275 14717
rect -693 14649 -607 14661
rect 195 14659 275 14661
rect -477 14601 -407 14613
rect 379 14601 459 14603
rect -477 14545 -465 14601
rect -409 14545 391 14601
rect 447 14545 459 14601
rect -477 14533 -407 14545
rect 379 14543 459 14545
rect 708 14601 788 14603
rect 975 14601 1045 14613
rect 708 14545 720 14601
rect 776 14545 977 14601
rect 1033 14545 1045 14601
rect 708 14543 788 14545
rect 975 14535 1045 14545
rect 563 14485 643 14487
rect -193 14429 575 14485
rect 631 14429 643 14485
rect -193 13698 -137 14429
rect 563 14427 643 14429
rect 195 14335 275 14349
rect -18 14313 28 14324
rect 195 14279 207 14335
rect 263 14279 275 14335
rect 379 14335 459 14349
rect 379 14279 391 14335
rect 447 14279 459 14335
rect 563 14335 643 14349
rect 563 14279 575 14335
rect 631 14279 643 14335
rect 810 14313 856 14324
rect 197 14276 208 14279
rect 262 14276 273 14279
rect 381 14276 392 14279
rect 446 14276 457 14279
rect 565 14276 576 14279
rect 630 14276 641 14279
rect 120 14230 166 14241
rect 28 14056 120 14230
rect 120 14045 166 14056
rect 304 14230 350 14241
rect 304 14045 350 14056
rect 488 14230 534 14241
rect 672 14230 718 14241
rect 655 14203 672 14205
rect 718 14203 735 14205
rect 655 14083 667 14203
rect 723 14083 735 14203
rect 655 14081 672 14083
rect 488 14045 534 14056
rect 718 14081 735 14083
rect 672 14045 718 14056
rect -18 13828 28 13973
rect 197 13964 208 14010
rect 262 13964 273 14010
rect 197 13931 273 13964
rect 381 13964 392 14010
rect 446 13964 457 14010
rect 381 13931 457 13964
rect 565 13964 576 14010
rect 630 13964 641 14010
rect 565 13931 641 13964
rect 810 13828 856 13973
rect -30 13816 50 13828
rect -30 13760 -18 13816
rect 38 13760 50 13816
rect -30 13748 50 13760
rect 788 13816 868 13828
rect 788 13760 800 13816
rect 856 13760 868 13816
rect 788 13748 868 13760
rect 1141 13698 1221 13708
rect -193 13642 1153 13698
rect 1209 13642 1221 13698
rect 1141 13640 1221 13642
rect 975 13589 1045 13591
rect -193 13588 1045 13589
rect -193 13534 977 13588
rect 1033 13534 1045 13588
rect -193 13533 1045 13534
rect -2085 13481 -1999 13485
rect -2085 13425 -2073 13481
rect -2017 13425 -1999 13481
rect -2085 13413 -1999 13425
rect -2574 13268 -2528 13279
rect -2359 13277 -2283 13310
rect -2359 13231 -2348 13277
rect -2294 13231 -2283 13277
rect -2175 13277 -2099 13310
rect -2175 13231 -2164 13277
rect -2110 13231 -2099 13277
rect -1991 13277 -1915 13310
rect -1991 13231 -1980 13277
rect -1926 13231 -1915 13277
rect -1746 13268 -1700 13279
rect -2436 13185 -2390 13196
rect -2453 13158 -2436 13160
rect -2252 13185 -2206 13196
rect -2390 13158 -2373 13160
rect -2528 13038 -2441 13158
rect -2385 13038 -2373 13158
rect -2453 13036 -2436 13038
rect -2528 12738 -2436 12858
rect -2390 13036 -2373 13038
rect -2269 12858 -2252 12860
rect -2068 13185 -2022 13196
rect -2085 13158 -2068 13160
rect -1884 13185 -1838 13196
rect -2022 13158 -2005 13160
rect -2085 13038 -2073 13158
rect -2017 13038 -2005 13158
rect -2085 13036 -2068 13038
rect -2206 12858 -2189 12860
rect -2269 12738 -2257 12858
rect -2201 12738 -2189 12858
rect -2269 12736 -2252 12738
rect -2436 12700 -2390 12711
rect -2206 12736 -2189 12738
rect -2252 12700 -2206 12711
rect -2022 13036 -2005 13038
rect -1901 12858 -1884 12860
rect -1763 13158 -1746 13160
rect -1700 13158 -1683 13160
rect -1763 13037 -1751 13158
rect -1695 13037 -1683 13158
rect -1763 13035 -1746 13037
rect -1838 12858 -1821 12860
rect -1901 12738 -1889 12858
rect -1833 12738 -1821 12858
rect -1901 12736 -1884 12738
rect -2068 12700 -2022 12711
rect -1838 12736 -1821 12738
rect -1884 12700 -1838 12711
rect -2359 12662 -2348 12665
rect -2294 12662 -2283 12665
rect -2175 12662 -2164 12665
rect -2110 12662 -2099 12665
rect -1991 12662 -1980 12665
rect -1926 12662 -1915 12665
rect -2574 12617 -2528 12628
rect -2361 12606 -2349 12662
rect -2293 12606 -2281 12662
rect -2361 12592 -2281 12606
rect -2177 12606 -2165 12662
rect -2109 12606 -2097 12662
rect -2177 12592 -2097 12606
rect -1993 12606 -1981 12662
rect -1925 12606 -1913 12662
rect -1700 13035 -1683 13037
rect -1746 12617 -1700 12628
rect -1993 12592 -1913 12606
rect -2361 12512 -2281 12514
rect -2749 12456 -2349 12512
rect -2293 12456 -2281 12512
rect -193 12512 -137 13533
rect 975 13525 1045 13533
rect 471 13481 557 13485
rect 471 13425 483 13481
rect 539 13425 557 13481
rect 471 13413 557 13425
rect -18 13268 28 13279
rect 197 13277 273 13310
rect 197 13231 208 13277
rect 262 13231 273 13277
rect 381 13277 457 13310
rect 381 13231 392 13277
rect 446 13231 457 13277
rect 565 13277 641 13310
rect 565 13231 576 13277
rect 630 13231 641 13277
rect 810 13268 856 13279
rect 120 13185 166 13196
rect 103 13158 120 13160
rect 304 13185 350 13196
rect 166 13158 183 13160
rect 28 13038 115 13158
rect 171 13038 183 13158
rect 103 13036 120 13038
rect 28 12738 120 12858
rect 166 13036 183 13038
rect 287 12858 304 12860
rect 488 13185 534 13196
rect 471 13158 488 13160
rect 672 13185 718 13196
rect 534 13158 551 13160
rect 471 13038 483 13158
rect 539 13038 551 13158
rect 471 13036 488 13038
rect 350 12858 367 12860
rect 287 12738 299 12858
rect 355 12738 367 12858
rect 287 12736 304 12738
rect 120 12700 166 12711
rect 350 12736 367 12738
rect 304 12700 350 12711
rect 534 13036 551 13038
rect 655 12858 672 12860
rect 793 13158 810 13160
rect 856 13158 873 13160
rect 793 13037 805 13158
rect 861 13037 873 13158
rect 793 13035 810 13037
rect 718 12858 735 12860
rect 655 12738 667 12858
rect 723 12738 735 12858
rect 655 12736 672 12738
rect 488 12700 534 12711
rect 718 12736 735 12738
rect 672 12700 718 12711
rect 197 12662 208 12665
rect 262 12662 273 12665
rect 381 12662 392 12665
rect 446 12662 457 12665
rect 565 12662 576 12665
rect 630 12662 641 12665
rect -18 12617 28 12628
rect 195 12606 207 12662
rect 263 12606 275 12662
rect 195 12592 275 12606
rect 379 12606 391 12662
rect 447 12606 459 12662
rect 379 12592 459 12606
rect 563 12606 575 12662
rect 631 12606 643 12662
rect 856 13035 873 13037
rect 810 12617 856 12628
rect 563 12592 643 12606
rect 195 12512 275 12514
rect -193 12456 207 12512
rect 263 12456 275 12512
rect 1293 12512 1349 15738
rect 3844 15738 5391 15794
rect 3349 14717 3435 14729
rect 3844 14717 3900 15738
rect 4513 15686 4599 15690
rect 4513 15630 4525 15686
rect 4581 15630 4599 15686
rect 4513 15618 4599 15630
rect 4024 15473 4070 15484
rect 4239 15482 4315 15515
rect 4239 15436 4250 15482
rect 4304 15436 4315 15482
rect 4423 15482 4499 15515
rect 4423 15436 4434 15482
rect 4488 15436 4499 15482
rect 4607 15482 4683 15515
rect 4607 15436 4618 15482
rect 4672 15436 4683 15482
rect 4852 15473 4898 15484
rect 4162 15390 4208 15401
rect 4145 15363 4162 15365
rect 4346 15390 4392 15401
rect 4208 15363 4225 15365
rect 4070 15243 4157 15363
rect 4213 15243 4225 15363
rect 4145 15241 4162 15243
rect 4070 14943 4162 15063
rect 4208 15241 4225 15243
rect 4329 15063 4346 15065
rect 4530 15390 4576 15401
rect 4513 15363 4530 15365
rect 4714 15390 4760 15401
rect 4576 15363 4593 15365
rect 4513 15243 4525 15363
rect 4581 15243 4593 15363
rect 4513 15241 4530 15243
rect 4392 15063 4409 15065
rect 4329 14943 4341 15063
rect 4397 14943 4409 15063
rect 4329 14941 4346 14943
rect 4162 14905 4208 14916
rect 4392 14941 4409 14943
rect 4346 14905 4392 14916
rect 4576 15241 4593 15243
rect 4697 15063 4714 15065
rect 4835 15363 4852 15365
rect 4898 15363 4915 15365
rect 4835 15242 4847 15363
rect 4903 15242 4915 15363
rect 4835 15240 4852 15242
rect 4760 15063 4777 15065
rect 4697 14943 4709 15063
rect 4765 14943 4777 15063
rect 4697 14941 4714 14943
rect 4530 14905 4576 14916
rect 4760 14941 4777 14943
rect 4714 14905 4760 14916
rect 4239 14867 4250 14870
rect 4304 14867 4315 14870
rect 4423 14867 4434 14870
rect 4488 14867 4499 14870
rect 4607 14867 4618 14870
rect 4672 14867 4683 14870
rect 4024 14822 4070 14833
rect 4237 14811 4249 14867
rect 4305 14811 4317 14867
rect 4237 14797 4317 14811
rect 4421 14811 4433 14867
rect 4489 14811 4501 14867
rect 4421 14797 4501 14811
rect 4605 14811 4617 14867
rect 4673 14811 4685 14867
rect 4898 15240 4915 15242
rect 4852 14822 4898 14833
rect 4605 14797 4685 14811
rect 4237 14717 4317 14719
rect 3349 14661 3361 14717
rect 3417 14661 4249 14717
rect 4305 14661 4317 14717
rect 3349 14649 3435 14661
rect 4237 14659 4317 14661
rect 3565 14601 3635 14613
rect 4421 14601 4501 14603
rect 3565 14545 3577 14601
rect 3633 14545 4433 14601
rect 4489 14545 4501 14601
rect 3565 14533 3635 14545
rect 4421 14543 4501 14545
rect 4750 14601 4830 14603
rect 5017 14601 5087 14613
rect 4750 14545 4762 14601
rect 4818 14545 5019 14601
rect 5075 14545 5087 14601
rect 4750 14543 4830 14545
rect 5017 14535 5087 14545
rect 4605 14485 4685 14487
rect 3849 14429 4617 14485
rect 4673 14429 4685 14485
rect 3849 13698 3905 14429
rect 4605 14427 4685 14429
rect 4237 14335 4317 14349
rect 4024 14313 4070 14324
rect 4237 14279 4249 14335
rect 4305 14279 4317 14335
rect 4421 14335 4501 14349
rect 4421 14279 4433 14335
rect 4489 14279 4501 14335
rect 4605 14335 4685 14349
rect 4605 14279 4617 14335
rect 4673 14279 4685 14335
rect 4852 14313 4898 14324
rect 4239 14276 4250 14279
rect 4304 14276 4315 14279
rect 4423 14276 4434 14279
rect 4488 14276 4499 14279
rect 4607 14276 4618 14279
rect 4672 14276 4683 14279
rect 4162 14230 4208 14241
rect 4070 14056 4162 14230
rect 4162 14045 4208 14056
rect 4346 14230 4392 14241
rect 4346 14045 4392 14056
rect 4530 14230 4576 14241
rect 4714 14230 4760 14241
rect 4697 14203 4714 14205
rect 4760 14203 4777 14205
rect 4697 14083 4709 14203
rect 4765 14083 4777 14203
rect 4697 14081 4714 14083
rect 4530 14045 4576 14056
rect 4760 14081 4777 14083
rect 4714 14045 4760 14056
rect 4024 13828 4070 13973
rect 4239 13964 4250 14010
rect 4304 13964 4315 14010
rect 4239 13931 4315 13964
rect 4423 13964 4434 14010
rect 4488 13964 4499 14010
rect 4423 13931 4499 13964
rect 4607 13964 4618 14010
rect 4672 13964 4683 14010
rect 4607 13931 4683 13964
rect 4852 13828 4898 13973
rect 4012 13816 4092 13828
rect 4012 13760 4024 13816
rect 4080 13760 4092 13816
rect 4012 13748 4092 13760
rect 4830 13816 4910 13828
rect 4830 13760 4842 13816
rect 4898 13760 4910 13816
rect 4830 13748 4910 13760
rect 5183 13698 5263 13708
rect 3849 13642 5195 13698
rect 5251 13642 5263 13698
rect 5183 13640 5263 13642
rect 5017 13589 5087 13591
rect 3849 13588 5087 13589
rect 3849 13534 5019 13588
rect 5075 13534 5087 13588
rect 3849 13533 5087 13534
rect 1957 13481 2043 13485
rect 1957 13425 1969 13481
rect 2025 13425 2043 13481
rect 1957 13413 2043 13425
rect 1468 13268 1514 13279
rect 1683 13277 1759 13310
rect 1683 13231 1694 13277
rect 1748 13231 1759 13277
rect 1867 13277 1943 13310
rect 1867 13231 1878 13277
rect 1932 13231 1943 13277
rect 2051 13277 2127 13310
rect 2051 13231 2062 13277
rect 2116 13231 2127 13277
rect 2296 13268 2342 13279
rect 1606 13185 1652 13196
rect 1589 13158 1606 13160
rect 1790 13185 1836 13196
rect 1652 13158 1669 13160
rect 1514 13038 1601 13158
rect 1657 13038 1669 13158
rect 1589 13036 1606 13038
rect 1514 12738 1606 12858
rect 1652 13036 1669 13038
rect 1773 12858 1790 12860
rect 1974 13185 2020 13196
rect 1957 13158 1974 13160
rect 2158 13185 2204 13196
rect 2020 13158 2037 13160
rect 1957 13038 1969 13158
rect 2025 13038 2037 13158
rect 1957 13036 1974 13038
rect 1836 12858 1853 12860
rect 1773 12738 1785 12858
rect 1841 12738 1853 12858
rect 1773 12736 1790 12738
rect 1606 12700 1652 12711
rect 1836 12736 1853 12738
rect 1790 12700 1836 12711
rect 2020 13036 2037 13038
rect 2141 12858 2158 12860
rect 2279 13158 2296 13160
rect 2342 13158 2359 13160
rect 2279 13037 2291 13158
rect 2347 13037 2359 13158
rect 2279 13035 2296 13037
rect 2204 12858 2221 12860
rect 2141 12738 2153 12858
rect 2209 12738 2221 12858
rect 2141 12736 2158 12738
rect 1974 12700 2020 12711
rect 2204 12736 2221 12738
rect 2158 12700 2204 12711
rect 1683 12662 1694 12665
rect 1748 12662 1759 12665
rect 1867 12662 1878 12665
rect 1932 12662 1943 12665
rect 2051 12662 2062 12665
rect 2116 12662 2127 12665
rect 1468 12617 1514 12628
rect 1681 12606 1693 12662
rect 1749 12606 1761 12662
rect 1681 12592 1761 12606
rect 1865 12606 1877 12662
rect 1933 12606 1945 12662
rect 1865 12592 1945 12606
rect 2049 12606 2061 12662
rect 2117 12606 2129 12662
rect 2342 13035 2359 13037
rect 2296 12617 2342 12628
rect 2049 12592 2129 12606
rect 1681 12512 1761 12514
rect 1293 12456 1693 12512
rect 1749 12456 1761 12512
rect 3849 12512 3905 13533
rect 5017 13525 5087 13533
rect 4513 13481 4599 13485
rect 4513 13425 4525 13481
rect 4581 13425 4599 13481
rect 4513 13413 4599 13425
rect 4024 13268 4070 13279
rect 4239 13277 4315 13310
rect 4239 13231 4250 13277
rect 4304 13231 4315 13277
rect 4423 13277 4499 13310
rect 4423 13231 4434 13277
rect 4488 13231 4499 13277
rect 4607 13277 4683 13310
rect 4607 13231 4618 13277
rect 4672 13231 4683 13277
rect 4852 13268 4898 13279
rect 4162 13185 4208 13196
rect 4145 13158 4162 13160
rect 4346 13185 4392 13196
rect 4208 13158 4225 13160
rect 4070 13038 4157 13158
rect 4213 13038 4225 13158
rect 4145 13036 4162 13038
rect 4070 12738 4162 12858
rect 4208 13036 4225 13038
rect 4329 12858 4346 12860
rect 4530 13185 4576 13196
rect 4513 13158 4530 13160
rect 4714 13185 4760 13196
rect 4576 13158 4593 13160
rect 4513 13038 4525 13158
rect 4581 13038 4593 13158
rect 4513 13036 4530 13038
rect 4392 12858 4409 12860
rect 4329 12738 4341 12858
rect 4397 12738 4409 12858
rect 4329 12736 4346 12738
rect 4162 12700 4208 12711
rect 4392 12736 4409 12738
rect 4346 12700 4392 12711
rect 4576 13036 4593 13038
rect 4697 12858 4714 12860
rect 4835 13158 4852 13160
rect 4898 13158 4915 13160
rect 4835 13037 4847 13158
rect 4903 13037 4915 13158
rect 4835 13035 4852 13037
rect 4760 12858 4777 12860
rect 4697 12738 4709 12858
rect 4765 12738 4777 12858
rect 4697 12736 4714 12738
rect 4530 12700 4576 12711
rect 4760 12736 4777 12738
rect 4714 12700 4760 12711
rect 4239 12662 4250 12665
rect 4304 12662 4315 12665
rect 4423 12662 4434 12665
rect 4488 12662 4499 12665
rect 4607 12662 4618 12665
rect 4672 12662 4683 12665
rect 4024 12617 4070 12628
rect 4237 12606 4249 12662
rect 4305 12606 4317 12662
rect 4237 12592 4317 12606
rect 4421 12606 4433 12662
rect 4489 12606 4501 12662
rect 4421 12592 4501 12606
rect 4605 12606 4617 12662
rect 4673 12606 4685 12662
rect 4898 13035 4915 13037
rect 4852 12617 4898 12628
rect 4605 12592 4685 12606
rect 4237 12512 4317 12514
rect 3849 12456 4249 12512
rect 4305 12456 4317 12512
rect 5335 12512 5391 15738
rect 7886 15738 9433 15794
rect 7391 14717 7477 14729
rect 7886 14717 7942 15738
rect 8555 15686 8641 15690
rect 8555 15630 8567 15686
rect 8623 15630 8641 15686
rect 8555 15618 8641 15630
rect 8066 15473 8112 15484
rect 8281 15482 8357 15515
rect 8281 15436 8292 15482
rect 8346 15436 8357 15482
rect 8465 15482 8541 15515
rect 8465 15436 8476 15482
rect 8530 15436 8541 15482
rect 8649 15482 8725 15515
rect 8649 15436 8660 15482
rect 8714 15436 8725 15482
rect 8894 15473 8940 15484
rect 8204 15390 8250 15401
rect 8187 15363 8204 15365
rect 8388 15390 8434 15401
rect 8250 15363 8267 15365
rect 8112 15243 8199 15363
rect 8255 15243 8267 15363
rect 8187 15241 8204 15243
rect 8112 14943 8204 15063
rect 8250 15241 8267 15243
rect 8371 15063 8388 15065
rect 8572 15390 8618 15401
rect 8555 15363 8572 15365
rect 8756 15390 8802 15401
rect 8618 15363 8635 15365
rect 8555 15243 8567 15363
rect 8623 15243 8635 15363
rect 8555 15241 8572 15243
rect 8434 15063 8451 15065
rect 8371 14943 8383 15063
rect 8439 14943 8451 15063
rect 8371 14941 8388 14943
rect 8204 14905 8250 14916
rect 8434 14941 8451 14943
rect 8388 14905 8434 14916
rect 8618 15241 8635 15243
rect 8739 15063 8756 15065
rect 8877 15363 8894 15365
rect 8940 15363 8957 15365
rect 8877 15242 8889 15363
rect 8945 15242 8957 15363
rect 8877 15240 8894 15242
rect 8802 15063 8819 15065
rect 8739 14943 8751 15063
rect 8807 14943 8819 15063
rect 8739 14941 8756 14943
rect 8572 14905 8618 14916
rect 8802 14941 8819 14943
rect 8756 14905 8802 14916
rect 8281 14867 8292 14870
rect 8346 14867 8357 14870
rect 8465 14867 8476 14870
rect 8530 14867 8541 14870
rect 8649 14867 8660 14870
rect 8714 14867 8725 14870
rect 8066 14822 8112 14833
rect 8279 14811 8291 14867
rect 8347 14811 8359 14867
rect 8279 14797 8359 14811
rect 8463 14811 8475 14867
rect 8531 14811 8543 14867
rect 8463 14797 8543 14811
rect 8647 14811 8659 14867
rect 8715 14811 8727 14867
rect 8940 15240 8957 15242
rect 8894 14822 8940 14833
rect 8647 14797 8727 14811
rect 8279 14717 8359 14719
rect 7391 14661 7403 14717
rect 7459 14661 8291 14717
rect 8347 14661 8359 14717
rect 7391 14649 7477 14661
rect 8279 14659 8359 14661
rect 7607 14601 7677 14613
rect 8463 14601 8543 14603
rect 7607 14545 7619 14601
rect 7675 14545 8475 14601
rect 8531 14545 8543 14601
rect 7607 14533 7677 14545
rect 8463 14543 8543 14545
rect 8792 14601 8872 14603
rect 9059 14601 9129 14613
rect 8792 14545 8804 14601
rect 8860 14545 9061 14601
rect 9117 14545 9129 14601
rect 8792 14543 8872 14545
rect 9059 14535 9129 14545
rect 8647 14485 8727 14487
rect 7891 14429 8659 14485
rect 8715 14429 8727 14485
rect 7891 13698 7947 14429
rect 8647 14427 8727 14429
rect 8279 14335 8359 14349
rect 8066 14313 8112 14324
rect 8279 14279 8291 14335
rect 8347 14279 8359 14335
rect 8463 14335 8543 14349
rect 8463 14279 8475 14335
rect 8531 14279 8543 14335
rect 8647 14335 8727 14349
rect 8647 14279 8659 14335
rect 8715 14279 8727 14335
rect 8894 14313 8940 14324
rect 8281 14276 8292 14279
rect 8346 14276 8357 14279
rect 8465 14276 8476 14279
rect 8530 14276 8541 14279
rect 8649 14276 8660 14279
rect 8714 14276 8725 14279
rect 8204 14230 8250 14241
rect 8112 14056 8204 14230
rect 8204 14045 8250 14056
rect 8388 14230 8434 14241
rect 8388 14045 8434 14056
rect 8572 14230 8618 14241
rect 8756 14230 8802 14241
rect 8739 14203 8756 14205
rect 8802 14203 8819 14205
rect 8739 14083 8751 14203
rect 8807 14083 8819 14203
rect 8739 14081 8756 14083
rect 8572 14045 8618 14056
rect 8802 14081 8819 14083
rect 8756 14045 8802 14056
rect 8066 13828 8112 13973
rect 8281 13964 8292 14010
rect 8346 13964 8357 14010
rect 8281 13931 8357 13964
rect 8465 13964 8476 14010
rect 8530 13964 8541 14010
rect 8465 13931 8541 13964
rect 8649 13964 8660 14010
rect 8714 13964 8725 14010
rect 8649 13931 8725 13964
rect 8894 13828 8940 13973
rect 8054 13816 8134 13828
rect 8054 13760 8066 13816
rect 8122 13760 8134 13816
rect 8054 13748 8134 13760
rect 8872 13816 8952 13828
rect 8872 13760 8884 13816
rect 8940 13760 8952 13816
rect 8872 13748 8952 13760
rect 9225 13698 9305 13708
rect 7891 13642 9237 13698
rect 9293 13642 9305 13698
rect 9225 13640 9305 13642
rect 9059 13589 9129 13591
rect 7891 13588 9129 13589
rect 7891 13534 9061 13588
rect 9117 13534 9129 13588
rect 7891 13533 9129 13534
rect 5999 13481 6085 13485
rect 5999 13425 6011 13481
rect 6067 13425 6085 13481
rect 5999 13413 6085 13425
rect 5510 13268 5556 13279
rect 5725 13277 5801 13310
rect 5725 13231 5736 13277
rect 5790 13231 5801 13277
rect 5909 13277 5985 13310
rect 5909 13231 5920 13277
rect 5974 13231 5985 13277
rect 6093 13277 6169 13310
rect 6093 13231 6104 13277
rect 6158 13231 6169 13277
rect 6338 13268 6384 13279
rect 5648 13185 5694 13196
rect 5631 13158 5648 13160
rect 5832 13185 5878 13196
rect 5694 13158 5711 13160
rect 5556 13038 5643 13158
rect 5699 13038 5711 13158
rect 5631 13036 5648 13038
rect 5556 12738 5648 12858
rect 5694 13036 5711 13038
rect 5815 12858 5832 12860
rect 6016 13185 6062 13196
rect 5999 13158 6016 13160
rect 6200 13185 6246 13196
rect 6062 13158 6079 13160
rect 5999 13038 6011 13158
rect 6067 13038 6079 13158
rect 5999 13036 6016 13038
rect 5878 12858 5895 12860
rect 5815 12738 5827 12858
rect 5883 12738 5895 12858
rect 5815 12736 5832 12738
rect 5648 12700 5694 12711
rect 5878 12736 5895 12738
rect 5832 12700 5878 12711
rect 6062 13036 6079 13038
rect 6183 12858 6200 12860
rect 6321 13158 6338 13160
rect 6384 13158 6401 13160
rect 6321 13037 6333 13158
rect 6389 13037 6401 13158
rect 6321 13035 6338 13037
rect 6246 12858 6263 12860
rect 6183 12738 6195 12858
rect 6251 12738 6263 12858
rect 6183 12736 6200 12738
rect 6016 12700 6062 12711
rect 6246 12736 6263 12738
rect 6200 12700 6246 12711
rect 5725 12662 5736 12665
rect 5790 12662 5801 12665
rect 5909 12662 5920 12665
rect 5974 12662 5985 12665
rect 6093 12662 6104 12665
rect 6158 12662 6169 12665
rect 5510 12617 5556 12628
rect 5723 12606 5735 12662
rect 5791 12606 5803 12662
rect 5723 12592 5803 12606
rect 5907 12606 5919 12662
rect 5975 12606 5987 12662
rect 5907 12592 5987 12606
rect 6091 12606 6103 12662
rect 6159 12606 6171 12662
rect 6384 13035 6401 13037
rect 6338 12617 6384 12628
rect 6091 12592 6171 12606
rect 5723 12512 5803 12514
rect 5335 12456 5735 12512
rect 5791 12456 5803 12512
rect 7891 12512 7947 13533
rect 9059 13525 9129 13533
rect 8555 13481 8641 13485
rect 8555 13425 8567 13481
rect 8623 13425 8641 13481
rect 8555 13413 8641 13425
rect 8066 13268 8112 13279
rect 8281 13277 8357 13310
rect 8281 13231 8292 13277
rect 8346 13231 8357 13277
rect 8465 13277 8541 13310
rect 8465 13231 8476 13277
rect 8530 13231 8541 13277
rect 8649 13277 8725 13310
rect 8649 13231 8660 13277
rect 8714 13231 8725 13277
rect 8894 13268 8940 13279
rect 8204 13185 8250 13196
rect 8187 13158 8204 13160
rect 8388 13185 8434 13196
rect 8250 13158 8267 13160
rect 8112 13038 8199 13158
rect 8255 13038 8267 13158
rect 8187 13036 8204 13038
rect 8112 12738 8204 12858
rect 8250 13036 8267 13038
rect 8371 12858 8388 12860
rect 8572 13185 8618 13196
rect 8555 13158 8572 13160
rect 8756 13185 8802 13196
rect 8618 13158 8635 13160
rect 8555 13038 8567 13158
rect 8623 13038 8635 13158
rect 8555 13036 8572 13038
rect 8434 12858 8451 12860
rect 8371 12738 8383 12858
rect 8439 12738 8451 12858
rect 8371 12736 8388 12738
rect 8204 12700 8250 12711
rect 8434 12736 8451 12738
rect 8388 12700 8434 12711
rect 8618 13036 8635 13038
rect 8739 12858 8756 12860
rect 8877 13158 8894 13160
rect 8940 13158 8957 13160
rect 8877 13037 8889 13158
rect 8945 13037 8957 13158
rect 8877 13035 8894 13037
rect 8802 12858 8819 12860
rect 8739 12738 8751 12858
rect 8807 12738 8819 12858
rect 8739 12736 8756 12738
rect 8572 12700 8618 12711
rect 8802 12736 8819 12738
rect 8756 12700 8802 12711
rect 8281 12662 8292 12665
rect 8346 12662 8357 12665
rect 8465 12662 8476 12665
rect 8530 12662 8541 12665
rect 8649 12662 8660 12665
rect 8714 12662 8725 12665
rect 8066 12617 8112 12628
rect 8279 12606 8291 12662
rect 8347 12606 8359 12662
rect 8279 12592 8359 12606
rect 8463 12606 8475 12662
rect 8531 12606 8543 12662
rect 8463 12592 8543 12606
rect 8647 12606 8659 12662
rect 8715 12606 8727 12662
rect 8940 13035 8957 13037
rect 8894 12617 8940 12628
rect 8647 12592 8727 12606
rect 8279 12512 8359 12514
rect 7891 12456 8291 12512
rect 8347 12456 8359 12512
rect 9377 12512 9433 15738
rect 11928 15738 13475 15794
rect 11433 14717 11519 14729
rect 11928 14717 11984 15738
rect 12597 15686 12683 15690
rect 12597 15630 12609 15686
rect 12665 15630 12683 15686
rect 12597 15618 12683 15630
rect 12108 15473 12154 15484
rect 12323 15482 12399 15515
rect 12323 15436 12334 15482
rect 12388 15436 12399 15482
rect 12507 15482 12583 15515
rect 12507 15436 12518 15482
rect 12572 15436 12583 15482
rect 12691 15482 12767 15515
rect 12691 15436 12702 15482
rect 12756 15436 12767 15482
rect 12936 15473 12982 15484
rect 12246 15390 12292 15401
rect 12229 15363 12246 15365
rect 12430 15390 12476 15401
rect 12292 15363 12309 15365
rect 12154 15243 12241 15363
rect 12297 15243 12309 15363
rect 12229 15241 12246 15243
rect 12154 14943 12246 15063
rect 12292 15241 12309 15243
rect 12413 15063 12430 15065
rect 12614 15390 12660 15401
rect 12597 15363 12614 15365
rect 12798 15390 12844 15401
rect 12660 15363 12677 15365
rect 12597 15243 12609 15363
rect 12665 15243 12677 15363
rect 12597 15241 12614 15243
rect 12476 15063 12493 15065
rect 12413 14943 12425 15063
rect 12481 14943 12493 15063
rect 12413 14941 12430 14943
rect 12246 14905 12292 14916
rect 12476 14941 12493 14943
rect 12430 14905 12476 14916
rect 12660 15241 12677 15243
rect 12781 15063 12798 15065
rect 12919 15363 12936 15365
rect 12982 15363 12999 15365
rect 12919 15242 12931 15363
rect 12987 15242 12999 15363
rect 12919 15240 12936 15242
rect 12844 15063 12861 15065
rect 12781 14943 12793 15063
rect 12849 14943 12861 15063
rect 12781 14941 12798 14943
rect 12614 14905 12660 14916
rect 12844 14941 12861 14943
rect 12798 14905 12844 14916
rect 12323 14867 12334 14870
rect 12388 14867 12399 14870
rect 12507 14867 12518 14870
rect 12572 14867 12583 14870
rect 12691 14867 12702 14870
rect 12756 14867 12767 14870
rect 12108 14822 12154 14833
rect 12321 14811 12333 14867
rect 12389 14811 12401 14867
rect 12321 14797 12401 14811
rect 12505 14811 12517 14867
rect 12573 14811 12585 14867
rect 12505 14797 12585 14811
rect 12689 14811 12701 14867
rect 12757 14811 12769 14867
rect 12982 15240 12999 15242
rect 12936 14822 12982 14833
rect 12689 14797 12769 14811
rect 12321 14717 12401 14719
rect 11433 14661 11445 14717
rect 11501 14661 12333 14717
rect 12389 14661 12401 14717
rect 11433 14649 11519 14661
rect 12321 14659 12401 14661
rect 11649 14601 11719 14613
rect 12505 14601 12585 14603
rect 11649 14545 11661 14601
rect 11717 14545 12517 14601
rect 12573 14545 12585 14601
rect 11649 14533 11719 14545
rect 12505 14543 12585 14545
rect 12834 14601 12914 14603
rect 13101 14601 13171 14613
rect 12834 14545 12846 14601
rect 12902 14545 13103 14601
rect 13159 14545 13171 14601
rect 12834 14543 12914 14545
rect 13101 14535 13171 14545
rect 12689 14485 12769 14487
rect 11933 14429 12701 14485
rect 12757 14429 12769 14485
rect 11933 13698 11989 14429
rect 12689 14427 12769 14429
rect 12321 14335 12401 14349
rect 12108 14313 12154 14324
rect 12321 14279 12333 14335
rect 12389 14279 12401 14335
rect 12505 14335 12585 14349
rect 12505 14279 12517 14335
rect 12573 14279 12585 14335
rect 12689 14335 12769 14349
rect 12689 14279 12701 14335
rect 12757 14279 12769 14335
rect 12936 14313 12982 14324
rect 12323 14276 12334 14279
rect 12388 14276 12399 14279
rect 12507 14276 12518 14279
rect 12572 14276 12583 14279
rect 12691 14276 12702 14279
rect 12756 14276 12767 14279
rect 12246 14230 12292 14241
rect 12154 14056 12246 14230
rect 12246 14045 12292 14056
rect 12430 14230 12476 14241
rect 12430 14045 12476 14056
rect 12614 14230 12660 14241
rect 12798 14230 12844 14241
rect 12781 14203 12798 14205
rect 12844 14203 12861 14205
rect 12781 14083 12793 14203
rect 12849 14083 12861 14203
rect 12781 14081 12798 14083
rect 12614 14045 12660 14056
rect 12844 14081 12861 14083
rect 12798 14045 12844 14056
rect 12108 13828 12154 13973
rect 12323 13964 12334 14010
rect 12388 13964 12399 14010
rect 12323 13931 12399 13964
rect 12507 13964 12518 14010
rect 12572 13964 12583 14010
rect 12507 13931 12583 13964
rect 12691 13964 12702 14010
rect 12756 13964 12767 14010
rect 12691 13931 12767 13964
rect 12936 13828 12982 13973
rect 12096 13816 12176 13828
rect 12096 13760 12108 13816
rect 12164 13760 12176 13816
rect 12096 13748 12176 13760
rect 12914 13816 12994 13828
rect 12914 13760 12926 13816
rect 12982 13760 12994 13816
rect 12914 13748 12994 13760
rect 13267 13698 13347 13708
rect 11933 13642 13279 13698
rect 13335 13642 13347 13698
rect 13267 13640 13347 13642
rect 13101 13589 13171 13591
rect 11933 13588 13171 13589
rect 11933 13534 13103 13588
rect 13159 13534 13171 13588
rect 11933 13533 13171 13534
rect 10041 13481 10127 13485
rect 10041 13425 10053 13481
rect 10109 13425 10127 13481
rect 10041 13413 10127 13425
rect 9552 13268 9598 13279
rect 9767 13277 9843 13310
rect 9767 13231 9778 13277
rect 9832 13231 9843 13277
rect 9951 13277 10027 13310
rect 9951 13231 9962 13277
rect 10016 13231 10027 13277
rect 10135 13277 10211 13310
rect 10135 13231 10146 13277
rect 10200 13231 10211 13277
rect 10380 13268 10426 13279
rect 9690 13185 9736 13196
rect 9673 13158 9690 13160
rect 9874 13185 9920 13196
rect 9736 13158 9753 13160
rect 9598 13038 9685 13158
rect 9741 13038 9753 13158
rect 9673 13036 9690 13038
rect 9598 12738 9690 12858
rect 9736 13036 9753 13038
rect 9857 12858 9874 12860
rect 10058 13185 10104 13196
rect 10041 13158 10058 13160
rect 10242 13185 10288 13196
rect 10104 13158 10121 13160
rect 10041 13038 10053 13158
rect 10109 13038 10121 13158
rect 10041 13036 10058 13038
rect 9920 12858 9937 12860
rect 9857 12738 9869 12858
rect 9925 12738 9937 12858
rect 9857 12736 9874 12738
rect 9690 12700 9736 12711
rect 9920 12736 9937 12738
rect 9874 12700 9920 12711
rect 10104 13036 10121 13038
rect 10225 12858 10242 12860
rect 10363 13158 10380 13160
rect 10426 13158 10443 13160
rect 10363 13037 10375 13158
rect 10431 13037 10443 13158
rect 10363 13035 10380 13037
rect 10288 12858 10305 12860
rect 10225 12738 10237 12858
rect 10293 12738 10305 12858
rect 10225 12736 10242 12738
rect 10058 12700 10104 12711
rect 10288 12736 10305 12738
rect 10242 12700 10288 12711
rect 9767 12662 9778 12665
rect 9832 12662 9843 12665
rect 9951 12662 9962 12665
rect 10016 12662 10027 12665
rect 10135 12662 10146 12665
rect 10200 12662 10211 12665
rect 9552 12617 9598 12628
rect 9765 12606 9777 12662
rect 9833 12606 9845 12662
rect 9765 12592 9845 12606
rect 9949 12606 9961 12662
rect 10017 12606 10029 12662
rect 9949 12592 10029 12606
rect 10133 12606 10145 12662
rect 10201 12606 10213 12662
rect 10426 13035 10443 13037
rect 10380 12617 10426 12628
rect 10133 12592 10213 12606
rect 9765 12512 9845 12514
rect 9377 12456 9777 12512
rect 9833 12456 9845 12512
rect 11933 12512 11989 13533
rect 13101 13525 13171 13533
rect 12597 13481 12683 13485
rect 12597 13425 12609 13481
rect 12665 13425 12683 13481
rect 12597 13413 12683 13425
rect 12108 13268 12154 13279
rect 12323 13277 12399 13310
rect 12323 13231 12334 13277
rect 12388 13231 12399 13277
rect 12507 13277 12583 13310
rect 12507 13231 12518 13277
rect 12572 13231 12583 13277
rect 12691 13277 12767 13310
rect 12691 13231 12702 13277
rect 12756 13231 12767 13277
rect 12936 13268 12982 13279
rect 12246 13185 12292 13196
rect 12229 13158 12246 13160
rect 12430 13185 12476 13196
rect 12292 13158 12309 13160
rect 12154 13038 12241 13158
rect 12297 13038 12309 13158
rect 12229 13036 12246 13038
rect 12154 12738 12246 12858
rect 12292 13036 12309 13038
rect 12413 12858 12430 12860
rect 12614 13185 12660 13196
rect 12597 13158 12614 13160
rect 12798 13185 12844 13196
rect 12660 13158 12677 13160
rect 12597 13038 12609 13158
rect 12665 13038 12677 13158
rect 12597 13036 12614 13038
rect 12476 12858 12493 12860
rect 12413 12738 12425 12858
rect 12481 12738 12493 12858
rect 12413 12736 12430 12738
rect 12246 12700 12292 12711
rect 12476 12736 12493 12738
rect 12430 12700 12476 12711
rect 12660 13036 12677 13038
rect 12781 12858 12798 12860
rect 12919 13158 12936 13160
rect 12982 13158 12999 13160
rect 12919 13037 12931 13158
rect 12987 13037 12999 13158
rect 12919 13035 12936 13037
rect 12844 12858 12861 12860
rect 12781 12738 12793 12858
rect 12849 12738 12861 12858
rect 12781 12736 12798 12738
rect 12614 12700 12660 12711
rect 12844 12736 12861 12738
rect 12798 12700 12844 12711
rect 12323 12662 12334 12665
rect 12388 12662 12399 12665
rect 12507 12662 12518 12665
rect 12572 12662 12583 12665
rect 12691 12662 12702 12665
rect 12756 12662 12767 12665
rect 12108 12617 12154 12628
rect 12321 12606 12333 12662
rect 12389 12606 12401 12662
rect 12321 12592 12401 12606
rect 12505 12606 12517 12662
rect 12573 12606 12585 12662
rect 12505 12592 12585 12606
rect 12689 12606 12701 12662
rect 12757 12606 12769 12662
rect 12982 13035 12999 13037
rect 12936 12617 12982 12628
rect 12689 12592 12769 12606
rect 12321 12512 12401 12514
rect 11933 12456 12333 12512
rect 12389 12456 12401 12512
rect 13419 12512 13475 15738
rect 14083 13481 14169 13485
rect 14083 13425 14095 13481
rect 14151 13425 14169 13481
rect 14083 13413 14169 13425
rect 13594 13268 13640 13279
rect 13809 13277 13885 13310
rect 13809 13231 13820 13277
rect 13874 13231 13885 13277
rect 13993 13277 14069 13310
rect 13993 13231 14004 13277
rect 14058 13231 14069 13277
rect 14177 13277 14253 13310
rect 14177 13231 14188 13277
rect 14242 13231 14253 13277
rect 14422 13268 14468 13279
rect 13732 13185 13778 13196
rect 13715 13158 13732 13160
rect 13916 13185 13962 13196
rect 13778 13158 13795 13160
rect 13640 13038 13727 13158
rect 13783 13038 13795 13158
rect 13715 13036 13732 13038
rect 13640 12738 13732 12858
rect 13778 13036 13795 13038
rect 13899 12858 13916 12860
rect 14100 13185 14146 13196
rect 14083 13158 14100 13160
rect 14284 13185 14330 13196
rect 14146 13158 14163 13160
rect 14083 13038 14095 13158
rect 14151 13038 14163 13158
rect 14083 13036 14100 13038
rect 13962 12858 13979 12860
rect 13899 12738 13911 12858
rect 13967 12738 13979 12858
rect 13899 12736 13916 12738
rect 13732 12700 13778 12711
rect 13962 12736 13979 12738
rect 13916 12700 13962 12711
rect 14146 13036 14163 13038
rect 14267 12858 14284 12860
rect 14405 13158 14422 13160
rect 14468 13158 14485 13160
rect 14405 13037 14417 13158
rect 14473 13037 14485 13158
rect 14405 13035 14422 13037
rect 14330 12858 14347 12860
rect 14267 12738 14279 12858
rect 14335 12738 14347 12858
rect 14267 12736 14284 12738
rect 14100 12700 14146 12711
rect 14330 12736 14347 12738
rect 14284 12700 14330 12711
rect 13809 12662 13820 12665
rect 13874 12662 13885 12665
rect 13993 12662 14004 12665
rect 14058 12662 14069 12665
rect 14177 12662 14188 12665
rect 14242 12662 14253 12665
rect 13594 12617 13640 12628
rect 13807 12606 13819 12662
rect 13875 12606 13887 12662
rect 13807 12592 13887 12606
rect 13991 12606 14003 12662
rect 14059 12606 14071 12662
rect 13991 12592 14071 12606
rect 14175 12606 14187 12662
rect 14243 12606 14255 12662
rect 14468 13035 14485 13037
rect 14422 12617 14468 12628
rect 14175 12592 14255 12606
rect 13807 12512 13887 12514
rect 13419 12456 13819 12512
rect 13875 12456 13887 12512
rect -11901 12454 -11821 12456
rect -10415 12454 -10335 12456
rect -7889 12454 -7809 12456
rect -6403 12454 -6323 12456
rect -3847 12454 -3767 12456
rect -2361 12454 -2281 12456
rect 195 12454 275 12456
rect 1681 12454 1761 12456
rect 4237 12454 4317 12456
rect 5723 12454 5803 12456
rect 8279 12454 8359 12456
rect 9765 12454 9845 12456
rect 12321 12454 12401 12456
rect 13807 12454 13887 12456
rect -12709 12396 -12639 12410
rect -11717 12396 -11637 12398
rect -12709 12340 -12697 12396
rect -12641 12340 -11705 12396
rect -11649 12340 -11637 12396
rect -12709 12328 -12639 12340
rect -11717 12338 -11637 12340
rect -11388 12396 -11308 12398
rect -10945 12396 -10885 12406
rect -10231 12396 -10151 12398
rect -11388 12340 -11376 12396
rect -11320 12340 -10943 12396
rect -10887 12340 -10219 12396
rect -10163 12340 -10151 12396
rect -11388 12338 -11308 12340
rect -10945 12328 -10885 12340
rect -10231 12338 -10151 12340
rect -9902 12396 -9822 12398
rect -9635 12396 -9565 12408
rect -8697 12396 -8627 12410
rect -7705 12396 -7625 12398
rect -9902 12340 -9890 12396
rect -9834 12340 -9633 12396
rect -9577 12340 -8765 12396
rect -9902 12338 -9822 12340
rect -9635 12330 -9565 12340
rect -11533 12280 -11453 12282
rect -10047 12280 -9967 12282
rect -12425 12224 -11521 12280
rect -11465 12224 -11453 12280
rect -13117 11494 -13047 11506
rect -12425 11494 -12369 12224
rect -11533 12222 -11453 12224
rect -10803 12224 -10035 12280
rect -9979 12224 -9967 12280
rect -11901 12130 -11821 12144
rect -12114 12108 -12068 12119
rect -11901 12074 -11889 12130
rect -11833 12074 -11821 12130
rect -11717 12130 -11637 12144
rect -11717 12074 -11705 12130
rect -11649 12074 -11637 12130
rect -11533 12130 -11453 12144
rect -11533 12074 -11521 12130
rect -11465 12074 -11453 12130
rect -11286 12108 -11240 12119
rect -11899 12071 -11888 12074
rect -11834 12071 -11823 12074
rect -11715 12071 -11704 12074
rect -11650 12071 -11639 12074
rect -11531 12071 -11520 12074
rect -11466 12071 -11455 12074
rect -11976 12025 -11930 12036
rect -12068 11851 -11976 12025
rect -11976 11840 -11930 11851
rect -11792 12025 -11746 12036
rect -11792 11840 -11746 11851
rect -11608 12025 -11562 12036
rect -11424 12025 -11378 12036
rect -11441 11998 -11424 12000
rect -11378 11998 -11361 12000
rect -11441 11878 -11429 11998
rect -11373 11878 -11361 11998
rect -11441 11876 -11424 11878
rect -11608 11840 -11562 11851
rect -11378 11876 -11361 11878
rect -11424 11840 -11378 11851
rect -12114 11623 -12068 11768
rect -11899 11759 -11888 11805
rect -11834 11759 -11823 11805
rect -11899 11726 -11823 11759
rect -11715 11759 -11704 11805
rect -11650 11759 -11639 11805
rect -11715 11726 -11639 11759
rect -11531 11759 -11520 11805
rect -11466 11759 -11455 11805
rect -11531 11726 -11455 11759
rect -11286 11623 -11240 11768
rect -12126 11611 -12046 11623
rect -12126 11555 -12114 11611
rect -12058 11555 -12046 11611
rect -12126 11543 -12046 11555
rect -11308 11611 -11230 11623
rect -11308 11555 -11296 11611
rect -11240 11555 -11230 11611
rect -11308 11543 -11230 11555
rect -13117 11438 -13105 11494
rect -13049 11438 -12369 11494
rect -10803 11494 -10747 12224
rect -10047 12222 -9967 12224
rect -8821 12218 -8765 12340
rect -8697 12340 -8685 12396
rect -8629 12340 -7693 12396
rect -7637 12340 -7625 12396
rect -8697 12328 -8627 12340
rect -7705 12338 -7625 12340
rect -7376 12396 -7296 12398
rect -6933 12396 -6873 12406
rect -6219 12396 -6139 12398
rect -7376 12340 -7364 12396
rect -7308 12340 -6931 12396
rect -6875 12340 -6207 12396
rect -6151 12340 -6139 12396
rect -7376 12338 -7296 12340
rect -6933 12328 -6873 12340
rect -6219 12338 -6139 12340
rect -5890 12396 -5810 12398
rect -5623 12396 -5553 12408
rect -4655 12396 -4585 12410
rect -3663 12396 -3583 12398
rect -5890 12340 -5878 12396
rect -5822 12340 -5621 12396
rect -5565 12340 -4753 12396
rect -5890 12338 -5810 12340
rect -5623 12330 -5553 12340
rect -7521 12280 -7441 12282
rect -6035 12280 -5955 12282
rect -8413 12224 -7509 12280
rect -7453 12224 -7441 12280
rect -8833 12208 -8753 12218
rect -8833 12152 -8821 12208
rect -8765 12152 -8753 12208
rect -8833 12150 -8753 12152
rect -10415 12130 -10335 12144
rect -10628 12108 -10582 12119
rect -10415 12074 -10403 12130
rect -10347 12074 -10335 12130
rect -10231 12130 -10151 12144
rect -10231 12074 -10219 12130
rect -10163 12074 -10151 12130
rect -10047 12130 -9967 12144
rect -10047 12074 -10035 12130
rect -9979 12074 -9967 12130
rect -9800 12108 -9754 12119
rect -10413 12071 -10402 12074
rect -10348 12071 -10337 12074
rect -10229 12071 -10218 12074
rect -10164 12071 -10153 12074
rect -10045 12071 -10034 12074
rect -9980 12071 -9969 12074
rect -10490 12025 -10444 12036
rect -10582 11851 -10490 12025
rect -10490 11840 -10444 11851
rect -10306 12025 -10260 12036
rect -10306 11840 -10260 11851
rect -10122 12025 -10076 12036
rect -9938 12025 -9892 12036
rect -9955 11998 -9938 12000
rect -9892 11998 -9875 12000
rect -9955 11878 -9943 11998
rect -9887 11878 -9875 11998
rect -9955 11876 -9938 11878
rect -10122 11840 -10076 11851
rect -9892 11876 -9875 11878
rect -9938 11840 -9892 11851
rect -10628 11623 -10582 11768
rect -10413 11759 -10402 11805
rect -10348 11759 -10337 11805
rect -10413 11726 -10337 11759
rect -10229 11759 -10218 11805
rect -10164 11759 -10153 11805
rect -10229 11726 -10153 11759
rect -10045 11759 -10034 11805
rect -9980 11759 -9969 11805
rect -10045 11726 -9969 11759
rect -9800 11623 -9754 11768
rect -10640 11611 -10560 11623
rect -10640 11555 -10628 11611
rect -10572 11555 -10560 11611
rect -10640 11543 -10560 11555
rect -9822 11611 -9744 11623
rect -9822 11555 -9810 11611
rect -9754 11555 -9744 11611
rect -9822 11543 -9744 11555
rect -9469 11494 -9389 11504
rect -10803 11438 -9457 11494
rect -9401 11438 -9389 11494
rect -13117 11426 -13047 11438
rect -12425 10191 -12369 11438
rect -9469 11436 -9389 11438
rect -9105 11494 -9035 11506
rect -8413 11494 -8357 12224
rect -7521 12222 -7441 12224
rect -6791 12224 -6023 12280
rect -5967 12224 -5955 12280
rect -7889 12130 -7809 12144
rect -8102 12108 -8056 12119
rect -7889 12074 -7877 12130
rect -7821 12074 -7809 12130
rect -7705 12130 -7625 12144
rect -7705 12074 -7693 12130
rect -7637 12074 -7625 12130
rect -7521 12130 -7441 12144
rect -7521 12074 -7509 12130
rect -7453 12074 -7441 12130
rect -7274 12108 -7228 12119
rect -7887 12071 -7876 12074
rect -7822 12071 -7811 12074
rect -7703 12071 -7692 12074
rect -7638 12071 -7627 12074
rect -7519 12071 -7508 12074
rect -7454 12071 -7443 12074
rect -7964 12025 -7918 12036
rect -8056 11851 -7964 12025
rect -7964 11840 -7918 11851
rect -7780 12025 -7734 12036
rect -7780 11840 -7734 11851
rect -7596 12025 -7550 12036
rect -7412 12025 -7366 12036
rect -7429 11998 -7412 12000
rect -7366 11998 -7349 12000
rect -7429 11878 -7417 11998
rect -7361 11878 -7349 11998
rect -7429 11876 -7412 11878
rect -7596 11840 -7550 11851
rect -7366 11876 -7349 11878
rect -7412 11840 -7366 11851
rect -8102 11623 -8056 11768
rect -7887 11759 -7876 11805
rect -7822 11759 -7811 11805
rect -7887 11726 -7811 11759
rect -7703 11759 -7692 11805
rect -7638 11759 -7627 11805
rect -7703 11726 -7627 11759
rect -7519 11759 -7508 11805
rect -7454 11759 -7443 11805
rect -7519 11726 -7443 11759
rect -7274 11623 -7228 11768
rect -8114 11611 -8034 11623
rect -8114 11555 -8102 11611
rect -8046 11555 -8034 11611
rect -8114 11543 -8034 11555
rect -7296 11611 -7218 11623
rect -7296 11555 -7284 11611
rect -7228 11555 -7218 11611
rect -7296 11543 -7218 11555
rect -9105 11438 -9093 11494
rect -9037 11438 -8357 11494
rect -6791 11494 -6735 12224
rect -6035 12222 -5955 12224
rect -4809 12218 -4753 12340
rect -4655 12340 -4643 12396
rect -4587 12340 -3651 12396
rect -3595 12340 -3583 12396
rect -4655 12328 -4585 12340
rect -3663 12338 -3583 12340
rect -3334 12396 -3254 12398
rect -2891 12396 -2831 12406
rect -2177 12396 -2097 12398
rect -3334 12340 -3322 12396
rect -3266 12340 -2889 12396
rect -2833 12340 -2165 12396
rect -2109 12340 -2097 12396
rect -3334 12338 -3254 12340
rect -2891 12328 -2831 12340
rect -2177 12338 -2097 12340
rect -1848 12396 -1768 12398
rect -1581 12396 -1511 12408
rect -613 12396 -543 12410
rect 379 12396 459 12398
rect -1848 12340 -1836 12396
rect -1780 12340 -1579 12396
rect -1523 12340 -711 12396
rect -1848 12338 -1768 12340
rect -1581 12330 -1511 12340
rect -3479 12280 -3399 12282
rect -1993 12280 -1913 12282
rect -4371 12224 -3467 12280
rect -3411 12224 -3399 12280
rect -4821 12208 -4741 12218
rect -4821 12152 -4809 12208
rect -4753 12152 -4741 12208
rect -4821 12150 -4741 12152
rect -6403 12130 -6323 12144
rect -6616 12108 -6570 12119
rect -6403 12074 -6391 12130
rect -6335 12074 -6323 12130
rect -6219 12130 -6139 12144
rect -6219 12074 -6207 12130
rect -6151 12074 -6139 12130
rect -6035 12130 -5955 12144
rect -6035 12074 -6023 12130
rect -5967 12074 -5955 12130
rect -5788 12108 -5742 12119
rect -6401 12071 -6390 12074
rect -6336 12071 -6325 12074
rect -6217 12071 -6206 12074
rect -6152 12071 -6141 12074
rect -6033 12071 -6022 12074
rect -5968 12071 -5957 12074
rect -6478 12025 -6432 12036
rect -6570 11851 -6478 12025
rect -6478 11840 -6432 11851
rect -6294 12025 -6248 12036
rect -6294 11840 -6248 11851
rect -6110 12025 -6064 12036
rect -5926 12025 -5880 12036
rect -5943 11998 -5926 12000
rect -5880 11998 -5863 12000
rect -5943 11878 -5931 11998
rect -5875 11878 -5863 11998
rect -5943 11876 -5926 11878
rect -6110 11840 -6064 11851
rect -5880 11876 -5863 11878
rect -5926 11840 -5880 11851
rect -6616 11623 -6570 11768
rect -6401 11759 -6390 11805
rect -6336 11759 -6325 11805
rect -6401 11726 -6325 11759
rect -6217 11759 -6206 11805
rect -6152 11759 -6141 11805
rect -6217 11726 -6141 11759
rect -6033 11759 -6022 11805
rect -5968 11759 -5957 11805
rect -6033 11726 -5957 11759
rect -5788 11623 -5742 11768
rect -6628 11611 -6548 11623
rect -6628 11555 -6616 11611
rect -6560 11555 -6548 11611
rect -6628 11543 -6548 11555
rect -5810 11611 -5732 11623
rect -5810 11555 -5798 11611
rect -5742 11555 -5732 11611
rect -5810 11543 -5732 11555
rect -5457 11494 -5377 11504
rect -6791 11438 -5445 11494
rect -5389 11438 -5377 11494
rect -9105 11426 -9035 11438
rect -10945 11383 -10875 11385
rect -9645 11384 -9565 11386
rect -12289 11327 -10943 11383
rect -10887 11327 -10875 11383
rect -12289 10307 -12233 11327
rect -10945 11315 -10875 11327
rect -10803 11328 -9633 11384
rect -9577 11328 -9565 11384
rect -11625 11276 -11539 11280
rect -11625 11220 -11613 11276
rect -11557 11220 -11539 11276
rect -11625 11208 -11539 11220
rect -12114 11063 -12068 11074
rect -11899 11072 -11823 11105
rect -11899 11026 -11888 11072
rect -11834 11026 -11823 11072
rect -11715 11072 -11639 11105
rect -11715 11026 -11704 11072
rect -11650 11026 -11639 11072
rect -11531 11072 -11455 11105
rect -11531 11026 -11520 11072
rect -11466 11026 -11455 11072
rect -11286 11063 -11240 11074
rect -11976 10980 -11930 10991
rect -11993 10953 -11976 10955
rect -11792 10980 -11746 10991
rect -11930 10953 -11913 10955
rect -12068 10833 -11981 10953
rect -11925 10833 -11913 10953
rect -11993 10831 -11976 10833
rect -12068 10533 -11976 10653
rect -11930 10831 -11913 10833
rect -11809 10653 -11792 10655
rect -11608 10980 -11562 10991
rect -11625 10953 -11608 10955
rect -11424 10980 -11378 10991
rect -11562 10953 -11545 10955
rect -11625 10833 -11613 10953
rect -11557 10833 -11545 10953
rect -11625 10831 -11608 10833
rect -11746 10653 -11729 10655
rect -11809 10533 -11797 10653
rect -11741 10533 -11729 10653
rect -11809 10531 -11792 10533
rect -11976 10495 -11930 10506
rect -11746 10531 -11729 10533
rect -11792 10495 -11746 10506
rect -11562 10831 -11545 10833
rect -11441 10653 -11424 10655
rect -11303 10953 -11286 10955
rect -11240 10953 -11223 10955
rect -11303 10832 -11291 10953
rect -11235 10832 -11223 10953
rect -11303 10830 -11286 10832
rect -11378 10653 -11361 10655
rect -11441 10533 -11429 10653
rect -11373 10533 -11361 10653
rect -11441 10531 -11424 10533
rect -11608 10495 -11562 10506
rect -11378 10531 -11361 10533
rect -11424 10495 -11378 10506
rect -11899 10457 -11888 10460
rect -11834 10457 -11823 10460
rect -11715 10457 -11704 10460
rect -11650 10457 -11639 10460
rect -11531 10457 -11520 10460
rect -11466 10457 -11455 10460
rect -12114 10412 -12068 10423
rect -11901 10401 -11889 10457
rect -11833 10401 -11821 10457
rect -11901 10387 -11821 10401
rect -11717 10401 -11705 10457
rect -11649 10401 -11637 10457
rect -11717 10387 -11637 10401
rect -11533 10401 -11521 10457
rect -11465 10401 -11453 10457
rect -11240 10830 -11223 10832
rect -11286 10412 -11240 10423
rect -11533 10387 -11453 10401
rect -11901 10307 -11821 10309
rect -12289 10251 -11889 10307
rect -11833 10251 -11821 10307
rect -10803 10308 -10747 11328
rect -9645 11316 -9565 11328
rect -10139 11277 -10053 11281
rect -10139 11221 -10127 11277
rect -10071 11221 -10053 11277
rect -10139 11209 -10053 11221
rect -10628 11064 -10582 11075
rect -10413 11073 -10337 11106
rect -10413 11027 -10402 11073
rect -10348 11027 -10337 11073
rect -10229 11073 -10153 11106
rect -10229 11027 -10218 11073
rect -10164 11027 -10153 11073
rect -10045 11073 -9969 11106
rect -10045 11027 -10034 11073
rect -9980 11027 -9969 11073
rect -9800 11064 -9754 11075
rect -10490 10981 -10444 10992
rect -10507 10954 -10490 10956
rect -10306 10981 -10260 10992
rect -10444 10954 -10427 10956
rect -10582 10834 -10495 10954
rect -10439 10834 -10427 10954
rect -10507 10832 -10490 10834
rect -10582 10534 -10490 10654
rect -10444 10832 -10427 10834
rect -10323 10654 -10306 10656
rect -10122 10981 -10076 10992
rect -10139 10954 -10122 10956
rect -9938 10981 -9892 10992
rect -10076 10954 -10059 10956
rect -10139 10834 -10127 10954
rect -10071 10834 -10059 10954
rect -10139 10832 -10122 10834
rect -10260 10654 -10243 10656
rect -10323 10534 -10311 10654
rect -10255 10534 -10243 10654
rect -10323 10532 -10306 10534
rect -10490 10496 -10444 10507
rect -10260 10532 -10243 10534
rect -10306 10496 -10260 10507
rect -10076 10832 -10059 10834
rect -9955 10654 -9938 10656
rect -9817 10954 -9800 10956
rect -9754 10954 -9737 10956
rect -9817 10833 -9805 10954
rect -9749 10833 -9737 10954
rect -9817 10831 -9800 10833
rect -9892 10654 -9875 10656
rect -9955 10534 -9943 10654
rect -9887 10534 -9875 10654
rect -9955 10532 -9938 10534
rect -10122 10496 -10076 10507
rect -9892 10532 -9875 10534
rect -9938 10496 -9892 10507
rect -10413 10458 -10402 10461
rect -10348 10458 -10337 10461
rect -10229 10458 -10218 10461
rect -10164 10458 -10153 10461
rect -10045 10458 -10034 10461
rect -9980 10458 -9969 10461
rect -10628 10413 -10582 10424
rect -10415 10402 -10403 10458
rect -10347 10402 -10335 10458
rect -10415 10388 -10335 10402
rect -10231 10402 -10219 10458
rect -10163 10402 -10151 10458
rect -10231 10388 -10151 10402
rect -10047 10402 -10035 10458
rect -9979 10402 -9967 10458
rect -9754 10831 -9737 10833
rect -9800 10413 -9754 10424
rect -10047 10388 -9967 10402
rect -10415 10308 -10335 10310
rect -10803 10252 -10403 10308
rect -10347 10252 -10335 10308
rect -11901 10249 -11821 10251
rect -10415 10250 -10335 10252
rect -11717 10191 -11637 10193
rect -12425 10135 -11705 10191
rect -11649 10135 -11637 10191
rect -11717 10133 -11637 10135
rect -11388 10191 -11308 10193
rect -11121 10192 -11051 10203
rect -10231 10192 -10151 10194
rect -11121 10191 -10219 10192
rect -11388 10135 -11376 10191
rect -11320 10135 -11119 10191
rect -11063 10136 -10219 10191
rect -10163 10136 -10151 10192
rect -11063 10135 -10803 10136
rect -11388 10133 -11308 10135
rect -11121 10125 -11051 10135
rect -10231 10134 -10151 10136
rect -9902 10192 -9822 10194
rect -9459 10192 -9389 10202
rect -9902 10136 -9890 10192
rect -9834 10136 -9457 10192
rect -9401 10136 -9389 10192
rect -9902 10134 -9822 10136
rect -9459 10124 -9389 10136
rect -8413 10191 -8357 11438
rect -5457 11436 -5377 11438
rect -5093 11494 -5023 11506
rect -4371 11494 -4315 12224
rect -3479 12222 -3399 12224
rect -2749 12224 -1981 12280
rect -1925 12224 -1913 12280
rect -3847 12130 -3767 12144
rect -4060 12108 -4014 12119
rect -3847 12074 -3835 12130
rect -3779 12074 -3767 12130
rect -3663 12130 -3583 12144
rect -3663 12074 -3651 12130
rect -3595 12074 -3583 12130
rect -3479 12130 -3399 12144
rect -3479 12074 -3467 12130
rect -3411 12074 -3399 12130
rect -3232 12108 -3186 12119
rect -3845 12071 -3834 12074
rect -3780 12071 -3769 12074
rect -3661 12071 -3650 12074
rect -3596 12071 -3585 12074
rect -3477 12071 -3466 12074
rect -3412 12071 -3401 12074
rect -3922 12025 -3876 12036
rect -4014 11851 -3922 12025
rect -3922 11840 -3876 11851
rect -3738 12025 -3692 12036
rect -3738 11840 -3692 11851
rect -3554 12025 -3508 12036
rect -3370 12025 -3324 12036
rect -3387 11998 -3370 12000
rect -3324 11998 -3307 12000
rect -3387 11878 -3375 11998
rect -3319 11878 -3307 11998
rect -3387 11876 -3370 11878
rect -3554 11840 -3508 11851
rect -3324 11876 -3307 11878
rect -3370 11840 -3324 11851
rect -4060 11623 -4014 11768
rect -3845 11759 -3834 11805
rect -3780 11759 -3769 11805
rect -3845 11726 -3769 11759
rect -3661 11759 -3650 11805
rect -3596 11759 -3585 11805
rect -3661 11726 -3585 11759
rect -3477 11759 -3466 11805
rect -3412 11759 -3401 11805
rect -3477 11726 -3401 11759
rect -3232 11623 -3186 11768
rect -4072 11611 -3992 11623
rect -4072 11555 -4060 11611
rect -4004 11555 -3992 11611
rect -4072 11543 -3992 11555
rect -3254 11611 -3176 11623
rect -3254 11555 -3242 11611
rect -3186 11555 -3176 11611
rect -3254 11543 -3176 11555
rect -5093 11438 -5081 11494
rect -5025 11438 -4315 11494
rect -2749 11494 -2693 12224
rect -1993 12222 -1913 12224
rect -767 12218 -711 12340
rect -613 12340 -601 12396
rect -545 12340 391 12396
rect 447 12340 459 12396
rect -613 12328 -543 12340
rect 379 12338 459 12340
rect 708 12396 788 12398
rect 1151 12396 1211 12406
rect 1865 12396 1945 12398
rect 708 12340 720 12396
rect 776 12340 1153 12396
rect 1209 12340 1877 12396
rect 1933 12340 1945 12396
rect 708 12338 788 12340
rect 1151 12328 1211 12340
rect 1865 12338 1945 12340
rect 2194 12396 2274 12398
rect 2461 12396 2531 12408
rect 3429 12396 3499 12410
rect 4421 12396 4501 12398
rect 2194 12340 2206 12396
rect 2262 12340 2463 12396
rect 2519 12340 3331 12396
rect 2194 12338 2274 12340
rect 2461 12330 2531 12340
rect 563 12280 643 12282
rect 2049 12280 2129 12282
rect -329 12224 575 12280
rect 631 12224 643 12280
rect -779 12208 -699 12218
rect -779 12152 -767 12208
rect -711 12152 -699 12208
rect -779 12150 -699 12152
rect -2361 12130 -2281 12144
rect -2574 12108 -2528 12119
rect -2361 12074 -2349 12130
rect -2293 12074 -2281 12130
rect -2177 12130 -2097 12144
rect -2177 12074 -2165 12130
rect -2109 12074 -2097 12130
rect -1993 12130 -1913 12144
rect -1993 12074 -1981 12130
rect -1925 12074 -1913 12130
rect -1746 12108 -1700 12119
rect -2359 12071 -2348 12074
rect -2294 12071 -2283 12074
rect -2175 12071 -2164 12074
rect -2110 12071 -2099 12074
rect -1991 12071 -1980 12074
rect -1926 12071 -1915 12074
rect -2436 12025 -2390 12036
rect -2528 11851 -2436 12025
rect -2436 11840 -2390 11851
rect -2252 12025 -2206 12036
rect -2252 11840 -2206 11851
rect -2068 12025 -2022 12036
rect -1884 12025 -1838 12036
rect -1901 11998 -1884 12000
rect -1838 11998 -1821 12000
rect -1901 11878 -1889 11998
rect -1833 11878 -1821 11998
rect -1901 11876 -1884 11878
rect -2068 11840 -2022 11851
rect -1838 11876 -1821 11878
rect -1884 11840 -1838 11851
rect -2574 11623 -2528 11768
rect -2359 11759 -2348 11805
rect -2294 11759 -2283 11805
rect -2359 11726 -2283 11759
rect -2175 11759 -2164 11805
rect -2110 11759 -2099 11805
rect -2175 11726 -2099 11759
rect -1991 11759 -1980 11805
rect -1926 11759 -1915 11805
rect -1991 11726 -1915 11759
rect -1746 11623 -1700 11768
rect -2586 11611 -2506 11623
rect -2586 11555 -2574 11611
rect -2518 11555 -2506 11611
rect -2586 11543 -2506 11555
rect -1768 11611 -1690 11623
rect -1768 11555 -1756 11611
rect -1700 11555 -1690 11611
rect -1768 11543 -1690 11555
rect -1415 11494 -1335 11504
rect -2749 11438 -1403 11494
rect -1347 11438 -1335 11494
rect -5093 11426 -5023 11438
rect -6933 11383 -6863 11385
rect -5633 11384 -5553 11386
rect -8277 11327 -6931 11383
rect -6875 11327 -6863 11383
rect -8277 10307 -8221 11327
rect -6933 11315 -6863 11327
rect -6791 11328 -5621 11384
rect -5565 11328 -5553 11384
rect -7613 11276 -7527 11280
rect -7613 11220 -7601 11276
rect -7545 11220 -7527 11276
rect -7613 11208 -7527 11220
rect -8102 11063 -8056 11074
rect -7887 11072 -7811 11105
rect -7887 11026 -7876 11072
rect -7822 11026 -7811 11072
rect -7703 11072 -7627 11105
rect -7703 11026 -7692 11072
rect -7638 11026 -7627 11072
rect -7519 11072 -7443 11105
rect -7519 11026 -7508 11072
rect -7454 11026 -7443 11072
rect -7274 11063 -7228 11074
rect -7964 10980 -7918 10991
rect -7981 10953 -7964 10955
rect -7780 10980 -7734 10991
rect -7918 10953 -7901 10955
rect -8056 10833 -7969 10953
rect -7913 10833 -7901 10953
rect -7981 10831 -7964 10833
rect -8056 10533 -7964 10653
rect -7918 10831 -7901 10833
rect -7797 10653 -7780 10655
rect -7596 10980 -7550 10991
rect -7613 10953 -7596 10955
rect -7412 10980 -7366 10991
rect -7550 10953 -7533 10955
rect -7613 10833 -7601 10953
rect -7545 10833 -7533 10953
rect -7613 10831 -7596 10833
rect -7734 10653 -7717 10655
rect -7797 10533 -7785 10653
rect -7729 10533 -7717 10653
rect -7797 10531 -7780 10533
rect -7964 10495 -7918 10506
rect -7734 10531 -7717 10533
rect -7780 10495 -7734 10506
rect -7550 10831 -7533 10833
rect -7429 10653 -7412 10655
rect -7291 10953 -7274 10955
rect -7228 10953 -7211 10955
rect -7291 10832 -7279 10953
rect -7223 10832 -7211 10953
rect -7291 10830 -7274 10832
rect -7366 10653 -7349 10655
rect -7429 10533 -7417 10653
rect -7361 10533 -7349 10653
rect -7429 10531 -7412 10533
rect -7596 10495 -7550 10506
rect -7366 10531 -7349 10533
rect -7412 10495 -7366 10506
rect -7887 10457 -7876 10460
rect -7822 10457 -7811 10460
rect -7703 10457 -7692 10460
rect -7638 10457 -7627 10460
rect -7519 10457 -7508 10460
rect -7454 10457 -7443 10460
rect -8102 10412 -8056 10423
rect -7889 10401 -7877 10457
rect -7821 10401 -7809 10457
rect -7889 10387 -7809 10401
rect -7705 10401 -7693 10457
rect -7637 10401 -7625 10457
rect -7705 10387 -7625 10401
rect -7521 10401 -7509 10457
rect -7453 10401 -7441 10457
rect -7228 10830 -7211 10832
rect -7274 10412 -7228 10423
rect -7521 10387 -7441 10401
rect -7889 10307 -7809 10309
rect -8277 10251 -7877 10307
rect -7821 10251 -7809 10307
rect -6791 10308 -6735 11328
rect -5633 11316 -5553 11328
rect -6127 11277 -6041 11281
rect -6127 11221 -6115 11277
rect -6059 11221 -6041 11277
rect -6127 11209 -6041 11221
rect -6616 11064 -6570 11075
rect -6401 11073 -6325 11106
rect -6401 11027 -6390 11073
rect -6336 11027 -6325 11073
rect -6217 11073 -6141 11106
rect -6217 11027 -6206 11073
rect -6152 11027 -6141 11073
rect -6033 11073 -5957 11106
rect -6033 11027 -6022 11073
rect -5968 11027 -5957 11073
rect -5788 11064 -5742 11075
rect -6478 10981 -6432 10992
rect -6495 10954 -6478 10956
rect -6294 10981 -6248 10992
rect -6432 10954 -6415 10956
rect -6570 10834 -6483 10954
rect -6427 10834 -6415 10954
rect -6495 10832 -6478 10834
rect -6570 10534 -6478 10654
rect -6432 10832 -6415 10834
rect -6311 10654 -6294 10656
rect -6110 10981 -6064 10992
rect -6127 10954 -6110 10956
rect -5926 10981 -5880 10992
rect -6064 10954 -6047 10956
rect -6127 10834 -6115 10954
rect -6059 10834 -6047 10954
rect -6127 10832 -6110 10834
rect -6248 10654 -6231 10656
rect -6311 10534 -6299 10654
rect -6243 10534 -6231 10654
rect -6311 10532 -6294 10534
rect -6478 10496 -6432 10507
rect -6248 10532 -6231 10534
rect -6294 10496 -6248 10507
rect -6064 10832 -6047 10834
rect -5943 10654 -5926 10656
rect -5805 10954 -5788 10956
rect -5742 10954 -5725 10956
rect -5805 10833 -5793 10954
rect -5737 10833 -5725 10954
rect -5805 10831 -5788 10833
rect -5880 10654 -5863 10656
rect -5943 10534 -5931 10654
rect -5875 10534 -5863 10654
rect -5943 10532 -5926 10534
rect -6110 10496 -6064 10507
rect -5880 10532 -5863 10534
rect -5926 10496 -5880 10507
rect -6401 10458 -6390 10461
rect -6336 10458 -6325 10461
rect -6217 10458 -6206 10461
rect -6152 10458 -6141 10461
rect -6033 10458 -6022 10461
rect -5968 10458 -5957 10461
rect -6616 10413 -6570 10424
rect -6403 10402 -6391 10458
rect -6335 10402 -6323 10458
rect -6403 10388 -6323 10402
rect -6219 10402 -6207 10458
rect -6151 10402 -6139 10458
rect -6219 10388 -6139 10402
rect -6035 10402 -6023 10458
rect -5967 10402 -5955 10458
rect -5742 10831 -5725 10833
rect -5788 10413 -5742 10424
rect -6035 10388 -5955 10402
rect -6403 10308 -6323 10310
rect -6791 10252 -6391 10308
rect -6335 10252 -6323 10308
rect -7889 10249 -7809 10251
rect -6403 10250 -6323 10252
rect -7705 10191 -7625 10193
rect -8413 10135 -7693 10191
rect -7637 10135 -7625 10191
rect -7705 10133 -7625 10135
rect -7376 10191 -7296 10193
rect -7109 10192 -7039 10203
rect -6219 10192 -6139 10194
rect -7109 10191 -6207 10192
rect -7376 10135 -7364 10191
rect -7308 10135 -7107 10191
rect -7051 10136 -6207 10191
rect -6151 10136 -6139 10192
rect -7051 10135 -6791 10136
rect -7376 10133 -7296 10135
rect -7109 10125 -7039 10135
rect -6219 10134 -6139 10136
rect -5890 10192 -5810 10194
rect -5447 10192 -5377 10202
rect -5890 10136 -5878 10192
rect -5822 10136 -5445 10192
rect -5389 10136 -5377 10192
rect -5890 10134 -5810 10136
rect -5447 10124 -5377 10136
rect -4371 10191 -4315 11438
rect -1415 11436 -1335 11438
rect -1051 11494 -981 11506
rect -329 11494 -273 12224
rect 563 12222 643 12224
rect 1293 12224 2061 12280
rect 2117 12224 2129 12280
rect 195 12130 275 12144
rect -18 12108 28 12119
rect 195 12074 207 12130
rect 263 12074 275 12130
rect 379 12130 459 12144
rect 379 12074 391 12130
rect 447 12074 459 12130
rect 563 12130 643 12144
rect 563 12074 575 12130
rect 631 12074 643 12130
rect 810 12108 856 12119
rect 197 12071 208 12074
rect 262 12071 273 12074
rect 381 12071 392 12074
rect 446 12071 457 12074
rect 565 12071 576 12074
rect 630 12071 641 12074
rect 120 12025 166 12036
rect 28 11851 120 12025
rect 120 11840 166 11851
rect 304 12025 350 12036
rect 304 11840 350 11851
rect 488 12025 534 12036
rect 672 12025 718 12036
rect 655 11998 672 12000
rect 718 11998 735 12000
rect 655 11878 667 11998
rect 723 11878 735 11998
rect 655 11876 672 11878
rect 488 11840 534 11851
rect 718 11876 735 11878
rect 672 11840 718 11851
rect -18 11623 28 11768
rect 197 11759 208 11805
rect 262 11759 273 11805
rect 197 11726 273 11759
rect 381 11759 392 11805
rect 446 11759 457 11805
rect 381 11726 457 11759
rect 565 11759 576 11805
rect 630 11759 641 11805
rect 565 11726 641 11759
rect 810 11623 856 11768
rect -30 11611 50 11623
rect -30 11555 -18 11611
rect 38 11555 50 11611
rect -30 11543 50 11555
rect 788 11611 866 11623
rect 788 11555 800 11611
rect 856 11555 866 11611
rect 788 11543 866 11555
rect -1051 11438 -1039 11494
rect -983 11438 -273 11494
rect 1293 11494 1349 12224
rect 2049 12222 2129 12224
rect 3275 12218 3331 12340
rect 3429 12340 3441 12396
rect 3497 12340 4433 12396
rect 4489 12340 4501 12396
rect 3429 12328 3499 12340
rect 4421 12338 4501 12340
rect 4750 12396 4830 12398
rect 5193 12396 5253 12406
rect 5907 12396 5987 12398
rect 4750 12340 4762 12396
rect 4818 12340 5195 12396
rect 5251 12340 5919 12396
rect 5975 12340 5987 12396
rect 4750 12338 4830 12340
rect 5193 12328 5253 12340
rect 5907 12338 5987 12340
rect 6236 12396 6316 12398
rect 6503 12396 6573 12408
rect 7471 12396 7541 12410
rect 8463 12396 8543 12398
rect 6236 12340 6248 12396
rect 6304 12340 6505 12396
rect 6561 12340 7373 12396
rect 6236 12338 6316 12340
rect 6503 12330 6573 12340
rect 4605 12280 4685 12282
rect 6091 12280 6171 12282
rect 3713 12224 4617 12280
rect 4673 12224 4685 12280
rect 3263 12208 3343 12218
rect 3263 12152 3275 12208
rect 3331 12152 3343 12208
rect 3263 12150 3343 12152
rect 1681 12130 1761 12144
rect 1468 12108 1514 12119
rect 1681 12074 1693 12130
rect 1749 12074 1761 12130
rect 1865 12130 1945 12144
rect 1865 12074 1877 12130
rect 1933 12074 1945 12130
rect 2049 12130 2129 12144
rect 2049 12074 2061 12130
rect 2117 12074 2129 12130
rect 2296 12108 2342 12119
rect 1683 12071 1694 12074
rect 1748 12071 1759 12074
rect 1867 12071 1878 12074
rect 1932 12071 1943 12074
rect 2051 12071 2062 12074
rect 2116 12071 2127 12074
rect 1606 12025 1652 12036
rect 1514 11851 1606 12025
rect 1606 11840 1652 11851
rect 1790 12025 1836 12036
rect 1790 11840 1836 11851
rect 1974 12025 2020 12036
rect 2158 12025 2204 12036
rect 2141 11998 2158 12000
rect 2204 11998 2221 12000
rect 2141 11878 2153 11998
rect 2209 11878 2221 11998
rect 2141 11876 2158 11878
rect 1974 11840 2020 11851
rect 2204 11876 2221 11878
rect 2158 11840 2204 11851
rect 1468 11623 1514 11768
rect 1683 11759 1694 11805
rect 1748 11759 1759 11805
rect 1683 11726 1759 11759
rect 1867 11759 1878 11805
rect 1932 11759 1943 11805
rect 1867 11726 1943 11759
rect 2051 11759 2062 11805
rect 2116 11759 2127 11805
rect 2051 11726 2127 11759
rect 2296 11623 2342 11768
rect 1456 11611 1536 11623
rect 1456 11555 1468 11611
rect 1524 11555 1536 11611
rect 1456 11543 1536 11555
rect 2274 11611 2352 11623
rect 2274 11555 2286 11611
rect 2342 11555 2352 11611
rect 2274 11543 2352 11555
rect 2627 11494 2707 11504
rect 1293 11438 2639 11494
rect 2695 11438 2707 11494
rect -1051 11426 -981 11438
rect -2891 11383 -2821 11385
rect -1591 11384 -1511 11386
rect -4235 11327 -2889 11383
rect -2833 11327 -2821 11383
rect -4235 10307 -4179 11327
rect -2891 11315 -2821 11327
rect -2749 11328 -1579 11384
rect -1523 11328 -1511 11384
rect -3571 11276 -3485 11280
rect -3571 11220 -3559 11276
rect -3503 11220 -3485 11276
rect -3571 11208 -3485 11220
rect -4060 11063 -4014 11074
rect -3845 11072 -3769 11105
rect -3845 11026 -3834 11072
rect -3780 11026 -3769 11072
rect -3661 11072 -3585 11105
rect -3661 11026 -3650 11072
rect -3596 11026 -3585 11072
rect -3477 11072 -3401 11105
rect -3477 11026 -3466 11072
rect -3412 11026 -3401 11072
rect -3232 11063 -3186 11074
rect -3922 10980 -3876 10991
rect -3939 10953 -3922 10955
rect -3738 10980 -3692 10991
rect -3876 10953 -3859 10955
rect -4014 10833 -3927 10953
rect -3871 10833 -3859 10953
rect -3939 10831 -3922 10833
rect -4014 10533 -3922 10653
rect -3876 10831 -3859 10833
rect -3755 10653 -3738 10655
rect -3554 10980 -3508 10991
rect -3571 10953 -3554 10955
rect -3370 10980 -3324 10991
rect -3508 10953 -3491 10955
rect -3571 10833 -3559 10953
rect -3503 10833 -3491 10953
rect -3571 10831 -3554 10833
rect -3692 10653 -3675 10655
rect -3755 10533 -3743 10653
rect -3687 10533 -3675 10653
rect -3755 10531 -3738 10533
rect -3922 10495 -3876 10506
rect -3692 10531 -3675 10533
rect -3738 10495 -3692 10506
rect -3508 10831 -3491 10833
rect -3387 10653 -3370 10655
rect -3249 10953 -3232 10955
rect -3186 10953 -3169 10955
rect -3249 10832 -3237 10953
rect -3181 10832 -3169 10953
rect -3249 10830 -3232 10832
rect -3324 10653 -3307 10655
rect -3387 10533 -3375 10653
rect -3319 10533 -3307 10653
rect -3387 10531 -3370 10533
rect -3554 10495 -3508 10506
rect -3324 10531 -3307 10533
rect -3370 10495 -3324 10506
rect -3845 10457 -3834 10460
rect -3780 10457 -3769 10460
rect -3661 10457 -3650 10460
rect -3596 10457 -3585 10460
rect -3477 10457 -3466 10460
rect -3412 10457 -3401 10460
rect -4060 10412 -4014 10423
rect -3847 10401 -3835 10457
rect -3779 10401 -3767 10457
rect -3847 10387 -3767 10401
rect -3663 10401 -3651 10457
rect -3595 10401 -3583 10457
rect -3663 10387 -3583 10401
rect -3479 10401 -3467 10457
rect -3411 10401 -3399 10457
rect -3186 10830 -3169 10832
rect -3232 10412 -3186 10423
rect -3479 10387 -3399 10401
rect -3847 10307 -3767 10309
rect -4235 10251 -3835 10307
rect -3779 10251 -3767 10307
rect -2749 10308 -2693 11328
rect -1591 11316 -1511 11328
rect -2085 11277 -1999 11281
rect -2085 11221 -2073 11277
rect -2017 11221 -1999 11277
rect -2085 11209 -1999 11221
rect -2574 11064 -2528 11075
rect -2359 11073 -2283 11106
rect -2359 11027 -2348 11073
rect -2294 11027 -2283 11073
rect -2175 11073 -2099 11106
rect -2175 11027 -2164 11073
rect -2110 11027 -2099 11073
rect -1991 11073 -1915 11106
rect -1991 11027 -1980 11073
rect -1926 11027 -1915 11073
rect -1746 11064 -1700 11075
rect -2436 10981 -2390 10992
rect -2453 10954 -2436 10956
rect -2252 10981 -2206 10992
rect -2390 10954 -2373 10956
rect -2528 10834 -2441 10954
rect -2385 10834 -2373 10954
rect -2453 10832 -2436 10834
rect -2528 10534 -2436 10654
rect -2390 10832 -2373 10834
rect -2269 10654 -2252 10656
rect -2068 10981 -2022 10992
rect -2085 10954 -2068 10956
rect -1884 10981 -1838 10992
rect -2022 10954 -2005 10956
rect -2085 10834 -2073 10954
rect -2017 10834 -2005 10954
rect -2085 10832 -2068 10834
rect -2206 10654 -2189 10656
rect -2269 10534 -2257 10654
rect -2201 10534 -2189 10654
rect -2269 10532 -2252 10534
rect -2436 10496 -2390 10507
rect -2206 10532 -2189 10534
rect -2252 10496 -2206 10507
rect -2022 10832 -2005 10834
rect -1901 10654 -1884 10656
rect -1763 10954 -1746 10956
rect -1700 10954 -1683 10956
rect -1763 10833 -1751 10954
rect -1695 10833 -1683 10954
rect -1763 10831 -1746 10833
rect -1838 10654 -1821 10656
rect -1901 10534 -1889 10654
rect -1833 10534 -1821 10654
rect -1901 10532 -1884 10534
rect -2068 10496 -2022 10507
rect -1838 10532 -1821 10534
rect -1884 10496 -1838 10507
rect -2359 10458 -2348 10461
rect -2294 10458 -2283 10461
rect -2175 10458 -2164 10461
rect -2110 10458 -2099 10461
rect -1991 10458 -1980 10461
rect -1926 10458 -1915 10461
rect -2574 10413 -2528 10424
rect -2361 10402 -2349 10458
rect -2293 10402 -2281 10458
rect -2361 10388 -2281 10402
rect -2177 10402 -2165 10458
rect -2109 10402 -2097 10458
rect -2177 10388 -2097 10402
rect -1993 10402 -1981 10458
rect -1925 10402 -1913 10458
rect -1700 10831 -1683 10833
rect -1746 10413 -1700 10424
rect -1993 10388 -1913 10402
rect -2361 10308 -2281 10310
rect -2749 10252 -2349 10308
rect -2293 10252 -2281 10308
rect -3847 10249 -3767 10251
rect -2361 10250 -2281 10252
rect -3663 10191 -3583 10193
rect -4371 10135 -3651 10191
rect -3595 10135 -3583 10191
rect -3663 10133 -3583 10135
rect -3334 10191 -3254 10193
rect -3067 10192 -2997 10203
rect -2177 10192 -2097 10194
rect -3067 10191 -2165 10192
rect -3334 10135 -3322 10191
rect -3266 10135 -3065 10191
rect -3009 10136 -2165 10191
rect -2109 10136 -2097 10192
rect -3009 10135 -2749 10136
rect -3334 10133 -3254 10135
rect -3067 10125 -2997 10135
rect -2177 10134 -2097 10136
rect -1848 10192 -1768 10194
rect -1405 10192 -1335 10202
rect -1848 10136 -1836 10192
rect -1780 10136 -1403 10192
rect -1347 10136 -1335 10192
rect -1848 10134 -1768 10136
rect -1405 10124 -1335 10136
rect -329 10191 -273 11438
rect 2627 11436 2707 11438
rect 2991 11494 3061 11506
rect 3713 11494 3769 12224
rect 4605 12222 4685 12224
rect 5335 12224 6103 12280
rect 6159 12224 6171 12280
rect 4237 12130 4317 12144
rect 4024 12108 4070 12119
rect 4237 12074 4249 12130
rect 4305 12074 4317 12130
rect 4421 12130 4501 12144
rect 4421 12074 4433 12130
rect 4489 12074 4501 12130
rect 4605 12130 4685 12144
rect 4605 12074 4617 12130
rect 4673 12074 4685 12130
rect 4852 12108 4898 12119
rect 4239 12071 4250 12074
rect 4304 12071 4315 12074
rect 4423 12071 4434 12074
rect 4488 12071 4499 12074
rect 4607 12071 4618 12074
rect 4672 12071 4683 12074
rect 4162 12025 4208 12036
rect 4070 11851 4162 12025
rect 4162 11840 4208 11851
rect 4346 12025 4392 12036
rect 4346 11840 4392 11851
rect 4530 12025 4576 12036
rect 4714 12025 4760 12036
rect 4697 11998 4714 12000
rect 4760 11998 4777 12000
rect 4697 11878 4709 11998
rect 4765 11878 4777 11998
rect 4697 11876 4714 11878
rect 4530 11840 4576 11851
rect 4760 11876 4777 11878
rect 4714 11840 4760 11851
rect 4024 11623 4070 11768
rect 4239 11759 4250 11805
rect 4304 11759 4315 11805
rect 4239 11726 4315 11759
rect 4423 11759 4434 11805
rect 4488 11759 4499 11805
rect 4423 11726 4499 11759
rect 4607 11759 4618 11805
rect 4672 11759 4683 11805
rect 4607 11726 4683 11759
rect 4852 11623 4898 11768
rect 4012 11611 4092 11623
rect 4012 11555 4024 11611
rect 4080 11555 4092 11611
rect 4012 11543 4092 11555
rect 4830 11611 4908 11623
rect 4830 11555 4842 11611
rect 4898 11555 4908 11611
rect 4830 11543 4908 11555
rect 2991 11438 3003 11494
rect 3059 11438 3769 11494
rect 5335 11494 5391 12224
rect 6091 12222 6171 12224
rect 7317 12218 7373 12340
rect 7471 12340 7483 12396
rect 7539 12340 8475 12396
rect 8531 12340 8543 12396
rect 7471 12328 7541 12340
rect 8463 12338 8543 12340
rect 8792 12396 8872 12398
rect 9235 12396 9295 12406
rect 9949 12396 10029 12398
rect 8792 12340 8804 12396
rect 8860 12340 9237 12396
rect 9293 12340 9961 12396
rect 10017 12340 10029 12396
rect 8792 12338 8872 12340
rect 9235 12328 9295 12340
rect 9949 12338 10029 12340
rect 10278 12396 10358 12398
rect 10545 12396 10615 12408
rect 11513 12396 11583 12410
rect 12505 12396 12585 12398
rect 10278 12340 10290 12396
rect 10346 12340 10547 12396
rect 10603 12340 11415 12396
rect 10278 12338 10358 12340
rect 10545 12330 10615 12340
rect 8647 12280 8727 12282
rect 10133 12280 10213 12282
rect 7755 12224 8659 12280
rect 8715 12224 8727 12280
rect 7305 12208 7385 12218
rect 7305 12152 7317 12208
rect 7373 12152 7385 12208
rect 7305 12150 7385 12152
rect 5723 12130 5803 12144
rect 5510 12108 5556 12119
rect 5723 12074 5735 12130
rect 5791 12074 5803 12130
rect 5907 12130 5987 12144
rect 5907 12074 5919 12130
rect 5975 12074 5987 12130
rect 6091 12130 6171 12144
rect 6091 12074 6103 12130
rect 6159 12074 6171 12130
rect 6338 12108 6384 12119
rect 5725 12071 5736 12074
rect 5790 12071 5801 12074
rect 5909 12071 5920 12074
rect 5974 12071 5985 12074
rect 6093 12071 6104 12074
rect 6158 12071 6169 12074
rect 5648 12025 5694 12036
rect 5556 11851 5648 12025
rect 5648 11840 5694 11851
rect 5832 12025 5878 12036
rect 5832 11840 5878 11851
rect 6016 12025 6062 12036
rect 6200 12025 6246 12036
rect 6183 11998 6200 12000
rect 6246 11998 6263 12000
rect 6183 11878 6195 11998
rect 6251 11878 6263 11998
rect 6183 11876 6200 11878
rect 6016 11840 6062 11851
rect 6246 11876 6263 11878
rect 6200 11840 6246 11851
rect 5510 11623 5556 11768
rect 5725 11759 5736 11805
rect 5790 11759 5801 11805
rect 5725 11726 5801 11759
rect 5909 11759 5920 11805
rect 5974 11759 5985 11805
rect 5909 11726 5985 11759
rect 6093 11759 6104 11805
rect 6158 11759 6169 11805
rect 6093 11726 6169 11759
rect 6338 11623 6384 11768
rect 5498 11611 5578 11623
rect 5498 11555 5510 11611
rect 5566 11555 5578 11611
rect 5498 11543 5578 11555
rect 6316 11611 6394 11623
rect 6316 11555 6328 11611
rect 6384 11555 6394 11611
rect 6316 11543 6394 11555
rect 6669 11494 6749 11504
rect 5335 11438 6681 11494
rect 6737 11438 6749 11494
rect 2991 11426 3061 11438
rect 1151 11383 1221 11385
rect 2451 11384 2531 11386
rect -193 11327 1153 11383
rect 1209 11327 1221 11383
rect -193 10307 -137 11327
rect 1151 11315 1221 11327
rect 1293 11328 2463 11384
rect 2519 11328 2531 11384
rect 471 11276 557 11280
rect 471 11220 483 11276
rect 539 11220 557 11276
rect 471 11208 557 11220
rect -18 11063 28 11074
rect 197 11072 273 11105
rect 197 11026 208 11072
rect 262 11026 273 11072
rect 381 11072 457 11105
rect 381 11026 392 11072
rect 446 11026 457 11072
rect 565 11072 641 11105
rect 565 11026 576 11072
rect 630 11026 641 11072
rect 810 11063 856 11074
rect 120 10980 166 10991
rect 103 10953 120 10955
rect 304 10980 350 10991
rect 166 10953 183 10955
rect 28 10833 115 10953
rect 171 10833 183 10953
rect 103 10831 120 10833
rect 28 10533 120 10653
rect 166 10831 183 10833
rect 287 10653 304 10655
rect 488 10980 534 10991
rect 471 10953 488 10955
rect 672 10980 718 10991
rect 534 10953 551 10955
rect 471 10833 483 10953
rect 539 10833 551 10953
rect 471 10831 488 10833
rect 350 10653 367 10655
rect 287 10533 299 10653
rect 355 10533 367 10653
rect 287 10531 304 10533
rect 120 10495 166 10506
rect 350 10531 367 10533
rect 304 10495 350 10506
rect 534 10831 551 10833
rect 655 10653 672 10655
rect 793 10953 810 10955
rect 856 10953 873 10955
rect 793 10832 805 10953
rect 861 10832 873 10953
rect 793 10830 810 10832
rect 718 10653 735 10655
rect 655 10533 667 10653
rect 723 10533 735 10653
rect 655 10531 672 10533
rect 488 10495 534 10506
rect 718 10531 735 10533
rect 672 10495 718 10506
rect 197 10457 208 10460
rect 262 10457 273 10460
rect 381 10457 392 10460
rect 446 10457 457 10460
rect 565 10457 576 10460
rect 630 10457 641 10460
rect -18 10412 28 10423
rect 195 10401 207 10457
rect 263 10401 275 10457
rect 195 10387 275 10401
rect 379 10401 391 10457
rect 447 10401 459 10457
rect 379 10387 459 10401
rect 563 10401 575 10457
rect 631 10401 643 10457
rect 856 10830 873 10832
rect 810 10412 856 10423
rect 563 10387 643 10401
rect 195 10307 275 10309
rect -193 10251 207 10307
rect 263 10251 275 10307
rect 1293 10308 1349 11328
rect 2451 11316 2531 11328
rect 1957 11277 2043 11281
rect 1957 11221 1969 11277
rect 2025 11221 2043 11277
rect 1957 11209 2043 11221
rect 1468 11064 1514 11075
rect 1683 11073 1759 11106
rect 1683 11027 1694 11073
rect 1748 11027 1759 11073
rect 1867 11073 1943 11106
rect 1867 11027 1878 11073
rect 1932 11027 1943 11073
rect 2051 11073 2127 11106
rect 2051 11027 2062 11073
rect 2116 11027 2127 11073
rect 2296 11064 2342 11075
rect 1606 10981 1652 10992
rect 1589 10954 1606 10956
rect 1790 10981 1836 10992
rect 1652 10954 1669 10956
rect 1514 10834 1601 10954
rect 1657 10834 1669 10954
rect 1589 10832 1606 10834
rect 1514 10534 1606 10654
rect 1652 10832 1669 10834
rect 1773 10654 1790 10656
rect 1974 10981 2020 10992
rect 1957 10954 1974 10956
rect 2158 10981 2204 10992
rect 2020 10954 2037 10956
rect 1957 10834 1969 10954
rect 2025 10834 2037 10954
rect 1957 10832 1974 10834
rect 1836 10654 1853 10656
rect 1773 10534 1785 10654
rect 1841 10534 1853 10654
rect 1773 10532 1790 10534
rect 1606 10496 1652 10507
rect 1836 10532 1853 10534
rect 1790 10496 1836 10507
rect 2020 10832 2037 10834
rect 2141 10654 2158 10656
rect 2279 10954 2296 10956
rect 2342 10954 2359 10956
rect 2279 10833 2291 10954
rect 2347 10833 2359 10954
rect 2279 10831 2296 10833
rect 2204 10654 2221 10656
rect 2141 10534 2153 10654
rect 2209 10534 2221 10654
rect 2141 10532 2158 10534
rect 1974 10496 2020 10507
rect 2204 10532 2221 10534
rect 2158 10496 2204 10507
rect 1683 10458 1694 10461
rect 1748 10458 1759 10461
rect 1867 10458 1878 10461
rect 1932 10458 1943 10461
rect 2051 10458 2062 10461
rect 2116 10458 2127 10461
rect 1468 10413 1514 10424
rect 1681 10402 1693 10458
rect 1749 10402 1761 10458
rect 1681 10388 1761 10402
rect 1865 10402 1877 10458
rect 1933 10402 1945 10458
rect 1865 10388 1945 10402
rect 2049 10402 2061 10458
rect 2117 10402 2129 10458
rect 2342 10831 2359 10833
rect 2296 10413 2342 10424
rect 2049 10388 2129 10402
rect 1681 10308 1761 10310
rect 1293 10252 1693 10308
rect 1749 10252 1761 10308
rect 195 10249 275 10251
rect 1681 10250 1761 10252
rect 379 10191 459 10193
rect -329 10135 391 10191
rect 447 10135 459 10191
rect 379 10133 459 10135
rect 708 10191 788 10193
rect 975 10192 1045 10203
rect 1865 10192 1945 10194
rect 975 10191 1877 10192
rect 708 10135 720 10191
rect 776 10135 977 10191
rect 1033 10136 1877 10191
rect 1933 10136 1945 10192
rect 1033 10135 1293 10136
rect 708 10133 788 10135
rect 975 10125 1045 10135
rect 1865 10134 1945 10136
rect 2194 10192 2274 10194
rect 2637 10192 2707 10202
rect 2194 10136 2206 10192
rect 2262 10136 2639 10192
rect 2695 10136 2707 10192
rect 2194 10134 2274 10136
rect 2637 10124 2707 10136
rect 3713 10191 3769 11438
rect 6669 11436 6749 11438
rect 7033 11494 7103 11506
rect 7755 11494 7811 12224
rect 8647 12222 8727 12224
rect 9377 12224 10145 12280
rect 10201 12224 10213 12280
rect 8279 12130 8359 12144
rect 8066 12108 8112 12119
rect 8279 12074 8291 12130
rect 8347 12074 8359 12130
rect 8463 12130 8543 12144
rect 8463 12074 8475 12130
rect 8531 12074 8543 12130
rect 8647 12130 8727 12144
rect 8647 12074 8659 12130
rect 8715 12074 8727 12130
rect 8894 12108 8940 12119
rect 8281 12071 8292 12074
rect 8346 12071 8357 12074
rect 8465 12071 8476 12074
rect 8530 12071 8541 12074
rect 8649 12071 8660 12074
rect 8714 12071 8725 12074
rect 8204 12025 8250 12036
rect 8112 11851 8204 12025
rect 8204 11840 8250 11851
rect 8388 12025 8434 12036
rect 8388 11840 8434 11851
rect 8572 12025 8618 12036
rect 8756 12025 8802 12036
rect 8739 11998 8756 12000
rect 8802 11998 8819 12000
rect 8739 11878 8751 11998
rect 8807 11878 8819 11998
rect 8739 11876 8756 11878
rect 8572 11840 8618 11851
rect 8802 11876 8819 11878
rect 8756 11840 8802 11851
rect 8066 11623 8112 11768
rect 8281 11759 8292 11805
rect 8346 11759 8357 11805
rect 8281 11726 8357 11759
rect 8465 11759 8476 11805
rect 8530 11759 8541 11805
rect 8465 11726 8541 11759
rect 8649 11759 8660 11805
rect 8714 11759 8725 11805
rect 8649 11726 8725 11759
rect 8894 11623 8940 11768
rect 8054 11611 8134 11623
rect 8054 11555 8066 11611
rect 8122 11555 8134 11611
rect 8054 11543 8134 11555
rect 8872 11611 8950 11623
rect 8872 11555 8884 11611
rect 8940 11555 8950 11611
rect 8872 11543 8950 11555
rect 7033 11438 7045 11494
rect 7101 11438 7811 11494
rect 9377 11494 9433 12224
rect 10133 12222 10213 12224
rect 11359 12218 11415 12340
rect 11513 12340 11525 12396
rect 11581 12340 12517 12396
rect 12573 12340 12585 12396
rect 11513 12328 11583 12340
rect 12505 12338 12585 12340
rect 12834 12396 12914 12398
rect 13277 12396 13337 12406
rect 13991 12396 14071 12398
rect 12834 12340 12846 12396
rect 12902 12340 13279 12396
rect 13335 12340 14003 12396
rect 14059 12340 14071 12396
rect 12834 12338 12914 12340
rect 13277 12328 13337 12340
rect 13991 12338 14071 12340
rect 14320 12396 14400 12398
rect 14587 12396 14657 12408
rect 14320 12340 14332 12396
rect 14388 12340 14589 12396
rect 14645 12340 14657 12396
rect 14320 12338 14400 12340
rect 14587 12330 14657 12340
rect 12689 12280 12769 12282
rect 14175 12280 14255 12282
rect 11797 12224 12701 12280
rect 12757 12224 12769 12280
rect 11347 12208 11427 12218
rect 11347 12152 11359 12208
rect 11415 12152 11427 12208
rect 11347 12150 11427 12152
rect 9765 12130 9845 12144
rect 9552 12108 9598 12119
rect 9765 12074 9777 12130
rect 9833 12074 9845 12130
rect 9949 12130 10029 12144
rect 9949 12074 9961 12130
rect 10017 12074 10029 12130
rect 10133 12130 10213 12144
rect 10133 12074 10145 12130
rect 10201 12074 10213 12130
rect 10380 12108 10426 12119
rect 9767 12071 9778 12074
rect 9832 12071 9843 12074
rect 9951 12071 9962 12074
rect 10016 12071 10027 12074
rect 10135 12071 10146 12074
rect 10200 12071 10211 12074
rect 9690 12025 9736 12036
rect 9598 11851 9690 12025
rect 9690 11840 9736 11851
rect 9874 12025 9920 12036
rect 9874 11840 9920 11851
rect 10058 12025 10104 12036
rect 10242 12025 10288 12036
rect 10225 11998 10242 12000
rect 10288 11998 10305 12000
rect 10225 11878 10237 11998
rect 10293 11878 10305 11998
rect 10225 11876 10242 11878
rect 10058 11840 10104 11851
rect 10288 11876 10305 11878
rect 10242 11840 10288 11851
rect 9552 11623 9598 11768
rect 9767 11759 9778 11805
rect 9832 11759 9843 11805
rect 9767 11726 9843 11759
rect 9951 11759 9962 11805
rect 10016 11759 10027 11805
rect 9951 11726 10027 11759
rect 10135 11759 10146 11805
rect 10200 11759 10211 11805
rect 10135 11726 10211 11759
rect 10380 11623 10426 11768
rect 9540 11611 9620 11623
rect 9540 11555 9552 11611
rect 9608 11555 9620 11611
rect 9540 11543 9620 11555
rect 10358 11611 10436 11623
rect 10358 11555 10370 11611
rect 10426 11555 10436 11611
rect 10358 11543 10436 11555
rect 10711 11494 10791 11504
rect 9377 11438 10723 11494
rect 10779 11438 10791 11494
rect 7033 11426 7103 11438
rect 5193 11383 5263 11385
rect 6493 11384 6573 11386
rect 3849 11327 5195 11383
rect 5251 11327 5263 11383
rect 3849 10307 3905 11327
rect 5193 11315 5263 11327
rect 5335 11328 6505 11384
rect 6561 11328 6573 11384
rect 4513 11276 4599 11280
rect 4513 11220 4525 11276
rect 4581 11220 4599 11276
rect 4513 11208 4599 11220
rect 4024 11063 4070 11074
rect 4239 11072 4315 11105
rect 4239 11026 4250 11072
rect 4304 11026 4315 11072
rect 4423 11072 4499 11105
rect 4423 11026 4434 11072
rect 4488 11026 4499 11072
rect 4607 11072 4683 11105
rect 4607 11026 4618 11072
rect 4672 11026 4683 11072
rect 4852 11063 4898 11074
rect 4162 10980 4208 10991
rect 4145 10953 4162 10955
rect 4346 10980 4392 10991
rect 4208 10953 4225 10955
rect 4070 10833 4157 10953
rect 4213 10833 4225 10953
rect 4145 10831 4162 10833
rect 4070 10533 4162 10653
rect 4208 10831 4225 10833
rect 4329 10653 4346 10655
rect 4530 10980 4576 10991
rect 4513 10953 4530 10955
rect 4714 10980 4760 10991
rect 4576 10953 4593 10955
rect 4513 10833 4525 10953
rect 4581 10833 4593 10953
rect 4513 10831 4530 10833
rect 4392 10653 4409 10655
rect 4329 10533 4341 10653
rect 4397 10533 4409 10653
rect 4329 10531 4346 10533
rect 4162 10495 4208 10506
rect 4392 10531 4409 10533
rect 4346 10495 4392 10506
rect 4576 10831 4593 10833
rect 4697 10653 4714 10655
rect 4835 10953 4852 10955
rect 4898 10953 4915 10955
rect 4835 10832 4847 10953
rect 4903 10832 4915 10953
rect 4835 10830 4852 10832
rect 4760 10653 4777 10655
rect 4697 10533 4709 10653
rect 4765 10533 4777 10653
rect 4697 10531 4714 10533
rect 4530 10495 4576 10506
rect 4760 10531 4777 10533
rect 4714 10495 4760 10506
rect 4239 10457 4250 10460
rect 4304 10457 4315 10460
rect 4423 10457 4434 10460
rect 4488 10457 4499 10460
rect 4607 10457 4618 10460
rect 4672 10457 4683 10460
rect 4024 10412 4070 10423
rect 4237 10401 4249 10457
rect 4305 10401 4317 10457
rect 4237 10387 4317 10401
rect 4421 10401 4433 10457
rect 4489 10401 4501 10457
rect 4421 10387 4501 10401
rect 4605 10401 4617 10457
rect 4673 10401 4685 10457
rect 4898 10830 4915 10832
rect 4852 10412 4898 10423
rect 4605 10387 4685 10401
rect 4237 10307 4317 10309
rect 3849 10251 4249 10307
rect 4305 10251 4317 10307
rect 5335 10308 5391 11328
rect 6493 11316 6573 11328
rect 5999 11277 6085 11281
rect 5999 11221 6011 11277
rect 6067 11221 6085 11277
rect 5999 11209 6085 11221
rect 5510 11064 5556 11075
rect 5725 11073 5801 11106
rect 5725 11027 5736 11073
rect 5790 11027 5801 11073
rect 5909 11073 5985 11106
rect 5909 11027 5920 11073
rect 5974 11027 5985 11073
rect 6093 11073 6169 11106
rect 6093 11027 6104 11073
rect 6158 11027 6169 11073
rect 6338 11064 6384 11075
rect 5648 10981 5694 10992
rect 5631 10954 5648 10956
rect 5832 10981 5878 10992
rect 5694 10954 5711 10956
rect 5556 10834 5643 10954
rect 5699 10834 5711 10954
rect 5631 10832 5648 10834
rect 5556 10534 5648 10654
rect 5694 10832 5711 10834
rect 5815 10654 5832 10656
rect 6016 10981 6062 10992
rect 5999 10954 6016 10956
rect 6200 10981 6246 10992
rect 6062 10954 6079 10956
rect 5999 10834 6011 10954
rect 6067 10834 6079 10954
rect 5999 10832 6016 10834
rect 5878 10654 5895 10656
rect 5815 10534 5827 10654
rect 5883 10534 5895 10654
rect 5815 10532 5832 10534
rect 5648 10496 5694 10507
rect 5878 10532 5895 10534
rect 5832 10496 5878 10507
rect 6062 10832 6079 10834
rect 6183 10654 6200 10656
rect 6321 10954 6338 10956
rect 6384 10954 6401 10956
rect 6321 10833 6333 10954
rect 6389 10833 6401 10954
rect 6321 10831 6338 10833
rect 6246 10654 6263 10656
rect 6183 10534 6195 10654
rect 6251 10534 6263 10654
rect 6183 10532 6200 10534
rect 6016 10496 6062 10507
rect 6246 10532 6263 10534
rect 6200 10496 6246 10507
rect 5725 10458 5736 10461
rect 5790 10458 5801 10461
rect 5909 10458 5920 10461
rect 5974 10458 5985 10461
rect 6093 10458 6104 10461
rect 6158 10458 6169 10461
rect 5510 10413 5556 10424
rect 5723 10402 5735 10458
rect 5791 10402 5803 10458
rect 5723 10388 5803 10402
rect 5907 10402 5919 10458
rect 5975 10402 5987 10458
rect 5907 10388 5987 10402
rect 6091 10402 6103 10458
rect 6159 10402 6171 10458
rect 6384 10831 6401 10833
rect 6338 10413 6384 10424
rect 6091 10388 6171 10402
rect 5723 10308 5803 10310
rect 5335 10252 5735 10308
rect 5791 10252 5803 10308
rect 4237 10249 4317 10251
rect 5723 10250 5803 10252
rect 4421 10191 4501 10193
rect 3713 10135 4433 10191
rect 4489 10135 4501 10191
rect 4421 10133 4501 10135
rect 4750 10191 4830 10193
rect 5017 10192 5087 10203
rect 5907 10192 5987 10194
rect 5017 10191 5919 10192
rect 4750 10135 4762 10191
rect 4818 10135 5019 10191
rect 5075 10136 5919 10191
rect 5975 10136 5987 10192
rect 5075 10135 5335 10136
rect 4750 10133 4830 10135
rect 5017 10125 5087 10135
rect 5907 10134 5987 10136
rect 6236 10192 6316 10194
rect 6679 10192 6749 10202
rect 6236 10136 6248 10192
rect 6304 10136 6681 10192
rect 6737 10136 6749 10192
rect 6236 10134 6316 10136
rect 6679 10124 6749 10136
rect 7755 10191 7811 11438
rect 10711 11436 10791 11438
rect 11075 11494 11145 11506
rect 11797 11494 11853 12224
rect 12689 12222 12769 12224
rect 13419 12224 14187 12280
rect 14243 12224 14255 12280
rect 12321 12130 12401 12144
rect 12108 12108 12154 12119
rect 12321 12074 12333 12130
rect 12389 12074 12401 12130
rect 12505 12130 12585 12144
rect 12505 12074 12517 12130
rect 12573 12074 12585 12130
rect 12689 12130 12769 12144
rect 12689 12074 12701 12130
rect 12757 12074 12769 12130
rect 12936 12108 12982 12119
rect 12323 12071 12334 12074
rect 12388 12071 12399 12074
rect 12507 12071 12518 12074
rect 12572 12071 12583 12074
rect 12691 12071 12702 12074
rect 12756 12071 12767 12074
rect 12246 12025 12292 12036
rect 12154 11851 12246 12025
rect 12246 11840 12292 11851
rect 12430 12025 12476 12036
rect 12430 11840 12476 11851
rect 12614 12025 12660 12036
rect 12798 12025 12844 12036
rect 12781 11998 12798 12000
rect 12844 11998 12861 12000
rect 12781 11878 12793 11998
rect 12849 11878 12861 11998
rect 12781 11876 12798 11878
rect 12614 11840 12660 11851
rect 12844 11876 12861 11878
rect 12798 11840 12844 11851
rect 12108 11623 12154 11768
rect 12323 11759 12334 11805
rect 12388 11759 12399 11805
rect 12323 11726 12399 11759
rect 12507 11759 12518 11805
rect 12572 11759 12583 11805
rect 12507 11726 12583 11759
rect 12691 11759 12702 11805
rect 12756 11759 12767 11805
rect 12691 11726 12767 11759
rect 12936 11623 12982 11768
rect 12096 11611 12176 11623
rect 12096 11555 12108 11611
rect 12164 11555 12176 11611
rect 12096 11543 12176 11555
rect 12914 11611 12992 11623
rect 12914 11555 12926 11611
rect 12982 11555 12992 11611
rect 12914 11543 12992 11555
rect 11075 11438 11087 11494
rect 11143 11438 11853 11494
rect 13419 11494 13475 12224
rect 14175 12222 14255 12224
rect 13807 12130 13887 12144
rect 13594 12108 13640 12119
rect 13807 12074 13819 12130
rect 13875 12074 13887 12130
rect 13991 12130 14071 12144
rect 13991 12074 14003 12130
rect 14059 12074 14071 12130
rect 14175 12130 14255 12144
rect 14175 12074 14187 12130
rect 14243 12074 14255 12130
rect 14422 12108 14468 12119
rect 13809 12071 13820 12074
rect 13874 12071 13885 12074
rect 13993 12071 14004 12074
rect 14058 12071 14069 12074
rect 14177 12071 14188 12074
rect 14242 12071 14253 12074
rect 13732 12025 13778 12036
rect 13640 11851 13732 12025
rect 13732 11840 13778 11851
rect 13916 12025 13962 12036
rect 13916 11840 13962 11851
rect 14100 12025 14146 12036
rect 14284 12025 14330 12036
rect 14267 11998 14284 12000
rect 14330 11998 14347 12000
rect 14267 11878 14279 11998
rect 14335 11878 14347 11998
rect 14267 11876 14284 11878
rect 14100 11840 14146 11851
rect 14330 11876 14347 11878
rect 14284 11840 14330 11851
rect 13594 11623 13640 11768
rect 13809 11759 13820 11805
rect 13874 11759 13885 11805
rect 13809 11726 13885 11759
rect 13993 11759 14004 11805
rect 14058 11759 14069 11805
rect 13993 11726 14069 11759
rect 14177 11759 14188 11805
rect 14242 11759 14253 11805
rect 14177 11726 14253 11759
rect 14422 11623 14468 11768
rect 13582 11611 13662 11623
rect 13582 11555 13594 11611
rect 13650 11555 13662 11611
rect 13582 11543 13662 11555
rect 14400 11611 14478 11623
rect 14400 11555 14412 11611
rect 14468 11555 14478 11611
rect 14400 11543 14478 11555
rect 14753 11494 14833 11504
rect 13419 11438 14765 11494
rect 14821 11438 14833 11494
rect 11075 11426 11145 11438
rect 9235 11383 9305 11385
rect 10535 11384 10615 11386
rect 7891 11327 9237 11383
rect 9293 11327 9305 11383
rect 7891 10307 7947 11327
rect 9235 11315 9305 11327
rect 9377 11328 10547 11384
rect 10603 11328 10615 11384
rect 8555 11276 8641 11280
rect 8555 11220 8567 11276
rect 8623 11220 8641 11276
rect 8555 11208 8641 11220
rect 8066 11063 8112 11074
rect 8281 11072 8357 11105
rect 8281 11026 8292 11072
rect 8346 11026 8357 11072
rect 8465 11072 8541 11105
rect 8465 11026 8476 11072
rect 8530 11026 8541 11072
rect 8649 11072 8725 11105
rect 8649 11026 8660 11072
rect 8714 11026 8725 11072
rect 8894 11063 8940 11074
rect 8204 10980 8250 10991
rect 8187 10953 8204 10955
rect 8388 10980 8434 10991
rect 8250 10953 8267 10955
rect 8112 10833 8199 10953
rect 8255 10833 8267 10953
rect 8187 10831 8204 10833
rect 8112 10533 8204 10653
rect 8250 10831 8267 10833
rect 8371 10653 8388 10655
rect 8572 10980 8618 10991
rect 8555 10953 8572 10955
rect 8756 10980 8802 10991
rect 8618 10953 8635 10955
rect 8555 10833 8567 10953
rect 8623 10833 8635 10953
rect 8555 10831 8572 10833
rect 8434 10653 8451 10655
rect 8371 10533 8383 10653
rect 8439 10533 8451 10653
rect 8371 10531 8388 10533
rect 8204 10495 8250 10506
rect 8434 10531 8451 10533
rect 8388 10495 8434 10506
rect 8618 10831 8635 10833
rect 8739 10653 8756 10655
rect 8877 10953 8894 10955
rect 8940 10953 8957 10955
rect 8877 10832 8889 10953
rect 8945 10832 8957 10953
rect 8877 10830 8894 10832
rect 8802 10653 8819 10655
rect 8739 10533 8751 10653
rect 8807 10533 8819 10653
rect 8739 10531 8756 10533
rect 8572 10495 8618 10506
rect 8802 10531 8819 10533
rect 8756 10495 8802 10506
rect 8281 10457 8292 10460
rect 8346 10457 8357 10460
rect 8465 10457 8476 10460
rect 8530 10457 8541 10460
rect 8649 10457 8660 10460
rect 8714 10457 8725 10460
rect 8066 10412 8112 10423
rect 8279 10401 8291 10457
rect 8347 10401 8359 10457
rect 8279 10387 8359 10401
rect 8463 10401 8475 10457
rect 8531 10401 8543 10457
rect 8463 10387 8543 10401
rect 8647 10401 8659 10457
rect 8715 10401 8727 10457
rect 8940 10830 8957 10832
rect 8894 10412 8940 10423
rect 8647 10387 8727 10401
rect 8279 10307 8359 10309
rect 7891 10251 8291 10307
rect 8347 10251 8359 10307
rect 9377 10308 9433 11328
rect 10535 11316 10615 11328
rect 10041 11277 10127 11281
rect 10041 11221 10053 11277
rect 10109 11221 10127 11277
rect 10041 11209 10127 11221
rect 9552 11064 9598 11075
rect 9767 11073 9843 11106
rect 9767 11027 9778 11073
rect 9832 11027 9843 11073
rect 9951 11073 10027 11106
rect 9951 11027 9962 11073
rect 10016 11027 10027 11073
rect 10135 11073 10211 11106
rect 10135 11027 10146 11073
rect 10200 11027 10211 11073
rect 10380 11064 10426 11075
rect 9690 10981 9736 10992
rect 9673 10954 9690 10956
rect 9874 10981 9920 10992
rect 9736 10954 9753 10956
rect 9598 10834 9685 10954
rect 9741 10834 9753 10954
rect 9673 10832 9690 10834
rect 9598 10534 9690 10654
rect 9736 10832 9753 10834
rect 9857 10654 9874 10656
rect 10058 10981 10104 10992
rect 10041 10954 10058 10956
rect 10242 10981 10288 10992
rect 10104 10954 10121 10956
rect 10041 10834 10053 10954
rect 10109 10834 10121 10954
rect 10041 10832 10058 10834
rect 9920 10654 9937 10656
rect 9857 10534 9869 10654
rect 9925 10534 9937 10654
rect 9857 10532 9874 10534
rect 9690 10496 9736 10507
rect 9920 10532 9937 10534
rect 9874 10496 9920 10507
rect 10104 10832 10121 10834
rect 10225 10654 10242 10656
rect 10363 10954 10380 10956
rect 10426 10954 10443 10956
rect 10363 10833 10375 10954
rect 10431 10833 10443 10954
rect 10363 10831 10380 10833
rect 10288 10654 10305 10656
rect 10225 10534 10237 10654
rect 10293 10534 10305 10654
rect 10225 10532 10242 10534
rect 10058 10496 10104 10507
rect 10288 10532 10305 10534
rect 10242 10496 10288 10507
rect 9767 10458 9778 10461
rect 9832 10458 9843 10461
rect 9951 10458 9962 10461
rect 10016 10458 10027 10461
rect 10135 10458 10146 10461
rect 10200 10458 10211 10461
rect 9552 10413 9598 10424
rect 9765 10402 9777 10458
rect 9833 10402 9845 10458
rect 9765 10388 9845 10402
rect 9949 10402 9961 10458
rect 10017 10402 10029 10458
rect 9949 10388 10029 10402
rect 10133 10402 10145 10458
rect 10201 10402 10213 10458
rect 10426 10831 10443 10833
rect 10380 10413 10426 10424
rect 10133 10388 10213 10402
rect 9765 10308 9845 10310
rect 9377 10252 9777 10308
rect 9833 10252 9845 10308
rect 8279 10249 8359 10251
rect 9765 10250 9845 10252
rect 8463 10191 8543 10193
rect 7755 10135 8475 10191
rect 8531 10135 8543 10191
rect 8463 10133 8543 10135
rect 8792 10191 8872 10193
rect 9059 10192 9129 10203
rect 9949 10192 10029 10194
rect 9059 10191 9961 10192
rect 8792 10135 8804 10191
rect 8860 10135 9061 10191
rect 9117 10136 9961 10191
rect 10017 10136 10029 10192
rect 9117 10135 9377 10136
rect 8792 10133 8872 10135
rect 9059 10125 9129 10135
rect 9949 10134 10029 10136
rect 10278 10192 10358 10194
rect 10721 10192 10791 10202
rect 10278 10136 10290 10192
rect 10346 10136 10723 10192
rect 10779 10136 10791 10192
rect 10278 10134 10358 10136
rect 10721 10124 10791 10136
rect 11797 10191 11853 11438
rect 14753 11436 14833 11438
rect 13277 11383 13347 11385
rect 14577 11384 14657 11386
rect 11933 11327 13279 11383
rect 13335 11327 13347 11383
rect 11933 10307 11989 11327
rect 13277 11315 13347 11327
rect 13419 11328 14589 11384
rect 14645 11328 14657 11384
rect 12597 11276 12683 11280
rect 12597 11220 12609 11276
rect 12665 11220 12683 11276
rect 12597 11208 12683 11220
rect 12108 11063 12154 11074
rect 12323 11072 12399 11105
rect 12323 11026 12334 11072
rect 12388 11026 12399 11072
rect 12507 11072 12583 11105
rect 12507 11026 12518 11072
rect 12572 11026 12583 11072
rect 12691 11072 12767 11105
rect 12691 11026 12702 11072
rect 12756 11026 12767 11072
rect 12936 11063 12982 11074
rect 12246 10980 12292 10991
rect 12229 10953 12246 10955
rect 12430 10980 12476 10991
rect 12292 10953 12309 10955
rect 12154 10833 12241 10953
rect 12297 10833 12309 10953
rect 12229 10831 12246 10833
rect 12154 10533 12246 10653
rect 12292 10831 12309 10833
rect 12413 10653 12430 10655
rect 12614 10980 12660 10991
rect 12597 10953 12614 10955
rect 12798 10980 12844 10991
rect 12660 10953 12677 10955
rect 12597 10833 12609 10953
rect 12665 10833 12677 10953
rect 12597 10831 12614 10833
rect 12476 10653 12493 10655
rect 12413 10533 12425 10653
rect 12481 10533 12493 10653
rect 12413 10531 12430 10533
rect 12246 10495 12292 10506
rect 12476 10531 12493 10533
rect 12430 10495 12476 10506
rect 12660 10831 12677 10833
rect 12781 10653 12798 10655
rect 12919 10953 12936 10955
rect 12982 10953 12999 10955
rect 12919 10832 12931 10953
rect 12987 10832 12999 10953
rect 12919 10830 12936 10832
rect 12844 10653 12861 10655
rect 12781 10533 12793 10653
rect 12849 10533 12861 10653
rect 12781 10531 12798 10533
rect 12614 10495 12660 10506
rect 12844 10531 12861 10533
rect 12798 10495 12844 10506
rect 12323 10457 12334 10460
rect 12388 10457 12399 10460
rect 12507 10457 12518 10460
rect 12572 10457 12583 10460
rect 12691 10457 12702 10460
rect 12756 10457 12767 10460
rect 12108 10412 12154 10423
rect 12321 10401 12333 10457
rect 12389 10401 12401 10457
rect 12321 10387 12401 10401
rect 12505 10401 12517 10457
rect 12573 10401 12585 10457
rect 12505 10387 12585 10401
rect 12689 10401 12701 10457
rect 12757 10401 12769 10457
rect 12982 10830 12999 10832
rect 12936 10412 12982 10423
rect 12689 10387 12769 10401
rect 12321 10307 12401 10309
rect 11933 10251 12333 10307
rect 12389 10251 12401 10307
rect 13419 10308 13475 11328
rect 14577 11316 14657 11328
rect 14083 11277 14169 11281
rect 14083 11221 14095 11277
rect 14151 11221 14169 11277
rect 14083 11209 14169 11221
rect 13594 11064 13640 11075
rect 13809 11073 13885 11106
rect 13809 11027 13820 11073
rect 13874 11027 13885 11073
rect 13993 11073 14069 11106
rect 13993 11027 14004 11073
rect 14058 11027 14069 11073
rect 14177 11073 14253 11106
rect 14177 11027 14188 11073
rect 14242 11027 14253 11073
rect 14422 11064 14468 11075
rect 13732 10981 13778 10992
rect 13715 10954 13732 10956
rect 13916 10981 13962 10992
rect 13778 10954 13795 10956
rect 13640 10834 13727 10954
rect 13783 10834 13795 10954
rect 13715 10832 13732 10834
rect 13640 10534 13732 10654
rect 13778 10832 13795 10834
rect 13899 10654 13916 10656
rect 14100 10981 14146 10992
rect 14083 10954 14100 10956
rect 14284 10981 14330 10992
rect 14146 10954 14163 10956
rect 14083 10834 14095 10954
rect 14151 10834 14163 10954
rect 14083 10832 14100 10834
rect 13962 10654 13979 10656
rect 13899 10534 13911 10654
rect 13967 10534 13979 10654
rect 13899 10532 13916 10534
rect 13732 10496 13778 10507
rect 13962 10532 13979 10534
rect 13916 10496 13962 10507
rect 14146 10832 14163 10834
rect 14267 10654 14284 10656
rect 14405 10954 14422 10956
rect 14468 10954 14485 10956
rect 14405 10833 14417 10954
rect 14473 10833 14485 10954
rect 14405 10831 14422 10833
rect 14330 10654 14347 10656
rect 14267 10534 14279 10654
rect 14335 10534 14347 10654
rect 14267 10532 14284 10534
rect 14100 10496 14146 10507
rect 14330 10532 14347 10534
rect 14284 10496 14330 10507
rect 13809 10458 13820 10461
rect 13874 10458 13885 10461
rect 13993 10458 14004 10461
rect 14058 10458 14069 10461
rect 14177 10458 14188 10461
rect 14242 10458 14253 10461
rect 13594 10413 13640 10424
rect 13807 10402 13819 10458
rect 13875 10402 13887 10458
rect 13807 10388 13887 10402
rect 13991 10402 14003 10458
rect 14059 10402 14071 10458
rect 13991 10388 14071 10402
rect 14175 10402 14187 10458
rect 14243 10402 14255 10458
rect 14468 10831 14485 10833
rect 14422 10413 14468 10424
rect 14175 10388 14255 10402
rect 13807 10308 13887 10310
rect 13419 10252 13819 10308
rect 13875 10252 13887 10308
rect 12321 10249 12401 10251
rect 13807 10250 13887 10252
rect 12505 10191 12585 10193
rect 11797 10135 12517 10191
rect 12573 10135 12585 10191
rect 12505 10133 12585 10135
rect 12834 10191 12914 10193
rect 13101 10192 13171 10203
rect 13991 10192 14071 10194
rect 13101 10191 14003 10192
rect 12834 10135 12846 10191
rect 12902 10135 13103 10191
rect 13159 10136 14003 10191
rect 14059 10136 14071 10192
rect 13159 10135 13419 10136
rect 12834 10133 12914 10135
rect 13101 10125 13171 10135
rect 13991 10134 14071 10136
rect 14320 10192 14400 10194
rect 14763 10192 14833 10202
rect 14320 10136 14332 10192
rect 14388 10136 14765 10192
rect 14821 10136 14833 10192
rect 14320 10134 14400 10136
rect 14763 10124 14833 10136
rect -12573 10075 -12503 10087
rect -11533 10075 -11453 10077
rect -10047 10076 -9967 10078
rect -12573 10019 -12561 10075
rect -12505 10019 -11521 10075
rect -11465 10019 -11453 10075
rect -12573 10007 -12503 10019
rect -12289 9288 -12233 10019
rect -11533 10017 -11453 10019
rect -10803 10020 -10035 10076
rect -9979 10020 -9967 10076
rect -11901 9925 -11821 9939
rect -12114 9903 -12068 9914
rect -11901 9869 -11889 9925
rect -11833 9869 -11821 9925
rect -11717 9925 -11637 9939
rect -11717 9869 -11705 9925
rect -11649 9869 -11637 9925
rect -11533 9925 -11453 9939
rect -11533 9869 -11521 9925
rect -11465 9869 -11453 9925
rect -11286 9903 -11240 9914
rect -11899 9866 -11888 9869
rect -11834 9866 -11823 9869
rect -11715 9866 -11704 9869
rect -11650 9866 -11639 9869
rect -11531 9866 -11520 9869
rect -11466 9866 -11455 9869
rect -11976 9820 -11930 9831
rect -12068 9646 -11976 9820
rect -11976 9635 -11930 9646
rect -11792 9820 -11746 9831
rect -11792 9635 -11746 9646
rect -11608 9820 -11562 9831
rect -11424 9820 -11378 9831
rect -11441 9793 -11424 9795
rect -11378 9793 -11361 9795
rect -11441 9673 -11429 9793
rect -11373 9673 -11361 9793
rect -11441 9671 -11424 9673
rect -11608 9635 -11562 9646
rect -11378 9671 -11361 9673
rect -11424 9635 -11378 9646
rect -12114 9418 -12068 9563
rect -11899 9554 -11888 9600
rect -11834 9554 -11823 9600
rect -11899 9521 -11823 9554
rect -11715 9554 -11704 9600
rect -11650 9554 -11639 9600
rect -11715 9521 -11639 9554
rect -11531 9554 -11520 9600
rect -11466 9554 -11455 9600
rect -11531 9521 -11455 9554
rect -11286 9418 -11240 9563
rect -12126 9406 -12046 9418
rect -12126 9350 -12114 9406
rect -12058 9350 -12046 9406
rect -12126 9338 -12046 9350
rect -11308 9406 -11230 9418
rect -11308 9350 -11296 9406
rect -11240 9350 -11230 9406
rect -11308 9338 -11230 9350
rect -10955 9288 -10875 9298
rect -12289 9232 -10943 9288
rect -10887 9232 -10875 9288
rect -10955 9230 -10875 9232
rect -11121 9179 -11051 9181
rect -12289 9178 -11051 9179
rect -12289 9124 -11119 9178
rect -11063 9124 -11051 9178
rect -12289 9123 -11051 9124
rect -12289 8102 -12233 9123
rect -11121 9115 -11051 9123
rect -11625 9071 -11539 9075
rect -11625 9015 -11613 9071
rect -11557 9015 -11539 9071
rect -11625 9003 -11539 9015
rect -12114 8858 -12068 8869
rect -11899 8867 -11823 8900
rect -11899 8821 -11888 8867
rect -11834 8821 -11823 8867
rect -11715 8867 -11639 8900
rect -11715 8821 -11704 8867
rect -11650 8821 -11639 8867
rect -11531 8867 -11455 8900
rect -11531 8821 -11520 8867
rect -11466 8821 -11455 8867
rect -11286 8858 -11240 8869
rect -11976 8775 -11930 8786
rect -11993 8748 -11976 8750
rect -11792 8775 -11746 8786
rect -11930 8748 -11913 8750
rect -12068 8628 -11981 8748
rect -11925 8628 -11913 8748
rect -11993 8626 -11976 8628
rect -12068 8328 -11976 8448
rect -11930 8626 -11913 8628
rect -11809 8448 -11792 8450
rect -11608 8775 -11562 8786
rect -11625 8748 -11608 8750
rect -11424 8775 -11378 8786
rect -11562 8748 -11545 8750
rect -11625 8628 -11613 8748
rect -11557 8628 -11545 8748
rect -11625 8626 -11608 8628
rect -11746 8448 -11729 8450
rect -11809 8328 -11797 8448
rect -11741 8328 -11729 8448
rect -11809 8326 -11792 8328
rect -11976 8290 -11930 8301
rect -11746 8326 -11729 8328
rect -11792 8290 -11746 8301
rect -11562 8626 -11545 8628
rect -11441 8448 -11424 8450
rect -11303 8748 -11286 8750
rect -11240 8748 -11223 8750
rect -11303 8627 -11291 8748
rect -11235 8627 -11223 8748
rect -11303 8625 -11286 8627
rect -11378 8448 -11361 8450
rect -11441 8328 -11429 8448
rect -11373 8328 -11361 8448
rect -11441 8326 -11424 8328
rect -11608 8290 -11562 8301
rect -11378 8326 -11361 8328
rect -11424 8290 -11378 8301
rect -11899 8252 -11888 8255
rect -11834 8252 -11823 8255
rect -11715 8252 -11704 8255
rect -11650 8252 -11639 8255
rect -11531 8252 -11520 8255
rect -11466 8252 -11455 8255
rect -12114 8207 -12068 8218
rect -11901 8196 -11889 8252
rect -11833 8196 -11821 8252
rect -11901 8182 -11821 8196
rect -11717 8196 -11705 8252
rect -11649 8196 -11637 8252
rect -11717 8182 -11637 8196
rect -11533 8196 -11521 8252
rect -11465 8196 -11453 8252
rect -11240 8625 -11223 8627
rect -11286 8207 -11240 8218
rect -11533 8182 -11453 8196
rect -11901 8102 -11821 8104
rect -12289 8046 -11889 8102
rect -11833 8046 -11821 8102
rect -11901 8044 -11821 8046
rect -12709 7986 -12639 8000
rect -11717 7986 -11637 7988
rect -12709 7930 -12697 7986
rect -12641 7930 -11705 7986
rect -11649 7930 -11637 7986
rect -12709 7918 -12639 7930
rect -11717 7928 -11637 7930
rect -11388 7986 -11308 7988
rect -10945 7986 -10885 7998
rect -11388 7930 -11376 7986
rect -11320 7930 -10943 7986
rect -10887 7930 -10885 7986
rect -11388 7928 -11308 7930
rect -10945 7918 -10885 7930
rect -12908 7870 -12828 7882
rect -11533 7870 -11453 7872
rect -12908 7814 -12896 7870
rect -12840 7814 -11521 7870
rect -11465 7814 -11453 7870
rect -12908 7802 -12828 7814
rect -11533 7812 -11453 7814
rect -11901 7720 -11821 7734
rect -12114 7698 -12068 7709
rect -11901 7664 -11889 7720
rect -11833 7664 -11821 7720
rect -11717 7720 -11637 7734
rect -11717 7664 -11705 7720
rect -11649 7664 -11637 7720
rect -11533 7720 -11453 7734
rect -11533 7664 -11521 7720
rect -11465 7664 -11453 7720
rect -11286 7698 -11240 7709
rect -11899 7661 -11888 7664
rect -11834 7661 -11823 7664
rect -11715 7661 -11704 7664
rect -11650 7661 -11639 7664
rect -11531 7661 -11520 7664
rect -11466 7661 -11455 7664
rect -11976 7615 -11930 7626
rect -12068 7441 -11976 7615
rect -11976 7430 -11930 7441
rect -11792 7615 -11746 7626
rect -11792 7430 -11746 7441
rect -11608 7615 -11562 7626
rect -11424 7615 -11378 7626
rect -11441 7588 -11424 7590
rect -11378 7588 -11361 7590
rect -11441 7468 -11429 7588
rect -11373 7468 -11361 7588
rect -11441 7466 -11424 7468
rect -11608 7430 -11562 7441
rect -11378 7466 -11361 7468
rect -11424 7430 -11378 7441
rect -12114 7213 -12068 7358
rect -11899 7349 -11888 7395
rect -11834 7349 -11823 7395
rect -11899 7316 -11823 7349
rect -11715 7349 -11704 7395
rect -11650 7349 -11639 7395
rect -11715 7316 -11639 7349
rect -11531 7349 -11520 7395
rect -11466 7349 -11455 7395
rect -11531 7316 -11455 7349
rect -11286 7213 -11240 7358
rect -12126 7201 -12046 7213
rect -12126 7145 -12114 7201
rect -12058 7145 -12046 7201
rect -12126 7133 -12046 7145
rect -11308 7201 -11228 7213
rect -11308 7145 -11296 7201
rect -11240 7145 -11228 7201
rect -11308 7133 -11228 7145
rect -12908 7083 -12822 7095
rect -12699 7083 -12639 7087
rect -10803 7083 -10747 10020
rect -10047 10018 -9967 10020
rect -8561 10075 -8491 10087
rect -7521 10075 -7441 10077
rect -6035 10076 -5955 10078
rect -8561 10019 -8549 10075
rect -8493 10019 -7509 10075
rect -7453 10019 -7441 10075
rect -8561 10007 -8491 10019
rect -10415 9926 -10335 9940
rect -10628 9904 -10582 9915
rect -10415 9870 -10403 9926
rect -10347 9870 -10335 9926
rect -10231 9926 -10151 9940
rect -10231 9870 -10219 9926
rect -10163 9870 -10151 9926
rect -10047 9926 -9967 9940
rect -10047 9870 -10035 9926
rect -9979 9870 -9967 9926
rect -9800 9904 -9754 9915
rect -10413 9867 -10402 9870
rect -10348 9867 -10337 9870
rect -10229 9867 -10218 9870
rect -10164 9867 -10153 9870
rect -10045 9867 -10034 9870
rect -9980 9867 -9969 9870
rect -10490 9821 -10444 9832
rect -10582 9647 -10490 9821
rect -10490 9636 -10444 9647
rect -10306 9821 -10260 9832
rect -10306 9636 -10260 9647
rect -10122 9821 -10076 9832
rect -9938 9821 -9892 9832
rect -9955 9794 -9938 9796
rect -9892 9794 -9875 9796
rect -9955 9674 -9943 9794
rect -9887 9674 -9875 9794
rect -9955 9672 -9938 9674
rect -10122 9636 -10076 9647
rect -9892 9672 -9875 9674
rect -9938 9636 -9892 9647
rect -10628 9419 -10582 9564
rect -10413 9555 -10402 9601
rect -10348 9555 -10337 9601
rect -10413 9522 -10337 9555
rect -10229 9555 -10218 9601
rect -10164 9555 -10153 9601
rect -10229 9522 -10153 9555
rect -10045 9555 -10034 9601
rect -9980 9555 -9969 9601
rect -10045 9522 -9969 9555
rect -9800 9419 -9754 9564
rect -10640 9407 -10560 9419
rect -10640 9351 -10628 9407
rect -10572 9351 -10560 9407
rect -10640 9339 -10560 9351
rect -9822 9407 -9744 9419
rect -9822 9351 -9810 9407
rect -9754 9351 -9744 9407
rect -9822 9339 -9744 9351
rect -8277 9288 -8221 10019
rect -7521 10017 -7441 10019
rect -6791 10020 -6023 10076
rect -5967 10020 -5955 10076
rect -7889 9925 -7809 9939
rect -8102 9903 -8056 9914
rect -7889 9869 -7877 9925
rect -7821 9869 -7809 9925
rect -7705 9925 -7625 9939
rect -7705 9869 -7693 9925
rect -7637 9869 -7625 9925
rect -7521 9925 -7441 9939
rect -7521 9869 -7509 9925
rect -7453 9869 -7441 9925
rect -7274 9903 -7228 9914
rect -7887 9866 -7876 9869
rect -7822 9866 -7811 9869
rect -7703 9866 -7692 9869
rect -7638 9866 -7627 9869
rect -7519 9866 -7508 9869
rect -7454 9866 -7443 9869
rect -7964 9820 -7918 9831
rect -8056 9646 -7964 9820
rect -7964 9635 -7918 9646
rect -7780 9820 -7734 9831
rect -7780 9635 -7734 9646
rect -7596 9820 -7550 9831
rect -7412 9820 -7366 9831
rect -7429 9793 -7412 9795
rect -7366 9793 -7349 9795
rect -7429 9673 -7417 9793
rect -7361 9673 -7349 9793
rect -7429 9671 -7412 9673
rect -7596 9635 -7550 9646
rect -7366 9671 -7349 9673
rect -7412 9635 -7366 9646
rect -8102 9418 -8056 9563
rect -7887 9554 -7876 9600
rect -7822 9554 -7811 9600
rect -7887 9521 -7811 9554
rect -7703 9554 -7692 9600
rect -7638 9554 -7627 9600
rect -7703 9521 -7627 9554
rect -7519 9554 -7508 9600
rect -7454 9554 -7443 9600
rect -7519 9521 -7443 9554
rect -7274 9418 -7228 9563
rect -8114 9406 -8034 9418
rect -8114 9350 -8102 9406
rect -8046 9350 -8034 9406
rect -8114 9338 -8034 9350
rect -7296 9406 -7218 9418
rect -7296 9350 -7284 9406
rect -7228 9350 -7218 9406
rect -7296 9338 -7218 9350
rect -6943 9288 -6863 9298
rect -8277 9232 -6931 9288
rect -6875 9232 -6863 9288
rect -6943 9230 -6863 9232
rect -7109 9179 -7039 9181
rect -8277 9178 -7039 9179
rect -8277 9124 -7107 9178
rect -7051 9124 -7039 9178
rect -8277 9123 -7039 9124
rect -8277 8102 -8221 9123
rect -7109 9115 -7039 9123
rect -7613 9071 -7527 9075
rect -7613 9015 -7601 9071
rect -7545 9015 -7527 9071
rect -7613 9003 -7527 9015
rect -8102 8858 -8056 8869
rect -7887 8867 -7811 8900
rect -7887 8821 -7876 8867
rect -7822 8821 -7811 8867
rect -7703 8867 -7627 8900
rect -7703 8821 -7692 8867
rect -7638 8821 -7627 8867
rect -7519 8867 -7443 8900
rect -7519 8821 -7508 8867
rect -7454 8821 -7443 8867
rect -7274 8858 -7228 8869
rect -7964 8775 -7918 8786
rect -7981 8748 -7964 8750
rect -7780 8775 -7734 8786
rect -7918 8748 -7901 8750
rect -8056 8628 -7969 8748
rect -7913 8628 -7901 8748
rect -7981 8626 -7964 8628
rect -8056 8328 -7964 8448
rect -7918 8626 -7901 8628
rect -7797 8448 -7780 8450
rect -7596 8775 -7550 8786
rect -7613 8748 -7596 8750
rect -7412 8775 -7366 8786
rect -7550 8748 -7533 8750
rect -7613 8628 -7601 8748
rect -7545 8628 -7533 8748
rect -7613 8626 -7596 8628
rect -7734 8448 -7717 8450
rect -7797 8328 -7785 8448
rect -7729 8328 -7717 8448
rect -7797 8326 -7780 8328
rect -7964 8290 -7918 8301
rect -7734 8326 -7717 8328
rect -7780 8290 -7734 8301
rect -7550 8626 -7533 8628
rect -7429 8448 -7412 8450
rect -7291 8748 -7274 8750
rect -7228 8748 -7211 8750
rect -7291 8627 -7279 8748
rect -7223 8627 -7211 8748
rect -7291 8625 -7274 8627
rect -7366 8448 -7349 8450
rect -7429 8328 -7417 8448
rect -7361 8328 -7349 8448
rect -7429 8326 -7412 8328
rect -7596 8290 -7550 8301
rect -7366 8326 -7349 8328
rect -7412 8290 -7366 8301
rect -7887 8252 -7876 8255
rect -7822 8252 -7811 8255
rect -7703 8252 -7692 8255
rect -7638 8252 -7627 8255
rect -7519 8252 -7508 8255
rect -7454 8252 -7443 8255
rect -8102 8207 -8056 8218
rect -7889 8196 -7877 8252
rect -7821 8196 -7809 8252
rect -7889 8182 -7809 8196
rect -7705 8196 -7693 8252
rect -7637 8196 -7625 8252
rect -7705 8182 -7625 8196
rect -7521 8196 -7509 8252
rect -7453 8196 -7441 8252
rect -7228 8625 -7211 8627
rect -7274 8207 -7228 8218
rect -7521 8182 -7441 8196
rect -7889 8102 -7809 8104
rect -8277 8046 -7877 8102
rect -7821 8046 -7809 8102
rect -7889 8044 -7809 8046
rect -8697 7986 -8627 8000
rect -7705 7986 -7625 7988
rect -8697 7930 -8685 7986
rect -8629 7930 -7693 7986
rect -7637 7930 -7625 7986
rect -8697 7918 -8627 7930
rect -7705 7928 -7625 7930
rect -7376 7986 -7296 7988
rect -6933 7986 -6873 7998
rect -7376 7930 -7364 7986
rect -7308 7930 -6931 7986
rect -6875 7930 -6873 7986
rect -7376 7928 -7296 7930
rect -6933 7918 -6873 7930
rect -8833 7870 -8763 7882
rect -7521 7870 -7441 7872
rect -8833 7814 -8821 7870
rect -8765 7814 -7509 7870
rect -7453 7814 -7441 7870
rect -8833 7802 -8763 7814
rect -7521 7812 -7441 7814
rect -7889 7720 -7809 7734
rect -8102 7698 -8056 7709
rect -7889 7664 -7877 7720
rect -7821 7664 -7809 7720
rect -7705 7720 -7625 7734
rect -7705 7664 -7693 7720
rect -7637 7664 -7625 7720
rect -7521 7720 -7441 7734
rect -7521 7664 -7509 7720
rect -7453 7664 -7441 7720
rect -7274 7698 -7228 7709
rect -7887 7661 -7876 7664
rect -7822 7661 -7811 7664
rect -7703 7661 -7692 7664
rect -7638 7661 -7627 7664
rect -7519 7661 -7508 7664
rect -7454 7661 -7443 7664
rect -7964 7615 -7918 7626
rect -8056 7441 -7964 7615
rect -7964 7430 -7918 7441
rect -7780 7615 -7734 7626
rect -7780 7430 -7734 7441
rect -7596 7615 -7550 7626
rect -7412 7615 -7366 7626
rect -7429 7588 -7412 7590
rect -7366 7588 -7349 7590
rect -7429 7468 -7417 7588
rect -7361 7468 -7349 7588
rect -7429 7466 -7412 7468
rect -7596 7430 -7550 7441
rect -7366 7466 -7349 7468
rect -7412 7430 -7366 7441
rect -8102 7213 -8056 7358
rect -7887 7349 -7876 7395
rect -7822 7349 -7811 7395
rect -7887 7316 -7811 7349
rect -7703 7349 -7692 7395
rect -7638 7349 -7627 7395
rect -7703 7316 -7627 7349
rect -7519 7349 -7508 7395
rect -7454 7349 -7443 7395
rect -7519 7316 -7443 7349
rect -7274 7213 -7228 7358
rect -8114 7201 -8034 7213
rect -8114 7145 -8102 7201
rect -8046 7145 -8034 7201
rect -8114 7133 -8034 7145
rect -7296 7201 -7216 7213
rect -7296 7145 -7284 7201
rect -7228 7145 -7216 7201
rect -7296 7133 -7216 7145
rect -12908 7027 -12896 7083
rect -12840 7027 -12697 7083
rect -12641 7027 -10747 7083
rect -8969 7083 -8899 7095
rect -8687 7083 -8627 7087
rect -6791 7083 -6735 10020
rect -6035 10018 -5955 10020
rect -4519 10075 -4449 10087
rect -3479 10075 -3399 10077
rect -1993 10076 -1913 10078
rect -4519 10019 -4507 10075
rect -4451 10019 -3467 10075
rect -3411 10019 -3399 10075
rect -4519 10007 -4449 10019
rect -6403 9926 -6323 9940
rect -6616 9904 -6570 9915
rect -6403 9870 -6391 9926
rect -6335 9870 -6323 9926
rect -6219 9926 -6139 9940
rect -6219 9870 -6207 9926
rect -6151 9870 -6139 9926
rect -6035 9926 -5955 9940
rect -6035 9870 -6023 9926
rect -5967 9870 -5955 9926
rect -5788 9904 -5742 9915
rect -6401 9867 -6390 9870
rect -6336 9867 -6325 9870
rect -6217 9867 -6206 9870
rect -6152 9867 -6141 9870
rect -6033 9867 -6022 9870
rect -5968 9867 -5957 9870
rect -6478 9821 -6432 9832
rect -6570 9647 -6478 9821
rect -6478 9636 -6432 9647
rect -6294 9821 -6248 9832
rect -6294 9636 -6248 9647
rect -6110 9821 -6064 9832
rect -5926 9821 -5880 9832
rect -5943 9794 -5926 9796
rect -5880 9794 -5863 9796
rect -5943 9674 -5931 9794
rect -5875 9674 -5863 9794
rect -5943 9672 -5926 9674
rect -6110 9636 -6064 9647
rect -5880 9672 -5863 9674
rect -5926 9636 -5880 9647
rect -6616 9419 -6570 9564
rect -6401 9555 -6390 9601
rect -6336 9555 -6325 9601
rect -6401 9522 -6325 9555
rect -6217 9555 -6206 9601
rect -6152 9555 -6141 9601
rect -6217 9522 -6141 9555
rect -6033 9555 -6022 9601
rect -5968 9555 -5957 9601
rect -6033 9522 -5957 9555
rect -5788 9419 -5742 9564
rect -6628 9407 -6548 9419
rect -6628 9351 -6616 9407
rect -6560 9351 -6548 9407
rect -6628 9339 -6548 9351
rect -5810 9407 -5732 9419
rect -5810 9351 -5798 9407
rect -5742 9351 -5732 9407
rect -5810 9339 -5732 9351
rect -4235 9288 -4179 10019
rect -3479 10017 -3399 10019
rect -2749 10020 -1981 10076
rect -1925 10020 -1913 10076
rect -3847 9925 -3767 9939
rect -4060 9903 -4014 9914
rect -3847 9869 -3835 9925
rect -3779 9869 -3767 9925
rect -3663 9925 -3583 9939
rect -3663 9869 -3651 9925
rect -3595 9869 -3583 9925
rect -3479 9925 -3399 9939
rect -3479 9869 -3467 9925
rect -3411 9869 -3399 9925
rect -3232 9903 -3186 9914
rect -3845 9866 -3834 9869
rect -3780 9866 -3769 9869
rect -3661 9866 -3650 9869
rect -3596 9866 -3585 9869
rect -3477 9866 -3466 9869
rect -3412 9866 -3401 9869
rect -3922 9820 -3876 9831
rect -4014 9646 -3922 9820
rect -3922 9635 -3876 9646
rect -3738 9820 -3692 9831
rect -3738 9635 -3692 9646
rect -3554 9820 -3508 9831
rect -3370 9820 -3324 9831
rect -3387 9793 -3370 9795
rect -3324 9793 -3307 9795
rect -3387 9673 -3375 9793
rect -3319 9673 -3307 9793
rect -3387 9671 -3370 9673
rect -3554 9635 -3508 9646
rect -3324 9671 -3307 9673
rect -3370 9635 -3324 9646
rect -4060 9418 -4014 9563
rect -3845 9554 -3834 9600
rect -3780 9554 -3769 9600
rect -3845 9521 -3769 9554
rect -3661 9554 -3650 9600
rect -3596 9554 -3585 9600
rect -3661 9521 -3585 9554
rect -3477 9554 -3466 9600
rect -3412 9554 -3401 9600
rect -3477 9521 -3401 9554
rect -3232 9418 -3186 9563
rect -4072 9406 -3992 9418
rect -4072 9350 -4060 9406
rect -4004 9350 -3992 9406
rect -4072 9338 -3992 9350
rect -3254 9406 -3176 9418
rect -3254 9350 -3242 9406
rect -3186 9350 -3176 9406
rect -3254 9338 -3176 9350
rect -2901 9288 -2821 9298
rect -4235 9232 -2889 9288
rect -2833 9232 -2821 9288
rect -2901 9230 -2821 9232
rect -3067 9179 -2997 9181
rect -4235 9178 -2997 9179
rect -4235 9124 -3065 9178
rect -3009 9124 -2997 9178
rect -4235 9123 -2997 9124
rect -4235 8102 -4179 9123
rect -3067 9115 -2997 9123
rect -3571 9071 -3485 9075
rect -3571 9015 -3559 9071
rect -3503 9015 -3485 9071
rect -3571 9003 -3485 9015
rect -4060 8858 -4014 8869
rect -3845 8867 -3769 8900
rect -3845 8821 -3834 8867
rect -3780 8821 -3769 8867
rect -3661 8867 -3585 8900
rect -3661 8821 -3650 8867
rect -3596 8821 -3585 8867
rect -3477 8867 -3401 8900
rect -3477 8821 -3466 8867
rect -3412 8821 -3401 8867
rect -3232 8858 -3186 8869
rect -3922 8775 -3876 8786
rect -3939 8748 -3922 8750
rect -3738 8775 -3692 8786
rect -3876 8748 -3859 8750
rect -4014 8628 -3927 8748
rect -3871 8628 -3859 8748
rect -3939 8626 -3922 8628
rect -4014 8328 -3922 8448
rect -3876 8626 -3859 8628
rect -3755 8448 -3738 8450
rect -3554 8775 -3508 8786
rect -3571 8748 -3554 8750
rect -3370 8775 -3324 8786
rect -3508 8748 -3491 8750
rect -3571 8628 -3559 8748
rect -3503 8628 -3491 8748
rect -3571 8626 -3554 8628
rect -3692 8448 -3675 8450
rect -3755 8328 -3743 8448
rect -3687 8328 -3675 8448
rect -3755 8326 -3738 8328
rect -3922 8290 -3876 8301
rect -3692 8326 -3675 8328
rect -3738 8290 -3692 8301
rect -3508 8626 -3491 8628
rect -3387 8448 -3370 8450
rect -3249 8748 -3232 8750
rect -3186 8748 -3169 8750
rect -3249 8627 -3237 8748
rect -3181 8627 -3169 8748
rect -3249 8625 -3232 8627
rect -3324 8448 -3307 8450
rect -3387 8328 -3375 8448
rect -3319 8328 -3307 8448
rect -3387 8326 -3370 8328
rect -3554 8290 -3508 8301
rect -3324 8326 -3307 8328
rect -3370 8290 -3324 8301
rect -3845 8252 -3834 8255
rect -3780 8252 -3769 8255
rect -3661 8252 -3650 8255
rect -3596 8252 -3585 8255
rect -3477 8252 -3466 8255
rect -3412 8252 -3401 8255
rect -4060 8207 -4014 8218
rect -3847 8196 -3835 8252
rect -3779 8196 -3767 8252
rect -3847 8182 -3767 8196
rect -3663 8196 -3651 8252
rect -3595 8196 -3583 8252
rect -3663 8182 -3583 8196
rect -3479 8196 -3467 8252
rect -3411 8196 -3399 8252
rect -3186 8625 -3169 8627
rect -3232 8207 -3186 8218
rect -3479 8182 -3399 8196
rect -3847 8102 -3767 8104
rect -4235 8046 -3835 8102
rect -3779 8046 -3767 8102
rect -3847 8044 -3767 8046
rect -4655 7986 -4585 8000
rect -3663 7986 -3583 7988
rect -4655 7930 -4643 7986
rect -4587 7930 -3651 7986
rect -3595 7930 -3583 7986
rect -4655 7918 -4585 7930
rect -3663 7928 -3583 7930
rect -3334 7986 -3254 7988
rect -2891 7986 -2831 7998
rect -3334 7930 -3322 7986
rect -3266 7930 -2889 7986
rect -2833 7930 -2831 7986
rect -3334 7928 -3254 7930
rect -2891 7918 -2831 7930
rect -4821 7870 -4741 7882
rect -3479 7870 -3399 7872
rect -4821 7814 -4809 7870
rect -4753 7814 -3467 7870
rect -3411 7814 -3399 7870
rect -4821 7802 -4741 7814
rect -3479 7812 -3399 7814
rect -3847 7720 -3767 7734
rect -4060 7698 -4014 7709
rect -3847 7664 -3835 7720
rect -3779 7664 -3767 7720
rect -3663 7720 -3583 7734
rect -3663 7664 -3651 7720
rect -3595 7664 -3583 7720
rect -3479 7720 -3399 7734
rect -3479 7664 -3467 7720
rect -3411 7664 -3399 7720
rect -3232 7698 -3186 7709
rect -3845 7661 -3834 7664
rect -3780 7661 -3769 7664
rect -3661 7661 -3650 7664
rect -3596 7661 -3585 7664
rect -3477 7661 -3466 7664
rect -3412 7661 -3401 7664
rect -3922 7615 -3876 7626
rect -4014 7441 -3922 7615
rect -3922 7430 -3876 7441
rect -3738 7615 -3692 7626
rect -3738 7430 -3692 7441
rect -3554 7615 -3508 7626
rect -3370 7615 -3324 7626
rect -3387 7588 -3370 7590
rect -3324 7588 -3307 7590
rect -3387 7468 -3375 7588
rect -3319 7468 -3307 7588
rect -3387 7466 -3370 7468
rect -3554 7430 -3508 7441
rect -3324 7466 -3307 7468
rect -3370 7430 -3324 7441
rect -4060 7213 -4014 7358
rect -3845 7349 -3834 7395
rect -3780 7349 -3769 7395
rect -3845 7316 -3769 7349
rect -3661 7349 -3650 7395
rect -3596 7349 -3585 7395
rect -3661 7316 -3585 7349
rect -3477 7349 -3466 7395
rect -3412 7349 -3401 7395
rect -3477 7316 -3401 7349
rect -3232 7213 -3186 7358
rect -4072 7201 -3992 7213
rect -4072 7145 -4060 7201
rect -4004 7145 -3992 7201
rect -4072 7133 -3992 7145
rect -3254 7201 -3174 7213
rect -3254 7145 -3242 7201
rect -3186 7145 -3174 7201
rect -3254 7133 -3174 7145
rect -8969 7027 -8957 7083
rect -8901 7027 -8685 7083
rect -8629 7027 -6735 7083
rect -4957 7083 -4887 7095
rect -4645 7083 -4585 7087
rect -2749 7083 -2693 10020
rect -1993 10018 -1913 10020
rect -477 10075 -407 10087
rect 563 10075 643 10077
rect 2049 10076 2129 10078
rect -477 10019 -465 10075
rect -409 10019 575 10075
rect 631 10019 643 10075
rect -477 10007 -407 10019
rect -2361 9926 -2281 9940
rect -2574 9904 -2528 9915
rect -2361 9870 -2349 9926
rect -2293 9870 -2281 9926
rect -2177 9926 -2097 9940
rect -2177 9870 -2165 9926
rect -2109 9870 -2097 9926
rect -1993 9926 -1913 9940
rect -1993 9870 -1981 9926
rect -1925 9870 -1913 9926
rect -1746 9904 -1700 9915
rect -2359 9867 -2348 9870
rect -2294 9867 -2283 9870
rect -2175 9867 -2164 9870
rect -2110 9867 -2099 9870
rect -1991 9867 -1980 9870
rect -1926 9867 -1915 9870
rect -2436 9821 -2390 9832
rect -2528 9647 -2436 9821
rect -2436 9636 -2390 9647
rect -2252 9821 -2206 9832
rect -2252 9636 -2206 9647
rect -2068 9821 -2022 9832
rect -1884 9821 -1838 9832
rect -1901 9794 -1884 9796
rect -1838 9794 -1821 9796
rect -1901 9674 -1889 9794
rect -1833 9674 -1821 9794
rect -1901 9672 -1884 9674
rect -2068 9636 -2022 9647
rect -1838 9672 -1821 9674
rect -1884 9636 -1838 9647
rect -2574 9419 -2528 9564
rect -2359 9555 -2348 9601
rect -2294 9555 -2283 9601
rect -2359 9522 -2283 9555
rect -2175 9555 -2164 9601
rect -2110 9555 -2099 9601
rect -2175 9522 -2099 9555
rect -1991 9555 -1980 9601
rect -1926 9555 -1915 9601
rect -1991 9522 -1915 9555
rect -1746 9419 -1700 9564
rect -2586 9407 -2506 9419
rect -2586 9351 -2574 9407
rect -2518 9351 -2506 9407
rect -2586 9339 -2506 9351
rect -1768 9407 -1690 9419
rect -1768 9351 -1756 9407
rect -1700 9351 -1690 9407
rect -1768 9339 -1690 9351
rect -193 9288 -137 10019
rect 563 10017 643 10019
rect 1293 10020 2061 10076
rect 2117 10020 2129 10076
rect 195 9925 275 9939
rect -18 9903 28 9914
rect 195 9869 207 9925
rect 263 9869 275 9925
rect 379 9925 459 9939
rect 379 9869 391 9925
rect 447 9869 459 9925
rect 563 9925 643 9939
rect 563 9869 575 9925
rect 631 9869 643 9925
rect 810 9903 856 9914
rect 197 9866 208 9869
rect 262 9866 273 9869
rect 381 9866 392 9869
rect 446 9866 457 9869
rect 565 9866 576 9869
rect 630 9866 641 9869
rect 120 9820 166 9831
rect 28 9646 120 9820
rect 120 9635 166 9646
rect 304 9820 350 9831
rect 304 9635 350 9646
rect 488 9820 534 9831
rect 672 9820 718 9831
rect 655 9793 672 9795
rect 718 9793 735 9795
rect 655 9673 667 9793
rect 723 9673 735 9793
rect 655 9671 672 9673
rect 488 9635 534 9646
rect 718 9671 735 9673
rect 672 9635 718 9646
rect -18 9418 28 9563
rect 197 9554 208 9600
rect 262 9554 273 9600
rect 197 9521 273 9554
rect 381 9554 392 9600
rect 446 9554 457 9600
rect 381 9521 457 9554
rect 565 9554 576 9600
rect 630 9554 641 9600
rect 565 9521 641 9554
rect 810 9418 856 9563
rect -30 9406 50 9418
rect -30 9350 -18 9406
rect 38 9350 50 9406
rect -30 9338 50 9350
rect 788 9406 866 9418
rect 788 9350 800 9406
rect 856 9350 866 9406
rect 788 9338 866 9350
rect 1141 9288 1221 9298
rect -193 9232 1153 9288
rect 1209 9232 1221 9288
rect 1141 9230 1221 9232
rect 975 9179 1045 9181
rect -193 9178 1045 9179
rect -193 9124 977 9178
rect 1033 9124 1045 9178
rect -193 9123 1045 9124
rect -193 8102 -137 9123
rect 975 9115 1045 9123
rect 471 9071 557 9075
rect 471 9015 483 9071
rect 539 9015 557 9071
rect 471 9003 557 9015
rect -18 8858 28 8869
rect 197 8867 273 8900
rect 197 8821 208 8867
rect 262 8821 273 8867
rect 381 8867 457 8900
rect 381 8821 392 8867
rect 446 8821 457 8867
rect 565 8867 641 8900
rect 565 8821 576 8867
rect 630 8821 641 8867
rect 810 8858 856 8869
rect 120 8775 166 8786
rect 103 8748 120 8750
rect 304 8775 350 8786
rect 166 8748 183 8750
rect 28 8628 115 8748
rect 171 8628 183 8748
rect 103 8626 120 8628
rect 28 8328 120 8448
rect 166 8626 183 8628
rect 287 8448 304 8450
rect 488 8775 534 8786
rect 471 8748 488 8750
rect 672 8775 718 8786
rect 534 8748 551 8750
rect 471 8628 483 8748
rect 539 8628 551 8748
rect 471 8626 488 8628
rect 350 8448 367 8450
rect 287 8328 299 8448
rect 355 8328 367 8448
rect 287 8326 304 8328
rect 120 8290 166 8301
rect 350 8326 367 8328
rect 304 8290 350 8301
rect 534 8626 551 8628
rect 655 8448 672 8450
rect 793 8748 810 8750
rect 856 8748 873 8750
rect 793 8627 805 8748
rect 861 8627 873 8748
rect 793 8625 810 8627
rect 718 8448 735 8450
rect 655 8328 667 8448
rect 723 8328 735 8448
rect 655 8326 672 8328
rect 488 8290 534 8301
rect 718 8326 735 8328
rect 672 8290 718 8301
rect 197 8252 208 8255
rect 262 8252 273 8255
rect 381 8252 392 8255
rect 446 8252 457 8255
rect 565 8252 576 8255
rect 630 8252 641 8255
rect -18 8207 28 8218
rect 195 8196 207 8252
rect 263 8196 275 8252
rect 195 8182 275 8196
rect 379 8196 391 8252
rect 447 8196 459 8252
rect 379 8182 459 8196
rect 563 8196 575 8252
rect 631 8196 643 8252
rect 856 8625 873 8627
rect 810 8207 856 8218
rect 563 8182 643 8196
rect 195 8102 275 8104
rect -193 8046 207 8102
rect 263 8046 275 8102
rect 195 8044 275 8046
rect -613 7986 -543 8000
rect 379 7986 459 7988
rect -613 7930 -601 7986
rect -545 7930 391 7986
rect 447 7930 459 7986
rect -613 7918 -543 7930
rect 379 7928 459 7930
rect 708 7986 788 7988
rect 1151 7986 1211 7998
rect 708 7930 720 7986
rect 776 7930 1153 7986
rect 1209 7930 1211 7986
rect 708 7928 788 7930
rect 1151 7918 1211 7930
rect -779 7870 -699 7882
rect 563 7870 643 7872
rect -779 7814 -767 7870
rect -711 7814 575 7870
rect 631 7814 643 7870
rect -779 7802 -699 7814
rect 563 7812 643 7814
rect 195 7720 275 7734
rect -18 7698 28 7709
rect 195 7664 207 7720
rect 263 7664 275 7720
rect 379 7720 459 7734
rect 379 7664 391 7720
rect 447 7664 459 7720
rect 563 7720 643 7734
rect 563 7664 575 7720
rect 631 7664 643 7720
rect 810 7698 856 7709
rect 197 7661 208 7664
rect 262 7661 273 7664
rect 381 7661 392 7664
rect 446 7661 457 7664
rect 565 7661 576 7664
rect 630 7661 641 7664
rect 120 7615 166 7626
rect 28 7441 120 7615
rect 120 7430 166 7441
rect 304 7615 350 7626
rect 304 7430 350 7441
rect 488 7615 534 7626
rect 672 7615 718 7626
rect 655 7588 672 7590
rect 718 7588 735 7590
rect 655 7468 667 7588
rect 723 7468 735 7588
rect 655 7466 672 7468
rect 488 7430 534 7441
rect 718 7466 735 7468
rect 672 7430 718 7441
rect -18 7213 28 7358
rect 197 7349 208 7395
rect 262 7349 273 7395
rect 197 7316 273 7349
rect 381 7349 392 7395
rect 446 7349 457 7395
rect 381 7316 457 7349
rect 565 7349 576 7395
rect 630 7349 641 7395
rect 565 7316 641 7349
rect 810 7213 856 7358
rect -30 7201 50 7213
rect -30 7145 -18 7201
rect 38 7145 50 7201
rect -30 7133 50 7145
rect 788 7201 868 7213
rect 788 7145 800 7201
rect 856 7145 868 7201
rect 788 7133 868 7145
rect -4957 7027 -4945 7083
rect -4889 7027 -4643 7083
rect -4587 7027 -2693 7083
rect -915 7083 -845 7095
rect -603 7083 -543 7087
rect 1293 7083 1349 10020
rect 2049 10018 2129 10020
rect 3565 10075 3635 10087
rect 4605 10075 4685 10077
rect 6091 10076 6171 10078
rect 3565 10019 3577 10075
rect 3633 10019 4617 10075
rect 4673 10019 4685 10075
rect 3565 10007 3635 10019
rect 1681 9926 1761 9940
rect 1468 9904 1514 9915
rect 1681 9870 1693 9926
rect 1749 9870 1761 9926
rect 1865 9926 1945 9940
rect 1865 9870 1877 9926
rect 1933 9870 1945 9926
rect 2049 9926 2129 9940
rect 2049 9870 2061 9926
rect 2117 9870 2129 9926
rect 2296 9904 2342 9915
rect 1683 9867 1694 9870
rect 1748 9867 1759 9870
rect 1867 9867 1878 9870
rect 1932 9867 1943 9870
rect 2051 9867 2062 9870
rect 2116 9867 2127 9870
rect 1606 9821 1652 9832
rect 1514 9647 1606 9821
rect 1606 9636 1652 9647
rect 1790 9821 1836 9832
rect 1790 9636 1836 9647
rect 1974 9821 2020 9832
rect 2158 9821 2204 9832
rect 2141 9794 2158 9796
rect 2204 9794 2221 9796
rect 2141 9674 2153 9794
rect 2209 9674 2221 9794
rect 2141 9672 2158 9674
rect 1974 9636 2020 9647
rect 2204 9672 2221 9674
rect 2158 9636 2204 9647
rect 1468 9419 1514 9564
rect 1683 9555 1694 9601
rect 1748 9555 1759 9601
rect 1683 9522 1759 9555
rect 1867 9555 1878 9601
rect 1932 9555 1943 9601
rect 1867 9522 1943 9555
rect 2051 9555 2062 9601
rect 2116 9555 2127 9601
rect 2051 9522 2127 9555
rect 2296 9419 2342 9564
rect 1456 9407 1536 9419
rect 1456 9351 1468 9407
rect 1524 9351 1536 9407
rect 1456 9339 1536 9351
rect 2274 9407 2352 9419
rect 2274 9351 2286 9407
rect 2342 9351 2352 9407
rect 2274 9339 2352 9351
rect 3849 9288 3905 10019
rect 4605 10017 4685 10019
rect 5335 10020 6103 10076
rect 6159 10020 6171 10076
rect 4237 9925 4317 9939
rect 4024 9903 4070 9914
rect 4237 9869 4249 9925
rect 4305 9869 4317 9925
rect 4421 9925 4501 9939
rect 4421 9869 4433 9925
rect 4489 9869 4501 9925
rect 4605 9925 4685 9939
rect 4605 9869 4617 9925
rect 4673 9869 4685 9925
rect 4852 9903 4898 9914
rect 4239 9866 4250 9869
rect 4304 9866 4315 9869
rect 4423 9866 4434 9869
rect 4488 9866 4499 9869
rect 4607 9866 4618 9869
rect 4672 9866 4683 9869
rect 4162 9820 4208 9831
rect 4070 9646 4162 9820
rect 4162 9635 4208 9646
rect 4346 9820 4392 9831
rect 4346 9635 4392 9646
rect 4530 9820 4576 9831
rect 4714 9820 4760 9831
rect 4697 9793 4714 9795
rect 4760 9793 4777 9795
rect 4697 9673 4709 9793
rect 4765 9673 4777 9793
rect 4697 9671 4714 9673
rect 4530 9635 4576 9646
rect 4760 9671 4777 9673
rect 4714 9635 4760 9646
rect 4024 9418 4070 9563
rect 4239 9554 4250 9600
rect 4304 9554 4315 9600
rect 4239 9521 4315 9554
rect 4423 9554 4434 9600
rect 4488 9554 4499 9600
rect 4423 9521 4499 9554
rect 4607 9554 4618 9600
rect 4672 9554 4683 9600
rect 4607 9521 4683 9554
rect 4852 9418 4898 9563
rect 4012 9406 4092 9418
rect 4012 9350 4024 9406
rect 4080 9350 4092 9406
rect 4012 9338 4092 9350
rect 4830 9406 4908 9418
rect 4830 9350 4842 9406
rect 4898 9350 4908 9406
rect 4830 9338 4908 9350
rect 5183 9288 5263 9298
rect 3849 9232 5195 9288
rect 5251 9232 5263 9288
rect 5183 9230 5263 9232
rect 5017 9179 5087 9181
rect 3849 9178 5087 9179
rect 3849 9124 5019 9178
rect 5075 9124 5087 9178
rect 3849 9123 5087 9124
rect 3849 8102 3905 9123
rect 5017 9115 5087 9123
rect 4513 9071 4599 9075
rect 4513 9015 4525 9071
rect 4581 9015 4599 9071
rect 4513 9003 4599 9015
rect 4024 8858 4070 8869
rect 4239 8867 4315 8900
rect 4239 8821 4250 8867
rect 4304 8821 4315 8867
rect 4423 8867 4499 8900
rect 4423 8821 4434 8867
rect 4488 8821 4499 8867
rect 4607 8867 4683 8900
rect 4607 8821 4618 8867
rect 4672 8821 4683 8867
rect 4852 8858 4898 8869
rect 4162 8775 4208 8786
rect 4145 8748 4162 8750
rect 4346 8775 4392 8786
rect 4208 8748 4225 8750
rect 4070 8628 4157 8748
rect 4213 8628 4225 8748
rect 4145 8626 4162 8628
rect 4070 8328 4162 8448
rect 4208 8626 4225 8628
rect 4329 8448 4346 8450
rect 4530 8775 4576 8786
rect 4513 8748 4530 8750
rect 4714 8775 4760 8786
rect 4576 8748 4593 8750
rect 4513 8628 4525 8748
rect 4581 8628 4593 8748
rect 4513 8626 4530 8628
rect 4392 8448 4409 8450
rect 4329 8328 4341 8448
rect 4397 8328 4409 8448
rect 4329 8326 4346 8328
rect 4162 8290 4208 8301
rect 4392 8326 4409 8328
rect 4346 8290 4392 8301
rect 4576 8626 4593 8628
rect 4697 8448 4714 8450
rect 4835 8748 4852 8750
rect 4898 8748 4915 8750
rect 4835 8627 4847 8748
rect 4903 8627 4915 8748
rect 4835 8625 4852 8627
rect 4760 8448 4777 8450
rect 4697 8328 4709 8448
rect 4765 8328 4777 8448
rect 4697 8326 4714 8328
rect 4530 8290 4576 8301
rect 4760 8326 4777 8328
rect 4714 8290 4760 8301
rect 4239 8252 4250 8255
rect 4304 8252 4315 8255
rect 4423 8252 4434 8255
rect 4488 8252 4499 8255
rect 4607 8252 4618 8255
rect 4672 8252 4683 8255
rect 4024 8207 4070 8218
rect 4237 8196 4249 8252
rect 4305 8196 4317 8252
rect 4237 8182 4317 8196
rect 4421 8196 4433 8252
rect 4489 8196 4501 8252
rect 4421 8182 4501 8196
rect 4605 8196 4617 8252
rect 4673 8196 4685 8252
rect 4898 8625 4915 8627
rect 4852 8207 4898 8218
rect 4605 8182 4685 8196
rect 4237 8102 4317 8104
rect 3849 8046 4249 8102
rect 4305 8046 4317 8102
rect 4237 8044 4317 8046
rect 3429 7986 3499 8000
rect 4421 7986 4501 7988
rect 3429 7930 3441 7986
rect 3497 7930 4433 7986
rect 4489 7930 4501 7986
rect 3429 7918 3499 7930
rect 4421 7928 4501 7930
rect 4750 7986 4830 7988
rect 5193 7986 5253 7998
rect 4750 7930 4762 7986
rect 4818 7930 5195 7986
rect 5251 7930 5253 7986
rect 4750 7928 4830 7930
rect 5193 7918 5253 7930
rect 3263 7870 3343 7882
rect 4605 7870 4685 7872
rect 3263 7814 3275 7870
rect 3331 7814 4617 7870
rect 4673 7814 4685 7870
rect 3263 7802 3343 7814
rect 4605 7812 4685 7814
rect 4237 7720 4317 7734
rect 4024 7698 4070 7709
rect 4237 7664 4249 7720
rect 4305 7664 4317 7720
rect 4421 7720 4501 7734
rect 4421 7664 4433 7720
rect 4489 7664 4501 7720
rect 4605 7720 4685 7734
rect 4605 7664 4617 7720
rect 4673 7664 4685 7720
rect 4852 7698 4898 7709
rect 4239 7661 4250 7664
rect 4304 7661 4315 7664
rect 4423 7661 4434 7664
rect 4488 7661 4499 7664
rect 4607 7661 4618 7664
rect 4672 7661 4683 7664
rect 4162 7615 4208 7626
rect 4070 7441 4162 7615
rect 4162 7430 4208 7441
rect 4346 7615 4392 7626
rect 4346 7430 4392 7441
rect 4530 7615 4576 7626
rect 4714 7615 4760 7626
rect 4697 7588 4714 7590
rect 4760 7588 4777 7590
rect 4697 7468 4709 7588
rect 4765 7468 4777 7588
rect 4697 7466 4714 7468
rect 4530 7430 4576 7441
rect 4760 7466 4777 7468
rect 4714 7430 4760 7441
rect 4024 7213 4070 7358
rect 4239 7349 4250 7395
rect 4304 7349 4315 7395
rect 4239 7316 4315 7349
rect 4423 7349 4434 7395
rect 4488 7349 4499 7395
rect 4423 7316 4499 7349
rect 4607 7349 4618 7395
rect 4672 7349 4683 7395
rect 4607 7316 4683 7349
rect 4852 7213 4898 7358
rect 4012 7201 4092 7213
rect 4012 7145 4024 7201
rect 4080 7145 4092 7201
rect 4012 7133 4092 7145
rect 4830 7201 4910 7213
rect 4830 7145 4842 7201
rect 4898 7145 4910 7201
rect 4830 7133 4910 7145
rect -915 7027 -903 7083
rect -847 7027 -601 7083
rect -545 7027 1349 7083
rect 3127 7083 3197 7095
rect 3439 7083 3499 7087
rect 5335 7083 5391 10020
rect 6091 10018 6171 10020
rect 7607 10075 7677 10087
rect 8647 10075 8727 10077
rect 10133 10076 10213 10078
rect 7607 10019 7619 10075
rect 7675 10019 8659 10075
rect 8715 10019 8727 10075
rect 7607 10007 7677 10019
rect 5723 9926 5803 9940
rect 5510 9904 5556 9915
rect 5723 9870 5735 9926
rect 5791 9870 5803 9926
rect 5907 9926 5987 9940
rect 5907 9870 5919 9926
rect 5975 9870 5987 9926
rect 6091 9926 6171 9940
rect 6091 9870 6103 9926
rect 6159 9870 6171 9926
rect 6338 9904 6384 9915
rect 5725 9867 5736 9870
rect 5790 9867 5801 9870
rect 5909 9867 5920 9870
rect 5974 9867 5985 9870
rect 6093 9867 6104 9870
rect 6158 9867 6169 9870
rect 5648 9821 5694 9832
rect 5556 9647 5648 9821
rect 5648 9636 5694 9647
rect 5832 9821 5878 9832
rect 5832 9636 5878 9647
rect 6016 9821 6062 9832
rect 6200 9821 6246 9832
rect 6183 9794 6200 9796
rect 6246 9794 6263 9796
rect 6183 9674 6195 9794
rect 6251 9674 6263 9794
rect 6183 9672 6200 9674
rect 6016 9636 6062 9647
rect 6246 9672 6263 9674
rect 6200 9636 6246 9647
rect 5510 9419 5556 9564
rect 5725 9555 5736 9601
rect 5790 9555 5801 9601
rect 5725 9522 5801 9555
rect 5909 9555 5920 9601
rect 5974 9555 5985 9601
rect 5909 9522 5985 9555
rect 6093 9555 6104 9601
rect 6158 9555 6169 9601
rect 6093 9522 6169 9555
rect 6338 9419 6384 9564
rect 5498 9407 5578 9419
rect 5498 9351 5510 9407
rect 5566 9351 5578 9407
rect 5498 9339 5578 9351
rect 6316 9407 6394 9419
rect 6316 9351 6328 9407
rect 6384 9351 6394 9407
rect 6316 9339 6394 9351
rect 7891 9288 7947 10019
rect 8647 10017 8727 10019
rect 9377 10020 10145 10076
rect 10201 10020 10213 10076
rect 8279 9925 8359 9939
rect 8066 9903 8112 9914
rect 8279 9869 8291 9925
rect 8347 9869 8359 9925
rect 8463 9925 8543 9939
rect 8463 9869 8475 9925
rect 8531 9869 8543 9925
rect 8647 9925 8727 9939
rect 8647 9869 8659 9925
rect 8715 9869 8727 9925
rect 8894 9903 8940 9914
rect 8281 9866 8292 9869
rect 8346 9866 8357 9869
rect 8465 9866 8476 9869
rect 8530 9866 8541 9869
rect 8649 9866 8660 9869
rect 8714 9866 8725 9869
rect 8204 9820 8250 9831
rect 8112 9646 8204 9820
rect 8204 9635 8250 9646
rect 8388 9820 8434 9831
rect 8388 9635 8434 9646
rect 8572 9820 8618 9831
rect 8756 9820 8802 9831
rect 8739 9793 8756 9795
rect 8802 9793 8819 9795
rect 8739 9673 8751 9793
rect 8807 9673 8819 9793
rect 8739 9671 8756 9673
rect 8572 9635 8618 9646
rect 8802 9671 8819 9673
rect 8756 9635 8802 9646
rect 8066 9418 8112 9563
rect 8281 9554 8292 9600
rect 8346 9554 8357 9600
rect 8281 9521 8357 9554
rect 8465 9554 8476 9600
rect 8530 9554 8541 9600
rect 8465 9521 8541 9554
rect 8649 9554 8660 9600
rect 8714 9554 8725 9600
rect 8649 9521 8725 9554
rect 8894 9418 8940 9563
rect 8054 9406 8134 9418
rect 8054 9350 8066 9406
rect 8122 9350 8134 9406
rect 8054 9338 8134 9350
rect 8872 9406 8950 9418
rect 8872 9350 8884 9406
rect 8940 9350 8950 9406
rect 8872 9338 8950 9350
rect 9225 9288 9305 9298
rect 7891 9232 9237 9288
rect 9293 9232 9305 9288
rect 9225 9230 9305 9232
rect 9059 9179 9129 9181
rect 7891 9178 9129 9179
rect 7891 9124 9061 9178
rect 9117 9124 9129 9178
rect 7891 9123 9129 9124
rect 7891 8102 7947 9123
rect 9059 9115 9129 9123
rect 8555 9071 8641 9075
rect 8555 9015 8567 9071
rect 8623 9015 8641 9071
rect 8555 9003 8641 9015
rect 8066 8858 8112 8869
rect 8281 8867 8357 8900
rect 8281 8821 8292 8867
rect 8346 8821 8357 8867
rect 8465 8867 8541 8900
rect 8465 8821 8476 8867
rect 8530 8821 8541 8867
rect 8649 8867 8725 8900
rect 8649 8821 8660 8867
rect 8714 8821 8725 8867
rect 8894 8858 8940 8869
rect 8204 8775 8250 8786
rect 8187 8748 8204 8750
rect 8388 8775 8434 8786
rect 8250 8748 8267 8750
rect 8112 8628 8199 8748
rect 8255 8628 8267 8748
rect 8187 8626 8204 8628
rect 8112 8328 8204 8448
rect 8250 8626 8267 8628
rect 8371 8448 8388 8450
rect 8572 8775 8618 8786
rect 8555 8748 8572 8750
rect 8756 8775 8802 8786
rect 8618 8748 8635 8750
rect 8555 8628 8567 8748
rect 8623 8628 8635 8748
rect 8555 8626 8572 8628
rect 8434 8448 8451 8450
rect 8371 8328 8383 8448
rect 8439 8328 8451 8448
rect 8371 8326 8388 8328
rect 8204 8290 8250 8301
rect 8434 8326 8451 8328
rect 8388 8290 8434 8301
rect 8618 8626 8635 8628
rect 8739 8448 8756 8450
rect 8877 8748 8894 8750
rect 8940 8748 8957 8750
rect 8877 8627 8889 8748
rect 8945 8627 8957 8748
rect 8877 8625 8894 8627
rect 8802 8448 8819 8450
rect 8739 8328 8751 8448
rect 8807 8328 8819 8448
rect 8739 8326 8756 8328
rect 8572 8290 8618 8301
rect 8802 8326 8819 8328
rect 8756 8290 8802 8301
rect 8281 8252 8292 8255
rect 8346 8252 8357 8255
rect 8465 8252 8476 8255
rect 8530 8252 8541 8255
rect 8649 8252 8660 8255
rect 8714 8252 8725 8255
rect 8066 8207 8112 8218
rect 8279 8196 8291 8252
rect 8347 8196 8359 8252
rect 8279 8182 8359 8196
rect 8463 8196 8475 8252
rect 8531 8196 8543 8252
rect 8463 8182 8543 8196
rect 8647 8196 8659 8252
rect 8715 8196 8727 8252
rect 8940 8625 8957 8627
rect 8894 8207 8940 8218
rect 8647 8182 8727 8196
rect 8279 8102 8359 8104
rect 7891 8046 8291 8102
rect 8347 8046 8359 8102
rect 8279 8044 8359 8046
rect 7471 7986 7541 8000
rect 8463 7986 8543 7988
rect 7471 7930 7483 7986
rect 7539 7930 8475 7986
rect 8531 7930 8543 7986
rect 7471 7918 7541 7930
rect 8463 7928 8543 7930
rect 8792 7986 8872 7988
rect 9235 7986 9295 7998
rect 8792 7930 8804 7986
rect 8860 7930 9237 7986
rect 9293 7930 9295 7986
rect 8792 7928 8872 7930
rect 9235 7918 9295 7930
rect 7305 7870 7385 7882
rect 8647 7870 8727 7872
rect 7305 7814 7317 7870
rect 7373 7814 8659 7870
rect 8715 7814 8727 7870
rect 7305 7802 7385 7814
rect 8647 7812 8727 7814
rect 8279 7720 8359 7734
rect 8066 7698 8112 7709
rect 8279 7664 8291 7720
rect 8347 7664 8359 7720
rect 8463 7720 8543 7734
rect 8463 7664 8475 7720
rect 8531 7664 8543 7720
rect 8647 7720 8727 7734
rect 8647 7664 8659 7720
rect 8715 7664 8727 7720
rect 8894 7698 8940 7709
rect 8281 7661 8292 7664
rect 8346 7661 8357 7664
rect 8465 7661 8476 7664
rect 8530 7661 8541 7664
rect 8649 7661 8660 7664
rect 8714 7661 8725 7664
rect 8204 7615 8250 7626
rect 8112 7441 8204 7615
rect 8204 7430 8250 7441
rect 8388 7615 8434 7626
rect 8388 7430 8434 7441
rect 8572 7615 8618 7626
rect 8756 7615 8802 7626
rect 8739 7588 8756 7590
rect 8802 7588 8819 7590
rect 8739 7468 8751 7588
rect 8807 7468 8819 7588
rect 8739 7466 8756 7468
rect 8572 7430 8618 7441
rect 8802 7466 8819 7468
rect 8756 7430 8802 7441
rect 8066 7213 8112 7358
rect 8281 7349 8292 7395
rect 8346 7349 8357 7395
rect 8281 7316 8357 7349
rect 8465 7349 8476 7395
rect 8530 7349 8541 7395
rect 8465 7316 8541 7349
rect 8649 7349 8660 7395
rect 8714 7349 8725 7395
rect 8649 7316 8725 7349
rect 8894 7213 8940 7358
rect 8054 7201 8134 7213
rect 8054 7145 8066 7201
rect 8122 7145 8134 7201
rect 8054 7133 8134 7145
rect 8872 7201 8952 7213
rect 8872 7145 8884 7201
rect 8940 7145 8952 7201
rect 8872 7133 8952 7145
rect 3127 7027 3139 7083
rect 3195 7027 3441 7083
rect 3497 7027 5391 7083
rect 7169 7083 7239 7095
rect 7481 7083 7541 7087
rect 9377 7083 9433 10020
rect 10133 10018 10213 10020
rect 11649 10075 11719 10087
rect 12689 10075 12769 10077
rect 14175 10076 14255 10078
rect 11649 10019 11661 10075
rect 11717 10019 12701 10075
rect 12757 10019 12769 10075
rect 11649 10007 11719 10019
rect 9765 9926 9845 9940
rect 9552 9904 9598 9915
rect 9765 9870 9777 9926
rect 9833 9870 9845 9926
rect 9949 9926 10029 9940
rect 9949 9870 9961 9926
rect 10017 9870 10029 9926
rect 10133 9926 10213 9940
rect 10133 9870 10145 9926
rect 10201 9870 10213 9926
rect 10380 9904 10426 9915
rect 9767 9867 9778 9870
rect 9832 9867 9843 9870
rect 9951 9867 9962 9870
rect 10016 9867 10027 9870
rect 10135 9867 10146 9870
rect 10200 9867 10211 9870
rect 9690 9821 9736 9832
rect 9598 9647 9690 9821
rect 9690 9636 9736 9647
rect 9874 9821 9920 9832
rect 9874 9636 9920 9647
rect 10058 9821 10104 9832
rect 10242 9821 10288 9832
rect 10225 9794 10242 9796
rect 10288 9794 10305 9796
rect 10225 9674 10237 9794
rect 10293 9674 10305 9794
rect 10225 9672 10242 9674
rect 10058 9636 10104 9647
rect 10288 9672 10305 9674
rect 10242 9636 10288 9647
rect 9552 9419 9598 9564
rect 9767 9555 9778 9601
rect 9832 9555 9843 9601
rect 9767 9522 9843 9555
rect 9951 9555 9962 9601
rect 10016 9555 10027 9601
rect 9951 9522 10027 9555
rect 10135 9555 10146 9601
rect 10200 9555 10211 9601
rect 10135 9522 10211 9555
rect 10380 9419 10426 9564
rect 9540 9407 9620 9419
rect 9540 9351 9552 9407
rect 9608 9351 9620 9407
rect 9540 9339 9620 9351
rect 10358 9407 10436 9419
rect 10358 9351 10370 9407
rect 10426 9351 10436 9407
rect 10358 9339 10436 9351
rect 11933 9288 11989 10019
rect 12689 10017 12769 10019
rect 13419 10020 14187 10076
rect 14243 10020 14255 10076
rect 12321 9925 12401 9939
rect 12108 9903 12154 9914
rect 12321 9869 12333 9925
rect 12389 9869 12401 9925
rect 12505 9925 12585 9939
rect 12505 9869 12517 9925
rect 12573 9869 12585 9925
rect 12689 9925 12769 9939
rect 12689 9869 12701 9925
rect 12757 9869 12769 9925
rect 12936 9903 12982 9914
rect 12323 9866 12334 9869
rect 12388 9866 12399 9869
rect 12507 9866 12518 9869
rect 12572 9866 12583 9869
rect 12691 9866 12702 9869
rect 12756 9866 12767 9869
rect 12246 9820 12292 9831
rect 12154 9646 12246 9820
rect 12246 9635 12292 9646
rect 12430 9820 12476 9831
rect 12430 9635 12476 9646
rect 12614 9820 12660 9831
rect 12798 9820 12844 9831
rect 12781 9793 12798 9795
rect 12844 9793 12861 9795
rect 12781 9673 12793 9793
rect 12849 9673 12861 9793
rect 12781 9671 12798 9673
rect 12614 9635 12660 9646
rect 12844 9671 12861 9673
rect 12798 9635 12844 9646
rect 12108 9418 12154 9563
rect 12323 9554 12334 9600
rect 12388 9554 12399 9600
rect 12323 9521 12399 9554
rect 12507 9554 12518 9600
rect 12572 9554 12583 9600
rect 12507 9521 12583 9554
rect 12691 9554 12702 9600
rect 12756 9554 12767 9600
rect 12691 9521 12767 9554
rect 12936 9418 12982 9563
rect 12096 9406 12176 9418
rect 12096 9350 12108 9406
rect 12164 9350 12176 9406
rect 12096 9338 12176 9350
rect 12914 9406 12992 9418
rect 12914 9350 12926 9406
rect 12982 9350 12992 9406
rect 12914 9338 12992 9350
rect 13267 9288 13347 9298
rect 11933 9232 13279 9288
rect 13335 9232 13347 9288
rect 13267 9230 13347 9232
rect 13101 9179 13171 9181
rect 11933 9178 13171 9179
rect 11933 9124 13103 9178
rect 13159 9124 13171 9178
rect 11933 9123 13171 9124
rect 11933 8102 11989 9123
rect 13101 9115 13171 9123
rect 12597 9071 12683 9075
rect 12597 9015 12609 9071
rect 12665 9015 12683 9071
rect 12597 9003 12683 9015
rect 12108 8858 12154 8869
rect 12323 8867 12399 8900
rect 12323 8821 12334 8867
rect 12388 8821 12399 8867
rect 12507 8867 12583 8900
rect 12507 8821 12518 8867
rect 12572 8821 12583 8867
rect 12691 8867 12767 8900
rect 12691 8821 12702 8867
rect 12756 8821 12767 8867
rect 12936 8858 12982 8869
rect 12246 8775 12292 8786
rect 12229 8748 12246 8750
rect 12430 8775 12476 8786
rect 12292 8748 12309 8750
rect 12154 8628 12241 8748
rect 12297 8628 12309 8748
rect 12229 8626 12246 8628
rect 12154 8328 12246 8448
rect 12292 8626 12309 8628
rect 12413 8448 12430 8450
rect 12614 8775 12660 8786
rect 12597 8748 12614 8750
rect 12798 8775 12844 8786
rect 12660 8748 12677 8750
rect 12597 8628 12609 8748
rect 12665 8628 12677 8748
rect 12597 8626 12614 8628
rect 12476 8448 12493 8450
rect 12413 8328 12425 8448
rect 12481 8328 12493 8448
rect 12413 8326 12430 8328
rect 12246 8290 12292 8301
rect 12476 8326 12493 8328
rect 12430 8290 12476 8301
rect 12660 8626 12677 8628
rect 12781 8448 12798 8450
rect 12919 8748 12936 8750
rect 12982 8748 12999 8750
rect 12919 8627 12931 8748
rect 12987 8627 12999 8748
rect 12919 8625 12936 8627
rect 12844 8448 12861 8450
rect 12781 8328 12793 8448
rect 12849 8328 12861 8448
rect 12781 8326 12798 8328
rect 12614 8290 12660 8301
rect 12844 8326 12861 8328
rect 12798 8290 12844 8301
rect 12323 8252 12334 8255
rect 12388 8252 12399 8255
rect 12507 8252 12518 8255
rect 12572 8252 12583 8255
rect 12691 8252 12702 8255
rect 12756 8252 12767 8255
rect 12108 8207 12154 8218
rect 12321 8196 12333 8252
rect 12389 8196 12401 8252
rect 12321 8182 12401 8196
rect 12505 8196 12517 8252
rect 12573 8196 12585 8252
rect 12505 8182 12585 8196
rect 12689 8196 12701 8252
rect 12757 8196 12769 8252
rect 12982 8625 12999 8627
rect 12936 8207 12982 8218
rect 12689 8182 12769 8196
rect 12321 8102 12401 8104
rect 11933 8046 12333 8102
rect 12389 8046 12401 8102
rect 12321 8044 12401 8046
rect 11513 7986 11583 8000
rect 12505 7986 12585 7988
rect 11513 7930 11525 7986
rect 11581 7930 12517 7986
rect 12573 7930 12585 7986
rect 11513 7918 11583 7930
rect 12505 7928 12585 7930
rect 12834 7986 12914 7988
rect 13277 7986 13337 7998
rect 12834 7930 12846 7986
rect 12902 7930 13279 7986
rect 13335 7930 13337 7986
rect 12834 7928 12914 7930
rect 13277 7918 13337 7930
rect 11347 7870 11427 7882
rect 12689 7870 12769 7872
rect 11347 7814 11359 7870
rect 11415 7814 12701 7870
rect 12757 7814 12769 7870
rect 11347 7802 11427 7814
rect 12689 7812 12769 7814
rect 12321 7720 12401 7734
rect 12108 7698 12154 7709
rect 12321 7664 12333 7720
rect 12389 7664 12401 7720
rect 12505 7720 12585 7734
rect 12505 7664 12517 7720
rect 12573 7664 12585 7720
rect 12689 7720 12769 7734
rect 12689 7664 12701 7720
rect 12757 7664 12769 7720
rect 12936 7698 12982 7709
rect 12323 7661 12334 7664
rect 12388 7661 12399 7664
rect 12507 7661 12518 7664
rect 12572 7661 12583 7664
rect 12691 7661 12702 7664
rect 12756 7661 12767 7664
rect 12246 7615 12292 7626
rect 12154 7441 12246 7615
rect 12246 7430 12292 7441
rect 12430 7615 12476 7626
rect 12430 7430 12476 7441
rect 12614 7615 12660 7626
rect 12798 7615 12844 7626
rect 12781 7588 12798 7590
rect 12844 7588 12861 7590
rect 12781 7468 12793 7588
rect 12849 7468 12861 7588
rect 12781 7466 12798 7468
rect 12614 7430 12660 7441
rect 12844 7466 12861 7468
rect 12798 7430 12844 7441
rect 12108 7213 12154 7358
rect 12323 7349 12334 7395
rect 12388 7349 12399 7395
rect 12323 7316 12399 7349
rect 12507 7349 12518 7395
rect 12572 7349 12583 7395
rect 12507 7316 12583 7349
rect 12691 7349 12702 7395
rect 12756 7349 12767 7395
rect 12691 7316 12767 7349
rect 12936 7213 12982 7358
rect 12096 7201 12176 7213
rect 12096 7145 12108 7201
rect 12164 7145 12176 7201
rect 12096 7133 12176 7145
rect 12914 7201 12994 7213
rect 12914 7145 12926 7201
rect 12982 7145 12994 7201
rect 12914 7133 12994 7145
rect 7169 7027 7181 7083
rect 7237 7027 7483 7083
rect 7539 7027 9433 7083
rect 11211 7083 11281 7095
rect 11523 7083 11583 7087
rect 13419 7083 13475 10020
rect 14175 10018 14255 10020
rect 13807 9926 13887 9940
rect 13594 9904 13640 9915
rect 13807 9870 13819 9926
rect 13875 9870 13887 9926
rect 13991 9926 14071 9940
rect 13991 9870 14003 9926
rect 14059 9870 14071 9926
rect 14175 9926 14255 9940
rect 14175 9870 14187 9926
rect 14243 9870 14255 9926
rect 14422 9904 14468 9915
rect 13809 9867 13820 9870
rect 13874 9867 13885 9870
rect 13993 9867 14004 9870
rect 14058 9867 14069 9870
rect 14177 9867 14188 9870
rect 14242 9867 14253 9870
rect 13732 9821 13778 9832
rect 13640 9647 13732 9821
rect 13732 9636 13778 9647
rect 13916 9821 13962 9832
rect 13916 9636 13962 9647
rect 14100 9821 14146 9832
rect 14284 9821 14330 9832
rect 14267 9794 14284 9796
rect 14330 9794 14347 9796
rect 14267 9674 14279 9794
rect 14335 9674 14347 9794
rect 14267 9672 14284 9674
rect 14100 9636 14146 9647
rect 14330 9672 14347 9674
rect 14284 9636 14330 9647
rect 13594 9419 13640 9564
rect 13809 9555 13820 9601
rect 13874 9555 13885 9601
rect 13809 9522 13885 9555
rect 13993 9555 14004 9601
rect 14058 9555 14069 9601
rect 13993 9522 14069 9555
rect 14177 9555 14188 9601
rect 14242 9555 14253 9601
rect 14177 9522 14253 9555
rect 14422 9419 14468 9564
rect 13582 9407 13662 9419
rect 13582 9351 13594 9407
rect 13650 9351 13662 9407
rect 13582 9339 13662 9351
rect 14400 9407 14478 9419
rect 14400 9351 14412 9407
rect 14468 9351 14478 9407
rect 14400 9339 14478 9351
rect 11211 7027 11223 7083
rect 11279 7027 11525 7083
rect 11581 7027 13475 7083
rect -12908 7015 -12822 7027
rect -12699 7015 -12639 7027
rect -8969 7015 -8899 7027
rect -8687 7015 -8627 7027
rect -4957 7015 -4887 7027
rect -4645 7015 -4585 7027
rect -915 7015 -845 7027
rect -603 7015 -543 7027
rect 3127 7015 3197 7027
rect 3439 7015 3499 7027
rect 7169 7015 7239 7027
rect 7481 7015 7541 7027
rect 11211 7015 11281 7027
rect 11523 7015 11583 7027
rect -12861 6434 -2430 6477
rect -12861 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -12861 6097 -2430 6134
rect -13680 4940 -13603 4954
rect -12380 4940 -12294 4954
rect -13680 4939 -12366 4940
rect -13680 4881 -13665 4939
rect -13607 4881 -12366 4939
rect -13680 4880 -12366 4881
rect -12306 4880 -12294 4940
rect -13680 4867 -13603 4880
rect -12380 4866 -12294 4880
rect -12085 3179 -12007 6097
rect -10476 5430 -10396 6097
rect -11031 5358 -9891 5430
rect -11031 5312 -10779 5358
rect -10733 5312 -10539 5358
rect -10493 5312 -10299 5358
rect -10253 5312 -10059 5358
rect -10013 5312 -9891 5358
rect -11031 5290 -9891 5312
rect -10911 5167 -10861 5290
rect -10911 4933 -10909 5167
rect -10863 4933 -10861 5167
rect -10741 5192 -10691 5220
rect -10741 4958 -10739 5192
rect -10693 4958 -10691 5192
rect -10741 4940 -10691 4958
rect -10571 5167 -10521 5290
rect -10911 4880 -10861 4933
rect -10771 4936 -10671 4940
rect -10771 4884 -10747 4936
rect -10695 4884 -10671 4936
rect -10771 4880 -10671 4884
rect -10571 4933 -10569 5167
rect -10523 4933 -10521 5167
rect -10571 4880 -10521 4933
rect -10401 5192 -10351 5220
rect -10401 4958 -10399 5192
rect -10353 4958 -10351 5192
rect -10741 4830 -10691 4880
rect -10401 4830 -10351 4958
rect -10231 5167 -10181 5290
rect -10231 4933 -10229 5167
rect -10183 4933 -10181 5167
rect -10231 4880 -10181 4933
rect -10061 5167 -10011 5220
rect -10061 4933 -10059 5167
rect -10013 4933 -10011 5167
rect -10061 4830 -10011 4933
rect -10741 4770 -10351 4830
rect -10301 4823 -10011 4830
rect -10301 4777 -10274 4823
rect -10228 4777 -10011 4823
rect -10301 4770 -10011 4777
rect -10741 4650 -10691 4770
rect -10401 4650 -10351 4770
rect -10741 4590 -10351 4650
rect -10211 4676 -10111 4680
rect -10211 4624 -10187 4676
rect -10135 4624 -10111 4676
rect -10211 4620 -10111 4624
rect -10911 4478 -10861 4540
rect -10911 4432 -10909 4478
rect -10863 4432 -10861 4478
rect -10911 4300 -10861 4432
rect -10741 4478 -10691 4590
rect -10741 4432 -10739 4478
rect -10693 4432 -10691 4478
rect -10741 4370 -10691 4432
rect -10571 4478 -10521 4540
rect -10571 4432 -10569 4478
rect -10523 4432 -10521 4478
rect -10571 4300 -10521 4432
rect -10401 4478 -10351 4590
rect -10401 4432 -10399 4478
rect -10353 4432 -10351 4478
rect -10401 4370 -10351 4432
rect -10231 4478 -10181 4540
rect -10231 4432 -10229 4478
rect -10183 4432 -10181 4478
rect -10231 4300 -10181 4432
rect -10061 4478 -10011 4770
rect -9396 4487 -9316 6097
rect -8216 5157 -8136 6097
rect -8644 5077 -7678 5157
rect -8644 4937 -8598 5077
rect -8429 4946 -8353 4979
rect -8429 4900 -8418 4946
rect -8364 4900 -8353 4946
rect -8184 4937 -8138 4948
rect -8506 4854 -8460 4865
rect -8598 4680 -8506 4854
rect -8322 4854 -8276 4865
rect -8339 4795 -8322 4805
rect -8276 4795 -8259 4805
rect -8339 4739 -8327 4795
rect -8271 4739 -8259 4795
rect -8339 4729 -8322 4739
rect -8506 4669 -8460 4680
rect -8276 4729 -8259 4739
rect -8322 4669 -8276 4680
rect -8644 4586 -8598 4597
rect -8429 4588 -8418 4634
rect -8364 4588 -8353 4634
rect -7969 4946 -7893 4979
rect -7969 4900 -7958 4946
rect -7904 4900 -7893 4946
rect -7724 4937 -7678 5077
rect -8046 4854 -8000 4865
rect -8063 4795 -8046 4805
rect -7862 4854 -7816 4865
rect -8000 4795 -7983 4805
rect -8063 4739 -8051 4795
rect -7995 4739 -7983 4795
rect -8063 4729 -8046 4739
rect -8000 4729 -7983 4739
rect -8046 4669 -8000 4680
rect -7816 4680 -7724 4854
rect -7862 4669 -7816 4680
rect -9522 4486 -9511 4487
rect -10061 4432 -10059 4478
rect -10013 4432 -10011 4478
rect -9593 4441 -9511 4486
rect -9211 4486 -9200 4487
rect -9211 4441 -9143 4486
rect -9593 4434 -9143 4441
rect -10061 4370 -10011 4432
rect -9585 4426 -9143 4434
rect -9485 4349 -9425 4426
rect -8419 4401 -8363 4588
rect -8184 4586 -8138 4597
rect -7969 4588 -7958 4634
rect -7904 4588 -7893 4634
rect -8201 4537 -8131 4539
rect -7959 4537 -7903 4588
rect -7724 4586 -7678 4597
rect -8201 4481 -8189 4537
rect -8133 4481 -7903 4537
rect -6996 4487 -6916 6097
rect -7122 4486 -7111 4487
rect -8201 4479 -8131 4481
rect -7179 4441 -7111 4486
rect -6811 4486 -6800 4487
rect -6811 4441 -6729 4486
rect -7179 4434 -6729 4441
rect -7179 4426 -6737 4434
rect -8419 4399 -8121 4401
rect -11031 4278 -9891 4300
rect -11031 4232 -10779 4278
rect -10733 4232 -10539 4278
rect -10493 4232 -10299 4278
rect -10253 4232 -10059 4278
rect -10013 4232 -9891 4278
rect -11031 4160 -9891 4232
rect -9485 4202 -9476 4349
rect -9430 4202 -9425 4349
rect -9292 4358 -9246 4360
rect -9292 4349 -9209 4358
rect -9476 3564 -9430 3575
rect -9246 3575 -9209 4349
rect -8419 4343 -8189 4399
rect -8133 4343 -8121 4399
rect -7076 4358 -7030 4360
rect -8419 4341 -8121 4343
rect -7113 4349 -7030 4358
rect -9292 3564 -9209 3575
rect -9399 3502 -9388 3529
rect -9401 3483 -9388 3502
rect -9334 3502 -9323 3529
rect -9334 3483 -9321 3502
rect -10531 3376 -10437 3388
rect -9401 3376 -9321 3483
rect -10531 3300 -10519 3376
rect -10439 3300 -9321 3376
rect -10531 3298 -10437 3300
rect -9401 3193 -9321 3300
rect -9401 3182 -9388 3193
rect -12086 2978 -12006 3179
rect -9399 3147 -9388 3182
rect -9334 3182 -9321 3193
rect -9273 3446 -9209 3564
rect -8644 4117 -8598 4128
rect -8429 4126 -8353 4159
rect -8429 4080 -8418 4126
rect -8364 4080 -8353 4126
rect -8184 4117 -8138 4128
rect -8506 4034 -8460 4045
rect -8598 3860 -8506 4034
rect -8322 4034 -8276 4045
rect -8339 3975 -8322 3985
rect -8276 3975 -8259 3985
rect -8339 3919 -8327 3975
rect -8271 3919 -8259 3975
rect -8339 3909 -8322 3919
rect -8506 3849 -8460 3860
rect -8276 3909 -8259 3919
rect -8322 3849 -8276 3860
rect -8429 3809 -8418 3814
rect -8644 3637 -8598 3777
rect -8431 3799 -8418 3809
rect -8364 3809 -8353 3814
rect -8364 3799 -8351 3809
rect -8431 3743 -8419 3799
rect -8363 3743 -8351 3799
rect -7969 4126 -7893 4159
rect -7969 4080 -7958 4126
rect -7904 4080 -7893 4126
rect -7724 4117 -7678 4128
rect -8046 4034 -8000 4045
rect -8063 3975 -8046 3985
rect -7862 4034 -7816 4045
rect -8000 3975 -7983 3985
rect -8063 3919 -8051 3975
rect -7995 3919 -7983 3975
rect -8063 3909 -8046 3919
rect -8000 3909 -7983 3919
rect -8046 3849 -8000 3860
rect -7816 3860 -7724 4034
rect -7862 3849 -7816 3860
rect -7969 3809 -7958 3814
rect -8184 3766 -8138 3777
rect -7971 3799 -7958 3809
rect -7904 3809 -7893 3814
rect -7904 3799 -7891 3809
rect -8431 3733 -8351 3743
rect -7971 3743 -7959 3799
rect -7903 3743 -7891 3799
rect -7971 3733 -7891 3743
rect -7724 3637 -7678 3777
rect -8644 3557 -7678 3637
rect -7113 3575 -7076 4349
rect -6897 4349 -6837 4426
rect -6897 4202 -6892 4349
rect -7113 3564 -7030 3575
rect -6846 4202 -6837 4349
rect -6892 3564 -6846 3575
rect -9273 3376 -9205 3446
rect -8421 3376 -8349 3378
rect -9273 3300 -8419 3376
rect -8363 3300 -8349 3376
rect -9334 3147 -9323 3182
rect -9273 3112 -9205 3300
rect -8421 3288 -8349 3300
rect -9476 3101 -9430 3112
rect -12103 2961 -11990 2978
rect -12103 2883 -12086 2961
rect -12006 2883 -11990 2961
rect -12103 2872 -11990 2883
rect -9477 2727 -9476 2810
rect -9292 3101 -9205 3112
rect -9430 2727 -9429 2810
rect -9477 2643 -9429 2727
rect -9246 2730 -9205 3101
rect -9292 2716 -9246 2727
rect -11227 2640 -8625 2643
rect -8205 2640 -8139 3557
rect -7113 3446 -7049 3564
rect -6999 3502 -6988 3529
rect -7973 3376 -7901 3378
rect -7117 3376 -7049 3446
rect -7973 3300 -7959 3376
rect -7903 3300 -7049 3376
rect -7973 3288 -7901 3300
rect -7117 3112 -7049 3300
rect -7001 3483 -6988 3502
rect -6934 3502 -6923 3529
rect -6934 3483 -6921 3502
rect -7001 3376 -6921 3483
rect -5895 3376 -5791 3388
rect -7001 3300 -5883 3376
rect -5803 3300 -5791 3376
rect -7001 3193 -6921 3300
rect -5895 3298 -5791 3300
rect -5675 3197 -5597 6097
rect -7001 3182 -6988 3193
rect -6999 3147 -6988 3182
rect -6934 3182 -6921 3193
rect -6934 3147 -6923 3182
rect -7117 3101 -7030 3112
rect -7117 2730 -7076 3101
rect -6892 3101 -6846 3112
rect -7076 2716 -7030 2727
rect -6893 2727 -6892 2810
rect -5676 3027 -5596 3197
rect -5696 2847 -5576 3027
rect -6846 2727 -6845 2810
rect -5696 2787 -5676 2847
rect -5596 2787 -5576 2847
rect -6893 2643 -6845 2727
rect -4791 2649 -4633 2664
rect -4791 2643 -4764 2649
rect -6914 2642 -4764 2643
rect -7131 2640 -4764 2642
rect -11700 2635 -4764 2640
rect -11700 2589 -9511 2635
rect -9211 2589 -7111 2635
rect -6811 2589 -4764 2635
rect -11700 2580 -4764 2589
rect -11700 2551 -11497 2580
rect -11227 2578 -4764 2580
rect -11700 2462 -11642 2551
rect -11551 2462 -11497 2551
rect -4791 2542 -4764 2578
rect -4655 2542 -4633 2649
rect -4791 2531 -4633 2542
rect -11700 2433 -11497 2462
rect -11391 2432 -11287 2446
rect -5035 2432 -4931 2444
rect -11391 2356 -11379 2432
rect -11299 2356 -5023 2432
rect -4943 2356 -4931 2432
rect -11391 2346 -11287 2356
rect -11162 1747 -11116 1758
rect -10947 1756 -10871 2356
rect -10947 1710 -10936 1756
rect -10882 1710 -10871 1756
rect -10702 1747 -10656 1758
rect -11024 1666 -10978 1675
rect -10840 1666 -10794 1675
rect -11116 1664 -10961 1666
rect -11116 1530 -11029 1664
rect -10973 1530 -10961 1664
rect -11116 1528 -10961 1530
rect -10857 1664 -10777 1666
rect -10857 1530 -10845 1664
rect -10789 1530 -10777 1664
rect -10857 1528 -10777 1530
rect -10719 1664 -10702 1666
rect -10302 1747 -10256 1758
rect -10656 1664 -10639 1666
rect -10719 1530 -10707 1664
rect -10651 1530 -10639 1664
rect -10719 1528 -10702 1530
rect -11024 1519 -10978 1528
rect -10840 1519 -10794 1528
rect -11162 1436 -11116 1447
rect -10947 1438 -10936 1484
rect -10882 1438 -10871 1484
rect -10947 1408 -10871 1438
rect -10656 1528 -10639 1530
rect -10702 1436 -10656 1447
rect -10087 1756 -10011 2356
rect -10087 1710 -10076 1756
rect -10022 1710 -10011 1756
rect -9842 1767 -9796 1778
rect -9323 1776 -8823 1832
rect -10164 1666 -10118 1675
rect -9980 1666 -9934 1675
rect -10256 1664 -10101 1666
rect -10256 1530 -10169 1664
rect -10113 1530 -10101 1664
rect -10256 1528 -10101 1530
rect -9997 1664 -9917 1666
rect -9997 1530 -9985 1664
rect -9929 1530 -9917 1664
rect -9997 1528 -9917 1530
rect -9859 1664 -9842 1666
rect -9627 1730 -9616 1776
rect -9442 1730 -9431 1776
rect -9323 1730 -9312 1776
rect -9138 1730 -9127 1776
rect -9019 1730 -9008 1776
rect -8834 1730 -8823 1776
rect -8715 1776 -8215 1832
rect -8715 1730 -8704 1776
rect -8530 1730 -8519 1776
rect -8411 1730 -8400 1776
rect -8226 1730 -8215 1776
rect -8107 1776 -7607 1832
rect -8107 1730 -8096 1776
rect -7922 1730 -7911 1776
rect -7803 1730 -7792 1776
rect -7618 1730 -7607 1776
rect -7499 1776 -6999 1832
rect -7499 1730 -7488 1776
rect -7314 1730 -7303 1776
rect -7195 1730 -7184 1776
rect -7010 1730 -6999 1776
rect -6891 1730 -6880 1776
rect -6706 1730 -6695 1776
rect -6526 1767 -6480 1778
rect -9704 1684 -9658 1695
rect -9796 1664 -9779 1666
rect -9859 1530 -9847 1664
rect -9791 1530 -9779 1664
rect -9859 1528 -9842 1530
rect -10164 1519 -10118 1528
rect -9980 1519 -9934 1528
rect -10302 1436 -10256 1447
rect -10087 1438 -10076 1484
rect -10022 1438 -10011 1484
rect -10087 1408 -10011 1438
rect -9796 1528 -9779 1530
rect -9400 1684 -9354 1695
rect -9417 1677 -9400 1679
rect -9096 1684 -9050 1695
rect -9354 1677 -9337 1679
rect -9417 1533 -9405 1677
rect -9349 1533 -9337 1677
rect -9417 1531 -9400 1533
rect -9704 1499 -9658 1510
rect -9354 1531 -9337 1533
rect -9113 1576 -9096 1586
rect -8792 1684 -8746 1695
rect -8809 1677 -8792 1679
rect -8488 1684 -8442 1695
rect -8746 1677 -8729 1679
rect -9050 1576 -9033 1586
rect -9113 1520 -9101 1576
rect -9045 1520 -9033 1576
rect -8809 1533 -8797 1677
rect -8741 1533 -8729 1677
rect -8809 1531 -8792 1533
rect -9113 1510 -9096 1520
rect -9050 1510 -9033 1520
rect -8746 1531 -8729 1533
rect -8505 1576 -8488 1586
rect -8184 1684 -8138 1695
rect -8201 1677 -8184 1679
rect -7880 1684 -7834 1695
rect -8138 1677 -8121 1679
rect -8442 1576 -8425 1586
rect -8505 1520 -8493 1576
rect -8437 1520 -8425 1576
rect -8201 1533 -8189 1677
rect -8133 1533 -8121 1677
rect -8201 1531 -8184 1533
rect -8505 1510 -8488 1520
rect -8442 1510 -8425 1520
rect -8138 1531 -8121 1533
rect -7897 1576 -7880 1586
rect -7576 1684 -7530 1695
rect -7593 1677 -7576 1679
rect -7272 1684 -7226 1695
rect -7530 1677 -7513 1679
rect -7834 1576 -7817 1586
rect -7897 1520 -7885 1576
rect -7829 1520 -7817 1576
rect -7593 1533 -7581 1677
rect -7525 1533 -7513 1677
rect -7593 1531 -7576 1533
rect -7897 1510 -7880 1520
rect -7834 1510 -7817 1520
rect -7530 1531 -7513 1533
rect -7289 1576 -7272 1586
rect -6968 1684 -6922 1695
rect -6985 1677 -6968 1679
rect -6664 1684 -6618 1695
rect -6922 1677 -6905 1679
rect -7226 1576 -7209 1586
rect -7289 1520 -7277 1576
rect -7221 1520 -7209 1576
rect -6985 1533 -6973 1677
rect -6917 1533 -6905 1677
rect -6985 1531 -6968 1533
rect -7289 1510 -7272 1520
rect -7226 1510 -7209 1520
rect -6922 1531 -6905 1533
rect -9400 1499 -9354 1510
rect -9096 1499 -9050 1510
rect -8792 1499 -8746 1510
rect -8488 1499 -8442 1510
rect -8184 1499 -8138 1510
rect -7880 1499 -7834 1510
rect -7576 1499 -7530 1510
rect -7272 1499 -7226 1510
rect -6968 1499 -6922 1510
rect -6543 1664 -6526 1666
rect -6311 1756 -6235 2356
rect -6311 1710 -6300 1756
rect -6246 1710 -6235 1756
rect -6066 1747 -6020 1758
rect -6388 1666 -6342 1675
rect -6204 1666 -6158 1675
rect -6480 1664 -6463 1666
rect -6543 1530 -6531 1664
rect -6475 1530 -6463 1664
rect -6543 1528 -6526 1530
rect -6664 1499 -6618 1510
rect -8310 1469 -8230 1479
rect -8310 1464 -8298 1469
rect -8242 1464 -8230 1469
rect -8092 1469 -8012 1479
rect -8092 1464 -8080 1469
rect -8024 1464 -8012 1469
rect -9842 1416 -9796 1427
rect -9627 1418 -9616 1464
rect -9442 1418 -9431 1464
rect -9323 1418 -9312 1464
rect -9138 1453 -9127 1464
rect -9019 1453 -9008 1464
rect -9138 1418 -9008 1453
rect -8834 1418 -8823 1464
rect -8715 1418 -8704 1464
rect -8530 1418 -8519 1464
rect -8411 1418 -8400 1464
rect -8226 1418 -8215 1464
rect -8107 1418 -8096 1464
rect -7922 1418 -7911 1464
rect -7803 1418 -7792 1464
rect -7618 1418 -7607 1464
rect -7499 1418 -7488 1464
rect -7314 1453 -7303 1464
rect -7195 1453 -7184 1464
rect -7314 1418 -7184 1453
rect -7010 1418 -6999 1464
rect -6891 1418 -6880 1464
rect -6706 1418 -6695 1464
rect -6480 1528 -6463 1530
rect -6405 1664 -6325 1666
rect -6405 1530 -6393 1664
rect -6337 1530 -6325 1664
rect -6405 1528 -6325 1530
rect -6221 1664 -6066 1666
rect -6221 1530 -6209 1664
rect -6153 1530 -6066 1664
rect -6221 1528 -6066 1530
rect -6388 1519 -6342 1528
rect -6204 1519 -6158 1528
rect -9263 1407 -8823 1418
rect -8310 1413 -8298 1418
rect -8242 1413 -8230 1418
rect -10531 1161 -10427 1173
rect -10009 1161 -9905 1171
rect -9263 1161 -9159 1407
rect -8310 1403 -8230 1413
rect -8092 1413 -8080 1418
rect -8024 1413 -8012 1418
rect -8092 1403 -8012 1413
rect -7499 1407 -7059 1418
rect -6526 1416 -6480 1427
rect -6311 1438 -6300 1484
rect -6246 1438 -6235 1484
rect -6311 1408 -6235 1438
rect -5666 1747 -5620 1758
rect -5683 1664 -5666 1666
rect -5451 1756 -5375 2356
rect -5035 2344 -4931 2356
rect -5451 1710 -5440 1756
rect -5386 1710 -5375 1756
rect -5206 1747 -5160 1758
rect -5528 1666 -5482 1675
rect -5344 1666 -5298 1675
rect -5620 1664 -5603 1666
rect -5683 1530 -5671 1664
rect -5615 1530 -5603 1664
rect -5683 1528 -5666 1530
rect -6066 1436 -6020 1447
rect -5620 1528 -5603 1530
rect -5545 1664 -5465 1666
rect -5545 1530 -5533 1664
rect -5477 1530 -5465 1664
rect -5545 1528 -5465 1530
rect -5361 1664 -5206 1666
rect -5361 1530 -5349 1664
rect -5293 1530 -5206 1664
rect -5361 1528 -5206 1530
rect -5528 1519 -5482 1528
rect -5344 1519 -5298 1528
rect -5666 1436 -5620 1447
rect -5451 1438 -5440 1484
rect -5386 1438 -5375 1484
rect -5451 1408 -5375 1438
rect -5206 1436 -5160 1447
rect -8655 1161 -8415 1169
rect -10531 1077 -10519 1161
rect -10439 1077 -9997 1161
rect -9917 1159 -8415 1161
rect -9917 1079 -9251 1159
rect -9171 1079 -8643 1159
rect -8563 1079 -8505 1159
rect -8425 1079 -8415 1159
rect -9917 1077 -8415 1079
rect -10531 1067 -10427 1077
rect -10009 1067 -9905 1077
rect -9263 1065 -9159 1077
rect -8655 1065 -8415 1077
rect -7909 1161 -7667 1169
rect -7163 1161 -7059 1407
rect -6417 1161 -6313 1171
rect -5895 1161 -5791 1171
rect -7909 1159 -6405 1161
rect -7909 1079 -7897 1159
rect -7817 1079 -7759 1159
rect -7679 1079 -7151 1159
rect -7071 1079 -6405 1159
rect -7909 1077 -6405 1079
rect -6325 1077 -5883 1161
rect -5803 1077 -5791 1161
rect -7909 1065 -7667 1077
rect -7163 1066 -7059 1077
rect -6417 1067 -6313 1077
rect -5895 1067 -5791 1077
rect -9461 865 -8657 880
rect -9980 811 -9934 822
rect -9461 820 -8842 865
rect -8762 820 -8657 865
rect -7665 865 -6861 880
rect -9997 415 -9980 425
rect -9765 774 -9754 820
rect -9580 774 -9569 820
rect -9461 774 -9450 820
rect -9276 774 -9265 820
rect -9157 774 -9146 820
rect -8972 774 -8961 820
rect -8853 774 -8842 820
rect -8668 774 -8657 820
rect -8549 774 -8538 820
rect -8364 774 -8353 820
rect -8184 811 -8138 822
rect -7665 820 -7560 865
rect -7480 820 -6861 865
rect -9842 728 -9796 739
rect -9934 415 -9917 425
rect -9997 271 -9985 415
rect -9929 271 -9917 415
rect -9538 728 -9492 739
rect -9555 505 -9538 507
rect -9234 728 -9188 739
rect -9251 721 -9234 723
rect -8930 728 -8884 739
rect -9188 721 -9171 723
rect -9251 577 -9239 721
rect -9183 577 -9171 721
rect -9251 575 -9234 577
rect -9492 505 -9475 507
rect -9555 361 -9543 505
rect -9487 361 -9475 505
rect -9555 359 -9538 361
rect -9842 343 -9796 354
rect -9492 359 -9475 361
rect -9538 343 -9492 354
rect -9188 575 -9171 577
rect -8947 505 -8930 507
rect -8626 728 -8580 739
rect -8643 721 -8626 723
rect -8322 728 -8276 739
rect -8580 721 -8563 723
rect -8643 577 -8631 721
rect -8575 577 -8563 721
rect -8643 575 -8626 577
rect -8884 505 -8867 507
rect -8947 361 -8935 505
rect -8879 361 -8867 505
rect -8947 359 -8930 361
rect -9234 343 -9188 354
rect -8884 359 -8867 361
rect -8930 343 -8884 354
rect -8580 575 -8563 577
rect -8626 343 -8580 354
rect -8322 343 -8276 354
rect -9997 260 -9917 271
rect -9765 262 -9754 308
rect -9580 262 -9569 308
rect -9461 262 -9450 308
rect -9276 262 -9265 308
rect -9157 262 -9146 308
rect -8972 262 -8961 308
rect -8853 262 -8842 308
rect -8668 262 -8657 308
rect -8549 262 -8538 308
rect -8364 262 -8353 308
rect -7969 774 -7958 820
rect -7784 774 -7773 820
rect -7665 774 -7654 820
rect -7480 774 -7469 820
rect -7361 774 -7350 820
rect -7176 774 -7165 820
rect -7057 774 -7046 820
rect -6872 774 -6861 820
rect -6753 774 -6742 820
rect -6568 774 -6557 820
rect -6388 811 -6342 822
rect -8046 728 -8000 739
rect -7742 728 -7696 739
rect -7759 721 -7742 723
rect -7438 728 -7392 739
rect -7696 721 -7679 723
rect -7759 577 -7747 721
rect -7691 577 -7679 721
rect -7759 575 -7742 577
rect -8046 343 -8000 354
rect -7696 575 -7679 577
rect -7455 505 -7438 507
rect -7134 728 -7088 739
rect -7151 721 -7134 723
rect -6830 728 -6784 739
rect -7088 721 -7071 723
rect -7151 577 -7139 721
rect -7083 577 -7071 721
rect -7151 575 -7134 577
rect -7392 505 -7375 507
rect -7455 361 -7443 505
rect -7387 361 -7375 505
rect -7455 359 -7438 361
rect -7742 343 -7696 354
rect -7392 359 -7375 361
rect -7438 343 -7392 354
rect -7088 575 -7071 577
rect -6847 505 -6830 507
rect -6526 728 -6480 739
rect -6784 505 -6767 507
rect -6847 361 -6835 505
rect -6779 361 -6767 505
rect -6847 359 -6830 361
rect -7134 343 -7088 354
rect -6784 359 -6767 361
rect -6830 343 -6784 354
rect -6526 343 -6480 354
rect -6405 415 -6388 425
rect -6342 415 -6325 425
rect -8184 260 -8138 271
rect -7969 262 -7958 308
rect -7784 262 -7773 308
rect -7665 262 -7654 308
rect -7480 262 -7469 308
rect -7361 262 -7350 308
rect -7176 262 -7165 308
rect -7057 262 -7046 308
rect -6872 262 -6861 308
rect -6753 262 -6742 308
rect -6568 262 -6557 308
rect -6405 271 -6393 415
rect -6337 271 -6325 415
rect -6405 260 -6325 271
rect -10869 -5 -10765 5
rect -9733 -5 -9629 7
rect -9567 -5 -9463 7
rect -8959 -5 -8855 7
rect -10869 -85 -10857 -5
rect -10777 -85 -9721 -5
rect -9641 -85 -9555 -5
rect -9475 -85 -8947 -5
rect -8867 -85 -8855 -5
rect -10869 -95 -10765 -85
rect -9733 -97 -9629 -85
rect -9567 -97 -9463 -85
rect -8959 -97 -8855 -85
rect -7467 -5 -7363 7
rect -6859 -5 -6755 7
rect -6693 -5 -6589 7
rect -5557 -5 -5453 5
rect -7467 -85 -7455 -5
rect -7375 -85 -6847 -5
rect -6767 -85 -6681 -5
rect -6601 -85 -5545 -5
rect -5465 -85 -5453 -5
rect -7467 -97 -7363 -85
rect -6859 -97 -6755 -85
rect -6693 -97 -6589 -85
rect -5557 -95 -5453 -85
rect -10315 -403 -10193 -392
rect -10315 -903 -10304 -403
rect -10204 -903 -10193 -403
rect -6129 -403 -6007 -392
rect -9931 -711 -9920 -665
rect -9746 -711 -9735 -665
rect -9627 -711 -9616 -665
rect -9442 -711 -9431 -665
rect -9323 -711 -9312 -665
rect -9138 -711 -9127 -665
rect -9019 -711 -9008 -665
rect -8834 -711 -8823 -665
rect -8715 -711 -8704 -665
rect -8530 -711 -8519 -665
rect -8411 -711 -8400 -665
rect -8226 -711 -8215 -665
rect -8107 -711 -8096 -665
rect -7922 -711 -7911 -665
rect -7803 -711 -7792 -665
rect -7618 -711 -7607 -665
rect -7499 -711 -7488 -665
rect -7314 -711 -7303 -665
rect -7195 -711 -7184 -665
rect -7010 -711 -6999 -665
rect -6891 -711 -6880 -665
rect -6706 -711 -6695 -665
rect -6587 -711 -6576 -665
rect -6402 -711 -6391 -665
rect -10315 -914 -10193 -903
rect -10008 -757 -9962 -746
rect -9704 -757 -9658 -746
rect -9721 -813 -9704 -803
rect -9400 -757 -9354 -746
rect -9658 -813 -9641 -803
rect -9721 -974 -9709 -813
rect -9653 -974 -9641 -813
rect -9721 -984 -9704 -974
rect -10008 -1042 -9962 -1031
rect -9658 -984 -9641 -974
rect -9417 -861 -9400 -851
rect -9096 -757 -9050 -746
rect -9113 -777 -9096 -767
rect -8792 -757 -8746 -746
rect -9050 -777 -9033 -767
rect -9354 -861 -9337 -851
rect -9704 -1042 -9658 -1031
rect -9417 -1022 -9405 -861
rect -9349 -1022 -9337 -861
rect -9113 -994 -9101 -777
rect -9045 -994 -9033 -777
rect -9113 -1002 -9096 -994
rect -9417 -1031 -9400 -1022
rect -9354 -1031 -9337 -1022
rect -9417 -1032 -9337 -1031
rect -9050 -1002 -9033 -994
rect -8809 -861 -8792 -851
rect -8488 -757 -8442 -746
rect -8505 -777 -8488 -767
rect -8184 -757 -8138 -746
rect -8442 -777 -8425 -767
rect -8505 -833 -8493 -777
rect -8437 -833 -8425 -777
rect -8505 -843 -8488 -833
rect -8746 -861 -8729 -851
rect -9400 -1042 -9354 -1032
rect -9096 -1042 -9050 -1031
rect -8809 -1022 -8797 -861
rect -8741 -1022 -8729 -861
rect -8809 -1031 -8792 -1022
rect -8746 -1031 -8729 -1022
rect -8809 -1032 -8729 -1031
rect -8442 -843 -8425 -833
rect -8792 -1042 -8746 -1032
rect -8488 -1042 -8442 -1031
rect -8201 -861 -8184 -851
rect -7880 -757 -7834 -746
rect -7897 -777 -7880 -767
rect -7576 -757 -7530 -746
rect -7834 -777 -7817 -767
rect -7897 -833 -7885 -777
rect -7829 -833 -7817 -777
rect -7897 -843 -7880 -833
rect -8138 -861 -8121 -851
rect -8201 -1022 -8189 -861
rect -8133 -1022 -8121 -861
rect -8201 -1031 -8184 -1022
rect -8138 -1031 -8121 -1022
rect -8201 -1032 -8121 -1031
rect -7834 -843 -7817 -833
rect -8184 -1042 -8138 -1032
rect -7880 -1042 -7834 -1031
rect -7593 -861 -7576 -851
rect -7272 -757 -7226 -746
rect -7289 -777 -7272 -767
rect -6968 -757 -6922 -746
rect -7226 -777 -7209 -767
rect -7530 -861 -7513 -851
rect -7593 -1022 -7581 -861
rect -7525 -1022 -7513 -861
rect -7593 -1031 -7576 -1022
rect -7530 -1031 -7513 -1022
rect -7593 -1032 -7513 -1031
rect -7289 -1022 -7277 -777
rect -7221 -1022 -7209 -777
rect -7289 -1031 -7272 -1022
rect -7226 -1031 -7209 -1022
rect -7289 -1032 -7209 -1031
rect -6985 -861 -6968 -851
rect -6664 -757 -6618 -746
rect -6681 -813 -6664 -803
rect -6360 -757 -6314 -746
rect -6618 -813 -6601 -803
rect -6922 -861 -6905 -851
rect -6985 -1022 -6973 -861
rect -6917 -1022 -6905 -861
rect -6681 -974 -6669 -813
rect -6613 -974 -6601 -813
rect -6681 -984 -6664 -974
rect -6985 -1031 -6968 -1022
rect -6922 -1031 -6905 -1022
rect -6985 -1032 -6905 -1031
rect -6618 -984 -6601 -974
rect -7576 -1042 -7530 -1032
rect -7272 -1042 -7226 -1032
rect -6968 -1042 -6922 -1032
rect -6664 -1042 -6618 -1031
rect -6129 -903 -6118 -403
rect -6018 -903 -6007 -403
rect -6129 -914 -6007 -903
rect -6360 -1042 -6314 -1031
rect -9276 -1077 -9261 -1068
rect -9191 -1077 -9176 -1068
rect -8971 -1077 -8956 -1068
rect -8886 -1077 -8871 -1068
rect -8061 -1077 -8046 -1068
rect -7976 -1077 -7961 -1068
rect -7756 -1077 -7741 -1068
rect -7671 -1077 -7656 -1068
rect -6841 -1077 -6826 -1068
rect -6756 -1077 -6741 -1068
rect -9931 -1123 -9920 -1077
rect -9746 -1123 -9735 -1077
rect -9627 -1123 -9616 -1077
rect -9442 -1123 -9431 -1077
rect -9323 -1123 -9312 -1077
rect -9138 -1123 -9127 -1077
rect -9019 -1123 -9008 -1077
rect -8834 -1123 -8823 -1077
rect -8715 -1123 -8704 -1077
rect -8530 -1123 -8519 -1077
rect -8411 -1123 -8400 -1077
rect -8226 -1123 -8215 -1077
rect -8107 -1123 -8096 -1077
rect -7922 -1123 -7911 -1077
rect -7803 -1123 -7792 -1077
rect -7618 -1123 -7607 -1077
rect -7499 -1123 -7488 -1077
rect -7314 -1123 -7303 -1077
rect -7195 -1123 -7184 -1077
rect -7010 -1123 -6999 -1077
rect -6891 -1123 -6880 -1077
rect -6706 -1123 -6695 -1077
rect -6587 -1123 -6576 -1077
rect -6402 -1123 -6391 -1077
rect -13722 -1178 -13632 -1166
rect -9626 -1178 -9431 -1123
rect -9321 -1128 -9261 -1123
rect -9191 -1128 -9136 -1123
rect -8971 -1128 -8956 -1123
rect -8886 -1128 -8871 -1123
rect -8716 -1178 -8521 -1123
rect -8411 -1178 -8216 -1123
rect -8061 -1128 -8046 -1123
rect -7976 -1128 -7961 -1123
rect -7756 -1128 -7741 -1123
rect -7671 -1128 -7656 -1123
rect -7496 -1178 -7301 -1123
rect -7196 -1178 -7001 -1123
rect -6841 -1128 -6826 -1123
rect -6756 -1128 -6741 -1123
rect -13722 -1179 -6031 -1178
rect -13722 -1252 -13707 -1179
rect -13634 -1193 -6031 -1179
rect -13634 -1226 -6511 -1193
rect -13634 -1252 -9254 -1226
rect -13722 -1253 -9254 -1252
rect -13722 -1266 -13632 -1253
rect -9266 -1282 -9254 -1253
rect -9198 -1253 -8039 -1226
rect -9198 -1282 -9186 -1253
rect -9266 -1292 -9186 -1282
rect -8051 -1282 -8039 -1253
rect -7983 -1253 -6511 -1226
rect -6451 -1253 -6031 -1193
rect -7983 -1282 -7971 -1253
rect -8051 -1292 -7971 -1282
rect -8961 -1474 -8881 -1464
rect -13717 -1503 -13627 -1491
rect -8961 -1503 -8949 -1474
rect -13717 -1504 -8949 -1503
rect -13717 -1577 -13704 -1504
rect -13631 -1530 -8949 -1504
rect -8893 -1503 -8881 -1474
rect -7746 -1474 -7666 -1464
rect -7746 -1503 -7734 -1474
rect -8893 -1530 -7734 -1503
rect -7678 -1503 -7666 -1474
rect -7678 -1530 -6251 -1503
rect -13631 -1563 -6251 -1530
rect -6191 -1563 -6031 -1503
rect -13631 -1577 -6031 -1563
rect -13717 -1578 -6031 -1577
rect -13717 -1591 -13627 -1578
rect -9626 -1628 -9431 -1578
rect -8716 -1628 -8521 -1578
rect -8411 -1628 -8216 -1578
rect -7501 -1628 -7306 -1578
rect -7196 -1628 -7001 -1578
rect -9931 -1674 -9920 -1628
rect -9746 -1674 -9735 -1628
rect -9627 -1674 -9616 -1628
rect -9442 -1674 -9431 -1628
rect -9323 -1674 -9312 -1628
rect -9138 -1674 -9127 -1628
rect -9019 -1674 -9008 -1628
rect -8834 -1674 -8823 -1628
rect -8715 -1674 -8704 -1628
rect -8530 -1674 -8519 -1628
rect -8411 -1674 -8400 -1628
rect -8226 -1674 -8215 -1628
rect -8107 -1674 -8096 -1628
rect -7922 -1674 -7911 -1628
rect -7803 -1674 -7792 -1628
rect -7618 -1674 -7607 -1628
rect -7499 -1674 -7488 -1628
rect -7314 -1674 -7303 -1628
rect -7195 -1674 -7184 -1628
rect -7010 -1674 -6999 -1628
rect -6891 -1674 -6880 -1628
rect -6706 -1674 -6695 -1628
rect -6587 -1674 -6576 -1628
rect -6402 -1674 -6391 -1628
rect -9276 -1688 -9261 -1674
rect -9191 -1688 -9176 -1674
rect -8971 -1688 -8956 -1674
rect -8886 -1688 -8871 -1674
rect -8061 -1688 -8046 -1674
rect -7976 -1688 -7961 -1674
rect -7756 -1688 -7741 -1674
rect -7671 -1688 -7656 -1674
rect -6841 -1688 -6826 -1674
rect -6756 -1688 -6741 -1674
rect -10008 -1720 -9962 -1709
rect -10315 -1848 -10193 -1837
rect -10315 -2348 -10304 -1848
rect -10204 -2348 -10193 -1848
rect -9704 -1720 -9658 -1709
rect -9721 -1921 -9704 -1911
rect -9400 -1720 -9354 -1709
rect -9417 -1732 -9400 -1722
rect -9096 -1720 -9050 -1709
rect -9354 -1732 -9337 -1722
rect -9417 -1893 -9405 -1732
rect -9349 -1893 -9337 -1732
rect -9417 -1903 -9400 -1893
rect -9658 -1921 -9641 -1911
rect -9721 -1977 -9709 -1921
rect -9653 -1977 -9641 -1921
rect -9721 -1987 -9704 -1977
rect -10008 -2005 -9962 -1994
rect -9658 -1987 -9641 -1977
rect -9704 -2005 -9658 -1994
rect -9354 -1903 -9337 -1893
rect -9113 -1766 -9096 -1756
rect -8792 -1720 -8746 -1709
rect -8809 -1732 -8792 -1722
rect -8488 -1720 -8442 -1709
rect -8746 -1732 -8729 -1722
rect -9050 -1766 -9033 -1756
rect -9113 -1977 -9101 -1766
rect -9045 -1977 -9033 -1766
rect -8809 -1893 -8797 -1732
rect -8741 -1893 -8729 -1732
rect -8809 -1903 -8792 -1893
rect -9113 -1987 -9096 -1977
rect -9400 -2005 -9354 -1994
rect -9050 -1987 -9033 -1977
rect -9096 -2005 -9050 -1994
rect -8746 -1903 -8729 -1893
rect -8505 -1732 -8488 -1722
rect -8184 -1720 -8138 -1709
rect -8442 -1732 -8425 -1722
rect -8505 -1977 -8493 -1732
rect -8437 -1977 -8425 -1732
rect -8201 -1732 -8184 -1722
rect -7880 -1720 -7834 -1709
rect -8138 -1732 -8121 -1722
rect -8201 -1893 -8189 -1732
rect -8133 -1893 -8121 -1732
rect -8201 -1903 -8184 -1893
rect -8505 -1987 -8488 -1977
rect -8792 -2005 -8746 -1994
rect -8442 -1987 -8425 -1977
rect -8488 -2005 -8442 -1994
rect -8138 -1903 -8121 -1893
rect -7897 -1766 -7880 -1756
rect -7576 -1720 -7530 -1709
rect -7593 -1732 -7576 -1722
rect -7272 -1720 -7226 -1709
rect -7530 -1732 -7513 -1722
rect -7834 -1766 -7817 -1756
rect -7897 -1977 -7885 -1766
rect -7829 -1977 -7817 -1766
rect -7593 -1893 -7581 -1732
rect -7525 -1893 -7513 -1732
rect -7593 -1903 -7576 -1893
rect -7897 -1987 -7880 -1977
rect -8184 -2005 -8138 -1994
rect -7834 -1987 -7817 -1977
rect -7880 -2005 -7834 -1994
rect -7530 -1903 -7513 -1893
rect -7289 -1732 -7272 -1722
rect -6968 -1720 -6922 -1709
rect -7226 -1732 -7209 -1722
rect -7289 -1977 -7277 -1732
rect -7221 -1977 -7209 -1732
rect -7289 -1987 -7272 -1977
rect -7576 -2005 -7530 -1994
rect -7226 -1987 -7209 -1977
rect -6985 -1732 -6968 -1722
rect -6664 -1720 -6618 -1709
rect -6922 -1732 -6905 -1722
rect -6985 -1977 -6973 -1732
rect -6917 -1977 -6905 -1732
rect -6985 -1987 -6968 -1977
rect -7272 -2005 -7226 -1994
rect -6922 -1987 -6905 -1977
rect -6681 -1920 -6664 -1910
rect -6360 -1720 -6314 -1709
rect -6618 -1920 -6601 -1910
rect -6681 -1977 -6669 -1920
rect -6613 -1977 -6601 -1920
rect -6681 -1987 -6664 -1977
rect -6968 -2005 -6922 -1994
rect -6618 -1987 -6601 -1977
rect -6664 -2005 -6618 -1994
rect -6360 -2005 -6314 -1994
rect -6129 -1848 -6007 -1837
rect -9931 -2086 -9920 -2040
rect -9746 -2086 -9735 -2040
rect -9627 -2086 -9616 -2040
rect -9442 -2086 -9431 -2040
rect -9323 -2086 -9312 -2040
rect -9138 -2086 -9127 -2040
rect -9019 -2086 -9008 -2040
rect -8834 -2086 -8823 -2040
rect -8715 -2086 -8704 -2040
rect -8530 -2086 -8519 -2040
rect -8411 -2086 -8400 -2040
rect -8226 -2086 -8215 -2040
rect -8107 -2086 -8096 -2040
rect -7922 -2086 -7911 -2040
rect -7803 -2086 -7792 -2040
rect -7618 -2086 -7607 -2040
rect -7499 -2086 -7488 -2040
rect -7314 -2086 -7303 -2040
rect -7195 -2086 -7184 -2040
rect -7010 -2086 -6999 -2040
rect -6891 -2086 -6880 -2040
rect -6706 -2086 -6695 -2040
rect -6587 -2086 -6576 -2040
rect -6402 -2086 -6391 -2040
rect -6129 -2144 -6118 -1848
rect -6143 -2160 -6118 -2144
rect -6018 -2144 -6007 -1848
rect -6143 -2297 -6129 -2160
rect -10315 -2359 -10193 -2348
rect -6144 -2370 -6129 -2297
rect -6018 -2308 -6002 -2144
rect -6018 -2348 -6007 -2308
rect -6024 -2370 -6007 -2348
rect -6144 -2388 -6007 -2370
rect -8598 -2563 -8552 -2552
rect -8615 -2652 -8598 -2650
rect -8383 -2554 -8307 -2524
rect -8383 -2600 -8372 -2554
rect -8318 -2600 -8307 -2554
rect -8199 -2554 -8123 -2524
rect -8199 -2600 -8188 -2554
rect -8134 -2600 -8123 -2554
rect -8015 -2554 -7939 -2524
rect -8015 -2600 -8004 -2554
rect -7950 -2600 -7939 -2554
rect -7770 -2563 -7724 -2552
rect -8460 -2646 -8414 -2635
rect -8552 -2652 -8535 -2650
rect -8615 -2774 -8603 -2652
rect -8547 -2774 -8535 -2652
rect -8615 -2776 -8598 -2774
rect -8552 -2776 -8535 -2774
rect -8276 -2646 -8230 -2635
rect -8293 -2652 -8276 -2650
rect -8092 -2646 -8046 -2635
rect -8230 -2652 -8213 -2650
rect -8293 -2774 -8281 -2652
rect -8225 -2774 -8213 -2652
rect -8293 -2776 -8276 -2774
rect -8460 -2791 -8414 -2780
rect -8230 -2776 -8213 -2774
rect -8109 -2652 -8092 -2650
rect -7908 -2646 -7862 -2635
rect -8046 -2652 -8029 -2650
rect -8109 -2774 -8097 -2652
rect -8041 -2774 -8029 -2652
rect -8109 -2776 -8092 -2774
rect -8276 -2791 -8230 -2780
rect -8046 -2776 -8029 -2774
rect -8092 -2791 -8046 -2780
rect -7908 -2791 -7862 -2780
rect -8598 -2874 -8552 -2863
rect -8383 -2872 -8372 -2826
rect -8318 -2872 -8307 -2826
rect -8383 -2902 -8307 -2872
rect -8199 -2872 -8188 -2826
rect -8134 -2872 -8123 -2826
rect -13382 -3003 -13286 -3000
rect -11391 -3003 -11287 -2993
rect -8199 -3003 -8123 -2872
rect -8015 -2872 -8004 -2826
rect -7950 -2872 -7939 -2826
rect -8015 -2902 -7939 -2872
rect -7770 -2874 -7724 -2863
rect -5035 -3003 -4931 -2993
rect -13382 -3004 -11379 -3003
rect -13382 -3082 -13368 -3004
rect -13290 -3082 -11379 -3004
rect -13382 -3083 -11379 -3082
rect -11299 -3083 -5023 -3003
rect -4943 -3083 -4931 -3003
rect -13382 -3096 -13286 -3083
rect -11391 -3093 -11287 -3083
rect -5035 -3093 -4931 -3083
rect -13302 -3363 -2407 -3321
rect -13302 -3375 -4454 -3363
rect -13302 -3376 -6132 -3375
rect -13302 -3443 -10639 -3376
rect -13302 -3530 -11640 -3443
rect -11555 -3463 -10639 -3443
rect -10550 -3381 -6132 -3376
rect -10550 -3463 -10083 -3381
rect -11555 -3530 -10083 -3463
rect -13302 -3592 -10083 -3530
rect -9728 -3578 -6132 -3381
rect -6018 -3429 -4454 -3375
rect -6018 -3531 -5654 -3429
rect -5550 -3451 -4454 -3429
rect -5550 -3531 -4764 -3451
rect -6018 -3558 -4764 -3531
rect -4655 -3558 -4454 -3451
rect -6018 -3578 -4454 -3558
rect -9728 -3592 -4454 -3578
rect -13302 -3663 -4454 -3592
rect -2454 -3663 -2407 -3363
rect -13302 -3701 -2407 -3663
<< via1 >>
rect 40739 39093 40957 39167
rect 40135 38547 40187 38599
rect 40695 38336 40747 38339
rect 40695 38290 40698 38336
rect 40698 38290 40744 38336
rect 40744 38290 40747 38336
rect 40695 38287 40747 38290
rect 40737 37749 40955 37823
rect -4343 37511 -4287 37567
rect -4711 37124 -4706 37244
rect -4706 37124 -4660 37244
rect -4660 37124 -4655 37244
rect -4343 37124 -4338 37244
rect -4338 37124 -4292 37244
rect -4292 37124 -4287 37244
rect -4527 36824 -4522 36944
rect -4522 36824 -4476 36944
rect -4476 36824 -4471 36944
rect -4021 37123 -4016 37244
rect -4016 37123 -3970 37244
rect -3970 37123 -3965 37244
rect -4159 36824 -4154 36944
rect -4154 36824 -4108 36944
rect -4108 36824 -4103 36944
rect -4619 36705 -4618 36748
rect -4618 36705 -4564 36748
rect -4564 36705 -4563 36748
rect -4619 36692 -4563 36705
rect -4435 36705 -4434 36748
rect -4434 36705 -4380 36748
rect -4380 36705 -4379 36748
rect -4435 36692 -4379 36705
rect -4251 36705 -4250 36748
rect -4250 36705 -4196 36748
rect -4196 36705 -4195 36748
rect -4251 36692 -4195 36705
rect -5507 36542 -5451 36598
rect -4619 36542 -4563 36598
rect -5291 36426 -5235 36482
rect -4435 36426 -4379 36482
rect -4106 36426 -4050 36482
rect -3849 36426 -3793 36482
rect -4251 36310 -4195 36366
rect -4619 36203 -4563 36216
rect -4619 36160 -4618 36203
rect -4618 36160 -4564 36203
rect -4564 36160 -4563 36203
rect -4435 36203 -4379 36216
rect -4435 36160 -4434 36203
rect -4434 36160 -4380 36203
rect -4380 36160 -4379 36203
rect -4251 36203 -4195 36216
rect -4251 36160 -4250 36203
rect -4250 36160 -4196 36203
rect -4196 36160 -4195 36203
rect -4159 35964 -4154 36084
rect -4154 35964 -4108 36084
rect -4108 35964 -4103 36084
rect -4844 35641 -4788 35697
rect -4026 35641 -3970 35697
rect -3673 35523 -3617 35579
rect -3849 35415 -3793 35469
rect -4343 35306 -4287 35362
rect -4711 34919 -4706 35039
rect -4706 34919 -4660 35039
rect -4660 34919 -4655 35039
rect -4343 34919 -4338 35039
rect -4338 34919 -4292 35039
rect -4292 34919 -4287 35039
rect -4527 34619 -4522 34739
rect -4522 34619 -4476 34739
rect -4476 34619 -4471 34739
rect -4021 34918 -4016 35039
rect -4016 34918 -3970 35039
rect -3970 34918 -3965 35039
rect -4159 34619 -4154 34739
rect -4154 34619 -4108 34739
rect -4108 34619 -4103 34739
rect -4619 34500 -4618 34543
rect -4618 34500 -4564 34543
rect -4564 34500 -4563 34543
rect -4619 34487 -4563 34500
rect -4435 34500 -4434 34543
rect -4434 34500 -4380 34543
rect -4380 34500 -4379 34543
rect -4435 34487 -4379 34500
rect -4251 34500 -4250 34543
rect -4250 34500 -4196 34543
rect -4196 34500 -4195 34543
rect -4251 34487 -4195 34500
rect -4619 34337 -4563 34393
rect 5129 37511 5185 37567
rect 4761 37124 4766 37244
rect 4766 37124 4812 37244
rect 4812 37124 4817 37244
rect 5129 37124 5134 37244
rect 5134 37124 5180 37244
rect 5180 37124 5185 37244
rect 4945 36824 4950 36944
rect 4950 36824 4996 36944
rect 4996 36824 5001 36944
rect 5451 37123 5456 37244
rect 5456 37123 5502 37244
rect 5502 37123 5507 37244
rect 5313 36824 5318 36944
rect 5318 36824 5364 36944
rect 5364 36824 5369 36944
rect 4853 36705 4854 36748
rect 4854 36705 4908 36748
rect 4908 36705 4909 36748
rect 4853 36692 4909 36705
rect 5037 36705 5038 36748
rect 5038 36705 5092 36748
rect 5092 36705 5093 36748
rect 5037 36692 5093 36705
rect 5221 36705 5222 36748
rect 5222 36705 5276 36748
rect 5276 36705 5277 36748
rect 5221 36692 5277 36705
rect 3965 36542 4021 36598
rect 4853 36542 4909 36598
rect 4181 36426 4237 36482
rect 5037 36426 5093 36482
rect 5366 36426 5422 36482
rect 5623 36426 5679 36482
rect 5221 36310 5277 36366
rect 4853 36203 4909 36216
rect 4853 36160 4854 36203
rect 4854 36160 4908 36203
rect 4908 36160 4909 36203
rect 5037 36203 5093 36216
rect 5037 36160 5038 36203
rect 5038 36160 5092 36203
rect 5092 36160 5093 36203
rect 5221 36203 5277 36216
rect 5221 36160 5222 36203
rect 5222 36160 5276 36203
rect 5276 36160 5277 36203
rect 5313 35964 5318 36084
rect 5318 35964 5364 36084
rect 5364 35964 5369 36084
rect 4628 35641 4684 35697
rect 5446 35641 5502 35697
rect 5799 35523 5855 35579
rect 5623 35415 5679 35469
rect -2857 35306 -2801 35362
rect -3225 34919 -3220 35039
rect -3220 34919 -3174 35039
rect -3174 34919 -3169 35039
rect -2857 34919 -2852 35039
rect -2852 34919 -2806 35039
rect -2806 34919 -2801 35039
rect -3041 34619 -3036 34739
rect -3036 34619 -2990 34739
rect -2990 34619 -2985 34739
rect -2535 34918 -2530 35039
rect -2530 34918 -2484 35039
rect -2484 34918 -2479 35039
rect -2673 34619 -2668 34739
rect -2668 34619 -2622 34739
rect -2622 34619 -2617 34739
rect -3133 34500 -3132 34543
rect -3132 34500 -3078 34543
rect -3078 34500 -3077 34543
rect -3133 34487 -3077 34500
rect -2949 34500 -2948 34543
rect -2948 34500 -2894 34543
rect -2894 34500 -2893 34543
rect -2949 34487 -2893 34500
rect -2765 34500 -2764 34543
rect -2764 34500 -2710 34543
rect -2710 34500 -2709 34543
rect -2765 34487 -2709 34500
rect -3133 34337 -3077 34393
rect 5129 35306 5185 35362
rect 4761 34919 4766 35039
rect 4766 34919 4812 35039
rect 4812 34919 4817 35039
rect 5129 34919 5134 35039
rect 5134 34919 5180 35039
rect 5180 34919 5185 35039
rect 4945 34619 4950 34739
rect 4950 34619 4996 34739
rect 4996 34619 5001 34739
rect 5451 34918 5456 35039
rect 5456 34918 5502 35039
rect 5502 34918 5507 35039
rect 5313 34619 5318 34739
rect 5318 34619 5364 34739
rect 5364 34619 5369 34739
rect 4853 34500 4854 34543
rect 4854 34500 4908 34543
rect 4908 34500 4909 34543
rect 4853 34487 4909 34500
rect 5037 34500 5038 34543
rect 5038 34500 5092 34543
rect 5092 34500 5093 34543
rect 5037 34487 5093 34500
rect 5221 34500 5222 34543
rect 5222 34500 5276 34543
rect 5276 34500 5277 34543
rect 5221 34487 5277 34500
rect 4853 34337 4909 34393
rect 14601 37512 14657 37568
rect 14233 37125 14238 37245
rect 14238 37125 14284 37245
rect 14284 37125 14289 37245
rect 14601 37125 14606 37245
rect 14606 37125 14652 37245
rect 14652 37125 14657 37245
rect 14417 36825 14422 36945
rect 14422 36825 14468 36945
rect 14468 36825 14473 36945
rect 14923 37124 14928 37245
rect 14928 37124 14974 37245
rect 14974 37124 14979 37245
rect 14785 36825 14790 36945
rect 14790 36825 14836 36945
rect 14836 36825 14841 36945
rect 14325 36706 14326 36749
rect 14326 36706 14380 36749
rect 14380 36706 14381 36749
rect 14325 36693 14381 36706
rect 14509 36706 14510 36749
rect 14510 36706 14564 36749
rect 14564 36706 14565 36749
rect 14509 36693 14565 36706
rect 14693 36706 14694 36749
rect 14694 36706 14748 36749
rect 14748 36706 14749 36749
rect 14693 36693 14749 36706
rect 13437 36543 13493 36599
rect 14325 36543 14381 36599
rect 13653 36427 13709 36483
rect 14509 36427 14565 36483
rect 14838 36427 14894 36483
rect 15095 36427 15151 36483
rect 14693 36311 14749 36367
rect 14325 36204 14381 36217
rect 14325 36161 14326 36204
rect 14326 36161 14380 36204
rect 14380 36161 14381 36204
rect 14509 36204 14565 36217
rect 14509 36161 14510 36204
rect 14510 36161 14564 36204
rect 14564 36161 14565 36204
rect 14693 36204 14749 36217
rect 14693 36161 14694 36204
rect 14694 36161 14748 36204
rect 14748 36161 14749 36204
rect 14785 35965 14790 36085
rect 14790 35965 14836 36085
rect 14836 35965 14841 36085
rect 14100 35642 14156 35698
rect 14918 35642 14974 35698
rect 15271 35524 15327 35580
rect 15095 35416 15151 35470
rect 6615 35306 6671 35362
rect 6247 34919 6252 35039
rect 6252 34919 6298 35039
rect 6298 34919 6303 35039
rect 6615 34919 6620 35039
rect 6620 34919 6666 35039
rect 6666 34919 6671 35039
rect 6431 34619 6436 34739
rect 6436 34619 6482 34739
rect 6482 34619 6487 34739
rect 6937 34918 6942 35039
rect 6942 34918 6988 35039
rect 6988 34918 6993 35039
rect 6799 34619 6804 34739
rect 6804 34619 6850 34739
rect 6850 34619 6855 34739
rect 6339 34500 6340 34543
rect 6340 34500 6394 34543
rect 6394 34500 6395 34543
rect 6339 34487 6395 34500
rect 6523 34500 6524 34543
rect 6524 34500 6578 34543
rect 6578 34500 6579 34543
rect 6523 34487 6579 34500
rect 6707 34500 6708 34543
rect 6708 34500 6762 34543
rect 6762 34500 6763 34543
rect 6707 34487 6763 34500
rect 6339 34337 6395 34393
rect 14601 35307 14657 35363
rect 14233 34920 14238 35040
rect 14238 34920 14284 35040
rect 14284 34920 14289 35040
rect 14601 34920 14606 35040
rect 14606 34920 14652 35040
rect 14652 34920 14657 35040
rect 14417 34620 14422 34740
rect 14422 34620 14468 34740
rect 14468 34620 14473 34740
rect 14923 34919 14928 35040
rect 14928 34919 14974 35040
rect 14974 34919 14979 35040
rect 14785 34620 14790 34740
rect 14790 34620 14836 34740
rect 14836 34620 14841 34740
rect 14325 34501 14326 34544
rect 14326 34501 14380 34544
rect 14380 34501 14381 34544
rect 14325 34488 14381 34501
rect 14509 34501 14510 34544
rect 14510 34501 14564 34544
rect 14564 34501 14565 34544
rect 14509 34488 14565 34501
rect 14693 34501 14694 34544
rect 14694 34501 14748 34544
rect 14748 34501 14749 34544
rect 14693 34488 14749 34501
rect 14325 34338 14381 34394
rect 24073 37512 24129 37568
rect 23705 37125 23710 37245
rect 23710 37125 23756 37245
rect 23756 37125 23761 37245
rect 24073 37125 24078 37245
rect 24078 37125 24124 37245
rect 24124 37125 24129 37245
rect 23889 36825 23894 36945
rect 23894 36825 23940 36945
rect 23940 36825 23945 36945
rect 24395 37124 24400 37245
rect 24400 37124 24446 37245
rect 24446 37124 24451 37245
rect 24257 36825 24262 36945
rect 24262 36825 24308 36945
rect 24308 36825 24313 36945
rect 23797 36706 23798 36749
rect 23798 36706 23852 36749
rect 23852 36706 23853 36749
rect 23797 36693 23853 36706
rect 23981 36706 23982 36749
rect 23982 36706 24036 36749
rect 24036 36706 24037 36749
rect 23981 36693 24037 36706
rect 24165 36706 24166 36749
rect 24166 36706 24220 36749
rect 24220 36706 24221 36749
rect 24165 36693 24221 36706
rect 22909 36543 22965 36599
rect 23797 36543 23853 36599
rect 23125 36427 23181 36483
rect 23981 36427 24037 36483
rect 24310 36427 24366 36483
rect 24567 36427 24623 36483
rect 24165 36311 24221 36367
rect 23797 36204 23853 36217
rect 23797 36161 23798 36204
rect 23798 36161 23852 36204
rect 23852 36161 23853 36204
rect 23981 36204 24037 36217
rect 23981 36161 23982 36204
rect 23982 36161 24036 36204
rect 24036 36161 24037 36204
rect 24165 36204 24221 36217
rect 24165 36161 24166 36204
rect 24166 36161 24220 36204
rect 24220 36161 24221 36204
rect 24257 35965 24262 36085
rect 24262 35965 24308 36085
rect 24308 35965 24313 36085
rect 23572 35642 23628 35698
rect 24390 35642 24446 35698
rect 24743 35524 24799 35580
rect 24567 35416 24623 35470
rect 16087 35307 16143 35363
rect 15719 34920 15724 35040
rect 15724 34920 15770 35040
rect 15770 34920 15775 35040
rect 16087 34920 16092 35040
rect 16092 34920 16138 35040
rect 16138 34920 16143 35040
rect 15903 34620 15908 34740
rect 15908 34620 15954 34740
rect 15954 34620 15959 34740
rect 16409 34919 16414 35040
rect 16414 34919 16460 35040
rect 16460 34919 16465 35040
rect 16271 34620 16276 34740
rect 16276 34620 16322 34740
rect 16322 34620 16327 34740
rect 15811 34501 15812 34544
rect 15812 34501 15866 34544
rect 15866 34501 15867 34544
rect 15811 34488 15867 34501
rect 15995 34501 15996 34544
rect 15996 34501 16050 34544
rect 16050 34501 16051 34544
rect 15995 34488 16051 34501
rect 16179 34501 16180 34544
rect 16180 34501 16234 34544
rect 16234 34501 16235 34544
rect 16179 34488 16235 34501
rect 15811 34338 15867 34394
rect 24073 35307 24129 35363
rect 23705 34920 23710 35040
rect 23710 34920 23756 35040
rect 23756 34920 23761 35040
rect 24073 34920 24078 35040
rect 24078 34920 24124 35040
rect 24124 34920 24129 35040
rect 23889 34620 23894 34740
rect 23894 34620 23940 34740
rect 23940 34620 23945 34740
rect 24395 34919 24400 35040
rect 24400 34919 24446 35040
rect 24446 34919 24451 35040
rect 24257 34620 24262 34740
rect 24262 34620 24308 34740
rect 24308 34620 24313 34740
rect 23797 34501 23798 34544
rect 23798 34501 23852 34544
rect 23852 34501 23853 34544
rect 23797 34488 23853 34501
rect 23981 34501 23982 34544
rect 23982 34501 24036 34544
rect 24036 34501 24037 34544
rect 23981 34488 24037 34501
rect 24165 34501 24166 34544
rect 24166 34501 24220 34544
rect 24220 34501 24221 34544
rect 24165 34488 24221 34501
rect 23797 34338 23853 34394
rect 33545 37512 33601 37568
rect 33177 37125 33182 37245
rect 33182 37125 33228 37245
rect 33228 37125 33233 37245
rect 33545 37125 33550 37245
rect 33550 37125 33596 37245
rect 33596 37125 33601 37245
rect 33361 36825 33366 36945
rect 33366 36825 33412 36945
rect 33412 36825 33417 36945
rect 33867 37124 33872 37245
rect 33872 37124 33918 37245
rect 33918 37124 33923 37245
rect 33729 36825 33734 36945
rect 33734 36825 33780 36945
rect 33780 36825 33785 36945
rect 33269 36706 33270 36749
rect 33270 36706 33324 36749
rect 33324 36706 33325 36749
rect 33269 36693 33325 36706
rect 33453 36706 33454 36749
rect 33454 36706 33508 36749
rect 33508 36706 33509 36749
rect 33453 36693 33509 36706
rect 33637 36706 33638 36749
rect 33638 36706 33692 36749
rect 33692 36706 33693 36749
rect 33637 36693 33693 36706
rect 32381 36543 32437 36599
rect 33269 36543 33325 36599
rect 32597 36427 32653 36483
rect 33453 36427 33509 36483
rect 33782 36427 33838 36483
rect 34039 36427 34095 36483
rect 33637 36311 33693 36367
rect 33269 36204 33325 36217
rect 33269 36161 33270 36204
rect 33270 36161 33324 36204
rect 33324 36161 33325 36204
rect 33453 36204 33509 36217
rect 33453 36161 33454 36204
rect 33454 36161 33508 36204
rect 33508 36161 33509 36204
rect 33637 36204 33693 36217
rect 33637 36161 33638 36204
rect 33638 36161 33692 36204
rect 33692 36161 33693 36204
rect 33729 35965 33734 36085
rect 33734 35965 33780 36085
rect 33780 35965 33785 36085
rect 33044 35642 33100 35698
rect 33862 35642 33918 35698
rect 34215 35524 34271 35580
rect 34039 35416 34095 35470
rect 25559 35307 25615 35363
rect 25191 34920 25196 35040
rect 25196 34920 25242 35040
rect 25242 34920 25247 35040
rect 25559 34920 25564 35040
rect 25564 34920 25610 35040
rect 25610 34920 25615 35040
rect 25375 34620 25380 34740
rect 25380 34620 25426 34740
rect 25426 34620 25431 34740
rect 25881 34919 25886 35040
rect 25886 34919 25932 35040
rect 25932 34919 25937 35040
rect 25743 34620 25748 34740
rect 25748 34620 25794 34740
rect 25794 34620 25799 34740
rect 25283 34501 25284 34544
rect 25284 34501 25338 34544
rect 25338 34501 25339 34544
rect 25283 34488 25339 34501
rect 25467 34501 25468 34544
rect 25468 34501 25522 34544
rect 25522 34501 25523 34544
rect 25467 34488 25523 34501
rect 25651 34501 25652 34544
rect 25652 34501 25706 34544
rect 25706 34501 25707 34544
rect 25651 34488 25707 34501
rect 25283 34338 25339 34394
rect 33545 35307 33601 35363
rect 33177 34920 33182 35040
rect 33182 34920 33228 35040
rect 33228 34920 33233 35040
rect 33545 34920 33550 35040
rect 33550 34920 33596 35040
rect 33596 34920 33601 35040
rect 33361 34620 33366 34740
rect 33366 34620 33412 34740
rect 33412 34620 33417 34740
rect 33867 34919 33872 35040
rect 33872 34919 33918 35040
rect 33918 34919 33923 35040
rect 33729 34620 33734 34740
rect 33734 34620 33780 34740
rect 33780 34620 33785 34740
rect 33269 34501 33270 34544
rect 33270 34501 33324 34544
rect 33324 34501 33325 34544
rect 33269 34488 33325 34501
rect 33453 34501 33454 34544
rect 33454 34501 33508 34544
rect 33508 34501 33509 34544
rect 33453 34488 33509 34501
rect 33637 34501 33638 34544
rect 33638 34501 33692 34544
rect 33692 34501 33693 34544
rect 33637 34488 33693 34501
rect 33269 34338 33325 34394
rect 43017 37512 43073 37568
rect 42649 37125 42654 37245
rect 42654 37125 42700 37245
rect 42700 37125 42705 37245
rect 43017 37125 43022 37245
rect 43022 37125 43068 37245
rect 43068 37125 43073 37245
rect 42833 36825 42838 36945
rect 42838 36825 42884 36945
rect 42884 36825 42889 36945
rect 43339 37124 43344 37245
rect 43344 37124 43390 37245
rect 43390 37124 43395 37245
rect 43201 36825 43206 36945
rect 43206 36825 43252 36945
rect 43252 36825 43257 36945
rect 42741 36706 42742 36749
rect 42742 36706 42796 36749
rect 42796 36706 42797 36749
rect 42741 36693 42797 36706
rect 42925 36706 42926 36749
rect 42926 36706 42980 36749
rect 42980 36706 42981 36749
rect 42925 36693 42981 36706
rect 43109 36706 43110 36749
rect 43110 36706 43164 36749
rect 43164 36706 43165 36749
rect 43109 36693 43165 36706
rect 41853 36543 41909 36599
rect 42741 36543 42797 36599
rect 42069 36427 42125 36483
rect 42925 36427 42981 36483
rect 43254 36427 43310 36483
rect 43511 36427 43567 36483
rect 43109 36311 43165 36367
rect 42741 36204 42797 36217
rect 42741 36161 42742 36204
rect 42742 36161 42796 36204
rect 42796 36161 42797 36204
rect 42925 36204 42981 36217
rect 42925 36161 42926 36204
rect 42926 36161 42980 36204
rect 42980 36161 42981 36204
rect 43109 36204 43165 36217
rect 43109 36161 43110 36204
rect 43110 36161 43164 36204
rect 43164 36161 43165 36204
rect 43201 35965 43206 36085
rect 43206 35965 43252 36085
rect 43252 35965 43257 36085
rect 42516 35642 42572 35698
rect 43334 35642 43390 35698
rect 43687 35524 43743 35580
rect 43511 35416 43567 35470
rect 35031 35307 35087 35363
rect 34663 34920 34668 35040
rect 34668 34920 34714 35040
rect 34714 34920 34719 35040
rect 35031 34920 35036 35040
rect 35036 34920 35082 35040
rect 35082 34920 35087 35040
rect 34847 34620 34852 34740
rect 34852 34620 34898 34740
rect 34898 34620 34903 34740
rect 35353 34919 35358 35040
rect 35358 34919 35404 35040
rect 35404 34919 35409 35040
rect 35215 34620 35220 34740
rect 35220 34620 35266 34740
rect 35266 34620 35271 34740
rect 34755 34501 34756 34544
rect 34756 34501 34810 34544
rect 34810 34501 34811 34544
rect 34755 34488 34811 34501
rect 34939 34501 34940 34544
rect 34940 34501 34994 34544
rect 34994 34501 34995 34544
rect 34939 34488 34995 34501
rect 35123 34501 35124 34544
rect 35124 34501 35178 34544
rect 35178 34501 35179 34544
rect 35123 34488 35179 34501
rect 34755 34338 34811 34394
rect 43017 35307 43073 35363
rect 42649 34920 42654 35040
rect 42654 34920 42700 35040
rect 42700 34920 42705 35040
rect 43017 34920 43022 35040
rect 43022 34920 43068 35040
rect 43068 34920 43073 35040
rect 42833 34620 42838 34740
rect 42838 34620 42884 34740
rect 42884 34620 42889 34740
rect 43339 34919 43344 35040
rect 43344 34919 43390 35040
rect 43390 34919 43395 35040
rect 43201 34620 43206 34740
rect 43206 34620 43252 34740
rect 43252 34620 43257 34740
rect 42741 34501 42742 34544
rect 42742 34501 42796 34544
rect 42796 34501 42797 34544
rect 42741 34488 42797 34501
rect 42925 34501 42926 34544
rect 42926 34501 42980 34544
rect 42980 34501 42981 34544
rect 42925 34488 42981 34501
rect 43109 34501 43110 34544
rect 43110 34501 43164 34544
rect 43164 34501 43165 34544
rect 43109 34488 43165 34501
rect 42741 34338 42797 34394
rect 44503 35307 44559 35363
rect 44135 34920 44140 35040
rect 44140 34920 44186 35040
rect 44186 34920 44191 35040
rect 44503 34920 44508 35040
rect 44508 34920 44554 35040
rect 44554 34920 44559 35040
rect 44319 34620 44324 34740
rect 44324 34620 44370 34740
rect 44370 34620 44375 34740
rect 44825 34919 44830 35040
rect 44830 34919 44876 35040
rect 44876 34919 44881 35040
rect 44687 34620 44692 34740
rect 44692 34620 44738 34740
rect 44738 34620 44743 34740
rect 44227 34501 44228 34544
rect 44228 34501 44282 34544
rect 44282 34501 44283 34544
rect 44227 34488 44283 34501
rect 44411 34501 44412 34544
rect 44412 34501 44466 34544
rect 44466 34501 44467 34544
rect 44411 34488 44467 34501
rect 44595 34501 44596 34544
rect 44596 34501 44650 34544
rect 44650 34501 44651 34544
rect 44595 34488 44651 34501
rect 44227 34338 44283 34394
rect -5427 34221 -5371 34277
rect -4435 34221 -4379 34277
rect -4106 34221 -4050 34277
rect -3673 34221 -3617 34277
rect -2949 34221 -2893 34277
rect -2620 34221 -2564 34277
rect -2363 34221 -2307 34277
rect 4045 34221 4101 34277
rect 5037 34221 5093 34277
rect 5366 34221 5422 34277
rect 5799 34221 5855 34277
rect 6523 34221 6579 34277
rect 6852 34221 6908 34277
rect 7109 34221 7165 34277
rect 13517 34222 13573 34278
rect 14509 34222 14565 34278
rect 14838 34222 14894 34278
rect 15271 34222 15327 34278
rect 15995 34222 16051 34278
rect 16324 34222 16380 34278
rect 16581 34222 16637 34278
rect 22989 34222 23045 34278
rect 23981 34222 24037 34278
rect 24310 34222 24366 34278
rect 24743 34222 24799 34278
rect 25467 34222 25523 34278
rect 25796 34222 25852 34278
rect 26053 34222 26109 34278
rect 32461 34222 32517 34278
rect 33453 34222 33509 34278
rect 33782 34222 33838 34278
rect 34215 34222 34271 34278
rect 34939 34222 34995 34278
rect 35268 34222 35324 34278
rect 35525 34222 35581 34278
rect 41933 34222 41989 34278
rect 42925 34222 42981 34278
rect 43254 34222 43310 34278
rect 43687 34222 43743 34278
rect 44411 34222 44467 34278
rect 44740 34222 44796 34278
rect 44997 34222 45053 34278
rect -4251 34105 -4195 34161
rect -2765 34105 -2709 34161
rect -4619 33998 -4563 34011
rect -4619 33955 -4618 33998
rect -4618 33955 -4564 33998
rect -4564 33955 -4563 33998
rect -4435 33998 -4379 34011
rect -4435 33955 -4434 33998
rect -4434 33955 -4380 33998
rect -4380 33955 -4379 33998
rect -4251 33998 -4195 34011
rect -4251 33955 -4250 33998
rect -4250 33955 -4196 33998
rect -4196 33955 -4195 33998
rect -4159 33759 -4154 33879
rect -4154 33759 -4108 33879
rect -4108 33759 -4103 33879
rect -4844 33436 -4788 33492
rect -4026 33436 -3970 33492
rect -5707 33319 -5651 33375
rect 5221 34105 5277 34161
rect -3133 33998 -3077 34011
rect -3133 33955 -3132 33998
rect -3132 33955 -3078 33998
rect -3078 33955 -3077 33998
rect -2949 33998 -2893 34011
rect -2949 33955 -2948 33998
rect -2948 33955 -2894 33998
rect -2894 33955 -2893 33998
rect -2765 33998 -2709 34011
rect -2765 33955 -2764 33998
rect -2764 33955 -2710 33998
rect -2710 33955 -2709 33998
rect -2673 33759 -2668 33879
rect -2668 33759 -2622 33879
rect -2622 33759 -2617 33879
rect -3358 33436 -3302 33492
rect -2540 33436 -2484 33492
rect -2187 33319 -2131 33375
rect 6707 34105 6763 34161
rect 4853 33998 4909 34011
rect 4853 33955 4854 33998
rect 4854 33955 4908 33998
rect 4908 33955 4909 33998
rect 5037 33998 5093 34011
rect 5037 33955 5038 33998
rect 5038 33955 5092 33998
rect 5092 33955 5093 33998
rect 5221 33998 5277 34011
rect 5221 33955 5222 33998
rect 5222 33955 5276 33998
rect 5276 33955 5277 33998
rect 5313 33759 5318 33879
rect 5318 33759 5364 33879
rect 5364 33759 5369 33879
rect 4628 33436 4684 33492
rect 5446 33436 5502 33492
rect 3765 33319 3821 33375
rect 14693 34106 14749 34162
rect 6339 33998 6395 34011
rect 6339 33955 6340 33998
rect 6340 33955 6394 33998
rect 6394 33955 6395 33998
rect 6523 33998 6579 34011
rect 6523 33955 6524 33998
rect 6524 33955 6578 33998
rect 6578 33955 6579 33998
rect 6707 33998 6763 34011
rect 6707 33955 6708 33998
rect 6708 33955 6762 33998
rect 6762 33955 6763 33998
rect 6799 33759 6804 33879
rect 6804 33759 6850 33879
rect 6850 33759 6855 33879
rect 6114 33436 6170 33492
rect 6932 33436 6988 33492
rect 7285 33319 7341 33375
rect -3673 33208 -3617 33264
rect -2363 33209 -2307 33265
rect -4343 33101 -4287 33157
rect -4711 32714 -4706 32834
rect -4706 32714 -4660 32834
rect -4660 32714 -4655 32834
rect -4343 32714 -4338 32834
rect -4338 32714 -4292 32834
rect -4292 32714 -4287 32834
rect -4527 32414 -4522 32534
rect -4522 32414 -4476 32534
rect -4476 32414 -4471 32534
rect -4021 32713 -4016 32834
rect -4016 32713 -3970 32834
rect -3970 32713 -3965 32834
rect -4159 32414 -4154 32534
rect -4154 32414 -4108 32534
rect -4108 32414 -4103 32534
rect -4619 32295 -4618 32338
rect -4618 32295 -4564 32338
rect -4564 32295 -4563 32338
rect -4619 32282 -4563 32295
rect -4435 32295 -4434 32338
rect -4434 32295 -4380 32338
rect -4380 32295 -4379 32338
rect -4435 32282 -4379 32295
rect -4251 32295 -4250 32338
rect -4250 32295 -4196 32338
rect -4196 32295 -4195 32338
rect -4251 32282 -4195 32295
rect -4619 32132 -4563 32188
rect -2857 33102 -2801 33158
rect -3225 32715 -3220 32835
rect -3220 32715 -3174 32835
rect -3174 32715 -3169 32835
rect -2857 32715 -2852 32835
rect -2852 32715 -2806 32835
rect -2806 32715 -2801 32835
rect -3041 32415 -3036 32535
rect -3036 32415 -2990 32535
rect -2990 32415 -2985 32535
rect -2535 32714 -2530 32835
rect -2530 32714 -2484 32835
rect -2484 32714 -2479 32835
rect -2673 32415 -2668 32535
rect -2668 32415 -2622 32535
rect -2622 32415 -2617 32535
rect -3133 32296 -3132 32339
rect -3132 32296 -3078 32339
rect -3078 32296 -3077 32339
rect -3133 32283 -3077 32296
rect -2949 32296 -2948 32339
rect -2948 32296 -2894 32339
rect -2894 32296 -2893 32339
rect -2949 32283 -2893 32296
rect -2765 32296 -2764 32339
rect -2764 32296 -2710 32339
rect -2710 32296 -2709 32339
rect -2765 32283 -2709 32296
rect -3133 32133 -3077 32189
rect -4435 32016 -4379 32072
rect -4106 32016 -4050 32072
rect -3849 32016 -3793 32072
rect -2949 32017 -2893 32073
rect -2620 32017 -2564 32073
rect -2187 32017 -2131 32073
rect -9853 31222 -9848 31462
rect -9848 31222 -9802 31462
rect -9802 31222 -9797 31462
rect -10199 30949 -10143 31005
rect -8761 31222 -8756 31462
rect -8756 31222 -8710 31462
rect -8710 31222 -8705 31462
rect -9751 30949 -9695 31005
rect -8281 31222 -8276 31462
rect -8276 31222 -8230 31462
rect -8230 31222 -8225 31462
rect -6327 31169 -6027 31969
rect 16179 34106 16235 34162
rect 14325 33999 14381 34012
rect 14325 33956 14326 33999
rect 14326 33956 14380 33999
rect 14380 33956 14381 33999
rect 14509 33999 14565 34012
rect 14509 33956 14510 33999
rect 14510 33956 14564 33999
rect 14564 33956 14565 33999
rect 14693 33999 14749 34012
rect 14693 33956 14694 33999
rect 14694 33956 14748 33999
rect 14748 33956 14749 33999
rect 14785 33760 14790 33880
rect 14790 33760 14836 33880
rect 14836 33760 14841 33880
rect 14100 33437 14156 33493
rect 14918 33437 14974 33493
rect 13237 33320 13293 33376
rect 24165 34106 24221 34162
rect 15811 33999 15867 34012
rect 15811 33956 15812 33999
rect 15812 33956 15866 33999
rect 15866 33956 15867 33999
rect 15995 33999 16051 34012
rect 15995 33956 15996 33999
rect 15996 33956 16050 33999
rect 16050 33956 16051 33999
rect 16179 33999 16235 34012
rect 16179 33956 16180 33999
rect 16180 33956 16234 33999
rect 16234 33956 16235 33999
rect 16271 33760 16276 33880
rect 16276 33760 16322 33880
rect 16322 33760 16327 33880
rect 15586 33437 15642 33493
rect 16404 33437 16460 33493
rect 16757 33320 16813 33376
rect 5799 33208 5855 33264
rect 7109 33209 7165 33265
rect 5129 33101 5185 33157
rect 4761 32714 4766 32834
rect 4766 32714 4812 32834
rect 4812 32714 4817 32834
rect 5129 32714 5134 32834
rect 5134 32714 5180 32834
rect 5180 32714 5185 32834
rect 4945 32414 4950 32534
rect 4950 32414 4996 32534
rect 4996 32414 5001 32534
rect 5451 32713 5456 32834
rect 5456 32713 5502 32834
rect 5502 32713 5507 32834
rect 5313 32414 5318 32534
rect 5318 32414 5364 32534
rect 5364 32414 5369 32534
rect 4853 32295 4854 32338
rect 4854 32295 4908 32338
rect 4908 32295 4909 32338
rect 4853 32282 4909 32295
rect 5037 32295 5038 32338
rect 5038 32295 5092 32338
rect 5092 32295 5093 32338
rect 5037 32282 5093 32295
rect 5221 32295 5222 32338
rect 5222 32295 5276 32338
rect 5276 32295 5277 32338
rect 5221 32282 5277 32295
rect 4853 32132 4909 32188
rect 6615 33102 6671 33158
rect 6247 32715 6252 32835
rect 6252 32715 6298 32835
rect 6298 32715 6303 32835
rect 6615 32715 6620 32835
rect 6620 32715 6666 32835
rect 6666 32715 6671 32835
rect 6431 32415 6436 32535
rect 6436 32415 6482 32535
rect 6482 32415 6487 32535
rect 6937 32714 6942 32835
rect 6942 32714 6988 32835
rect 6988 32714 6993 32835
rect 6799 32415 6804 32535
rect 6804 32415 6850 32535
rect 6850 32415 6855 32535
rect 6339 32296 6340 32339
rect 6340 32296 6394 32339
rect 6394 32296 6395 32339
rect 6339 32283 6395 32296
rect 6523 32296 6524 32339
rect 6524 32296 6578 32339
rect 6578 32296 6579 32339
rect 6523 32283 6579 32296
rect 6707 32296 6708 32339
rect 6708 32296 6762 32339
rect 6762 32296 6763 32339
rect 6707 32283 6763 32296
rect 6339 32133 6395 32189
rect 5037 32016 5093 32072
rect 5366 32016 5422 32072
rect 5623 32016 5679 32072
rect 6523 32017 6579 32073
rect 6852 32017 6908 32073
rect 7285 32017 7341 32073
rect -5291 31900 -5235 31956
rect -4251 31900 -4195 31956
rect -8459 30871 -8403 30927
rect -8939 30793 -8883 30849
rect -10543 29802 -10538 30042
rect -10538 29802 -10492 30042
rect -10492 29802 -10487 30042
rect -9649 30511 -9644 30567
rect -9644 30511 -9598 30567
rect -9598 30511 -9593 30567
rect -9169 30511 -9164 30567
rect -9164 30511 -9118 30567
rect -9118 30511 -9113 30567
rect -8965 30511 -8960 30567
rect -8960 30511 -8914 30567
rect -8914 30511 -8909 30567
rect -8761 30511 -8756 30567
rect -8756 30511 -8710 30567
rect -8710 30511 -8705 30567
rect -2765 31901 -2709 31957
rect -4619 31793 -4563 31806
rect -4619 31750 -4618 31793
rect -4618 31750 -4564 31793
rect -4564 31750 -4563 31793
rect -4435 31793 -4379 31806
rect -4435 31750 -4434 31793
rect -4434 31750 -4380 31793
rect -4380 31750 -4379 31793
rect -4251 31793 -4195 31806
rect -4251 31750 -4250 31793
rect -4250 31750 -4196 31793
rect -4196 31750 -4195 31793
rect -4159 31554 -4154 31674
rect -4154 31554 -4108 31674
rect -4108 31554 -4103 31674
rect -4844 31231 -4788 31287
rect -4026 31231 -3970 31287
rect -3673 31113 -3617 31169
rect -7695 30833 -5927 30973
rect -3849 31005 -3793 31059
rect -8281 30511 -8276 30567
rect -8276 30511 -8230 30567
rect -8230 30511 -8225 30567
rect -9985 30090 -9905 30166
rect -8755 30059 -8155 30199
rect -7421 30330 -7416 30570
rect -7416 30330 -7370 30570
rect -7370 30330 -7365 30570
rect -6737 30330 -6732 30570
rect -6732 30330 -6686 30570
rect -6686 30330 -6681 30570
rect -6941 29996 -6936 30236
rect -6936 29996 -6890 30236
rect -6890 29996 -6885 30236
rect -6533 29996 -6528 30236
rect -6528 29996 -6482 30236
rect -6482 29996 -6477 30236
rect -6053 30046 -6048 30286
rect -6048 30046 -6002 30286
rect -6002 30046 -5997 30286
rect -8755 29659 -8155 29799
rect -7523 29773 -7467 29829
rect -10721 29451 -10665 29507
rect -10543 29091 -10538 29147
rect -10538 29091 -10492 29147
rect -10492 29091 -10487 29147
rect -12256 27872 -12251 28112
rect -12251 27872 -12205 28112
rect -12205 27872 -12200 28112
rect -9853 28882 -9848 29122
rect -9848 28882 -9802 29122
rect -9802 28882 -9797 29122
rect -8761 28882 -8756 29122
rect -8756 28882 -8710 29122
rect -8710 28882 -8705 29122
rect -9751 28609 -9695 28665
rect -8281 28882 -8276 29122
rect -8276 28882 -8230 29122
rect -8230 28882 -8225 29122
rect -4343 30896 -4287 30952
rect -4711 30509 -4706 30629
rect -4706 30509 -4660 30629
rect -4660 30509 -4655 30629
rect -4343 30509 -4338 30629
rect -4338 30509 -4292 30629
rect -4292 30509 -4287 30629
rect -4527 30209 -4522 30329
rect -4522 30209 -4476 30329
rect -4476 30209 -4471 30329
rect -4021 30508 -4016 30629
rect -4016 30508 -3970 30629
rect -3970 30508 -3965 30629
rect -4159 30209 -4154 30329
rect -4154 30209 -4108 30329
rect -4108 30209 -4103 30329
rect -4619 30090 -4618 30133
rect -4618 30090 -4564 30133
rect -4564 30090 -4563 30133
rect -4619 30077 -4563 30090
rect -4435 30090 -4434 30133
rect -4434 30090 -4380 30133
rect -4380 30090 -4379 30133
rect -4435 30077 -4379 30090
rect -4251 30090 -4250 30133
rect -4250 30090 -4196 30133
rect -4196 30090 -4195 30133
rect -4251 30077 -4195 30090
rect -4619 29927 -4563 29983
rect -5427 29811 -5371 29867
rect -4435 29811 -4379 29867
rect -4106 29811 -4050 29867
rect -3673 29811 -3617 29867
rect -6231 29695 -6175 29751
rect -5661 29696 -5607 29750
rect -4251 29695 -4195 29751
rect -6839 29617 -6783 29673
rect -7625 29335 -7620 29391
rect -7620 29335 -7574 29391
rect -7574 29335 -7569 29391
rect -6737 29335 -6732 29391
rect -6732 29335 -6686 29391
rect -6686 29335 -6681 29391
rect -6053 29335 -6048 29391
rect -6048 29335 -6002 29391
rect -6002 29335 -5997 29391
rect -4619 29588 -4563 29601
rect -4619 29545 -4618 29588
rect -4618 29545 -4564 29588
rect -4564 29545 -4563 29588
rect -4435 29588 -4379 29601
rect -4435 29545 -4434 29588
rect -4434 29545 -4380 29588
rect -4380 29545 -4379 29588
rect -4251 29588 -4195 29601
rect -4251 29545 -4250 29588
rect -4250 29545 -4196 29588
rect -4196 29545 -4195 29588
rect -4159 29349 -4154 29469
rect -4154 29349 -4108 29469
rect -4108 29349 -4103 29469
rect -4844 29026 -4788 29082
rect -4026 29026 -3970 29082
rect -7695 28873 -5927 29013
rect -3133 31794 -3077 31807
rect -3133 31751 -3132 31794
rect -3132 31751 -3078 31794
rect -3078 31751 -3077 31794
rect -2949 31794 -2893 31807
rect -2949 31751 -2948 31794
rect -2948 31751 -2894 31794
rect -2894 31751 -2893 31794
rect -2765 31794 -2709 31807
rect -2765 31751 -2764 31794
rect -2764 31751 -2710 31794
rect -2710 31751 -2709 31794
rect -2673 31555 -2668 31675
rect -2668 31555 -2622 31675
rect -2622 31555 -2617 31675
rect -3358 31232 -3302 31288
rect -2540 31232 -2484 31288
rect -1245 31169 -1045 31969
rect -381 31222 -376 31462
rect -376 31222 -330 31462
rect -330 31222 -325 31462
rect 711 31222 716 31462
rect 716 31222 762 31462
rect 762 31222 767 31462
rect -279 30949 -223 31005
rect 1191 31222 1196 31462
rect 1196 31222 1242 31462
rect 1242 31222 1247 31462
rect 3145 31169 3445 31969
rect 25651 34106 25707 34162
rect 23797 33999 23853 34012
rect 23797 33956 23798 33999
rect 23798 33956 23852 33999
rect 23852 33956 23853 33999
rect 23981 33999 24037 34012
rect 23981 33956 23982 33999
rect 23982 33956 24036 33999
rect 24036 33956 24037 33999
rect 24165 33999 24221 34012
rect 24165 33956 24166 33999
rect 24166 33956 24220 33999
rect 24220 33956 24221 33999
rect 24257 33760 24262 33880
rect 24262 33760 24308 33880
rect 24308 33760 24313 33880
rect 23572 33437 23628 33493
rect 24390 33437 24446 33493
rect 22709 33320 22765 33376
rect 33637 34106 33693 34162
rect 25283 33999 25339 34012
rect 25283 33956 25284 33999
rect 25284 33956 25338 33999
rect 25338 33956 25339 33999
rect 25467 33999 25523 34012
rect 25467 33956 25468 33999
rect 25468 33956 25522 33999
rect 25522 33956 25523 33999
rect 25651 33999 25707 34012
rect 25651 33956 25652 33999
rect 25652 33956 25706 33999
rect 25706 33956 25707 33999
rect 25743 33760 25748 33880
rect 25748 33760 25794 33880
rect 25794 33760 25799 33880
rect 25058 33437 25114 33493
rect 25876 33437 25932 33493
rect 26229 33320 26285 33376
rect 15271 33209 15327 33265
rect 16581 33210 16637 33266
rect 14601 33102 14657 33158
rect 14233 32715 14238 32835
rect 14238 32715 14284 32835
rect 14284 32715 14289 32835
rect 14601 32715 14606 32835
rect 14606 32715 14652 32835
rect 14652 32715 14657 32835
rect 14417 32415 14422 32535
rect 14422 32415 14468 32535
rect 14468 32415 14473 32535
rect 14923 32714 14928 32835
rect 14928 32714 14974 32835
rect 14974 32714 14979 32835
rect 14785 32415 14790 32535
rect 14790 32415 14836 32535
rect 14836 32415 14841 32535
rect 14325 32296 14326 32339
rect 14326 32296 14380 32339
rect 14380 32296 14381 32339
rect 14325 32283 14381 32296
rect 14509 32296 14510 32339
rect 14510 32296 14564 32339
rect 14564 32296 14565 32339
rect 14509 32283 14565 32296
rect 14693 32296 14694 32339
rect 14694 32296 14748 32339
rect 14748 32296 14749 32339
rect 14693 32283 14749 32296
rect 14325 32133 14381 32189
rect 16087 33103 16143 33159
rect 15719 32716 15724 32836
rect 15724 32716 15770 32836
rect 15770 32716 15775 32836
rect 16087 32716 16092 32836
rect 16092 32716 16138 32836
rect 16138 32716 16143 32836
rect 15903 32416 15908 32536
rect 15908 32416 15954 32536
rect 15954 32416 15959 32536
rect 16409 32715 16414 32836
rect 16414 32715 16460 32836
rect 16460 32715 16465 32836
rect 16271 32416 16276 32536
rect 16276 32416 16322 32536
rect 16322 32416 16327 32536
rect 15811 32297 15812 32340
rect 15812 32297 15866 32340
rect 15866 32297 15867 32340
rect 15811 32284 15867 32297
rect 15995 32297 15996 32340
rect 15996 32297 16050 32340
rect 16050 32297 16051 32340
rect 15995 32284 16051 32297
rect 16179 32297 16180 32340
rect 16180 32297 16234 32340
rect 16234 32297 16235 32340
rect 16179 32284 16235 32297
rect 15811 32134 15867 32190
rect 14509 32017 14565 32073
rect 14838 32017 14894 32073
rect 15095 32017 15151 32073
rect 15995 32018 16051 32074
rect 16324 32018 16380 32074
rect 16757 32018 16813 32074
rect 4181 31900 4237 31956
rect 5221 31900 5277 31956
rect 1013 30871 1069 30927
rect 533 30793 589 30849
rect -1071 29802 -1066 30042
rect -1066 29802 -1020 30042
rect -1020 29802 -1015 30042
rect -177 30511 -172 30567
rect -172 30511 -126 30567
rect -126 30511 -121 30567
rect 303 30511 308 30567
rect 308 30511 354 30567
rect 354 30511 359 30567
rect 507 30511 512 30567
rect 512 30511 558 30567
rect 558 30511 563 30567
rect 711 30511 716 30567
rect 716 30511 762 30567
rect 762 30511 767 30567
rect 6707 31901 6763 31957
rect 4853 31793 4909 31806
rect 4853 31750 4854 31793
rect 4854 31750 4908 31793
rect 4908 31750 4909 31793
rect 5037 31793 5093 31806
rect 5037 31750 5038 31793
rect 5038 31750 5092 31793
rect 5092 31750 5093 31793
rect 5221 31793 5277 31806
rect 5221 31750 5222 31793
rect 5222 31750 5276 31793
rect 5276 31750 5277 31793
rect 5313 31554 5318 31674
rect 5318 31554 5364 31674
rect 5364 31554 5369 31674
rect 4628 31231 4684 31287
rect 5446 31231 5502 31287
rect 5799 31113 5855 31169
rect 1777 30833 3545 30973
rect 5623 31005 5679 31059
rect 1191 30511 1196 30567
rect 1196 30511 1242 30567
rect 1242 30511 1247 30567
rect 717 30059 1317 30199
rect 2051 30330 2056 30570
rect 2056 30330 2102 30570
rect 2102 30330 2107 30570
rect 2735 30330 2740 30570
rect 2740 30330 2786 30570
rect 2786 30330 2791 30570
rect 2531 29996 2536 30236
rect 2536 29996 2582 30236
rect 2582 29996 2587 30236
rect 2939 29996 2944 30236
rect 2944 29996 2990 30236
rect 2990 29996 2995 30236
rect 3419 30046 3424 30286
rect 3424 30046 3470 30286
rect 3470 30046 3475 30286
rect 717 29659 1317 29799
rect 1949 29773 2005 29829
rect -1249 29451 -1193 29507
rect -5610 28908 -5554 28964
rect -5427 28908 -5371 28964
rect -1071 29091 -1066 29147
rect -1066 29091 -1020 29147
rect -1020 29091 -1015 29147
rect -8459 28531 -8403 28587
rect -8939 28453 -8883 28509
rect -9649 28171 -9644 28227
rect -9644 28171 -9598 28227
rect -9598 28171 -9593 28227
rect -9169 28171 -9164 28227
rect -9164 28171 -9118 28227
rect -9118 28171 -9113 28227
rect -8965 28171 -8960 28227
rect -8960 28171 -8914 28227
rect -8914 28171 -8909 28227
rect -8761 28171 -8756 28227
rect -8756 28171 -8710 28227
rect -8710 28171 -8705 28227
rect -8281 28171 -8276 28227
rect -8276 28171 -8230 28227
rect -8230 28171 -8225 28227
rect -6327 27889 -6027 28689
rect -381 28882 -376 29122
rect -376 28882 -330 29122
rect -330 28882 -325 29122
rect 711 28882 716 29122
rect 716 28882 762 29122
rect 762 28882 767 29122
rect -279 28609 -223 28665
rect 1191 28882 1196 29122
rect 1196 28882 1242 29122
rect 1242 28882 1247 29122
rect 5129 30896 5185 30952
rect 4761 30509 4766 30629
rect 4766 30509 4812 30629
rect 4812 30509 4817 30629
rect 5129 30509 5134 30629
rect 5134 30509 5180 30629
rect 5180 30509 5185 30629
rect 4945 30209 4950 30329
rect 4950 30209 4996 30329
rect 4996 30209 5001 30329
rect 5451 30508 5456 30629
rect 5456 30508 5502 30629
rect 5502 30508 5507 30629
rect 5313 30209 5318 30329
rect 5318 30209 5364 30329
rect 5364 30209 5369 30329
rect 4853 30090 4854 30133
rect 4854 30090 4908 30133
rect 4908 30090 4909 30133
rect 4853 30077 4909 30090
rect 5037 30090 5038 30133
rect 5038 30090 5092 30133
rect 5092 30090 5093 30133
rect 5037 30077 5093 30090
rect 5221 30090 5222 30133
rect 5222 30090 5276 30133
rect 5276 30090 5277 30133
rect 5221 30077 5277 30090
rect 4853 29927 4909 29983
rect 4045 29811 4101 29867
rect 5037 29811 5093 29867
rect 5366 29811 5422 29867
rect 5799 29811 5855 29867
rect 3241 29695 3297 29751
rect 3811 29696 3865 29750
rect 5221 29695 5277 29751
rect 2633 29617 2689 29673
rect 1847 29335 1852 29391
rect 1852 29335 1898 29391
rect 1898 29335 1903 29391
rect 2735 29335 2740 29391
rect 2740 29335 2786 29391
rect 2786 29335 2791 29391
rect 3419 29335 3424 29391
rect 3424 29335 3470 29391
rect 3470 29335 3475 29391
rect 4853 29588 4909 29601
rect 4853 29545 4854 29588
rect 4854 29545 4908 29588
rect 4908 29545 4909 29588
rect 5037 29588 5093 29601
rect 5037 29545 5038 29588
rect 5038 29545 5092 29588
rect 5092 29545 5093 29588
rect 5221 29588 5277 29601
rect 5221 29545 5222 29588
rect 5222 29545 5276 29588
rect 5276 29545 5277 29588
rect 5313 29349 5318 29469
rect 5318 29349 5364 29469
rect 5364 29349 5369 29469
rect 4628 29026 4684 29082
rect 5446 29026 5502 29082
rect 1777 28873 3545 29013
rect 6339 31794 6395 31807
rect 6339 31751 6340 31794
rect 6340 31751 6394 31794
rect 6394 31751 6395 31794
rect 6523 31794 6579 31807
rect 6523 31751 6524 31794
rect 6524 31751 6578 31794
rect 6578 31751 6579 31794
rect 6707 31794 6763 31807
rect 6707 31751 6708 31794
rect 6708 31751 6762 31794
rect 6762 31751 6763 31794
rect 6799 31555 6804 31675
rect 6804 31555 6850 31675
rect 6850 31555 6855 31675
rect 6114 31232 6170 31288
rect 6932 31232 6988 31288
rect 8227 31170 8427 31970
rect 9091 31223 9096 31463
rect 9096 31223 9142 31463
rect 9142 31223 9147 31463
rect 10183 31223 10188 31463
rect 10188 31223 10234 31463
rect 10234 31223 10239 31463
rect 9193 30950 9249 31006
rect 10663 31223 10668 31463
rect 10668 31223 10714 31463
rect 10714 31223 10719 31463
rect 12617 31170 12917 31970
rect 35123 34106 35179 34162
rect 33269 33999 33325 34012
rect 33269 33956 33270 33999
rect 33270 33956 33324 33999
rect 33324 33956 33325 33999
rect 33453 33999 33509 34012
rect 33453 33956 33454 33999
rect 33454 33956 33508 33999
rect 33508 33956 33509 33999
rect 33637 33999 33693 34012
rect 33637 33956 33638 33999
rect 33638 33956 33692 33999
rect 33692 33956 33693 33999
rect 33729 33760 33734 33880
rect 33734 33760 33780 33880
rect 33780 33760 33785 33880
rect 33044 33437 33100 33493
rect 33862 33437 33918 33493
rect 32181 33320 32237 33376
rect 43109 34106 43165 34162
rect 34755 33999 34811 34012
rect 34755 33956 34756 33999
rect 34756 33956 34810 33999
rect 34810 33956 34811 33999
rect 34939 33999 34995 34012
rect 34939 33956 34940 33999
rect 34940 33956 34994 33999
rect 34994 33956 34995 33999
rect 35123 33999 35179 34012
rect 35123 33956 35124 33999
rect 35124 33956 35178 33999
rect 35178 33956 35179 33999
rect 35215 33760 35220 33880
rect 35220 33760 35266 33880
rect 35266 33760 35271 33880
rect 34530 33437 34586 33493
rect 35348 33437 35404 33493
rect 35701 33320 35757 33376
rect 24743 33209 24799 33265
rect 26053 33210 26109 33266
rect 24073 33102 24129 33158
rect 23705 32715 23710 32835
rect 23710 32715 23756 32835
rect 23756 32715 23761 32835
rect 24073 32715 24078 32835
rect 24078 32715 24124 32835
rect 24124 32715 24129 32835
rect 23889 32415 23894 32535
rect 23894 32415 23940 32535
rect 23940 32415 23945 32535
rect 24395 32714 24400 32835
rect 24400 32714 24446 32835
rect 24446 32714 24451 32835
rect 24257 32415 24262 32535
rect 24262 32415 24308 32535
rect 24308 32415 24313 32535
rect 23797 32296 23798 32339
rect 23798 32296 23852 32339
rect 23852 32296 23853 32339
rect 23797 32283 23853 32296
rect 23981 32296 23982 32339
rect 23982 32296 24036 32339
rect 24036 32296 24037 32339
rect 23981 32283 24037 32296
rect 24165 32296 24166 32339
rect 24166 32296 24220 32339
rect 24220 32296 24221 32339
rect 24165 32283 24221 32296
rect 23797 32133 23853 32189
rect 25559 33103 25615 33159
rect 25191 32716 25196 32836
rect 25196 32716 25242 32836
rect 25242 32716 25247 32836
rect 25559 32716 25564 32836
rect 25564 32716 25610 32836
rect 25610 32716 25615 32836
rect 25375 32416 25380 32536
rect 25380 32416 25426 32536
rect 25426 32416 25431 32536
rect 25881 32715 25886 32836
rect 25886 32715 25932 32836
rect 25932 32715 25937 32836
rect 25743 32416 25748 32536
rect 25748 32416 25794 32536
rect 25794 32416 25799 32536
rect 25283 32297 25284 32340
rect 25284 32297 25338 32340
rect 25338 32297 25339 32340
rect 25283 32284 25339 32297
rect 25467 32297 25468 32340
rect 25468 32297 25522 32340
rect 25522 32297 25523 32340
rect 25467 32284 25523 32297
rect 25651 32297 25652 32340
rect 25652 32297 25706 32340
rect 25706 32297 25707 32340
rect 25651 32284 25707 32297
rect 25283 32134 25339 32190
rect 23981 32017 24037 32073
rect 24310 32017 24366 32073
rect 24567 32017 24623 32073
rect 25467 32018 25523 32074
rect 25796 32018 25852 32074
rect 26229 32018 26285 32074
rect 13653 31901 13709 31957
rect 14693 31901 14749 31957
rect 10485 30872 10541 30928
rect 10005 30794 10061 30850
rect 8401 29803 8406 30043
rect 8406 29803 8452 30043
rect 8452 29803 8457 30043
rect 9295 30512 9300 30568
rect 9300 30512 9346 30568
rect 9346 30512 9351 30568
rect 9775 30512 9780 30568
rect 9780 30512 9826 30568
rect 9826 30512 9831 30568
rect 9979 30512 9984 30568
rect 9984 30512 10030 30568
rect 10030 30512 10035 30568
rect 10183 30512 10188 30568
rect 10188 30512 10234 30568
rect 10234 30512 10239 30568
rect 16179 31902 16235 31958
rect 14325 31794 14381 31807
rect 14325 31751 14326 31794
rect 14326 31751 14380 31794
rect 14380 31751 14381 31794
rect 14509 31794 14565 31807
rect 14509 31751 14510 31794
rect 14510 31751 14564 31794
rect 14564 31751 14565 31794
rect 14693 31794 14749 31807
rect 14693 31751 14694 31794
rect 14694 31751 14748 31794
rect 14748 31751 14749 31794
rect 14785 31555 14790 31675
rect 14790 31555 14836 31675
rect 14836 31555 14841 31675
rect 14100 31232 14156 31288
rect 14918 31232 14974 31288
rect 15271 31114 15327 31170
rect 11249 30834 13017 30974
rect 15095 31006 15151 31060
rect 10663 30512 10668 30568
rect 10668 30512 10714 30568
rect 10714 30512 10719 30568
rect 10189 30060 10789 30200
rect 11523 30331 11528 30571
rect 11528 30331 11574 30571
rect 11574 30331 11579 30571
rect 12207 30331 12212 30571
rect 12212 30331 12258 30571
rect 12258 30331 12263 30571
rect 12003 29997 12008 30237
rect 12008 29997 12054 30237
rect 12054 29997 12059 30237
rect 12411 29997 12416 30237
rect 12416 29997 12462 30237
rect 12462 29997 12467 30237
rect 12891 30047 12896 30287
rect 12896 30047 12942 30287
rect 12942 30047 12947 30287
rect 10189 29660 10789 29800
rect 11421 29774 11477 29830
rect 8223 29452 8279 29508
rect 3862 28908 3918 28964
rect 4045 28908 4101 28964
rect 8401 29092 8406 29148
rect 8406 29092 8452 29148
rect 8452 29092 8457 29148
rect 1013 28531 1069 28587
rect 533 28453 589 28509
rect -177 28171 -172 28227
rect -172 28171 -126 28227
rect -126 28171 -121 28227
rect 303 28171 308 28227
rect 308 28171 354 28227
rect 354 28171 359 28227
rect 507 28171 512 28227
rect 512 28171 558 28227
rect 558 28171 563 28227
rect 711 28171 716 28227
rect 716 28171 762 28227
rect 762 28171 767 28227
rect 1191 28171 1196 28227
rect 1196 28171 1242 28227
rect 1242 28171 1247 28227
rect 3145 27889 3445 28689
rect 9091 28883 9096 29123
rect 9096 28883 9142 29123
rect 9142 28883 9147 29123
rect 10183 28883 10188 29123
rect 10188 28883 10234 29123
rect 10234 28883 10239 29123
rect 9193 28610 9249 28666
rect 10663 28883 10668 29123
rect 10668 28883 10714 29123
rect 10714 28883 10719 29123
rect 14601 30897 14657 30953
rect 14233 30510 14238 30630
rect 14238 30510 14284 30630
rect 14284 30510 14289 30630
rect 14601 30510 14606 30630
rect 14606 30510 14652 30630
rect 14652 30510 14657 30630
rect 14417 30210 14422 30330
rect 14422 30210 14468 30330
rect 14468 30210 14473 30330
rect 14923 30509 14928 30630
rect 14928 30509 14974 30630
rect 14974 30509 14979 30630
rect 14785 30210 14790 30330
rect 14790 30210 14836 30330
rect 14836 30210 14841 30330
rect 14325 30091 14326 30134
rect 14326 30091 14380 30134
rect 14380 30091 14381 30134
rect 14325 30078 14381 30091
rect 14509 30091 14510 30134
rect 14510 30091 14564 30134
rect 14564 30091 14565 30134
rect 14509 30078 14565 30091
rect 14693 30091 14694 30134
rect 14694 30091 14748 30134
rect 14748 30091 14749 30134
rect 14693 30078 14749 30091
rect 14325 29928 14381 29984
rect 13517 29812 13573 29868
rect 14509 29812 14565 29868
rect 14838 29812 14894 29868
rect 15271 29812 15327 29868
rect 12713 29696 12769 29752
rect 13283 29697 13337 29751
rect 14693 29696 14749 29752
rect 12105 29618 12161 29674
rect 11319 29336 11324 29392
rect 11324 29336 11370 29392
rect 11370 29336 11375 29392
rect 12207 29336 12212 29392
rect 12212 29336 12258 29392
rect 12258 29336 12263 29392
rect 12891 29336 12896 29392
rect 12896 29336 12942 29392
rect 12942 29336 12947 29392
rect 14325 29589 14381 29602
rect 14325 29546 14326 29589
rect 14326 29546 14380 29589
rect 14380 29546 14381 29589
rect 14509 29589 14565 29602
rect 14509 29546 14510 29589
rect 14510 29546 14564 29589
rect 14564 29546 14565 29589
rect 14693 29589 14749 29602
rect 14693 29546 14694 29589
rect 14694 29546 14748 29589
rect 14748 29546 14749 29589
rect 14785 29350 14790 29470
rect 14790 29350 14836 29470
rect 14836 29350 14841 29470
rect 14100 29027 14156 29083
rect 14918 29027 14974 29083
rect 11249 28874 13017 29014
rect 15811 31795 15867 31808
rect 15811 31752 15812 31795
rect 15812 31752 15866 31795
rect 15866 31752 15867 31795
rect 15995 31795 16051 31808
rect 15995 31752 15996 31795
rect 15996 31752 16050 31795
rect 16050 31752 16051 31795
rect 16179 31795 16235 31808
rect 16179 31752 16180 31795
rect 16180 31752 16234 31795
rect 16234 31752 16235 31795
rect 16271 31556 16276 31676
rect 16276 31556 16322 31676
rect 16322 31556 16327 31676
rect 15586 31233 15642 31289
rect 16404 31233 16460 31289
rect 17699 31170 17899 31970
rect 18563 31223 18568 31463
rect 18568 31223 18614 31463
rect 18614 31223 18619 31463
rect 19655 31223 19660 31463
rect 19660 31223 19706 31463
rect 19706 31223 19711 31463
rect 18665 30950 18721 31006
rect 20135 31223 20140 31463
rect 20140 31223 20186 31463
rect 20186 31223 20191 31463
rect 22089 31170 22389 31970
rect 44595 34106 44651 34162
rect 42741 33999 42797 34012
rect 42741 33956 42742 33999
rect 42742 33956 42796 33999
rect 42796 33956 42797 33999
rect 42925 33999 42981 34012
rect 42925 33956 42926 33999
rect 42926 33956 42980 33999
rect 42980 33956 42981 33999
rect 43109 33999 43165 34012
rect 43109 33956 43110 33999
rect 43110 33956 43164 33999
rect 43164 33956 43165 33999
rect 43201 33760 43206 33880
rect 43206 33760 43252 33880
rect 43252 33760 43257 33880
rect 42516 33437 42572 33493
rect 43334 33437 43390 33493
rect 41653 33320 41709 33376
rect 44227 33999 44283 34012
rect 44227 33956 44228 33999
rect 44228 33956 44282 33999
rect 44282 33956 44283 33999
rect 44411 33999 44467 34012
rect 44411 33956 44412 33999
rect 44412 33956 44466 33999
rect 44466 33956 44467 33999
rect 44595 33999 44651 34012
rect 44595 33956 44596 33999
rect 44596 33956 44650 33999
rect 44650 33956 44651 33999
rect 44687 33760 44692 33880
rect 44692 33760 44738 33880
rect 44738 33760 44743 33880
rect 44002 33437 44058 33493
rect 44820 33437 44876 33493
rect 45173 33320 45229 33376
rect 34215 33209 34271 33265
rect 35525 33210 35581 33266
rect 33545 33102 33601 33158
rect 33177 32715 33182 32835
rect 33182 32715 33228 32835
rect 33228 32715 33233 32835
rect 33545 32715 33550 32835
rect 33550 32715 33596 32835
rect 33596 32715 33601 32835
rect 33361 32415 33366 32535
rect 33366 32415 33412 32535
rect 33412 32415 33417 32535
rect 33867 32714 33872 32835
rect 33872 32714 33918 32835
rect 33918 32714 33923 32835
rect 33729 32415 33734 32535
rect 33734 32415 33780 32535
rect 33780 32415 33785 32535
rect 33269 32296 33270 32339
rect 33270 32296 33324 32339
rect 33324 32296 33325 32339
rect 33269 32283 33325 32296
rect 33453 32296 33454 32339
rect 33454 32296 33508 32339
rect 33508 32296 33509 32339
rect 33453 32283 33509 32296
rect 33637 32296 33638 32339
rect 33638 32296 33692 32339
rect 33692 32296 33693 32339
rect 33637 32283 33693 32296
rect 33269 32133 33325 32189
rect 35031 33103 35087 33159
rect 34663 32716 34668 32836
rect 34668 32716 34714 32836
rect 34714 32716 34719 32836
rect 35031 32716 35036 32836
rect 35036 32716 35082 32836
rect 35082 32716 35087 32836
rect 34847 32416 34852 32536
rect 34852 32416 34898 32536
rect 34898 32416 34903 32536
rect 35353 32715 35358 32836
rect 35358 32715 35404 32836
rect 35404 32715 35409 32836
rect 35215 32416 35220 32536
rect 35220 32416 35266 32536
rect 35266 32416 35271 32536
rect 34755 32297 34756 32340
rect 34756 32297 34810 32340
rect 34810 32297 34811 32340
rect 34755 32284 34811 32297
rect 34939 32297 34940 32340
rect 34940 32297 34994 32340
rect 34994 32297 34995 32340
rect 34939 32284 34995 32297
rect 35123 32297 35124 32340
rect 35124 32297 35178 32340
rect 35178 32297 35179 32340
rect 35123 32284 35179 32297
rect 34755 32134 34811 32190
rect 33453 32017 33509 32073
rect 33782 32017 33838 32073
rect 34039 32017 34095 32073
rect 34939 32018 34995 32074
rect 35268 32018 35324 32074
rect 35701 32018 35757 32074
rect 23125 31901 23181 31957
rect 24165 31901 24221 31957
rect 19957 30872 20013 30928
rect 19477 30794 19533 30850
rect 17873 29803 17878 30043
rect 17878 29803 17924 30043
rect 17924 29803 17929 30043
rect 18767 30512 18772 30568
rect 18772 30512 18818 30568
rect 18818 30512 18823 30568
rect 19247 30512 19252 30568
rect 19252 30512 19298 30568
rect 19298 30512 19303 30568
rect 19451 30512 19456 30568
rect 19456 30512 19502 30568
rect 19502 30512 19507 30568
rect 19655 30512 19660 30568
rect 19660 30512 19706 30568
rect 19706 30512 19711 30568
rect 25651 31902 25707 31958
rect 23797 31794 23853 31807
rect 23797 31751 23798 31794
rect 23798 31751 23852 31794
rect 23852 31751 23853 31794
rect 23981 31794 24037 31807
rect 23981 31751 23982 31794
rect 23982 31751 24036 31794
rect 24036 31751 24037 31794
rect 24165 31794 24221 31807
rect 24165 31751 24166 31794
rect 24166 31751 24220 31794
rect 24220 31751 24221 31794
rect 24257 31555 24262 31675
rect 24262 31555 24308 31675
rect 24308 31555 24313 31675
rect 23572 31232 23628 31288
rect 24390 31232 24446 31288
rect 24743 31114 24799 31170
rect 20721 30834 22489 30974
rect 24567 31006 24623 31060
rect 20135 30512 20140 30568
rect 20140 30512 20186 30568
rect 20186 30512 20191 30568
rect 19661 30060 20261 30200
rect 20995 30331 21000 30571
rect 21000 30331 21046 30571
rect 21046 30331 21051 30571
rect 21679 30331 21684 30571
rect 21684 30331 21730 30571
rect 21730 30331 21735 30571
rect 21475 29997 21480 30237
rect 21480 29997 21526 30237
rect 21526 29997 21531 30237
rect 21883 29997 21888 30237
rect 21888 29997 21934 30237
rect 21934 29997 21939 30237
rect 22363 30047 22368 30287
rect 22368 30047 22414 30287
rect 22414 30047 22419 30287
rect 19661 29660 20261 29800
rect 20893 29774 20949 29830
rect 17695 29452 17751 29508
rect 13334 28909 13390 28965
rect 13517 28909 13573 28965
rect 17873 29092 17878 29148
rect 17878 29092 17924 29148
rect 17924 29092 17929 29148
rect 10485 28532 10541 28588
rect 10005 28454 10061 28510
rect 9295 28172 9300 28228
rect 9300 28172 9346 28228
rect 9346 28172 9351 28228
rect 9775 28172 9780 28228
rect 9780 28172 9826 28228
rect 9826 28172 9831 28228
rect 9979 28172 9984 28228
rect 9984 28172 10030 28228
rect 10030 28172 10035 28228
rect 10183 28172 10188 28228
rect 10188 28172 10234 28228
rect 10234 28172 10239 28228
rect 10663 28172 10668 28228
rect 10668 28172 10714 28228
rect 10714 28172 10719 28228
rect 12617 27890 12917 28690
rect 18563 28883 18568 29123
rect 18568 28883 18614 29123
rect 18614 28883 18619 29123
rect 19655 28883 19660 29123
rect 19660 28883 19706 29123
rect 19706 28883 19711 29123
rect 18665 28610 18721 28666
rect 20135 28883 20140 29123
rect 20140 28883 20186 29123
rect 20186 28883 20191 29123
rect 24073 30897 24129 30953
rect 23705 30510 23710 30630
rect 23710 30510 23756 30630
rect 23756 30510 23761 30630
rect 24073 30510 24078 30630
rect 24078 30510 24124 30630
rect 24124 30510 24129 30630
rect 23889 30210 23894 30330
rect 23894 30210 23940 30330
rect 23940 30210 23945 30330
rect 24395 30509 24400 30630
rect 24400 30509 24446 30630
rect 24446 30509 24451 30630
rect 24257 30210 24262 30330
rect 24262 30210 24308 30330
rect 24308 30210 24313 30330
rect 23797 30091 23798 30134
rect 23798 30091 23852 30134
rect 23852 30091 23853 30134
rect 23797 30078 23853 30091
rect 23981 30091 23982 30134
rect 23982 30091 24036 30134
rect 24036 30091 24037 30134
rect 23981 30078 24037 30091
rect 24165 30091 24166 30134
rect 24166 30091 24220 30134
rect 24220 30091 24221 30134
rect 24165 30078 24221 30091
rect 23797 29928 23853 29984
rect 22989 29812 23045 29868
rect 23981 29812 24037 29868
rect 24310 29812 24366 29868
rect 24743 29812 24799 29868
rect 22185 29696 22241 29752
rect 22755 29697 22809 29751
rect 24165 29696 24221 29752
rect 21577 29618 21633 29674
rect 20791 29336 20796 29392
rect 20796 29336 20842 29392
rect 20842 29336 20847 29392
rect 21679 29336 21684 29392
rect 21684 29336 21730 29392
rect 21730 29336 21735 29392
rect 22363 29336 22368 29392
rect 22368 29336 22414 29392
rect 22414 29336 22419 29392
rect 23797 29589 23853 29602
rect 23797 29546 23798 29589
rect 23798 29546 23852 29589
rect 23852 29546 23853 29589
rect 23981 29589 24037 29602
rect 23981 29546 23982 29589
rect 23982 29546 24036 29589
rect 24036 29546 24037 29589
rect 24165 29589 24221 29602
rect 24165 29546 24166 29589
rect 24166 29546 24220 29589
rect 24220 29546 24221 29589
rect 24257 29350 24262 29470
rect 24262 29350 24308 29470
rect 24308 29350 24313 29470
rect 23572 29027 23628 29083
rect 24390 29027 24446 29083
rect 20721 28874 22489 29014
rect 25283 31795 25339 31808
rect 25283 31752 25284 31795
rect 25284 31752 25338 31795
rect 25338 31752 25339 31795
rect 25467 31795 25523 31808
rect 25467 31752 25468 31795
rect 25468 31752 25522 31795
rect 25522 31752 25523 31795
rect 25651 31795 25707 31808
rect 25651 31752 25652 31795
rect 25652 31752 25706 31795
rect 25706 31752 25707 31795
rect 25743 31556 25748 31676
rect 25748 31556 25794 31676
rect 25794 31556 25799 31676
rect 25058 31233 25114 31289
rect 25876 31233 25932 31289
rect 27171 31170 27371 31970
rect 28035 31223 28040 31463
rect 28040 31223 28086 31463
rect 28086 31223 28091 31463
rect 29127 31223 29132 31463
rect 29132 31223 29178 31463
rect 29178 31223 29183 31463
rect 28137 30950 28193 31006
rect 29607 31223 29612 31463
rect 29612 31223 29658 31463
rect 29658 31223 29663 31463
rect 31561 31170 31861 31970
rect 43687 33209 43743 33265
rect 44997 33210 45053 33266
rect 43017 33102 43073 33158
rect 42649 32715 42654 32835
rect 42654 32715 42700 32835
rect 42700 32715 42705 32835
rect 43017 32715 43022 32835
rect 43022 32715 43068 32835
rect 43068 32715 43073 32835
rect 42833 32415 42838 32535
rect 42838 32415 42884 32535
rect 42884 32415 42889 32535
rect 43339 32714 43344 32835
rect 43344 32714 43390 32835
rect 43390 32714 43395 32835
rect 43201 32415 43206 32535
rect 43206 32415 43252 32535
rect 43252 32415 43257 32535
rect 42741 32296 42742 32339
rect 42742 32296 42796 32339
rect 42796 32296 42797 32339
rect 42741 32283 42797 32296
rect 42925 32296 42926 32339
rect 42926 32296 42980 32339
rect 42980 32296 42981 32339
rect 42925 32283 42981 32296
rect 43109 32296 43110 32339
rect 43110 32296 43164 32339
rect 43164 32296 43165 32339
rect 43109 32283 43165 32296
rect 42741 32133 42797 32189
rect 44503 33103 44559 33159
rect 44135 32716 44140 32836
rect 44140 32716 44186 32836
rect 44186 32716 44191 32836
rect 44503 32716 44508 32836
rect 44508 32716 44554 32836
rect 44554 32716 44559 32836
rect 44319 32416 44324 32536
rect 44324 32416 44370 32536
rect 44370 32416 44375 32536
rect 44825 32715 44830 32836
rect 44830 32715 44876 32836
rect 44876 32715 44881 32836
rect 44687 32416 44692 32536
rect 44692 32416 44738 32536
rect 44738 32416 44743 32536
rect 44227 32297 44228 32340
rect 44228 32297 44282 32340
rect 44282 32297 44283 32340
rect 44227 32284 44283 32297
rect 44411 32297 44412 32340
rect 44412 32297 44466 32340
rect 44466 32297 44467 32340
rect 44411 32284 44467 32297
rect 44595 32297 44596 32340
rect 44596 32297 44650 32340
rect 44650 32297 44651 32340
rect 44595 32284 44651 32297
rect 44227 32134 44283 32190
rect 42925 32017 42981 32073
rect 43254 32017 43310 32073
rect 43511 32017 43567 32073
rect 44411 32018 44467 32074
rect 44740 32018 44796 32074
rect 45173 32018 45229 32074
rect 32597 31901 32653 31957
rect 33637 31901 33693 31957
rect 29429 30872 29485 30928
rect 28949 30794 29005 30850
rect 27345 29803 27350 30043
rect 27350 29803 27396 30043
rect 27396 29803 27401 30043
rect 28239 30512 28244 30568
rect 28244 30512 28290 30568
rect 28290 30512 28295 30568
rect 28719 30512 28724 30568
rect 28724 30512 28770 30568
rect 28770 30512 28775 30568
rect 28923 30512 28928 30568
rect 28928 30512 28974 30568
rect 28974 30512 28979 30568
rect 29127 30512 29132 30568
rect 29132 30512 29178 30568
rect 29178 30512 29183 30568
rect 35123 31902 35179 31958
rect 33269 31794 33325 31807
rect 33269 31751 33270 31794
rect 33270 31751 33324 31794
rect 33324 31751 33325 31794
rect 33453 31794 33509 31807
rect 33453 31751 33454 31794
rect 33454 31751 33508 31794
rect 33508 31751 33509 31794
rect 33637 31794 33693 31807
rect 33637 31751 33638 31794
rect 33638 31751 33692 31794
rect 33692 31751 33693 31794
rect 33729 31555 33734 31675
rect 33734 31555 33780 31675
rect 33780 31555 33785 31675
rect 33044 31232 33100 31288
rect 33862 31232 33918 31288
rect 34215 31114 34271 31170
rect 30193 30834 31961 30974
rect 34039 31006 34095 31060
rect 29607 30512 29612 30568
rect 29612 30512 29658 30568
rect 29658 30512 29663 30568
rect 29133 30060 29733 30200
rect 30467 30331 30472 30571
rect 30472 30331 30518 30571
rect 30518 30331 30523 30571
rect 31151 30331 31156 30571
rect 31156 30331 31202 30571
rect 31202 30331 31207 30571
rect 30947 29997 30952 30237
rect 30952 29997 30998 30237
rect 30998 29997 31003 30237
rect 31355 29997 31360 30237
rect 31360 29997 31406 30237
rect 31406 29997 31411 30237
rect 31835 30047 31840 30287
rect 31840 30047 31886 30287
rect 31886 30047 31891 30287
rect 29133 29660 29733 29800
rect 30365 29774 30421 29830
rect 27167 29452 27223 29508
rect 22806 28909 22862 28965
rect 22989 28909 23045 28965
rect 27345 29092 27350 29148
rect 27350 29092 27396 29148
rect 27396 29092 27401 29148
rect 19957 28532 20013 28588
rect 19477 28454 19533 28510
rect 18767 28172 18772 28228
rect 18772 28172 18818 28228
rect 18818 28172 18823 28228
rect 19247 28172 19252 28228
rect 19252 28172 19298 28228
rect 19298 28172 19303 28228
rect 19451 28172 19456 28228
rect 19456 28172 19502 28228
rect 19502 28172 19507 28228
rect 19655 28172 19660 28228
rect 19660 28172 19706 28228
rect 19706 28172 19711 28228
rect 20135 28172 20140 28228
rect 20140 28172 20186 28228
rect 20186 28172 20191 28228
rect 22089 27890 22389 28690
rect 28035 28883 28040 29123
rect 28040 28883 28086 29123
rect 28086 28883 28091 29123
rect 29127 28883 29132 29123
rect 29132 28883 29178 29123
rect 29178 28883 29183 29123
rect 28137 28610 28193 28666
rect 29607 28883 29612 29123
rect 29612 28883 29658 29123
rect 29658 28883 29663 29123
rect 33545 30897 33601 30953
rect 33177 30510 33182 30630
rect 33182 30510 33228 30630
rect 33228 30510 33233 30630
rect 33545 30510 33550 30630
rect 33550 30510 33596 30630
rect 33596 30510 33601 30630
rect 33361 30210 33366 30330
rect 33366 30210 33412 30330
rect 33412 30210 33417 30330
rect 33867 30509 33872 30630
rect 33872 30509 33918 30630
rect 33918 30509 33923 30630
rect 33729 30210 33734 30330
rect 33734 30210 33780 30330
rect 33780 30210 33785 30330
rect 33269 30091 33270 30134
rect 33270 30091 33324 30134
rect 33324 30091 33325 30134
rect 33269 30078 33325 30091
rect 33453 30091 33454 30134
rect 33454 30091 33508 30134
rect 33508 30091 33509 30134
rect 33453 30078 33509 30091
rect 33637 30091 33638 30134
rect 33638 30091 33692 30134
rect 33692 30091 33693 30134
rect 33637 30078 33693 30091
rect 33269 29928 33325 29984
rect 32461 29812 32517 29868
rect 33453 29812 33509 29868
rect 33782 29812 33838 29868
rect 34215 29812 34271 29868
rect 31657 29696 31713 29752
rect 32227 29697 32281 29751
rect 33637 29696 33693 29752
rect 31049 29618 31105 29674
rect 30263 29336 30268 29392
rect 30268 29336 30314 29392
rect 30314 29336 30319 29392
rect 31151 29336 31156 29392
rect 31156 29336 31202 29392
rect 31202 29336 31207 29392
rect 31835 29336 31840 29392
rect 31840 29336 31886 29392
rect 31886 29336 31891 29392
rect 33269 29589 33325 29602
rect 33269 29546 33270 29589
rect 33270 29546 33324 29589
rect 33324 29546 33325 29589
rect 33453 29589 33509 29602
rect 33453 29546 33454 29589
rect 33454 29546 33508 29589
rect 33508 29546 33509 29589
rect 33637 29589 33693 29602
rect 33637 29546 33638 29589
rect 33638 29546 33692 29589
rect 33692 29546 33693 29589
rect 33729 29350 33734 29470
rect 33734 29350 33780 29470
rect 33780 29350 33785 29470
rect 33044 29027 33100 29083
rect 33862 29027 33918 29083
rect 30193 28874 31961 29014
rect 34755 31795 34811 31808
rect 34755 31752 34756 31795
rect 34756 31752 34810 31795
rect 34810 31752 34811 31795
rect 34939 31795 34995 31808
rect 34939 31752 34940 31795
rect 34940 31752 34994 31795
rect 34994 31752 34995 31795
rect 35123 31795 35179 31808
rect 35123 31752 35124 31795
rect 35124 31752 35178 31795
rect 35178 31752 35179 31795
rect 35215 31556 35220 31676
rect 35220 31556 35266 31676
rect 35266 31556 35271 31676
rect 34530 31233 34586 31289
rect 35348 31233 35404 31289
rect 36643 31170 36843 31970
rect 37507 31223 37512 31463
rect 37512 31223 37558 31463
rect 37558 31223 37563 31463
rect 38599 31223 38604 31463
rect 38604 31223 38650 31463
rect 38650 31223 38655 31463
rect 37609 30950 37665 31006
rect 39079 31223 39084 31463
rect 39084 31223 39130 31463
rect 39130 31223 39135 31463
rect 41033 31170 41333 31970
rect 42069 31901 42125 31957
rect 43109 31901 43165 31957
rect 38901 30872 38957 30928
rect 38421 30794 38477 30850
rect 36817 29803 36822 30043
rect 36822 29803 36868 30043
rect 36868 29803 36873 30043
rect 37711 30512 37716 30568
rect 37716 30512 37762 30568
rect 37762 30512 37767 30568
rect 38191 30512 38196 30568
rect 38196 30512 38242 30568
rect 38242 30512 38247 30568
rect 38395 30512 38400 30568
rect 38400 30512 38446 30568
rect 38446 30512 38451 30568
rect 38599 30512 38604 30568
rect 38604 30512 38650 30568
rect 38650 30512 38655 30568
rect 44595 31902 44651 31958
rect 42741 31794 42797 31807
rect 42741 31751 42742 31794
rect 42742 31751 42796 31794
rect 42796 31751 42797 31794
rect 42925 31794 42981 31807
rect 42925 31751 42926 31794
rect 42926 31751 42980 31794
rect 42980 31751 42981 31794
rect 43109 31794 43165 31807
rect 43109 31751 43110 31794
rect 43110 31751 43164 31794
rect 43164 31751 43165 31794
rect 43201 31555 43206 31675
rect 43206 31555 43252 31675
rect 43252 31555 43257 31675
rect 42516 31232 42572 31288
rect 43334 31232 43390 31288
rect 43687 31114 43743 31170
rect 39665 30834 41433 30974
rect 43511 31006 43567 31060
rect 39079 30512 39084 30568
rect 39084 30512 39130 30568
rect 39130 30512 39135 30568
rect 38605 30060 39205 30200
rect 39939 30331 39944 30571
rect 39944 30331 39990 30571
rect 39990 30331 39995 30571
rect 40623 30331 40628 30571
rect 40628 30331 40674 30571
rect 40674 30331 40679 30571
rect 40419 29997 40424 30237
rect 40424 29997 40470 30237
rect 40470 29997 40475 30237
rect 40827 29997 40832 30237
rect 40832 29997 40878 30237
rect 40878 29997 40883 30237
rect 41307 30047 41312 30287
rect 41312 30047 41358 30287
rect 41358 30047 41363 30287
rect 38605 29660 39205 29800
rect 39837 29774 39893 29830
rect 36639 29452 36695 29508
rect 32278 28909 32334 28965
rect 32461 28909 32517 28965
rect 36817 29092 36822 29148
rect 36822 29092 36868 29148
rect 36868 29092 36873 29148
rect 29429 28532 29485 28588
rect 28949 28454 29005 28510
rect 28239 28172 28244 28228
rect 28244 28172 28290 28228
rect 28290 28172 28295 28228
rect 28719 28172 28724 28228
rect 28724 28172 28770 28228
rect 28770 28172 28775 28228
rect 28923 28172 28928 28228
rect 28928 28172 28974 28228
rect 28974 28172 28979 28228
rect 29127 28172 29132 28228
rect 29132 28172 29178 28228
rect 29178 28172 29183 28228
rect 29607 28172 29612 28228
rect 29612 28172 29658 28228
rect 29658 28172 29663 28228
rect 31561 27890 31861 28690
rect 37507 28883 37512 29123
rect 37512 28883 37558 29123
rect 37558 28883 37563 29123
rect 38599 28883 38604 29123
rect 38604 28883 38650 29123
rect 38650 28883 38655 29123
rect 37609 28610 37665 28666
rect 39079 28883 39084 29123
rect 39084 28883 39130 29123
rect 39130 28883 39135 29123
rect 43017 30897 43073 30953
rect 42649 30510 42654 30630
rect 42654 30510 42700 30630
rect 42700 30510 42705 30630
rect 43017 30510 43022 30630
rect 43022 30510 43068 30630
rect 43068 30510 43073 30630
rect 42833 30210 42838 30330
rect 42838 30210 42884 30330
rect 42884 30210 42889 30330
rect 43339 30509 43344 30630
rect 43344 30509 43390 30630
rect 43390 30509 43395 30630
rect 43201 30210 43206 30330
rect 43206 30210 43252 30330
rect 43252 30210 43257 30330
rect 42741 30091 42742 30134
rect 42742 30091 42796 30134
rect 42796 30091 42797 30134
rect 42741 30078 42797 30091
rect 42925 30091 42926 30134
rect 42926 30091 42980 30134
rect 42980 30091 42981 30134
rect 42925 30078 42981 30091
rect 43109 30091 43110 30134
rect 43110 30091 43164 30134
rect 43164 30091 43165 30134
rect 43109 30078 43165 30091
rect 42741 29928 42797 29984
rect 41933 29812 41989 29868
rect 42925 29812 42981 29868
rect 43254 29812 43310 29868
rect 43687 29812 43743 29868
rect 41129 29696 41185 29752
rect 41699 29697 41753 29751
rect 43109 29696 43165 29752
rect 40521 29618 40577 29674
rect 39735 29336 39740 29392
rect 39740 29336 39786 29392
rect 39786 29336 39791 29392
rect 40623 29336 40628 29392
rect 40628 29336 40674 29392
rect 40674 29336 40679 29392
rect 41307 29336 41312 29392
rect 41312 29336 41358 29392
rect 41358 29336 41363 29392
rect 42741 29589 42797 29602
rect 42741 29546 42742 29589
rect 42742 29546 42796 29589
rect 42796 29546 42797 29589
rect 42925 29589 42981 29602
rect 42925 29546 42926 29589
rect 42926 29546 42980 29589
rect 42980 29546 42981 29589
rect 43109 29589 43165 29602
rect 43109 29546 43110 29589
rect 43110 29546 43164 29589
rect 43164 29546 43165 29589
rect 43201 29350 43206 29470
rect 43206 29350 43252 29470
rect 43252 29350 43257 29470
rect 42516 29027 42572 29083
rect 43334 29027 43390 29083
rect 39665 28874 41433 29014
rect 44227 31795 44283 31808
rect 44227 31752 44228 31795
rect 44228 31752 44282 31795
rect 44282 31752 44283 31795
rect 44411 31795 44467 31808
rect 44411 31752 44412 31795
rect 44412 31752 44466 31795
rect 44466 31752 44467 31795
rect 44595 31795 44651 31808
rect 44595 31752 44596 31795
rect 44596 31752 44650 31795
rect 44650 31752 44651 31795
rect 44687 31556 44692 31676
rect 44692 31556 44738 31676
rect 44738 31556 44743 31676
rect 44002 31233 44058 31289
rect 44820 31233 44876 31289
rect 41750 28909 41806 28965
rect 41933 28909 41989 28965
rect 38901 28532 38957 28588
rect 38421 28454 38477 28510
rect 37711 28172 37716 28228
rect 37716 28172 37762 28228
rect 37762 28172 37767 28228
rect 38191 28172 38196 28228
rect 38196 28172 38242 28228
rect 38242 28172 38247 28228
rect 38395 28172 38400 28228
rect 38400 28172 38446 28228
rect 38446 28172 38451 28228
rect 38599 28172 38604 28228
rect 38604 28172 38650 28228
rect 38650 28172 38655 28228
rect 39079 28172 39084 28228
rect 39084 28172 39130 28228
rect 39130 28172 39135 28228
rect 41033 27890 41333 28690
rect -12434 27521 -12378 27577
rect -12256 27161 -12251 27217
rect -12251 27161 -12205 27217
rect -12205 27161 -12200 27217
rect -737 26018 -681 26074
rect 7111 26018 7167 26074
rect 3305 25842 3361 25898
rect 11153 25842 11209 25898
rect -8875 25666 -8819 25722
rect -1027 25666 -971 25722
rect 7347 25666 7403 25722
rect 15195 25666 15251 25722
rect -4779 25490 -4723 25546
rect 3069 25490 3125 25546
rect 11389 25490 11445 25546
rect 19237 25490 19293 25546
rect -7601 25209 -7545 25265
rect -7969 24822 -7964 24942
rect -7964 24822 -7918 24942
rect -7918 24822 -7913 24942
rect -7601 24822 -7596 24942
rect -7596 24822 -7550 24942
rect -7550 24822 -7545 24942
rect -7785 24522 -7780 24642
rect -7780 24522 -7734 24642
rect -7734 24522 -7729 24642
rect -7279 24821 -7274 24942
rect -7274 24821 -7228 24942
rect -7228 24821 -7223 24942
rect -7417 24522 -7412 24642
rect -7412 24522 -7366 24642
rect -7366 24522 -7361 24642
rect -7877 24403 -7876 24446
rect -7876 24403 -7822 24446
rect -7822 24403 -7821 24446
rect -7877 24390 -7821 24403
rect -7693 24403 -7692 24446
rect -7692 24403 -7638 24446
rect -7638 24403 -7637 24446
rect -7693 24390 -7637 24403
rect -7509 24403 -7508 24446
rect -7508 24403 -7454 24446
rect -7454 24403 -7453 24446
rect -7509 24390 -7453 24403
rect -9229 24240 -9173 24296
rect -7877 24240 -7821 24296
rect -8549 24124 -8493 24180
rect -7693 24124 -7637 24180
rect -7364 24124 -7308 24180
rect -7107 24124 -7051 24180
rect -7509 24008 -7453 24064
rect -7877 23901 -7821 23914
rect -7877 23858 -7876 23901
rect -7876 23858 -7822 23901
rect -7822 23858 -7821 23901
rect -7693 23901 -7637 23914
rect -7693 23858 -7692 23901
rect -7692 23858 -7638 23901
rect -7638 23858 -7637 23901
rect -7509 23901 -7453 23914
rect -7509 23858 -7508 23901
rect -7508 23858 -7454 23901
rect -7454 23858 -7453 23901
rect -7417 23662 -7412 23782
rect -7412 23662 -7366 23782
rect -7366 23662 -7361 23782
rect -8102 23339 -8046 23395
rect -7284 23339 -7228 23395
rect -6931 23221 -6875 23277
rect -7107 23113 -7051 23167
rect -7601 23004 -7545 23060
rect -7969 22617 -7964 22737
rect -7964 22617 -7918 22737
rect -7918 22617 -7913 22737
rect -7601 22617 -7596 22737
rect -7596 22617 -7550 22737
rect -7550 22617 -7545 22737
rect -7785 22317 -7780 22437
rect -7780 22317 -7734 22437
rect -7734 22317 -7729 22437
rect -7279 22616 -7274 22737
rect -7274 22616 -7228 22737
rect -7228 22616 -7223 22737
rect -7417 22317 -7412 22437
rect -7412 22317 -7366 22437
rect -7366 22317 -7361 22437
rect -7877 22198 -7876 22241
rect -7876 22198 -7822 22241
rect -7822 22198 -7821 22241
rect -7877 22185 -7821 22198
rect -7693 22198 -7692 22241
rect -7692 22198 -7638 22241
rect -7638 22198 -7637 22241
rect -7693 22185 -7637 22198
rect -7509 22198 -7508 22241
rect -7508 22198 -7454 22241
rect -7454 22198 -7453 22241
rect -7509 22185 -7453 22198
rect -7877 22035 -7821 22091
rect -3559 25206 -3503 25262
rect -3927 24819 -3922 24939
rect -3922 24819 -3876 24939
rect -3876 24819 -3871 24939
rect -3559 24819 -3554 24939
rect -3554 24819 -3508 24939
rect -3508 24819 -3503 24939
rect -3743 24519 -3738 24639
rect -3738 24519 -3692 24639
rect -3692 24519 -3687 24639
rect -3237 24818 -3232 24939
rect -3232 24818 -3186 24939
rect -3186 24818 -3181 24939
rect -3375 24519 -3370 24639
rect -3370 24519 -3324 24639
rect -3324 24519 -3319 24639
rect -3835 24400 -3834 24443
rect -3834 24400 -3780 24443
rect -3780 24400 -3779 24443
rect -3835 24387 -3779 24400
rect -3651 24400 -3650 24443
rect -3650 24400 -3596 24443
rect -3596 24400 -3595 24443
rect -3651 24387 -3595 24400
rect -3467 24400 -3466 24443
rect -3466 24400 -3412 24443
rect -3412 24400 -3411 24443
rect -3467 24387 -3411 24400
rect -5217 24237 -5161 24293
rect -3835 24237 -3779 24293
rect -4507 24121 -4451 24177
rect -3651 24121 -3595 24177
rect -3322 24121 -3266 24177
rect -3065 24121 -3009 24177
rect -3467 24005 -3411 24061
rect -3835 23898 -3779 23911
rect -3835 23855 -3834 23898
rect -3834 23855 -3780 23898
rect -3780 23855 -3779 23898
rect -3651 23898 -3595 23911
rect -3651 23855 -3650 23898
rect -3650 23855 -3596 23898
rect -3596 23855 -3595 23898
rect -3467 23898 -3411 23911
rect -3467 23855 -3466 23898
rect -3466 23855 -3412 23898
rect -3412 23855 -3411 23898
rect -3375 23659 -3370 23779
rect -3370 23659 -3324 23779
rect -3324 23659 -3319 23779
rect -4060 23336 -4004 23392
rect -3242 23336 -3186 23392
rect -2889 23218 -2833 23274
rect -3065 23110 -3009 23164
rect -6115 23004 -6059 23060
rect -6483 22617 -6478 22737
rect -6478 22617 -6432 22737
rect -6432 22617 -6427 22737
rect -6115 22617 -6110 22737
rect -6110 22617 -6064 22737
rect -6064 22617 -6059 22737
rect -6299 22317 -6294 22437
rect -6294 22317 -6248 22437
rect -6248 22317 -6243 22437
rect -5793 22616 -5788 22737
rect -5788 22616 -5742 22737
rect -5742 22616 -5737 22737
rect -5931 22317 -5926 22437
rect -5926 22317 -5880 22437
rect -5880 22317 -5875 22437
rect -6391 22198 -6390 22241
rect -6390 22198 -6336 22241
rect -6336 22198 -6335 22241
rect -6391 22185 -6335 22198
rect -6207 22198 -6206 22241
rect -6206 22198 -6152 22241
rect -6152 22198 -6151 22241
rect -6207 22185 -6151 22198
rect -6023 22198 -6022 22241
rect -6022 22198 -5968 22241
rect -5968 22198 -5967 22241
rect -6023 22185 -5967 22198
rect -6391 22035 -6335 22091
rect -3559 23001 -3503 23057
rect -3927 22614 -3922 22734
rect -3922 22614 -3876 22734
rect -3876 22614 -3871 22734
rect -3559 22614 -3554 22734
rect -3554 22614 -3508 22734
rect -3508 22614 -3503 22734
rect -3743 22314 -3738 22434
rect -3738 22314 -3692 22434
rect -3692 22314 -3687 22434
rect -3237 22613 -3232 22734
rect -3232 22613 -3186 22734
rect -3186 22613 -3181 22734
rect -3375 22314 -3370 22434
rect -3370 22314 -3324 22434
rect -3324 22314 -3319 22434
rect -3835 22195 -3834 22238
rect -3834 22195 -3780 22238
rect -3780 22195 -3779 22238
rect -3835 22182 -3779 22195
rect -3651 22195 -3650 22238
rect -3650 22195 -3596 22238
rect -3596 22195 -3595 22238
rect -3651 22182 -3595 22195
rect -3467 22195 -3466 22238
rect -3466 22195 -3412 22238
rect -3412 22195 -3411 22238
rect -3467 22182 -3411 22195
rect -3835 22032 -3779 22088
rect 483 25206 539 25262
rect 115 24819 120 24939
rect 120 24819 166 24939
rect 166 24819 171 24939
rect 483 24819 488 24939
rect 488 24819 534 24939
rect 534 24819 539 24939
rect 299 24519 304 24639
rect 304 24519 350 24639
rect 350 24519 355 24639
rect 805 24818 810 24939
rect 810 24818 856 24939
rect 856 24818 861 24939
rect 667 24519 672 24639
rect 672 24519 718 24639
rect 718 24519 723 24639
rect 207 24400 208 24443
rect 208 24400 262 24443
rect 262 24400 263 24443
rect 207 24387 263 24400
rect 391 24400 392 24443
rect 392 24400 446 24443
rect 446 24400 447 24443
rect 391 24387 447 24400
rect 575 24400 576 24443
rect 576 24400 630 24443
rect 630 24400 631 24443
rect 575 24387 631 24400
rect -1175 24237 -1119 24293
rect 207 24237 263 24293
rect -465 24121 -409 24177
rect 391 24121 447 24177
rect 720 24121 776 24177
rect 977 24121 1033 24177
rect 575 24005 631 24061
rect 207 23898 263 23911
rect 207 23855 208 23898
rect 208 23855 262 23898
rect 262 23855 263 23898
rect 391 23898 447 23911
rect 391 23855 392 23898
rect 392 23855 446 23898
rect 446 23855 447 23898
rect 575 23898 631 23911
rect 575 23855 576 23898
rect 576 23855 630 23898
rect 630 23855 631 23898
rect 667 23659 672 23779
rect 672 23659 718 23779
rect 718 23659 723 23779
rect -18 23336 38 23392
rect 800 23336 856 23392
rect 1153 23218 1209 23274
rect 977 23110 1033 23164
rect -2073 23001 -2017 23057
rect -2441 22614 -2436 22734
rect -2436 22614 -2390 22734
rect -2390 22614 -2385 22734
rect -2073 22614 -2068 22734
rect -2068 22614 -2022 22734
rect -2022 22614 -2017 22734
rect -2257 22314 -2252 22434
rect -2252 22314 -2206 22434
rect -2206 22314 -2201 22434
rect -1751 22613 -1746 22734
rect -1746 22613 -1700 22734
rect -1700 22613 -1695 22734
rect -1889 22314 -1884 22434
rect -1884 22314 -1838 22434
rect -1838 22314 -1833 22434
rect -2349 22195 -2348 22238
rect -2348 22195 -2294 22238
rect -2294 22195 -2293 22238
rect -2349 22182 -2293 22195
rect -2165 22195 -2164 22238
rect -2164 22195 -2110 22238
rect -2110 22195 -2109 22238
rect -2165 22182 -2109 22195
rect -1981 22195 -1980 22238
rect -1980 22195 -1926 22238
rect -1926 22195 -1925 22238
rect -1981 22182 -1925 22195
rect -2349 22032 -2293 22088
rect 483 23001 539 23057
rect 115 22614 120 22734
rect 120 22614 166 22734
rect 166 22614 171 22734
rect 483 22614 488 22734
rect 488 22614 534 22734
rect 534 22614 539 22734
rect 299 22314 304 22434
rect 304 22314 350 22434
rect 350 22314 355 22434
rect 805 22613 810 22734
rect 810 22613 856 22734
rect 856 22613 861 22734
rect 667 22314 672 22434
rect 672 22314 718 22434
rect 718 22314 723 22434
rect 207 22195 208 22238
rect 208 22195 262 22238
rect 262 22195 263 22238
rect 207 22182 263 22195
rect 391 22195 392 22238
rect 392 22195 446 22238
rect 446 22195 447 22238
rect 391 22182 447 22195
rect 575 22195 576 22238
rect 576 22195 630 22238
rect 630 22195 631 22238
rect 575 22182 631 22195
rect 207 22032 263 22088
rect 4525 25206 4581 25262
rect 4157 24819 4162 24939
rect 4162 24819 4208 24939
rect 4208 24819 4213 24939
rect 4525 24819 4530 24939
rect 4530 24819 4576 24939
rect 4576 24819 4581 24939
rect 4341 24519 4346 24639
rect 4346 24519 4392 24639
rect 4392 24519 4397 24639
rect 4847 24818 4852 24939
rect 4852 24818 4898 24939
rect 4898 24818 4903 24939
rect 4709 24519 4714 24639
rect 4714 24519 4760 24639
rect 4760 24519 4765 24639
rect 4249 24400 4250 24443
rect 4250 24400 4304 24443
rect 4304 24400 4305 24443
rect 4249 24387 4305 24400
rect 4433 24400 4434 24443
rect 4434 24400 4488 24443
rect 4488 24400 4489 24443
rect 4433 24387 4489 24400
rect 4617 24400 4618 24443
rect 4618 24400 4672 24443
rect 4672 24400 4673 24443
rect 4617 24387 4673 24400
rect 2867 24237 2923 24293
rect 4249 24237 4305 24293
rect 3577 24121 3633 24177
rect 4433 24121 4489 24177
rect 4762 24121 4818 24177
rect 5019 24121 5075 24177
rect 4617 24005 4673 24061
rect 4249 23898 4305 23911
rect 4249 23855 4250 23898
rect 4250 23855 4304 23898
rect 4304 23855 4305 23898
rect 4433 23898 4489 23911
rect 4433 23855 4434 23898
rect 4434 23855 4488 23898
rect 4488 23855 4489 23898
rect 4617 23898 4673 23911
rect 4617 23855 4618 23898
rect 4618 23855 4672 23898
rect 4672 23855 4673 23898
rect 4709 23659 4714 23779
rect 4714 23659 4760 23779
rect 4760 23659 4765 23779
rect 4024 23336 4080 23392
rect 4842 23336 4898 23392
rect 5195 23218 5251 23274
rect 5019 23110 5075 23164
rect 1969 23001 2025 23057
rect 1601 22614 1606 22734
rect 1606 22614 1652 22734
rect 1652 22614 1657 22734
rect 1969 22614 1974 22734
rect 1974 22614 2020 22734
rect 2020 22614 2025 22734
rect 1785 22314 1790 22434
rect 1790 22314 1836 22434
rect 1836 22314 1841 22434
rect 2291 22613 2296 22734
rect 2296 22613 2342 22734
rect 2342 22613 2347 22734
rect 2153 22314 2158 22434
rect 2158 22314 2204 22434
rect 2204 22314 2209 22434
rect 1693 22195 1694 22238
rect 1694 22195 1748 22238
rect 1748 22195 1749 22238
rect 1693 22182 1749 22195
rect 1877 22195 1878 22238
rect 1878 22195 1932 22238
rect 1932 22195 1933 22238
rect 1877 22182 1933 22195
rect 2061 22195 2062 22238
rect 2062 22195 2116 22238
rect 2116 22195 2117 22238
rect 2061 22182 2117 22195
rect 1693 22032 1749 22088
rect 4525 23001 4581 23057
rect 4157 22614 4162 22734
rect 4162 22614 4208 22734
rect 4208 22614 4213 22734
rect 4525 22614 4530 22734
rect 4530 22614 4576 22734
rect 4576 22614 4581 22734
rect 4341 22314 4346 22434
rect 4346 22314 4392 22434
rect 4392 22314 4397 22434
rect 4847 22613 4852 22734
rect 4852 22613 4898 22734
rect 4898 22613 4903 22734
rect 4709 22314 4714 22434
rect 4714 22314 4760 22434
rect 4760 22314 4765 22434
rect 4249 22195 4250 22238
rect 4250 22195 4304 22238
rect 4304 22195 4305 22238
rect 4249 22182 4305 22195
rect 4433 22195 4434 22238
rect 4434 22195 4488 22238
rect 4488 22195 4489 22238
rect 4433 22182 4489 22195
rect 4617 22195 4618 22238
rect 4618 22195 4672 22238
rect 4672 22195 4673 22238
rect 4617 22182 4673 22195
rect 4249 22032 4305 22088
rect 8567 25206 8623 25262
rect 8199 24819 8204 24939
rect 8204 24819 8250 24939
rect 8250 24819 8255 24939
rect 8567 24819 8572 24939
rect 8572 24819 8618 24939
rect 8618 24819 8623 24939
rect 8383 24519 8388 24639
rect 8388 24519 8434 24639
rect 8434 24519 8439 24639
rect 8889 24818 8894 24939
rect 8894 24818 8940 24939
rect 8940 24818 8945 24939
rect 8751 24519 8756 24639
rect 8756 24519 8802 24639
rect 8802 24519 8807 24639
rect 8291 24400 8292 24443
rect 8292 24400 8346 24443
rect 8346 24400 8347 24443
rect 8291 24387 8347 24400
rect 8475 24400 8476 24443
rect 8476 24400 8530 24443
rect 8530 24400 8531 24443
rect 8475 24387 8531 24400
rect 8659 24400 8660 24443
rect 8660 24400 8714 24443
rect 8714 24400 8715 24443
rect 8659 24387 8715 24400
rect 6909 24237 6965 24293
rect 8291 24237 8347 24293
rect 7619 24121 7675 24177
rect 8475 24121 8531 24177
rect 8804 24121 8860 24177
rect 9061 24121 9117 24177
rect 8659 24005 8715 24061
rect 8291 23898 8347 23911
rect 8291 23855 8292 23898
rect 8292 23855 8346 23898
rect 8346 23855 8347 23898
rect 8475 23898 8531 23911
rect 8475 23855 8476 23898
rect 8476 23855 8530 23898
rect 8530 23855 8531 23898
rect 8659 23898 8715 23911
rect 8659 23855 8660 23898
rect 8660 23855 8714 23898
rect 8714 23855 8715 23898
rect 8751 23659 8756 23779
rect 8756 23659 8802 23779
rect 8802 23659 8807 23779
rect 8066 23336 8122 23392
rect 8884 23336 8940 23392
rect 9237 23218 9293 23274
rect 9061 23110 9117 23164
rect 6011 23001 6067 23057
rect 5643 22614 5648 22734
rect 5648 22614 5694 22734
rect 5694 22614 5699 22734
rect 6011 22614 6016 22734
rect 6016 22614 6062 22734
rect 6062 22614 6067 22734
rect 5827 22314 5832 22434
rect 5832 22314 5878 22434
rect 5878 22314 5883 22434
rect 6333 22613 6338 22734
rect 6338 22613 6384 22734
rect 6384 22613 6389 22734
rect 6195 22314 6200 22434
rect 6200 22314 6246 22434
rect 6246 22314 6251 22434
rect 5735 22195 5736 22238
rect 5736 22195 5790 22238
rect 5790 22195 5791 22238
rect 5735 22182 5791 22195
rect 5919 22195 5920 22238
rect 5920 22195 5974 22238
rect 5974 22195 5975 22238
rect 5919 22182 5975 22195
rect 6103 22195 6104 22238
rect 6104 22195 6158 22238
rect 6158 22195 6159 22238
rect 6103 22182 6159 22195
rect 5735 22032 5791 22088
rect 8567 23001 8623 23057
rect 8199 22614 8204 22734
rect 8204 22614 8250 22734
rect 8250 22614 8255 22734
rect 8567 22614 8572 22734
rect 8572 22614 8618 22734
rect 8618 22614 8623 22734
rect 8383 22314 8388 22434
rect 8388 22314 8434 22434
rect 8434 22314 8439 22434
rect 8889 22613 8894 22734
rect 8894 22613 8940 22734
rect 8940 22613 8945 22734
rect 8751 22314 8756 22434
rect 8756 22314 8802 22434
rect 8802 22314 8807 22434
rect 8291 22195 8292 22238
rect 8292 22195 8346 22238
rect 8346 22195 8347 22238
rect 8291 22182 8347 22195
rect 8475 22195 8476 22238
rect 8476 22195 8530 22238
rect 8530 22195 8531 22238
rect 8475 22182 8531 22195
rect 8659 22195 8660 22238
rect 8660 22195 8714 22238
rect 8714 22195 8715 22238
rect 8659 22182 8715 22195
rect 8291 22032 8347 22088
rect 12609 25206 12665 25262
rect 12241 24819 12246 24939
rect 12246 24819 12292 24939
rect 12292 24819 12297 24939
rect 12609 24819 12614 24939
rect 12614 24819 12660 24939
rect 12660 24819 12665 24939
rect 12425 24519 12430 24639
rect 12430 24519 12476 24639
rect 12476 24519 12481 24639
rect 12931 24818 12936 24939
rect 12936 24818 12982 24939
rect 12982 24818 12987 24939
rect 12793 24519 12798 24639
rect 12798 24519 12844 24639
rect 12844 24519 12849 24639
rect 12333 24400 12334 24443
rect 12334 24400 12388 24443
rect 12388 24400 12389 24443
rect 12333 24387 12389 24400
rect 12517 24400 12518 24443
rect 12518 24400 12572 24443
rect 12572 24400 12573 24443
rect 12517 24387 12573 24400
rect 12701 24400 12702 24443
rect 12702 24400 12756 24443
rect 12756 24400 12757 24443
rect 12701 24387 12757 24400
rect 10951 24237 11007 24293
rect 12333 24237 12389 24293
rect 11661 24121 11717 24177
rect 12517 24121 12573 24177
rect 12846 24121 12902 24177
rect 13103 24121 13159 24177
rect 12701 24005 12757 24061
rect 12333 23898 12389 23911
rect 12333 23855 12334 23898
rect 12334 23855 12388 23898
rect 12388 23855 12389 23898
rect 12517 23898 12573 23911
rect 12517 23855 12518 23898
rect 12518 23855 12572 23898
rect 12572 23855 12573 23898
rect 12701 23898 12757 23911
rect 12701 23855 12702 23898
rect 12702 23855 12756 23898
rect 12756 23855 12757 23898
rect 12793 23659 12798 23779
rect 12798 23659 12844 23779
rect 12844 23659 12849 23779
rect 12108 23336 12164 23392
rect 12926 23336 12982 23392
rect 13279 23218 13335 23274
rect 13103 23110 13159 23164
rect 10053 23001 10109 23057
rect 9685 22614 9690 22734
rect 9690 22614 9736 22734
rect 9736 22614 9741 22734
rect 10053 22614 10058 22734
rect 10058 22614 10104 22734
rect 10104 22614 10109 22734
rect 9869 22314 9874 22434
rect 9874 22314 9920 22434
rect 9920 22314 9925 22434
rect 10375 22613 10380 22734
rect 10380 22613 10426 22734
rect 10426 22613 10431 22734
rect 10237 22314 10242 22434
rect 10242 22314 10288 22434
rect 10288 22314 10293 22434
rect 9777 22195 9778 22238
rect 9778 22195 9832 22238
rect 9832 22195 9833 22238
rect 9777 22182 9833 22195
rect 9961 22195 9962 22238
rect 9962 22195 10016 22238
rect 10016 22195 10017 22238
rect 9961 22182 10017 22195
rect 10145 22195 10146 22238
rect 10146 22195 10200 22238
rect 10200 22195 10201 22238
rect 10145 22182 10201 22195
rect 9777 22032 9833 22088
rect 12609 23001 12665 23057
rect 12241 22614 12246 22734
rect 12246 22614 12292 22734
rect 12292 22614 12297 22734
rect 12609 22614 12614 22734
rect 12614 22614 12660 22734
rect 12660 22614 12665 22734
rect 12425 22314 12430 22434
rect 12430 22314 12476 22434
rect 12476 22314 12481 22434
rect 12931 22613 12936 22734
rect 12936 22613 12982 22734
rect 12982 22613 12987 22734
rect 12793 22314 12798 22434
rect 12798 22314 12844 22434
rect 12844 22314 12849 22434
rect 12333 22195 12334 22238
rect 12334 22195 12388 22238
rect 12388 22195 12389 22238
rect 12333 22182 12389 22195
rect 12517 22195 12518 22238
rect 12518 22195 12572 22238
rect 12572 22195 12573 22238
rect 12517 22182 12573 22195
rect 12701 22195 12702 22238
rect 12702 22195 12756 22238
rect 12756 22195 12757 22238
rect 12701 22182 12757 22195
rect 12333 22032 12389 22088
rect 16651 25206 16707 25262
rect 16283 24819 16288 24939
rect 16288 24819 16334 24939
rect 16334 24819 16339 24939
rect 16651 24819 16656 24939
rect 16656 24819 16702 24939
rect 16702 24819 16707 24939
rect 16467 24519 16472 24639
rect 16472 24519 16518 24639
rect 16518 24519 16523 24639
rect 16973 24818 16978 24939
rect 16978 24818 17024 24939
rect 17024 24818 17029 24939
rect 16835 24519 16840 24639
rect 16840 24519 16886 24639
rect 16886 24519 16891 24639
rect 16375 24400 16376 24443
rect 16376 24400 16430 24443
rect 16430 24400 16431 24443
rect 16375 24387 16431 24400
rect 16559 24400 16560 24443
rect 16560 24400 16614 24443
rect 16614 24400 16615 24443
rect 16559 24387 16615 24400
rect 16743 24400 16744 24443
rect 16744 24400 16798 24443
rect 16798 24400 16799 24443
rect 16743 24387 16799 24400
rect 14993 24237 15049 24293
rect 16375 24237 16431 24293
rect 15703 24121 15759 24177
rect 16559 24121 16615 24177
rect 16888 24121 16944 24177
rect 17145 24121 17201 24177
rect 16743 24005 16799 24061
rect 16375 23898 16431 23911
rect 16375 23855 16376 23898
rect 16376 23855 16430 23898
rect 16430 23855 16431 23898
rect 16559 23898 16615 23911
rect 16559 23855 16560 23898
rect 16560 23855 16614 23898
rect 16614 23855 16615 23898
rect 16743 23898 16799 23911
rect 16743 23855 16744 23898
rect 16744 23855 16798 23898
rect 16798 23855 16799 23898
rect 16835 23659 16840 23779
rect 16840 23659 16886 23779
rect 16886 23659 16891 23779
rect 16150 23336 16206 23392
rect 16968 23336 17024 23392
rect 17321 23218 17377 23274
rect 17145 23110 17201 23164
rect 14095 23001 14151 23057
rect 13727 22614 13732 22734
rect 13732 22614 13778 22734
rect 13778 22614 13783 22734
rect 14095 22614 14100 22734
rect 14100 22614 14146 22734
rect 14146 22614 14151 22734
rect 13911 22314 13916 22434
rect 13916 22314 13962 22434
rect 13962 22314 13967 22434
rect 14417 22613 14422 22734
rect 14422 22613 14468 22734
rect 14468 22613 14473 22734
rect 14279 22314 14284 22434
rect 14284 22314 14330 22434
rect 14330 22314 14335 22434
rect 13819 22195 13820 22238
rect 13820 22195 13874 22238
rect 13874 22195 13875 22238
rect 13819 22182 13875 22195
rect 14003 22195 14004 22238
rect 14004 22195 14058 22238
rect 14058 22195 14059 22238
rect 14003 22182 14059 22195
rect 14187 22195 14188 22238
rect 14188 22195 14242 22238
rect 14242 22195 14243 22238
rect 14187 22182 14243 22195
rect 13819 22032 13875 22088
rect 16651 23001 16707 23057
rect 16283 22614 16288 22734
rect 16288 22614 16334 22734
rect 16334 22614 16339 22734
rect 16651 22614 16656 22734
rect 16656 22614 16702 22734
rect 16702 22614 16707 22734
rect 16467 22314 16472 22434
rect 16472 22314 16518 22434
rect 16518 22314 16523 22434
rect 16973 22613 16978 22734
rect 16978 22613 17024 22734
rect 17024 22613 17029 22734
rect 16835 22314 16840 22434
rect 16840 22314 16886 22434
rect 16886 22314 16891 22434
rect 16375 22195 16376 22238
rect 16376 22195 16430 22238
rect 16430 22195 16431 22238
rect 16375 22182 16431 22195
rect 16559 22195 16560 22238
rect 16560 22195 16614 22238
rect 16614 22195 16615 22238
rect 16559 22182 16615 22195
rect 16743 22195 16744 22238
rect 16744 22195 16798 22238
rect 16798 22195 16799 22238
rect 16743 22182 16799 22195
rect 16375 22032 16431 22088
rect 18137 23001 18193 23057
rect 17769 22614 17774 22734
rect 17774 22614 17820 22734
rect 17820 22614 17825 22734
rect 18137 22614 18142 22734
rect 18142 22614 18188 22734
rect 18188 22614 18193 22734
rect 17953 22314 17958 22434
rect 17958 22314 18004 22434
rect 18004 22314 18009 22434
rect 18459 22613 18464 22734
rect 18464 22613 18510 22734
rect 18510 22613 18515 22734
rect 18321 22314 18326 22434
rect 18326 22314 18372 22434
rect 18372 22314 18377 22434
rect 17861 22195 17862 22238
rect 17862 22195 17916 22238
rect 17916 22195 17917 22238
rect 17861 22182 17917 22195
rect 18045 22195 18046 22238
rect 18046 22195 18100 22238
rect 18100 22195 18101 22238
rect 18045 22182 18101 22195
rect 18229 22195 18230 22238
rect 18230 22195 18284 22238
rect 18284 22195 18285 22238
rect 18229 22182 18285 22195
rect 17861 22032 17917 22088
rect -8685 21919 -8629 21975
rect -7693 21919 -7637 21975
rect -7364 21919 -7308 21975
rect -6931 21919 -6875 21975
rect -6207 21919 -6151 21975
rect -5878 21919 -5822 21975
rect -5621 21919 -5565 21975
rect -5081 21919 -5025 21975
rect -4643 21916 -4587 21972
rect -3651 21916 -3595 21972
rect -3322 21916 -3266 21972
rect -2889 21916 -2833 21972
rect -2165 21916 -2109 21972
rect -1836 21916 -1780 21972
rect -1579 21916 -1523 21972
rect -1027 21916 -971 21972
rect -601 21916 -545 21972
rect 391 21916 447 21972
rect 720 21916 776 21972
rect 1153 21916 1209 21972
rect 1877 21916 1933 21972
rect 2206 21916 2262 21972
rect 2463 21916 2519 21972
rect 3069 21916 3125 21972
rect 3441 21916 3497 21972
rect 4433 21916 4489 21972
rect 4762 21916 4818 21972
rect 5195 21916 5251 21972
rect 5919 21916 5975 21972
rect 6248 21916 6304 21972
rect 6505 21916 6561 21972
rect 7111 21916 7167 21972
rect 7483 21916 7539 21972
rect 8475 21916 8531 21972
rect 8804 21916 8860 21972
rect 9237 21916 9293 21972
rect 9961 21916 10017 21972
rect 10290 21916 10346 21972
rect 10547 21916 10603 21972
rect 11153 21916 11209 21972
rect 11525 21916 11581 21972
rect 12517 21916 12573 21972
rect 12846 21916 12902 21972
rect 13279 21916 13335 21972
rect 14003 21916 14059 21972
rect 14332 21916 14388 21972
rect 14589 21916 14645 21972
rect 15195 21916 15251 21972
rect 15567 21916 15623 21972
rect 16559 21916 16615 21972
rect 16888 21916 16944 21972
rect 17321 21916 17377 21972
rect 18045 21916 18101 21972
rect 18374 21916 18430 21972
rect 18631 21916 18687 21972
rect 19237 21916 19293 21972
rect -7509 21803 -7453 21859
rect -6023 21803 -5967 21859
rect -7877 21696 -7821 21709
rect -7877 21653 -7876 21696
rect -7876 21653 -7822 21696
rect -7822 21653 -7821 21696
rect -7693 21696 -7637 21709
rect -7693 21653 -7692 21696
rect -7692 21653 -7638 21696
rect -7638 21653 -7637 21696
rect -7509 21696 -7453 21709
rect -7509 21653 -7508 21696
rect -7508 21653 -7454 21696
rect -7454 21653 -7453 21696
rect -7417 21457 -7412 21577
rect -7412 21457 -7366 21577
rect -7366 21457 -7361 21577
rect -8102 21134 -8046 21190
rect -7284 21134 -7228 21190
rect -8875 21017 -8819 21073
rect -3467 21800 -3411 21856
rect -6391 21696 -6335 21709
rect -6391 21653 -6390 21696
rect -6390 21653 -6336 21696
rect -6336 21653 -6335 21696
rect -6207 21696 -6151 21709
rect -6207 21653 -6206 21696
rect -6206 21653 -6152 21696
rect -6152 21653 -6151 21696
rect -6023 21696 -5967 21709
rect -6023 21653 -6022 21696
rect -6022 21653 -5968 21696
rect -5968 21653 -5967 21696
rect -5931 21457 -5926 21577
rect -5926 21457 -5880 21577
rect -5880 21457 -5875 21577
rect -6616 21134 -6560 21190
rect -5798 21134 -5742 21190
rect -5445 21017 -5389 21073
rect -1981 21800 -1925 21856
rect -3835 21693 -3779 21706
rect -3835 21650 -3834 21693
rect -3834 21650 -3780 21693
rect -3780 21650 -3779 21693
rect -3651 21693 -3595 21706
rect -3651 21650 -3650 21693
rect -3650 21650 -3596 21693
rect -3596 21650 -3595 21693
rect -3467 21693 -3411 21706
rect -3467 21650 -3466 21693
rect -3466 21650 -3412 21693
rect -3412 21650 -3411 21693
rect -3375 21454 -3370 21574
rect -3370 21454 -3324 21574
rect -3324 21454 -3319 21574
rect -4060 21131 -4004 21187
rect -3242 21131 -3186 21187
rect -4779 21014 -4723 21070
rect 575 21800 631 21856
rect -2349 21693 -2293 21706
rect -2349 21650 -2348 21693
rect -2348 21650 -2294 21693
rect -2294 21650 -2293 21693
rect -2165 21693 -2109 21706
rect -2165 21650 -2164 21693
rect -2164 21650 -2110 21693
rect -2110 21650 -2109 21693
rect -1981 21693 -1925 21706
rect -1981 21650 -1980 21693
rect -1980 21650 -1926 21693
rect -1926 21650 -1925 21693
rect -1889 21454 -1884 21574
rect -1884 21454 -1838 21574
rect -1838 21454 -1833 21574
rect -2574 21131 -2518 21187
rect -1756 21131 -1700 21187
rect -1403 21014 -1347 21070
rect -6931 20906 -6875 20962
rect -5621 20907 -5565 20963
rect -7601 20799 -7545 20855
rect -7969 20412 -7964 20532
rect -7964 20412 -7918 20532
rect -7918 20412 -7913 20532
rect -7601 20412 -7596 20532
rect -7596 20412 -7550 20532
rect -7550 20412 -7545 20532
rect -7785 20112 -7780 20232
rect -7780 20112 -7734 20232
rect -7734 20112 -7729 20232
rect -7279 20411 -7274 20532
rect -7274 20411 -7228 20532
rect -7228 20411 -7223 20532
rect -7417 20112 -7412 20232
rect -7412 20112 -7366 20232
rect -7366 20112 -7361 20232
rect -7877 19993 -7876 20036
rect -7876 19993 -7822 20036
rect -7822 19993 -7821 20036
rect -7877 19980 -7821 19993
rect -7693 19993 -7692 20036
rect -7692 19993 -7638 20036
rect -7638 19993 -7637 20036
rect -7693 19980 -7637 19993
rect -7509 19993 -7508 20036
rect -7508 19993 -7454 20036
rect -7454 19993 -7453 20036
rect -7509 19980 -7453 19993
rect -7877 19830 -7821 19886
rect -6115 20800 -6059 20856
rect -6483 20413 -6478 20533
rect -6478 20413 -6432 20533
rect -6432 20413 -6427 20533
rect -6115 20413 -6110 20533
rect -6110 20413 -6064 20533
rect -6064 20413 -6059 20533
rect -6299 20113 -6294 20233
rect -6294 20113 -6248 20233
rect -6248 20113 -6243 20233
rect -5793 20412 -5788 20533
rect -5788 20412 -5742 20533
rect -5742 20412 -5737 20533
rect -5931 20113 -5926 20233
rect -5926 20113 -5880 20233
rect -5880 20113 -5875 20233
rect -6391 19994 -6390 20037
rect -6390 19994 -6336 20037
rect -6336 19994 -6335 20037
rect -6391 19981 -6335 19994
rect -6207 19994 -6206 20037
rect -6206 19994 -6152 20037
rect -6152 19994 -6151 20037
rect -6207 19981 -6151 19994
rect -6023 19994 -6022 20037
rect -6022 19994 -5968 20037
rect -5968 19994 -5967 20037
rect -6023 19981 -5967 19994
rect -6391 19831 -6335 19887
rect -7693 19714 -7637 19770
rect -7364 19714 -7308 19770
rect -7107 19714 -7051 19770
rect -6207 19715 -6151 19771
rect -5878 19715 -5822 19771
rect -5445 19715 -5389 19771
rect 2061 21800 2117 21856
rect 207 21693 263 21706
rect 207 21650 208 21693
rect 208 21650 262 21693
rect 262 21650 263 21693
rect 391 21693 447 21706
rect 391 21650 392 21693
rect 392 21650 446 21693
rect 446 21650 447 21693
rect 575 21693 631 21706
rect 575 21650 576 21693
rect 576 21650 630 21693
rect 630 21650 631 21693
rect 667 21454 672 21574
rect 672 21454 718 21574
rect 718 21454 723 21574
rect -18 21131 38 21187
rect 800 21131 856 21187
rect -737 21014 -681 21070
rect 4617 21800 4673 21856
rect 1693 21693 1749 21706
rect 1693 21650 1694 21693
rect 1694 21650 1748 21693
rect 1748 21650 1749 21693
rect 1877 21693 1933 21706
rect 1877 21650 1878 21693
rect 1878 21650 1932 21693
rect 1932 21650 1933 21693
rect 2061 21693 2117 21706
rect 2061 21650 2062 21693
rect 2062 21650 2116 21693
rect 2116 21650 2117 21693
rect 2153 21454 2158 21574
rect 2158 21454 2204 21574
rect 2204 21454 2209 21574
rect 1468 21131 1524 21187
rect 2286 21131 2342 21187
rect 2639 21014 2695 21070
rect -2889 20903 -2833 20959
rect -1579 20904 -1523 20960
rect -3559 20796 -3503 20852
rect -3927 20409 -3922 20529
rect -3922 20409 -3876 20529
rect -3876 20409 -3871 20529
rect -3559 20409 -3554 20529
rect -3554 20409 -3508 20529
rect -3508 20409 -3503 20529
rect -3743 20109 -3738 20229
rect -3738 20109 -3692 20229
rect -3692 20109 -3687 20229
rect -3237 20408 -3232 20529
rect -3232 20408 -3186 20529
rect -3186 20408 -3181 20529
rect -3375 20109 -3370 20229
rect -3370 20109 -3324 20229
rect -3324 20109 -3319 20229
rect -3835 19990 -3834 20033
rect -3834 19990 -3780 20033
rect -3780 19990 -3779 20033
rect -3835 19977 -3779 19990
rect -3651 19990 -3650 20033
rect -3650 19990 -3596 20033
rect -3596 19990 -3595 20033
rect -3651 19977 -3595 19990
rect -3467 19990 -3466 20033
rect -3466 19990 -3412 20033
rect -3412 19990 -3411 20033
rect -3467 19977 -3411 19990
rect -3835 19827 -3779 19883
rect -2073 20797 -2017 20853
rect -2441 20410 -2436 20530
rect -2436 20410 -2390 20530
rect -2390 20410 -2385 20530
rect -2073 20410 -2068 20530
rect -2068 20410 -2022 20530
rect -2022 20410 -2017 20530
rect -2257 20110 -2252 20230
rect -2252 20110 -2206 20230
rect -2206 20110 -2201 20230
rect -1751 20409 -1746 20530
rect -1746 20409 -1700 20530
rect -1700 20409 -1695 20530
rect -1889 20110 -1884 20230
rect -1884 20110 -1838 20230
rect -1838 20110 -1833 20230
rect -2349 19991 -2348 20034
rect -2348 19991 -2294 20034
rect -2294 19991 -2293 20034
rect -2349 19978 -2293 19991
rect -2165 19991 -2164 20034
rect -2164 19991 -2110 20034
rect -2110 19991 -2109 20034
rect -2165 19978 -2109 19991
rect -1981 19991 -1980 20034
rect -1980 19991 -1926 20034
rect -1926 19991 -1925 20034
rect -1981 19978 -1925 19991
rect -2349 19828 -2293 19884
rect -3651 19711 -3595 19767
rect -3322 19711 -3266 19767
rect -3065 19711 -3009 19767
rect -2165 19712 -2109 19768
rect -1836 19712 -1780 19768
rect -1403 19712 -1347 19768
rect 6103 21800 6159 21856
rect 4249 21693 4305 21706
rect 4249 21650 4250 21693
rect 4250 21650 4304 21693
rect 4304 21650 4305 21693
rect 4433 21693 4489 21706
rect 4433 21650 4434 21693
rect 4434 21650 4488 21693
rect 4488 21650 4489 21693
rect 4617 21693 4673 21706
rect 4617 21650 4618 21693
rect 4618 21650 4672 21693
rect 4672 21650 4673 21693
rect 4709 21454 4714 21574
rect 4714 21454 4760 21574
rect 4760 21454 4765 21574
rect 4024 21131 4080 21187
rect 4842 21131 4898 21187
rect 3305 21014 3361 21070
rect 8659 21800 8715 21856
rect 5735 21693 5791 21706
rect 5735 21650 5736 21693
rect 5736 21650 5790 21693
rect 5790 21650 5791 21693
rect 5919 21693 5975 21706
rect 5919 21650 5920 21693
rect 5920 21650 5974 21693
rect 5974 21650 5975 21693
rect 6103 21693 6159 21706
rect 6103 21650 6104 21693
rect 6104 21650 6158 21693
rect 6158 21650 6159 21693
rect 6195 21454 6200 21574
rect 6200 21454 6246 21574
rect 6246 21454 6251 21574
rect 5510 21131 5566 21187
rect 6328 21131 6384 21187
rect 6681 21014 6737 21070
rect 1153 20903 1209 20959
rect 2463 20904 2519 20960
rect 483 20796 539 20852
rect 115 20409 120 20529
rect 120 20409 166 20529
rect 166 20409 171 20529
rect 483 20409 488 20529
rect 488 20409 534 20529
rect 534 20409 539 20529
rect 299 20109 304 20229
rect 304 20109 350 20229
rect 350 20109 355 20229
rect 805 20408 810 20529
rect 810 20408 856 20529
rect 856 20408 861 20529
rect 667 20109 672 20229
rect 672 20109 718 20229
rect 718 20109 723 20229
rect 207 19990 208 20033
rect 208 19990 262 20033
rect 262 19990 263 20033
rect 207 19977 263 19990
rect 391 19990 392 20033
rect 392 19990 446 20033
rect 446 19990 447 20033
rect 391 19977 447 19990
rect 575 19990 576 20033
rect 576 19990 630 20033
rect 630 19990 631 20033
rect 575 19977 631 19990
rect 207 19827 263 19883
rect 1969 20797 2025 20853
rect 1601 20410 1606 20530
rect 1606 20410 1652 20530
rect 1652 20410 1657 20530
rect 1969 20410 1974 20530
rect 1974 20410 2020 20530
rect 2020 20410 2025 20530
rect 1785 20110 1790 20230
rect 1790 20110 1836 20230
rect 1836 20110 1841 20230
rect 2291 20409 2296 20530
rect 2296 20409 2342 20530
rect 2342 20409 2347 20530
rect 2153 20110 2158 20230
rect 2158 20110 2204 20230
rect 2204 20110 2209 20230
rect 1693 19991 1694 20034
rect 1694 19991 1748 20034
rect 1748 19991 1749 20034
rect 1693 19978 1749 19991
rect 1877 19991 1878 20034
rect 1878 19991 1932 20034
rect 1932 19991 1933 20034
rect 1877 19978 1933 19991
rect 2061 19991 2062 20034
rect 2062 19991 2116 20034
rect 2116 19991 2117 20034
rect 2061 19978 2117 19991
rect 1693 19828 1749 19884
rect 391 19711 447 19767
rect 720 19711 776 19767
rect 977 19711 1033 19767
rect 1877 19712 1933 19768
rect 2206 19712 2262 19768
rect 2639 19712 2695 19768
rect 10145 21800 10201 21856
rect 8291 21693 8347 21706
rect 8291 21650 8292 21693
rect 8292 21650 8346 21693
rect 8346 21650 8347 21693
rect 8475 21693 8531 21706
rect 8475 21650 8476 21693
rect 8476 21650 8530 21693
rect 8530 21650 8531 21693
rect 8659 21693 8715 21706
rect 8659 21650 8660 21693
rect 8660 21650 8714 21693
rect 8714 21650 8715 21693
rect 8751 21454 8756 21574
rect 8756 21454 8802 21574
rect 8802 21454 8807 21574
rect 8066 21131 8122 21187
rect 8884 21131 8940 21187
rect 7347 21014 7403 21070
rect 12701 21800 12757 21856
rect 9777 21693 9833 21706
rect 9777 21650 9778 21693
rect 9778 21650 9832 21693
rect 9832 21650 9833 21693
rect 9961 21693 10017 21706
rect 9961 21650 9962 21693
rect 9962 21650 10016 21693
rect 10016 21650 10017 21693
rect 10145 21693 10201 21706
rect 10145 21650 10146 21693
rect 10146 21650 10200 21693
rect 10200 21650 10201 21693
rect 10237 21454 10242 21574
rect 10242 21454 10288 21574
rect 10288 21454 10293 21574
rect 9552 21131 9608 21187
rect 10370 21131 10426 21187
rect 10723 21014 10779 21070
rect 5195 20903 5251 20959
rect 6505 20904 6561 20960
rect 4525 20796 4581 20852
rect 4157 20409 4162 20529
rect 4162 20409 4208 20529
rect 4208 20409 4213 20529
rect 4525 20409 4530 20529
rect 4530 20409 4576 20529
rect 4576 20409 4581 20529
rect 4341 20109 4346 20229
rect 4346 20109 4392 20229
rect 4392 20109 4397 20229
rect 4847 20408 4852 20529
rect 4852 20408 4898 20529
rect 4898 20408 4903 20529
rect 4709 20109 4714 20229
rect 4714 20109 4760 20229
rect 4760 20109 4765 20229
rect 4249 19990 4250 20033
rect 4250 19990 4304 20033
rect 4304 19990 4305 20033
rect 4249 19977 4305 19990
rect 4433 19990 4434 20033
rect 4434 19990 4488 20033
rect 4488 19990 4489 20033
rect 4433 19977 4489 19990
rect 4617 19990 4618 20033
rect 4618 19990 4672 20033
rect 4672 19990 4673 20033
rect 4617 19977 4673 19990
rect 4249 19827 4305 19883
rect 6011 20797 6067 20853
rect 5643 20410 5648 20530
rect 5648 20410 5694 20530
rect 5694 20410 5699 20530
rect 6011 20410 6016 20530
rect 6016 20410 6062 20530
rect 6062 20410 6067 20530
rect 5827 20110 5832 20230
rect 5832 20110 5878 20230
rect 5878 20110 5883 20230
rect 6333 20409 6338 20530
rect 6338 20409 6384 20530
rect 6384 20409 6389 20530
rect 6195 20110 6200 20230
rect 6200 20110 6246 20230
rect 6246 20110 6251 20230
rect 5735 19991 5736 20034
rect 5736 19991 5790 20034
rect 5790 19991 5791 20034
rect 5735 19978 5791 19991
rect 5919 19991 5920 20034
rect 5920 19991 5974 20034
rect 5974 19991 5975 20034
rect 5919 19978 5975 19991
rect 6103 19991 6104 20034
rect 6104 19991 6158 20034
rect 6158 19991 6159 20034
rect 6103 19978 6159 19991
rect 5735 19828 5791 19884
rect 4433 19711 4489 19767
rect 4762 19711 4818 19767
rect 5019 19711 5075 19767
rect 5919 19712 5975 19768
rect 6248 19712 6304 19768
rect 6681 19712 6737 19768
rect 14187 21800 14243 21856
rect 12333 21693 12389 21706
rect 12333 21650 12334 21693
rect 12334 21650 12388 21693
rect 12388 21650 12389 21693
rect 12517 21693 12573 21706
rect 12517 21650 12518 21693
rect 12518 21650 12572 21693
rect 12572 21650 12573 21693
rect 12701 21693 12757 21706
rect 12701 21650 12702 21693
rect 12702 21650 12756 21693
rect 12756 21650 12757 21693
rect 12793 21454 12798 21574
rect 12798 21454 12844 21574
rect 12844 21454 12849 21574
rect 12108 21131 12164 21187
rect 12926 21131 12982 21187
rect 11389 21014 11445 21070
rect 16743 21800 16799 21856
rect 13819 21693 13875 21706
rect 13819 21650 13820 21693
rect 13820 21650 13874 21693
rect 13874 21650 13875 21693
rect 14003 21693 14059 21706
rect 14003 21650 14004 21693
rect 14004 21650 14058 21693
rect 14058 21650 14059 21693
rect 14187 21693 14243 21706
rect 14187 21650 14188 21693
rect 14188 21650 14242 21693
rect 14242 21650 14243 21693
rect 14279 21454 14284 21574
rect 14284 21454 14330 21574
rect 14330 21454 14335 21574
rect 13594 21131 13650 21187
rect 14412 21131 14468 21187
rect 14765 21014 14821 21070
rect 9237 20903 9293 20959
rect 10547 20904 10603 20960
rect 8567 20796 8623 20852
rect 8199 20409 8204 20529
rect 8204 20409 8250 20529
rect 8250 20409 8255 20529
rect 8567 20409 8572 20529
rect 8572 20409 8618 20529
rect 8618 20409 8623 20529
rect 8383 20109 8388 20229
rect 8388 20109 8434 20229
rect 8434 20109 8439 20229
rect 8889 20408 8894 20529
rect 8894 20408 8940 20529
rect 8940 20408 8945 20529
rect 8751 20109 8756 20229
rect 8756 20109 8802 20229
rect 8802 20109 8807 20229
rect 8291 19990 8292 20033
rect 8292 19990 8346 20033
rect 8346 19990 8347 20033
rect 8291 19977 8347 19990
rect 8475 19990 8476 20033
rect 8476 19990 8530 20033
rect 8530 19990 8531 20033
rect 8475 19977 8531 19990
rect 8659 19990 8660 20033
rect 8660 19990 8714 20033
rect 8714 19990 8715 20033
rect 8659 19977 8715 19990
rect 8291 19827 8347 19883
rect 10053 20797 10109 20853
rect 9685 20410 9690 20530
rect 9690 20410 9736 20530
rect 9736 20410 9741 20530
rect 10053 20410 10058 20530
rect 10058 20410 10104 20530
rect 10104 20410 10109 20530
rect 9869 20110 9874 20230
rect 9874 20110 9920 20230
rect 9920 20110 9925 20230
rect 10375 20409 10380 20530
rect 10380 20409 10426 20530
rect 10426 20409 10431 20530
rect 10237 20110 10242 20230
rect 10242 20110 10288 20230
rect 10288 20110 10293 20230
rect 9777 19991 9778 20034
rect 9778 19991 9832 20034
rect 9832 19991 9833 20034
rect 9777 19978 9833 19991
rect 9961 19991 9962 20034
rect 9962 19991 10016 20034
rect 10016 19991 10017 20034
rect 9961 19978 10017 19991
rect 10145 19991 10146 20034
rect 10146 19991 10200 20034
rect 10200 19991 10201 20034
rect 10145 19978 10201 19991
rect 9777 19828 9833 19884
rect 8475 19711 8531 19767
rect 8804 19711 8860 19767
rect 9061 19711 9117 19767
rect 9961 19712 10017 19768
rect 10290 19712 10346 19768
rect 10723 19712 10779 19768
rect 18229 21800 18285 21856
rect 16375 21693 16431 21706
rect 16375 21650 16376 21693
rect 16376 21650 16430 21693
rect 16430 21650 16431 21693
rect 16559 21693 16615 21706
rect 16559 21650 16560 21693
rect 16560 21650 16614 21693
rect 16614 21650 16615 21693
rect 16743 21693 16799 21706
rect 16743 21650 16744 21693
rect 16744 21650 16798 21693
rect 16798 21650 16799 21693
rect 16835 21454 16840 21574
rect 16840 21454 16886 21574
rect 16886 21454 16891 21574
rect 16150 21131 16206 21187
rect 16968 21131 17024 21187
rect 15386 21014 15442 21070
rect 17861 21693 17917 21706
rect 17861 21650 17862 21693
rect 17862 21650 17916 21693
rect 17916 21650 17917 21693
rect 18045 21693 18101 21706
rect 18045 21650 18046 21693
rect 18046 21650 18100 21693
rect 18100 21650 18101 21693
rect 18229 21693 18285 21706
rect 18229 21650 18230 21693
rect 18230 21650 18284 21693
rect 18284 21650 18285 21693
rect 18321 21454 18326 21574
rect 18326 21454 18372 21574
rect 18372 21454 18377 21574
rect 17636 21131 17692 21187
rect 18454 21131 18510 21187
rect 18807 21014 18863 21070
rect 13279 20903 13335 20959
rect 14589 20904 14645 20960
rect 12609 20796 12665 20852
rect 12241 20409 12246 20529
rect 12246 20409 12292 20529
rect 12292 20409 12297 20529
rect 12609 20409 12614 20529
rect 12614 20409 12660 20529
rect 12660 20409 12665 20529
rect 12425 20109 12430 20229
rect 12430 20109 12476 20229
rect 12476 20109 12481 20229
rect 12931 20408 12936 20529
rect 12936 20408 12982 20529
rect 12982 20408 12987 20529
rect 12793 20109 12798 20229
rect 12798 20109 12844 20229
rect 12844 20109 12849 20229
rect 12333 19990 12334 20033
rect 12334 19990 12388 20033
rect 12388 19990 12389 20033
rect 12333 19977 12389 19990
rect 12517 19990 12518 20033
rect 12518 19990 12572 20033
rect 12572 19990 12573 20033
rect 12517 19977 12573 19990
rect 12701 19990 12702 20033
rect 12702 19990 12756 20033
rect 12756 19990 12757 20033
rect 12701 19977 12757 19990
rect 12333 19827 12389 19883
rect 14095 20797 14151 20853
rect 13727 20410 13732 20530
rect 13732 20410 13778 20530
rect 13778 20410 13783 20530
rect 14095 20410 14100 20530
rect 14100 20410 14146 20530
rect 14146 20410 14151 20530
rect 13911 20110 13916 20230
rect 13916 20110 13962 20230
rect 13962 20110 13967 20230
rect 14417 20409 14422 20530
rect 14422 20409 14468 20530
rect 14468 20409 14473 20530
rect 14279 20110 14284 20230
rect 14284 20110 14330 20230
rect 14330 20110 14335 20230
rect 13819 19991 13820 20034
rect 13820 19991 13874 20034
rect 13874 19991 13875 20034
rect 13819 19978 13875 19991
rect 14003 19991 14004 20034
rect 14004 19991 14058 20034
rect 14058 19991 14059 20034
rect 14003 19978 14059 19991
rect 14187 19991 14188 20034
rect 14188 19991 14242 20034
rect 14242 19991 14243 20034
rect 14187 19978 14243 19991
rect 13819 19828 13875 19884
rect 12517 19711 12573 19767
rect 12846 19711 12902 19767
rect 13103 19711 13159 19767
rect 14003 19712 14059 19768
rect 14332 19712 14388 19768
rect 14765 19712 14821 19768
rect 17321 20903 17377 20959
rect 18631 20904 18687 20960
rect 16651 20796 16707 20852
rect 16283 20409 16288 20529
rect 16288 20409 16334 20529
rect 16334 20409 16339 20529
rect 16651 20409 16656 20529
rect 16656 20409 16702 20529
rect 16702 20409 16707 20529
rect 16467 20109 16472 20229
rect 16472 20109 16518 20229
rect 16518 20109 16523 20229
rect 16973 20408 16978 20529
rect 16978 20408 17024 20529
rect 17024 20408 17029 20529
rect 16835 20109 16840 20229
rect 16840 20109 16886 20229
rect 16886 20109 16891 20229
rect 16375 19990 16376 20033
rect 16376 19990 16430 20033
rect 16430 19990 16431 20033
rect 16375 19977 16431 19990
rect 16559 19990 16560 20033
rect 16560 19990 16614 20033
rect 16614 19990 16615 20033
rect 16559 19977 16615 19990
rect 16743 19990 16744 20033
rect 16744 19990 16798 20033
rect 16798 19990 16799 20033
rect 16743 19977 16799 19990
rect 16375 19827 16431 19883
rect 18137 20797 18193 20853
rect 17769 20410 17774 20530
rect 17774 20410 17820 20530
rect 17820 20410 17825 20530
rect 18137 20410 18142 20530
rect 18142 20410 18188 20530
rect 18188 20410 18193 20530
rect 17953 20110 17958 20230
rect 17958 20110 18004 20230
rect 18004 20110 18009 20230
rect 18459 20409 18464 20530
rect 18464 20409 18510 20530
rect 18510 20409 18515 20530
rect 18321 20110 18326 20230
rect 18326 20110 18372 20230
rect 18372 20110 18377 20230
rect 17861 19991 17862 20034
rect 17862 19991 17916 20034
rect 17916 19991 17917 20034
rect 17861 19978 17917 19991
rect 18045 19991 18046 20034
rect 18046 19991 18100 20034
rect 18100 19991 18101 20034
rect 18045 19978 18101 19991
rect 18229 19991 18230 20034
rect 18230 19991 18284 20034
rect 18284 19991 18285 20034
rect 18229 19978 18285 19991
rect 17861 19828 17917 19884
rect 16559 19711 16615 19767
rect 16888 19711 16944 19767
rect 17145 19711 17201 19767
rect 18045 19712 18101 19768
rect 18374 19712 18430 19768
rect 18807 19712 18863 19768
rect -8549 19598 -8493 19654
rect -7509 19598 -7453 19654
rect -6023 19599 -5967 19655
rect -7877 19491 -7821 19504
rect -7877 19448 -7876 19491
rect -7876 19448 -7822 19491
rect -7822 19448 -7821 19491
rect -7693 19491 -7637 19504
rect -7693 19448 -7692 19491
rect -7692 19448 -7638 19491
rect -7638 19448 -7637 19491
rect -7509 19491 -7453 19504
rect -7509 19448 -7508 19491
rect -7508 19448 -7454 19491
rect -7454 19448 -7453 19491
rect -7417 19252 -7412 19372
rect -7412 19252 -7366 19372
rect -7366 19252 -7361 19372
rect -8102 18929 -8046 18985
rect -7284 18929 -7228 18985
rect -6931 18811 -6875 18867
rect -7107 18703 -7051 18757
rect -7601 18594 -7545 18650
rect -7969 18207 -7964 18327
rect -7964 18207 -7918 18327
rect -7918 18207 -7913 18327
rect -7601 18207 -7596 18327
rect -7596 18207 -7550 18327
rect -7550 18207 -7545 18327
rect -7785 17907 -7780 18027
rect -7780 17907 -7734 18027
rect -7734 17907 -7729 18027
rect -7279 18206 -7274 18327
rect -7274 18206 -7228 18327
rect -7228 18206 -7223 18327
rect -7417 17907 -7412 18027
rect -7412 17907 -7366 18027
rect -7366 17907 -7361 18027
rect -7877 17788 -7876 17831
rect -7876 17788 -7822 17831
rect -7822 17788 -7821 17831
rect -7877 17775 -7821 17788
rect -7693 17788 -7692 17831
rect -7692 17788 -7638 17831
rect -7638 17788 -7637 17831
rect -7693 17775 -7637 17788
rect -7509 17788 -7508 17831
rect -7508 17788 -7454 17831
rect -7454 17788 -7453 17831
rect -7509 17775 -7453 17788
rect -7877 17625 -7821 17681
rect -8685 17509 -8629 17565
rect -7693 17509 -7637 17565
rect -7364 17509 -7308 17565
rect -6931 17509 -6875 17565
rect -9501 17393 -9445 17449
rect -7509 17393 -7453 17449
rect -7877 17286 -7821 17299
rect -7877 17243 -7876 17286
rect -7876 17243 -7822 17286
rect -7822 17243 -7821 17286
rect -7693 17286 -7637 17299
rect -7693 17243 -7692 17286
rect -7692 17243 -7638 17286
rect -7638 17243 -7637 17286
rect -7509 17286 -7453 17299
rect -7509 17243 -7508 17286
rect -7508 17243 -7454 17286
rect -7454 17243 -7453 17286
rect -7417 17047 -7412 17167
rect -7412 17047 -7366 17167
rect -7366 17047 -7361 17167
rect -8102 16724 -8046 16780
rect -7284 16724 -7228 16780
rect -4507 19595 -4451 19651
rect -3467 19595 -3411 19651
rect -6391 19492 -6335 19505
rect -6391 19449 -6390 19492
rect -6390 19449 -6336 19492
rect -6336 19449 -6335 19492
rect -6207 19492 -6151 19505
rect -6207 19449 -6206 19492
rect -6206 19449 -6152 19492
rect -6152 19449 -6151 19492
rect -6023 19492 -5967 19505
rect -6023 19449 -6022 19492
rect -6022 19449 -5968 19492
rect -5968 19449 -5967 19492
rect -5931 19253 -5926 19373
rect -5926 19253 -5880 19373
rect -5880 19253 -5875 19373
rect -6616 18930 -6560 18986
rect -5798 18930 -5742 18986
rect -1981 19596 -1925 19652
rect -3835 19488 -3779 19501
rect -3835 19445 -3834 19488
rect -3834 19445 -3780 19488
rect -3780 19445 -3779 19488
rect -3651 19488 -3595 19501
rect -3651 19445 -3650 19488
rect -3650 19445 -3596 19488
rect -3596 19445 -3595 19488
rect -3467 19488 -3411 19501
rect -3467 19445 -3466 19488
rect -3466 19445 -3412 19488
rect -3412 19445 -3411 19488
rect -3375 19249 -3370 19369
rect -3370 19249 -3324 19369
rect -3324 19249 -3319 19369
rect -4060 18926 -4004 18982
rect -3242 18926 -3186 18982
rect -2889 18808 -2833 18864
rect -3065 18700 -3009 18754
rect -3559 18591 -3503 18647
rect -3927 18204 -3922 18324
rect -3922 18204 -3876 18324
rect -3876 18204 -3871 18324
rect -3559 18204 -3554 18324
rect -3554 18204 -3508 18324
rect -3508 18204 -3503 18324
rect -3743 17904 -3738 18024
rect -3738 17904 -3692 18024
rect -3692 17904 -3687 18024
rect -3237 18203 -3232 18324
rect -3232 18203 -3186 18324
rect -3186 18203 -3181 18324
rect -3375 17904 -3370 18024
rect -3370 17904 -3324 18024
rect -3324 17904 -3319 18024
rect -3835 17785 -3834 17828
rect -3834 17785 -3780 17828
rect -3780 17785 -3779 17828
rect -3835 17772 -3779 17785
rect -3651 17785 -3650 17828
rect -3650 17785 -3596 17828
rect -3596 17785 -3595 17828
rect -3651 17772 -3595 17785
rect -3467 17785 -3466 17828
rect -3466 17785 -3412 17828
rect -3412 17785 -3411 17828
rect -3467 17772 -3411 17785
rect -3835 17622 -3779 17678
rect -4643 17506 -4587 17562
rect -3651 17506 -3595 17562
rect -3322 17506 -3266 17562
rect -2889 17506 -2833 17562
rect -5489 17390 -5433 17446
rect -3467 17390 -3411 17446
rect -3835 17283 -3779 17296
rect -3835 17240 -3834 17283
rect -3834 17240 -3780 17283
rect -3780 17240 -3779 17283
rect -3651 17283 -3595 17296
rect -3651 17240 -3650 17283
rect -3650 17240 -3596 17283
rect -3596 17240 -3595 17283
rect -3467 17283 -3411 17296
rect -3467 17240 -3466 17283
rect -3466 17240 -3412 17283
rect -3412 17240 -3411 17283
rect -3375 17044 -3370 17164
rect -3370 17044 -3324 17164
rect -3324 17044 -3319 17164
rect -4060 16721 -4004 16777
rect -3242 16721 -3186 16777
rect -8957 16606 -8901 16662
rect -8685 16606 -8629 16662
rect -465 19595 -409 19651
rect 575 19595 631 19651
rect -2349 19489 -2293 19502
rect -2349 19446 -2348 19489
rect -2348 19446 -2294 19489
rect -2294 19446 -2293 19489
rect -2165 19489 -2109 19502
rect -2165 19446 -2164 19489
rect -2164 19446 -2110 19489
rect -2110 19446 -2109 19489
rect -1981 19489 -1925 19502
rect -1981 19446 -1980 19489
rect -1980 19446 -1926 19489
rect -1926 19446 -1925 19489
rect -1889 19250 -1884 19370
rect -1884 19250 -1838 19370
rect -1838 19250 -1833 19370
rect -2574 18927 -2518 18983
rect -1756 18927 -1700 18983
rect 2061 19596 2117 19652
rect 207 19488 263 19501
rect 207 19445 208 19488
rect 208 19445 262 19488
rect 262 19445 263 19488
rect 391 19488 447 19501
rect 391 19445 392 19488
rect 392 19445 446 19488
rect 446 19445 447 19488
rect 575 19488 631 19501
rect 575 19445 576 19488
rect 576 19445 630 19488
rect 630 19445 631 19488
rect 667 19249 672 19369
rect 672 19249 718 19369
rect 718 19249 723 19369
rect -18 18926 38 18982
rect 800 18926 856 18982
rect 1153 18808 1209 18864
rect 977 18700 1033 18754
rect 483 18591 539 18647
rect 115 18204 120 18324
rect 120 18204 166 18324
rect 166 18204 171 18324
rect 483 18204 488 18324
rect 488 18204 534 18324
rect 534 18204 539 18324
rect 299 17904 304 18024
rect 304 17904 350 18024
rect 350 17904 355 18024
rect 805 18203 810 18324
rect 810 18203 856 18324
rect 856 18203 861 18324
rect 667 17904 672 18024
rect 672 17904 718 18024
rect 718 17904 723 18024
rect 207 17785 208 17828
rect 208 17785 262 17828
rect 262 17785 263 17828
rect 207 17772 263 17785
rect 391 17785 392 17828
rect 392 17785 446 17828
rect 446 17785 447 17828
rect 391 17772 447 17785
rect 575 17785 576 17828
rect 576 17785 630 17828
rect 630 17785 631 17828
rect 575 17772 631 17785
rect 207 17622 263 17678
rect -601 17506 -545 17562
rect 391 17506 447 17562
rect 720 17506 776 17562
rect 1153 17506 1209 17562
rect -1447 17390 -1391 17446
rect 575 17390 631 17446
rect 207 17283 263 17296
rect 207 17240 208 17283
rect 208 17240 262 17283
rect 262 17240 263 17283
rect 391 17283 447 17296
rect 391 17240 392 17283
rect 392 17240 446 17283
rect 446 17240 447 17283
rect 575 17283 631 17296
rect 575 17240 576 17283
rect 576 17240 630 17283
rect 630 17240 631 17283
rect 667 17044 672 17164
rect 672 17044 718 17164
rect 718 17044 723 17164
rect -18 16721 38 16777
rect 800 16721 856 16777
rect -4945 16603 -4889 16659
rect -4643 16603 -4587 16659
rect 3577 19595 3633 19651
rect 4617 19595 4673 19651
rect 1693 19489 1749 19502
rect 1693 19446 1694 19489
rect 1694 19446 1748 19489
rect 1748 19446 1749 19489
rect 1877 19489 1933 19502
rect 1877 19446 1878 19489
rect 1878 19446 1932 19489
rect 1932 19446 1933 19489
rect 2061 19489 2117 19502
rect 2061 19446 2062 19489
rect 2062 19446 2116 19489
rect 2116 19446 2117 19489
rect 2153 19250 2158 19370
rect 2158 19250 2204 19370
rect 2204 19250 2209 19370
rect 1468 18927 1524 18983
rect 2286 18927 2342 18983
rect 6103 19596 6159 19652
rect 4249 19488 4305 19501
rect 4249 19445 4250 19488
rect 4250 19445 4304 19488
rect 4304 19445 4305 19488
rect 4433 19488 4489 19501
rect 4433 19445 4434 19488
rect 4434 19445 4488 19488
rect 4488 19445 4489 19488
rect 4617 19488 4673 19501
rect 4617 19445 4618 19488
rect 4618 19445 4672 19488
rect 4672 19445 4673 19488
rect 4709 19249 4714 19369
rect 4714 19249 4760 19369
rect 4760 19249 4765 19369
rect 4024 18926 4080 18982
rect 4842 18926 4898 18982
rect 5195 18808 5251 18864
rect 5019 18700 5075 18754
rect 4525 18591 4581 18647
rect 4157 18204 4162 18324
rect 4162 18204 4208 18324
rect 4208 18204 4213 18324
rect 4525 18204 4530 18324
rect 4530 18204 4576 18324
rect 4576 18204 4581 18324
rect 4341 17904 4346 18024
rect 4346 17904 4392 18024
rect 4392 17904 4397 18024
rect 4847 18203 4852 18324
rect 4852 18203 4898 18324
rect 4898 18203 4903 18324
rect 4709 17904 4714 18024
rect 4714 17904 4760 18024
rect 4760 17904 4765 18024
rect 4249 17785 4250 17828
rect 4250 17785 4304 17828
rect 4304 17785 4305 17828
rect 4249 17772 4305 17785
rect 4433 17785 4434 17828
rect 4434 17785 4488 17828
rect 4488 17785 4489 17828
rect 4433 17772 4489 17785
rect 4617 17785 4618 17828
rect 4618 17785 4672 17828
rect 4672 17785 4673 17828
rect 4617 17772 4673 17785
rect 4249 17622 4305 17678
rect 3441 17506 3497 17562
rect 4433 17506 4489 17562
rect 4762 17506 4818 17562
rect 5195 17506 5251 17562
rect 2595 17390 2651 17446
rect 4617 17390 4673 17446
rect 4249 17283 4305 17296
rect 4249 17240 4250 17283
rect 4250 17240 4304 17283
rect 4304 17240 4305 17283
rect 4433 17283 4489 17296
rect 4433 17240 4434 17283
rect 4434 17240 4488 17283
rect 4488 17240 4489 17283
rect 4617 17283 4673 17296
rect 4617 17240 4618 17283
rect 4618 17240 4672 17283
rect 4672 17240 4673 17283
rect 4709 17044 4714 17164
rect 4714 17044 4760 17164
rect 4760 17044 4765 17164
rect 4024 16721 4080 16777
rect 4842 16721 4898 16777
rect -903 16603 -847 16659
rect -601 16603 -545 16659
rect 7619 19595 7675 19651
rect 8659 19595 8715 19651
rect 5735 19489 5791 19502
rect 5735 19446 5736 19489
rect 5736 19446 5790 19489
rect 5790 19446 5791 19489
rect 5919 19489 5975 19502
rect 5919 19446 5920 19489
rect 5920 19446 5974 19489
rect 5974 19446 5975 19489
rect 6103 19489 6159 19502
rect 6103 19446 6104 19489
rect 6104 19446 6158 19489
rect 6158 19446 6159 19489
rect 6195 19250 6200 19370
rect 6200 19250 6246 19370
rect 6246 19250 6251 19370
rect 5510 18927 5566 18983
rect 6328 18927 6384 18983
rect 10145 19596 10201 19652
rect 8291 19488 8347 19501
rect 8291 19445 8292 19488
rect 8292 19445 8346 19488
rect 8346 19445 8347 19488
rect 8475 19488 8531 19501
rect 8475 19445 8476 19488
rect 8476 19445 8530 19488
rect 8530 19445 8531 19488
rect 8659 19488 8715 19501
rect 8659 19445 8660 19488
rect 8660 19445 8714 19488
rect 8714 19445 8715 19488
rect 8751 19249 8756 19369
rect 8756 19249 8802 19369
rect 8802 19249 8807 19369
rect 8066 18926 8122 18982
rect 8884 18926 8940 18982
rect 9237 18808 9293 18864
rect 9061 18700 9117 18754
rect 8567 18591 8623 18647
rect 8199 18204 8204 18324
rect 8204 18204 8250 18324
rect 8250 18204 8255 18324
rect 8567 18204 8572 18324
rect 8572 18204 8618 18324
rect 8618 18204 8623 18324
rect 8383 17904 8388 18024
rect 8388 17904 8434 18024
rect 8434 17904 8439 18024
rect 8889 18203 8894 18324
rect 8894 18203 8940 18324
rect 8940 18203 8945 18324
rect 8751 17904 8756 18024
rect 8756 17904 8802 18024
rect 8802 17904 8807 18024
rect 8291 17785 8292 17828
rect 8292 17785 8346 17828
rect 8346 17785 8347 17828
rect 8291 17772 8347 17785
rect 8475 17785 8476 17828
rect 8476 17785 8530 17828
rect 8530 17785 8531 17828
rect 8475 17772 8531 17785
rect 8659 17785 8660 17828
rect 8660 17785 8714 17828
rect 8714 17785 8715 17828
rect 8659 17772 8715 17785
rect 8291 17622 8347 17678
rect 7483 17506 7539 17562
rect 8475 17506 8531 17562
rect 8804 17506 8860 17562
rect 9237 17506 9293 17562
rect 6637 17390 6693 17446
rect 8659 17390 8715 17446
rect 8291 17283 8347 17296
rect 8291 17240 8292 17283
rect 8292 17240 8346 17283
rect 8346 17240 8347 17283
rect 8475 17283 8531 17296
rect 8475 17240 8476 17283
rect 8476 17240 8530 17283
rect 8530 17240 8531 17283
rect 8659 17283 8715 17296
rect 8659 17240 8660 17283
rect 8660 17240 8714 17283
rect 8714 17240 8715 17283
rect 8751 17044 8756 17164
rect 8756 17044 8802 17164
rect 8802 17044 8807 17164
rect 8066 16721 8122 16777
rect 8884 16721 8940 16777
rect 3139 16603 3195 16659
rect 3441 16603 3497 16659
rect 11661 19595 11717 19651
rect 12701 19595 12757 19651
rect 9777 19489 9833 19502
rect 9777 19446 9778 19489
rect 9778 19446 9832 19489
rect 9832 19446 9833 19489
rect 9961 19489 10017 19502
rect 9961 19446 9962 19489
rect 9962 19446 10016 19489
rect 10016 19446 10017 19489
rect 10145 19489 10201 19502
rect 10145 19446 10146 19489
rect 10146 19446 10200 19489
rect 10200 19446 10201 19489
rect 10237 19250 10242 19370
rect 10242 19250 10288 19370
rect 10288 19250 10293 19370
rect 9552 18927 9608 18983
rect 10370 18927 10426 18983
rect 14187 19596 14243 19652
rect 12333 19488 12389 19501
rect 12333 19445 12334 19488
rect 12334 19445 12388 19488
rect 12388 19445 12389 19488
rect 12517 19488 12573 19501
rect 12517 19445 12518 19488
rect 12518 19445 12572 19488
rect 12572 19445 12573 19488
rect 12701 19488 12757 19501
rect 12701 19445 12702 19488
rect 12702 19445 12756 19488
rect 12756 19445 12757 19488
rect 12793 19249 12798 19369
rect 12798 19249 12844 19369
rect 12844 19249 12849 19369
rect 12108 18926 12164 18982
rect 12926 18926 12982 18982
rect 13279 18808 13335 18864
rect 13103 18700 13159 18754
rect 12609 18591 12665 18647
rect 12241 18204 12246 18324
rect 12246 18204 12292 18324
rect 12292 18204 12297 18324
rect 12609 18204 12614 18324
rect 12614 18204 12660 18324
rect 12660 18204 12665 18324
rect 12425 17904 12430 18024
rect 12430 17904 12476 18024
rect 12476 17904 12481 18024
rect 12931 18203 12936 18324
rect 12936 18203 12982 18324
rect 12982 18203 12987 18324
rect 12793 17904 12798 18024
rect 12798 17904 12844 18024
rect 12844 17904 12849 18024
rect 12333 17785 12334 17828
rect 12334 17785 12388 17828
rect 12388 17785 12389 17828
rect 12333 17772 12389 17785
rect 12517 17785 12518 17828
rect 12518 17785 12572 17828
rect 12572 17785 12573 17828
rect 12517 17772 12573 17785
rect 12701 17785 12702 17828
rect 12702 17785 12756 17828
rect 12756 17785 12757 17828
rect 12701 17772 12757 17785
rect 12333 17622 12389 17678
rect 11525 17506 11581 17562
rect 12517 17506 12573 17562
rect 12846 17506 12902 17562
rect 13279 17506 13335 17562
rect 10679 17390 10735 17446
rect 12701 17390 12757 17446
rect 12333 17283 12389 17296
rect 12333 17240 12334 17283
rect 12334 17240 12388 17283
rect 12388 17240 12389 17283
rect 12517 17283 12573 17296
rect 12517 17240 12518 17283
rect 12518 17240 12572 17283
rect 12572 17240 12573 17283
rect 12701 17283 12757 17296
rect 12701 17240 12702 17283
rect 12702 17240 12756 17283
rect 12756 17240 12757 17283
rect 12793 17044 12798 17164
rect 12798 17044 12844 17164
rect 12844 17044 12849 17164
rect 12108 16721 12164 16777
rect 12926 16721 12982 16777
rect 7181 16603 7237 16659
rect 7483 16603 7539 16659
rect 15703 19595 15759 19651
rect 16743 19595 16799 19651
rect 13819 19489 13875 19502
rect 13819 19446 13820 19489
rect 13820 19446 13874 19489
rect 13874 19446 13875 19489
rect 14003 19489 14059 19502
rect 14003 19446 14004 19489
rect 14004 19446 14058 19489
rect 14058 19446 14059 19489
rect 14187 19489 14243 19502
rect 14187 19446 14188 19489
rect 14188 19446 14242 19489
rect 14242 19446 14243 19489
rect 14279 19250 14284 19370
rect 14284 19250 14330 19370
rect 14330 19250 14335 19370
rect 13594 18927 13650 18983
rect 14412 18927 14468 18983
rect 18229 19596 18285 19652
rect 16375 19488 16431 19501
rect 16375 19445 16376 19488
rect 16376 19445 16430 19488
rect 16430 19445 16431 19488
rect 16559 19488 16615 19501
rect 16559 19445 16560 19488
rect 16560 19445 16614 19488
rect 16614 19445 16615 19488
rect 16743 19488 16799 19501
rect 16743 19445 16744 19488
rect 16744 19445 16798 19488
rect 16798 19445 16799 19488
rect 16835 19249 16840 19369
rect 16840 19249 16886 19369
rect 16886 19249 16891 19369
rect 16150 18926 16206 18982
rect 16968 18926 17024 18982
rect 17321 18808 17377 18864
rect 17145 18700 17201 18754
rect 16651 18591 16707 18647
rect 16283 18204 16288 18324
rect 16288 18204 16334 18324
rect 16334 18204 16339 18324
rect 16651 18204 16656 18324
rect 16656 18204 16702 18324
rect 16702 18204 16707 18324
rect 16467 17904 16472 18024
rect 16472 17904 16518 18024
rect 16518 17904 16523 18024
rect 16973 18203 16978 18324
rect 16978 18203 17024 18324
rect 17024 18203 17029 18324
rect 16835 17904 16840 18024
rect 16840 17904 16886 18024
rect 16886 17904 16891 18024
rect 16375 17785 16376 17828
rect 16376 17785 16430 17828
rect 16430 17785 16431 17828
rect 16375 17772 16431 17785
rect 16559 17785 16560 17828
rect 16560 17785 16614 17828
rect 16614 17785 16615 17828
rect 16559 17772 16615 17785
rect 16743 17785 16744 17828
rect 16744 17785 16798 17828
rect 16798 17785 16799 17828
rect 16743 17772 16799 17785
rect 16375 17622 16431 17678
rect 15567 17506 15623 17562
rect 16559 17506 16615 17562
rect 16888 17506 16944 17562
rect 17321 17506 17377 17562
rect 15386 17390 15442 17446
rect 16743 17390 16799 17446
rect 16375 17283 16431 17296
rect 16375 17240 16376 17283
rect 16376 17240 16430 17283
rect 16430 17240 16431 17283
rect 16559 17283 16615 17296
rect 16559 17240 16560 17283
rect 16560 17240 16614 17283
rect 16614 17240 16615 17283
rect 16743 17283 16799 17296
rect 16743 17240 16744 17283
rect 16744 17240 16798 17283
rect 16798 17240 16799 17283
rect 16835 17044 16840 17164
rect 16840 17044 16886 17164
rect 16886 17044 16891 17164
rect 16150 16721 16206 16777
rect 16968 16721 17024 16777
rect 11223 16603 11279 16659
rect 11525 16603 11581 16659
rect 17861 19489 17917 19502
rect 17861 19446 17862 19489
rect 17862 19446 17916 19489
rect 17916 19446 17917 19489
rect 18045 19489 18101 19502
rect 18045 19446 18046 19489
rect 18046 19446 18100 19489
rect 18100 19446 18101 19489
rect 18229 19489 18285 19502
rect 18229 19446 18230 19489
rect 18230 19446 18284 19489
rect 18284 19446 18285 19489
rect 18321 19250 18326 19370
rect 18326 19250 18372 19370
rect 18372 19250 18377 19370
rect 17636 18927 17692 18983
rect 18454 18927 18510 18983
rect 15265 16603 15321 16659
rect 15567 16603 15623 16659
rect -11613 15630 -11557 15686
rect -11981 15243 -11976 15363
rect -11976 15243 -11930 15363
rect -11930 15243 -11925 15363
rect -11613 15243 -11608 15363
rect -11608 15243 -11562 15363
rect -11562 15243 -11557 15363
rect -11797 14943 -11792 15063
rect -11792 14943 -11746 15063
rect -11746 14943 -11741 15063
rect -11291 15242 -11286 15363
rect -11286 15242 -11240 15363
rect -11240 15242 -11235 15363
rect -11429 14943 -11424 15063
rect -11424 14943 -11378 15063
rect -11378 14943 -11373 15063
rect -11889 14824 -11888 14867
rect -11888 14824 -11834 14867
rect -11834 14824 -11833 14867
rect -11889 14811 -11833 14824
rect -11705 14824 -11704 14867
rect -11704 14824 -11650 14867
rect -11650 14824 -11649 14867
rect -11705 14811 -11649 14824
rect -11521 14824 -11520 14867
rect -11520 14824 -11466 14867
rect -11466 14824 -11465 14867
rect -11521 14811 -11465 14824
rect -12833 14661 -12777 14717
rect -11889 14661 -11833 14717
rect -12561 14545 -12505 14601
rect -11705 14545 -11649 14601
rect -11376 14545 -11320 14601
rect -11119 14545 -11063 14601
rect -11521 14429 -11465 14485
rect -11889 14322 -11833 14335
rect -11889 14279 -11888 14322
rect -11888 14279 -11834 14322
rect -11834 14279 -11833 14322
rect -11705 14322 -11649 14335
rect -11705 14279 -11704 14322
rect -11704 14279 -11650 14322
rect -11650 14279 -11649 14322
rect -11521 14322 -11465 14335
rect -11521 14279 -11520 14322
rect -11520 14279 -11466 14322
rect -11466 14279 -11465 14322
rect -11429 14083 -11424 14203
rect -11424 14083 -11378 14203
rect -11378 14083 -11373 14203
rect -12114 13760 -12058 13816
rect -11296 13760 -11240 13816
rect -10943 13642 -10887 13698
rect -11119 13534 -11063 13588
rect -11613 13425 -11557 13481
rect -11981 13038 -11976 13158
rect -11976 13038 -11930 13158
rect -11930 13038 -11925 13158
rect -11613 13038 -11608 13158
rect -11608 13038 -11562 13158
rect -11562 13038 -11557 13158
rect -11797 12738 -11792 12858
rect -11792 12738 -11746 12858
rect -11746 12738 -11741 12858
rect -11291 13037 -11286 13158
rect -11286 13037 -11240 13158
rect -11240 13037 -11235 13158
rect -11429 12738 -11424 12858
rect -11424 12738 -11378 12858
rect -11378 12738 -11373 12858
rect -11889 12619 -11888 12662
rect -11888 12619 -11834 12662
rect -11834 12619 -11833 12662
rect -11889 12606 -11833 12619
rect -11705 12619 -11704 12662
rect -11704 12619 -11650 12662
rect -11650 12619 -11649 12662
rect -11705 12606 -11649 12619
rect -11521 12619 -11520 12662
rect -11520 12619 -11466 12662
rect -11466 12619 -11465 12662
rect -11521 12606 -11465 12619
rect -11889 12456 -11833 12512
rect -7601 15630 -7545 15686
rect -7969 15243 -7964 15363
rect -7964 15243 -7918 15363
rect -7918 15243 -7913 15363
rect -7601 15243 -7596 15363
rect -7596 15243 -7550 15363
rect -7550 15243 -7545 15363
rect -7785 14943 -7780 15063
rect -7780 14943 -7734 15063
rect -7734 14943 -7729 15063
rect -7279 15242 -7274 15363
rect -7274 15242 -7228 15363
rect -7228 15242 -7223 15363
rect -7417 14943 -7412 15063
rect -7412 14943 -7366 15063
rect -7366 14943 -7361 15063
rect -7877 14824 -7876 14867
rect -7876 14824 -7822 14867
rect -7822 14824 -7821 14867
rect -7877 14811 -7821 14824
rect -7693 14824 -7692 14867
rect -7692 14824 -7638 14867
rect -7638 14824 -7637 14867
rect -7693 14811 -7637 14824
rect -7509 14824 -7508 14867
rect -7508 14824 -7454 14867
rect -7454 14824 -7453 14867
rect -7509 14811 -7453 14824
rect -8765 14661 -8709 14717
rect -7877 14661 -7821 14717
rect -8549 14545 -8493 14601
rect -7693 14545 -7637 14601
rect -7364 14545 -7308 14601
rect -7107 14545 -7051 14601
rect -7509 14429 -7453 14485
rect -7877 14322 -7821 14335
rect -7877 14279 -7876 14322
rect -7876 14279 -7822 14322
rect -7822 14279 -7821 14322
rect -7693 14322 -7637 14335
rect -7693 14279 -7692 14322
rect -7692 14279 -7638 14322
rect -7638 14279 -7637 14322
rect -7509 14322 -7453 14335
rect -7509 14279 -7508 14322
rect -7508 14279 -7454 14322
rect -7454 14279 -7453 14322
rect -7417 14083 -7412 14203
rect -7412 14083 -7366 14203
rect -7366 14083 -7361 14203
rect -8102 13760 -8046 13816
rect -7284 13760 -7228 13816
rect -6931 13642 -6875 13698
rect -7107 13534 -7051 13588
rect -10127 13425 -10071 13481
rect -10495 13038 -10490 13158
rect -10490 13038 -10444 13158
rect -10444 13038 -10439 13158
rect -10127 13038 -10122 13158
rect -10122 13038 -10076 13158
rect -10076 13038 -10071 13158
rect -10311 12738 -10306 12858
rect -10306 12738 -10260 12858
rect -10260 12738 -10255 12858
rect -9805 13037 -9800 13158
rect -9800 13037 -9754 13158
rect -9754 13037 -9749 13158
rect -9943 12738 -9938 12858
rect -9938 12738 -9892 12858
rect -9892 12738 -9887 12858
rect -10403 12619 -10402 12662
rect -10402 12619 -10348 12662
rect -10348 12619 -10347 12662
rect -10403 12606 -10347 12619
rect -10219 12619 -10218 12662
rect -10218 12619 -10164 12662
rect -10164 12619 -10163 12662
rect -10219 12606 -10163 12619
rect -10035 12619 -10034 12662
rect -10034 12619 -9980 12662
rect -9980 12619 -9979 12662
rect -10035 12606 -9979 12619
rect -10403 12456 -10347 12512
rect -7601 13425 -7545 13481
rect -7969 13038 -7964 13158
rect -7964 13038 -7918 13158
rect -7918 13038 -7913 13158
rect -7601 13038 -7596 13158
rect -7596 13038 -7550 13158
rect -7550 13038 -7545 13158
rect -7785 12738 -7780 12858
rect -7780 12738 -7734 12858
rect -7734 12738 -7729 12858
rect -7279 13037 -7274 13158
rect -7274 13037 -7228 13158
rect -7228 13037 -7223 13158
rect -7417 12738 -7412 12858
rect -7412 12738 -7366 12858
rect -7366 12738 -7361 12858
rect -7877 12619 -7876 12662
rect -7876 12619 -7822 12662
rect -7822 12619 -7821 12662
rect -7877 12606 -7821 12619
rect -7693 12619 -7692 12662
rect -7692 12619 -7638 12662
rect -7638 12619 -7637 12662
rect -7693 12606 -7637 12619
rect -7509 12619 -7508 12662
rect -7508 12619 -7454 12662
rect -7454 12619 -7453 12662
rect -7509 12606 -7453 12619
rect -7877 12456 -7821 12512
rect -3559 15630 -3503 15686
rect -3927 15243 -3922 15363
rect -3922 15243 -3876 15363
rect -3876 15243 -3871 15363
rect -3559 15243 -3554 15363
rect -3554 15243 -3508 15363
rect -3508 15243 -3503 15363
rect -3743 14943 -3738 15063
rect -3738 14943 -3692 15063
rect -3692 14943 -3687 15063
rect -3237 15242 -3232 15363
rect -3232 15242 -3186 15363
rect -3186 15242 -3181 15363
rect -3375 14943 -3370 15063
rect -3370 14943 -3324 15063
rect -3324 14943 -3319 15063
rect -3835 14824 -3834 14867
rect -3834 14824 -3780 14867
rect -3780 14824 -3779 14867
rect -3835 14811 -3779 14824
rect -3651 14824 -3650 14867
rect -3650 14824 -3596 14867
rect -3596 14824 -3595 14867
rect -3651 14811 -3595 14824
rect -3467 14824 -3466 14867
rect -3466 14824 -3412 14867
rect -3412 14824 -3411 14867
rect -3467 14811 -3411 14824
rect -4723 14661 -4667 14717
rect -3835 14661 -3779 14717
rect -4507 14545 -4451 14601
rect -3651 14545 -3595 14601
rect -3322 14545 -3266 14601
rect -3065 14545 -3009 14601
rect -3467 14429 -3411 14485
rect -3835 14322 -3779 14335
rect -3835 14279 -3834 14322
rect -3834 14279 -3780 14322
rect -3780 14279 -3779 14322
rect -3651 14322 -3595 14335
rect -3651 14279 -3650 14322
rect -3650 14279 -3596 14322
rect -3596 14279 -3595 14322
rect -3467 14322 -3411 14335
rect -3467 14279 -3466 14322
rect -3466 14279 -3412 14322
rect -3412 14279 -3411 14322
rect -3375 14083 -3370 14203
rect -3370 14083 -3324 14203
rect -3324 14083 -3319 14203
rect -4060 13760 -4004 13816
rect -3242 13760 -3186 13816
rect -2889 13642 -2833 13698
rect -3065 13534 -3009 13588
rect -6115 13425 -6059 13481
rect -6483 13038 -6478 13158
rect -6478 13038 -6432 13158
rect -6432 13038 -6427 13158
rect -6115 13038 -6110 13158
rect -6110 13038 -6064 13158
rect -6064 13038 -6059 13158
rect -6299 12738 -6294 12858
rect -6294 12738 -6248 12858
rect -6248 12738 -6243 12858
rect -5793 13037 -5788 13158
rect -5788 13037 -5742 13158
rect -5742 13037 -5737 13158
rect -5931 12738 -5926 12858
rect -5926 12738 -5880 12858
rect -5880 12738 -5875 12858
rect -6391 12619 -6390 12662
rect -6390 12619 -6336 12662
rect -6336 12619 -6335 12662
rect -6391 12606 -6335 12619
rect -6207 12619 -6206 12662
rect -6206 12619 -6152 12662
rect -6152 12619 -6151 12662
rect -6207 12606 -6151 12619
rect -6023 12619 -6022 12662
rect -6022 12619 -5968 12662
rect -5968 12619 -5967 12662
rect -6023 12606 -5967 12619
rect -6391 12456 -6335 12512
rect -3559 13425 -3503 13481
rect -3927 13038 -3922 13158
rect -3922 13038 -3876 13158
rect -3876 13038 -3871 13158
rect -3559 13038 -3554 13158
rect -3554 13038 -3508 13158
rect -3508 13038 -3503 13158
rect -3743 12738 -3738 12858
rect -3738 12738 -3692 12858
rect -3692 12738 -3687 12858
rect -3237 13037 -3232 13158
rect -3232 13037 -3186 13158
rect -3186 13037 -3181 13158
rect -3375 12738 -3370 12858
rect -3370 12738 -3324 12858
rect -3324 12738 -3319 12858
rect -3835 12619 -3834 12662
rect -3834 12619 -3780 12662
rect -3780 12619 -3779 12662
rect -3835 12606 -3779 12619
rect -3651 12619 -3650 12662
rect -3650 12619 -3596 12662
rect -3596 12619 -3595 12662
rect -3651 12606 -3595 12619
rect -3467 12619 -3466 12662
rect -3466 12619 -3412 12662
rect -3412 12619 -3411 12662
rect -3467 12606 -3411 12619
rect -3835 12456 -3779 12512
rect 483 15630 539 15686
rect 115 15243 120 15363
rect 120 15243 166 15363
rect 166 15243 171 15363
rect 483 15243 488 15363
rect 488 15243 534 15363
rect 534 15243 539 15363
rect 299 14943 304 15063
rect 304 14943 350 15063
rect 350 14943 355 15063
rect 805 15242 810 15363
rect 810 15242 856 15363
rect 856 15242 861 15363
rect 667 14943 672 15063
rect 672 14943 718 15063
rect 718 14943 723 15063
rect 207 14824 208 14867
rect 208 14824 262 14867
rect 262 14824 263 14867
rect 207 14811 263 14824
rect 391 14824 392 14867
rect 392 14824 446 14867
rect 446 14824 447 14867
rect 391 14811 447 14824
rect 575 14824 576 14867
rect 576 14824 630 14867
rect 630 14824 631 14867
rect 575 14811 631 14824
rect -681 14661 -625 14717
rect 207 14661 263 14717
rect -465 14545 -409 14601
rect 391 14545 447 14601
rect 720 14545 776 14601
rect 977 14545 1033 14601
rect 575 14429 631 14485
rect 207 14322 263 14335
rect 207 14279 208 14322
rect 208 14279 262 14322
rect 262 14279 263 14322
rect 391 14322 447 14335
rect 391 14279 392 14322
rect 392 14279 446 14322
rect 446 14279 447 14322
rect 575 14322 631 14335
rect 575 14279 576 14322
rect 576 14279 630 14322
rect 630 14279 631 14322
rect 667 14083 672 14203
rect 672 14083 718 14203
rect 718 14083 723 14203
rect -18 13760 38 13816
rect 800 13760 856 13816
rect 1153 13642 1209 13698
rect 977 13534 1033 13588
rect -2073 13425 -2017 13481
rect -2441 13038 -2436 13158
rect -2436 13038 -2390 13158
rect -2390 13038 -2385 13158
rect -2073 13038 -2068 13158
rect -2068 13038 -2022 13158
rect -2022 13038 -2017 13158
rect -2257 12738 -2252 12858
rect -2252 12738 -2206 12858
rect -2206 12738 -2201 12858
rect -1751 13037 -1746 13158
rect -1746 13037 -1700 13158
rect -1700 13037 -1695 13158
rect -1889 12738 -1884 12858
rect -1884 12738 -1838 12858
rect -1838 12738 -1833 12858
rect -2349 12619 -2348 12662
rect -2348 12619 -2294 12662
rect -2294 12619 -2293 12662
rect -2349 12606 -2293 12619
rect -2165 12619 -2164 12662
rect -2164 12619 -2110 12662
rect -2110 12619 -2109 12662
rect -2165 12606 -2109 12619
rect -1981 12619 -1980 12662
rect -1980 12619 -1926 12662
rect -1926 12619 -1925 12662
rect -1981 12606 -1925 12619
rect -2349 12456 -2293 12512
rect 483 13425 539 13481
rect 115 13038 120 13158
rect 120 13038 166 13158
rect 166 13038 171 13158
rect 483 13038 488 13158
rect 488 13038 534 13158
rect 534 13038 539 13158
rect 299 12738 304 12858
rect 304 12738 350 12858
rect 350 12738 355 12858
rect 805 13037 810 13158
rect 810 13037 856 13158
rect 856 13037 861 13158
rect 667 12738 672 12858
rect 672 12738 718 12858
rect 718 12738 723 12858
rect 207 12619 208 12662
rect 208 12619 262 12662
rect 262 12619 263 12662
rect 207 12606 263 12619
rect 391 12619 392 12662
rect 392 12619 446 12662
rect 446 12619 447 12662
rect 391 12606 447 12619
rect 575 12619 576 12662
rect 576 12619 630 12662
rect 630 12619 631 12662
rect 575 12606 631 12619
rect 207 12456 263 12512
rect 4525 15630 4581 15686
rect 4157 15243 4162 15363
rect 4162 15243 4208 15363
rect 4208 15243 4213 15363
rect 4525 15243 4530 15363
rect 4530 15243 4576 15363
rect 4576 15243 4581 15363
rect 4341 14943 4346 15063
rect 4346 14943 4392 15063
rect 4392 14943 4397 15063
rect 4847 15242 4852 15363
rect 4852 15242 4898 15363
rect 4898 15242 4903 15363
rect 4709 14943 4714 15063
rect 4714 14943 4760 15063
rect 4760 14943 4765 15063
rect 4249 14824 4250 14867
rect 4250 14824 4304 14867
rect 4304 14824 4305 14867
rect 4249 14811 4305 14824
rect 4433 14824 4434 14867
rect 4434 14824 4488 14867
rect 4488 14824 4489 14867
rect 4433 14811 4489 14824
rect 4617 14824 4618 14867
rect 4618 14824 4672 14867
rect 4672 14824 4673 14867
rect 4617 14811 4673 14824
rect 3361 14661 3417 14717
rect 4249 14661 4305 14717
rect 3577 14545 3633 14601
rect 4433 14545 4489 14601
rect 4762 14545 4818 14601
rect 5019 14545 5075 14601
rect 4617 14429 4673 14485
rect 4249 14322 4305 14335
rect 4249 14279 4250 14322
rect 4250 14279 4304 14322
rect 4304 14279 4305 14322
rect 4433 14322 4489 14335
rect 4433 14279 4434 14322
rect 4434 14279 4488 14322
rect 4488 14279 4489 14322
rect 4617 14322 4673 14335
rect 4617 14279 4618 14322
rect 4618 14279 4672 14322
rect 4672 14279 4673 14322
rect 4709 14083 4714 14203
rect 4714 14083 4760 14203
rect 4760 14083 4765 14203
rect 4024 13760 4080 13816
rect 4842 13760 4898 13816
rect 5195 13642 5251 13698
rect 5019 13534 5075 13588
rect 1969 13425 2025 13481
rect 1601 13038 1606 13158
rect 1606 13038 1652 13158
rect 1652 13038 1657 13158
rect 1969 13038 1974 13158
rect 1974 13038 2020 13158
rect 2020 13038 2025 13158
rect 1785 12738 1790 12858
rect 1790 12738 1836 12858
rect 1836 12738 1841 12858
rect 2291 13037 2296 13158
rect 2296 13037 2342 13158
rect 2342 13037 2347 13158
rect 2153 12738 2158 12858
rect 2158 12738 2204 12858
rect 2204 12738 2209 12858
rect 1693 12619 1694 12662
rect 1694 12619 1748 12662
rect 1748 12619 1749 12662
rect 1693 12606 1749 12619
rect 1877 12619 1878 12662
rect 1878 12619 1932 12662
rect 1932 12619 1933 12662
rect 1877 12606 1933 12619
rect 2061 12619 2062 12662
rect 2062 12619 2116 12662
rect 2116 12619 2117 12662
rect 2061 12606 2117 12619
rect 1693 12456 1749 12512
rect 4525 13425 4581 13481
rect 4157 13038 4162 13158
rect 4162 13038 4208 13158
rect 4208 13038 4213 13158
rect 4525 13038 4530 13158
rect 4530 13038 4576 13158
rect 4576 13038 4581 13158
rect 4341 12738 4346 12858
rect 4346 12738 4392 12858
rect 4392 12738 4397 12858
rect 4847 13037 4852 13158
rect 4852 13037 4898 13158
rect 4898 13037 4903 13158
rect 4709 12738 4714 12858
rect 4714 12738 4760 12858
rect 4760 12738 4765 12858
rect 4249 12619 4250 12662
rect 4250 12619 4304 12662
rect 4304 12619 4305 12662
rect 4249 12606 4305 12619
rect 4433 12619 4434 12662
rect 4434 12619 4488 12662
rect 4488 12619 4489 12662
rect 4433 12606 4489 12619
rect 4617 12619 4618 12662
rect 4618 12619 4672 12662
rect 4672 12619 4673 12662
rect 4617 12606 4673 12619
rect 4249 12456 4305 12512
rect 8567 15630 8623 15686
rect 8199 15243 8204 15363
rect 8204 15243 8250 15363
rect 8250 15243 8255 15363
rect 8567 15243 8572 15363
rect 8572 15243 8618 15363
rect 8618 15243 8623 15363
rect 8383 14943 8388 15063
rect 8388 14943 8434 15063
rect 8434 14943 8439 15063
rect 8889 15242 8894 15363
rect 8894 15242 8940 15363
rect 8940 15242 8945 15363
rect 8751 14943 8756 15063
rect 8756 14943 8802 15063
rect 8802 14943 8807 15063
rect 8291 14824 8292 14867
rect 8292 14824 8346 14867
rect 8346 14824 8347 14867
rect 8291 14811 8347 14824
rect 8475 14824 8476 14867
rect 8476 14824 8530 14867
rect 8530 14824 8531 14867
rect 8475 14811 8531 14824
rect 8659 14824 8660 14867
rect 8660 14824 8714 14867
rect 8714 14824 8715 14867
rect 8659 14811 8715 14824
rect 7403 14661 7459 14717
rect 8291 14661 8347 14717
rect 7619 14545 7675 14601
rect 8475 14545 8531 14601
rect 8804 14545 8860 14601
rect 9061 14545 9117 14601
rect 8659 14429 8715 14485
rect 8291 14322 8347 14335
rect 8291 14279 8292 14322
rect 8292 14279 8346 14322
rect 8346 14279 8347 14322
rect 8475 14322 8531 14335
rect 8475 14279 8476 14322
rect 8476 14279 8530 14322
rect 8530 14279 8531 14322
rect 8659 14322 8715 14335
rect 8659 14279 8660 14322
rect 8660 14279 8714 14322
rect 8714 14279 8715 14322
rect 8751 14083 8756 14203
rect 8756 14083 8802 14203
rect 8802 14083 8807 14203
rect 8066 13760 8122 13816
rect 8884 13760 8940 13816
rect 9237 13642 9293 13698
rect 9061 13534 9117 13588
rect 6011 13425 6067 13481
rect 5643 13038 5648 13158
rect 5648 13038 5694 13158
rect 5694 13038 5699 13158
rect 6011 13038 6016 13158
rect 6016 13038 6062 13158
rect 6062 13038 6067 13158
rect 5827 12738 5832 12858
rect 5832 12738 5878 12858
rect 5878 12738 5883 12858
rect 6333 13037 6338 13158
rect 6338 13037 6384 13158
rect 6384 13037 6389 13158
rect 6195 12738 6200 12858
rect 6200 12738 6246 12858
rect 6246 12738 6251 12858
rect 5735 12619 5736 12662
rect 5736 12619 5790 12662
rect 5790 12619 5791 12662
rect 5735 12606 5791 12619
rect 5919 12619 5920 12662
rect 5920 12619 5974 12662
rect 5974 12619 5975 12662
rect 5919 12606 5975 12619
rect 6103 12619 6104 12662
rect 6104 12619 6158 12662
rect 6158 12619 6159 12662
rect 6103 12606 6159 12619
rect 5735 12456 5791 12512
rect 8567 13425 8623 13481
rect 8199 13038 8204 13158
rect 8204 13038 8250 13158
rect 8250 13038 8255 13158
rect 8567 13038 8572 13158
rect 8572 13038 8618 13158
rect 8618 13038 8623 13158
rect 8383 12738 8388 12858
rect 8388 12738 8434 12858
rect 8434 12738 8439 12858
rect 8889 13037 8894 13158
rect 8894 13037 8940 13158
rect 8940 13037 8945 13158
rect 8751 12738 8756 12858
rect 8756 12738 8802 12858
rect 8802 12738 8807 12858
rect 8291 12619 8292 12662
rect 8292 12619 8346 12662
rect 8346 12619 8347 12662
rect 8291 12606 8347 12619
rect 8475 12619 8476 12662
rect 8476 12619 8530 12662
rect 8530 12619 8531 12662
rect 8475 12606 8531 12619
rect 8659 12619 8660 12662
rect 8660 12619 8714 12662
rect 8714 12619 8715 12662
rect 8659 12606 8715 12619
rect 8291 12456 8347 12512
rect 12609 15630 12665 15686
rect 12241 15243 12246 15363
rect 12246 15243 12292 15363
rect 12292 15243 12297 15363
rect 12609 15243 12614 15363
rect 12614 15243 12660 15363
rect 12660 15243 12665 15363
rect 12425 14943 12430 15063
rect 12430 14943 12476 15063
rect 12476 14943 12481 15063
rect 12931 15242 12936 15363
rect 12936 15242 12982 15363
rect 12982 15242 12987 15363
rect 12793 14943 12798 15063
rect 12798 14943 12844 15063
rect 12844 14943 12849 15063
rect 12333 14824 12334 14867
rect 12334 14824 12388 14867
rect 12388 14824 12389 14867
rect 12333 14811 12389 14824
rect 12517 14824 12518 14867
rect 12518 14824 12572 14867
rect 12572 14824 12573 14867
rect 12517 14811 12573 14824
rect 12701 14824 12702 14867
rect 12702 14824 12756 14867
rect 12756 14824 12757 14867
rect 12701 14811 12757 14824
rect 11445 14661 11501 14717
rect 12333 14661 12389 14717
rect 11661 14545 11717 14601
rect 12517 14545 12573 14601
rect 12846 14545 12902 14601
rect 13103 14545 13159 14601
rect 12701 14429 12757 14485
rect 12333 14322 12389 14335
rect 12333 14279 12334 14322
rect 12334 14279 12388 14322
rect 12388 14279 12389 14322
rect 12517 14322 12573 14335
rect 12517 14279 12518 14322
rect 12518 14279 12572 14322
rect 12572 14279 12573 14322
rect 12701 14322 12757 14335
rect 12701 14279 12702 14322
rect 12702 14279 12756 14322
rect 12756 14279 12757 14322
rect 12793 14083 12798 14203
rect 12798 14083 12844 14203
rect 12844 14083 12849 14203
rect 12108 13760 12164 13816
rect 12926 13760 12982 13816
rect 13279 13642 13335 13698
rect 13103 13534 13159 13588
rect 10053 13425 10109 13481
rect 9685 13038 9690 13158
rect 9690 13038 9736 13158
rect 9736 13038 9741 13158
rect 10053 13038 10058 13158
rect 10058 13038 10104 13158
rect 10104 13038 10109 13158
rect 9869 12738 9874 12858
rect 9874 12738 9920 12858
rect 9920 12738 9925 12858
rect 10375 13037 10380 13158
rect 10380 13037 10426 13158
rect 10426 13037 10431 13158
rect 10237 12738 10242 12858
rect 10242 12738 10288 12858
rect 10288 12738 10293 12858
rect 9777 12619 9778 12662
rect 9778 12619 9832 12662
rect 9832 12619 9833 12662
rect 9777 12606 9833 12619
rect 9961 12619 9962 12662
rect 9962 12619 10016 12662
rect 10016 12619 10017 12662
rect 9961 12606 10017 12619
rect 10145 12619 10146 12662
rect 10146 12619 10200 12662
rect 10200 12619 10201 12662
rect 10145 12606 10201 12619
rect 9777 12456 9833 12512
rect 12609 13425 12665 13481
rect 12241 13038 12246 13158
rect 12246 13038 12292 13158
rect 12292 13038 12297 13158
rect 12609 13038 12614 13158
rect 12614 13038 12660 13158
rect 12660 13038 12665 13158
rect 12425 12738 12430 12858
rect 12430 12738 12476 12858
rect 12476 12738 12481 12858
rect 12931 13037 12936 13158
rect 12936 13037 12982 13158
rect 12982 13037 12987 13158
rect 12793 12738 12798 12858
rect 12798 12738 12844 12858
rect 12844 12738 12849 12858
rect 12333 12619 12334 12662
rect 12334 12619 12388 12662
rect 12388 12619 12389 12662
rect 12333 12606 12389 12619
rect 12517 12619 12518 12662
rect 12518 12619 12572 12662
rect 12572 12619 12573 12662
rect 12517 12606 12573 12619
rect 12701 12619 12702 12662
rect 12702 12619 12756 12662
rect 12756 12619 12757 12662
rect 12701 12606 12757 12619
rect 12333 12456 12389 12512
rect 14095 13425 14151 13481
rect 13727 13038 13732 13158
rect 13732 13038 13778 13158
rect 13778 13038 13783 13158
rect 14095 13038 14100 13158
rect 14100 13038 14146 13158
rect 14146 13038 14151 13158
rect 13911 12738 13916 12858
rect 13916 12738 13962 12858
rect 13962 12738 13967 12858
rect 14417 13037 14422 13158
rect 14422 13037 14468 13158
rect 14468 13037 14473 13158
rect 14279 12738 14284 12858
rect 14284 12738 14330 12858
rect 14330 12738 14335 12858
rect 13819 12619 13820 12662
rect 13820 12619 13874 12662
rect 13874 12619 13875 12662
rect 13819 12606 13875 12619
rect 14003 12619 14004 12662
rect 14004 12619 14058 12662
rect 14058 12619 14059 12662
rect 14003 12606 14059 12619
rect 14187 12619 14188 12662
rect 14188 12619 14242 12662
rect 14242 12619 14243 12662
rect 14187 12606 14243 12619
rect 13819 12456 13875 12512
rect -12697 12340 -12641 12396
rect -11705 12340 -11649 12396
rect -11376 12340 -11320 12396
rect -10943 12340 -10887 12396
rect -10219 12340 -10163 12396
rect -9890 12340 -9834 12396
rect -9633 12340 -9577 12396
rect -11521 12224 -11465 12280
rect -10035 12224 -9979 12280
rect -11889 12117 -11833 12130
rect -11889 12074 -11888 12117
rect -11888 12074 -11834 12117
rect -11834 12074 -11833 12117
rect -11705 12117 -11649 12130
rect -11705 12074 -11704 12117
rect -11704 12074 -11650 12117
rect -11650 12074 -11649 12117
rect -11521 12117 -11465 12130
rect -11521 12074 -11520 12117
rect -11520 12074 -11466 12117
rect -11466 12074 -11465 12117
rect -11429 11878 -11424 11998
rect -11424 11878 -11378 11998
rect -11378 11878 -11373 11998
rect -12114 11555 -12058 11611
rect -11296 11555 -11240 11611
rect -13105 11438 -13049 11494
rect -8685 12340 -8629 12396
rect -7693 12340 -7637 12396
rect -7364 12340 -7308 12396
rect -6931 12340 -6875 12396
rect -6207 12340 -6151 12396
rect -5878 12340 -5822 12396
rect -5621 12340 -5565 12396
rect -7509 12224 -7453 12280
rect -8821 12152 -8765 12208
rect -10403 12117 -10347 12130
rect -10403 12074 -10402 12117
rect -10402 12074 -10348 12117
rect -10348 12074 -10347 12117
rect -10219 12117 -10163 12130
rect -10219 12074 -10218 12117
rect -10218 12074 -10164 12117
rect -10164 12074 -10163 12117
rect -10035 12117 -9979 12130
rect -10035 12074 -10034 12117
rect -10034 12074 -9980 12117
rect -9980 12074 -9979 12117
rect -9943 11878 -9938 11998
rect -9938 11878 -9892 11998
rect -9892 11878 -9887 11998
rect -10628 11555 -10572 11611
rect -9810 11555 -9754 11611
rect -9457 11438 -9401 11494
rect -6023 12224 -5967 12280
rect -7877 12117 -7821 12130
rect -7877 12074 -7876 12117
rect -7876 12074 -7822 12117
rect -7822 12074 -7821 12117
rect -7693 12117 -7637 12130
rect -7693 12074 -7692 12117
rect -7692 12074 -7638 12117
rect -7638 12074 -7637 12117
rect -7509 12117 -7453 12130
rect -7509 12074 -7508 12117
rect -7508 12074 -7454 12117
rect -7454 12074 -7453 12117
rect -7417 11878 -7412 11998
rect -7412 11878 -7366 11998
rect -7366 11878 -7361 11998
rect -8102 11555 -8046 11611
rect -7284 11555 -7228 11611
rect -9093 11438 -9037 11494
rect -4643 12340 -4587 12396
rect -3651 12340 -3595 12396
rect -3322 12340 -3266 12396
rect -2889 12340 -2833 12396
rect -2165 12340 -2109 12396
rect -1836 12340 -1780 12396
rect -1579 12340 -1523 12396
rect -3467 12224 -3411 12280
rect -4809 12152 -4753 12208
rect -6391 12117 -6335 12130
rect -6391 12074 -6390 12117
rect -6390 12074 -6336 12117
rect -6336 12074 -6335 12117
rect -6207 12117 -6151 12130
rect -6207 12074 -6206 12117
rect -6206 12074 -6152 12117
rect -6152 12074 -6151 12117
rect -6023 12117 -5967 12130
rect -6023 12074 -6022 12117
rect -6022 12074 -5968 12117
rect -5968 12074 -5967 12117
rect -5931 11878 -5926 11998
rect -5926 11878 -5880 11998
rect -5880 11878 -5875 11998
rect -6616 11555 -6560 11611
rect -5798 11555 -5742 11611
rect -5445 11438 -5389 11494
rect -10943 11327 -10887 11383
rect -9633 11328 -9577 11384
rect -11613 11220 -11557 11276
rect -11981 10833 -11976 10953
rect -11976 10833 -11930 10953
rect -11930 10833 -11925 10953
rect -11613 10833 -11608 10953
rect -11608 10833 -11562 10953
rect -11562 10833 -11557 10953
rect -11797 10533 -11792 10653
rect -11792 10533 -11746 10653
rect -11746 10533 -11741 10653
rect -11291 10832 -11286 10953
rect -11286 10832 -11240 10953
rect -11240 10832 -11235 10953
rect -11429 10533 -11424 10653
rect -11424 10533 -11378 10653
rect -11378 10533 -11373 10653
rect -11889 10414 -11888 10457
rect -11888 10414 -11834 10457
rect -11834 10414 -11833 10457
rect -11889 10401 -11833 10414
rect -11705 10414 -11704 10457
rect -11704 10414 -11650 10457
rect -11650 10414 -11649 10457
rect -11705 10401 -11649 10414
rect -11521 10414 -11520 10457
rect -11520 10414 -11466 10457
rect -11466 10414 -11465 10457
rect -11521 10401 -11465 10414
rect -11889 10251 -11833 10307
rect -10127 11221 -10071 11277
rect -10495 10834 -10490 10954
rect -10490 10834 -10444 10954
rect -10444 10834 -10439 10954
rect -10127 10834 -10122 10954
rect -10122 10834 -10076 10954
rect -10076 10834 -10071 10954
rect -10311 10534 -10306 10654
rect -10306 10534 -10260 10654
rect -10260 10534 -10255 10654
rect -9805 10833 -9800 10954
rect -9800 10833 -9754 10954
rect -9754 10833 -9749 10954
rect -9943 10534 -9938 10654
rect -9938 10534 -9892 10654
rect -9892 10534 -9887 10654
rect -10403 10415 -10402 10458
rect -10402 10415 -10348 10458
rect -10348 10415 -10347 10458
rect -10403 10402 -10347 10415
rect -10219 10415 -10218 10458
rect -10218 10415 -10164 10458
rect -10164 10415 -10163 10458
rect -10219 10402 -10163 10415
rect -10035 10415 -10034 10458
rect -10034 10415 -9980 10458
rect -9980 10415 -9979 10458
rect -10035 10402 -9979 10415
rect -10403 10252 -10347 10308
rect -11705 10135 -11649 10191
rect -11376 10135 -11320 10191
rect -11119 10135 -11063 10191
rect -10219 10136 -10163 10192
rect -9890 10136 -9834 10192
rect -9457 10136 -9401 10192
rect -1981 12224 -1925 12280
rect -3835 12117 -3779 12130
rect -3835 12074 -3834 12117
rect -3834 12074 -3780 12117
rect -3780 12074 -3779 12117
rect -3651 12117 -3595 12130
rect -3651 12074 -3650 12117
rect -3650 12074 -3596 12117
rect -3596 12074 -3595 12117
rect -3467 12117 -3411 12130
rect -3467 12074 -3466 12117
rect -3466 12074 -3412 12117
rect -3412 12074 -3411 12117
rect -3375 11878 -3370 11998
rect -3370 11878 -3324 11998
rect -3324 11878 -3319 11998
rect -4060 11555 -4004 11611
rect -3242 11555 -3186 11611
rect -5081 11438 -5025 11494
rect -601 12340 -545 12396
rect 391 12340 447 12396
rect 720 12340 776 12396
rect 1153 12340 1209 12396
rect 1877 12340 1933 12396
rect 2206 12340 2262 12396
rect 2463 12340 2519 12396
rect 575 12224 631 12280
rect -767 12152 -711 12208
rect -2349 12117 -2293 12130
rect -2349 12074 -2348 12117
rect -2348 12074 -2294 12117
rect -2294 12074 -2293 12117
rect -2165 12117 -2109 12130
rect -2165 12074 -2164 12117
rect -2164 12074 -2110 12117
rect -2110 12074 -2109 12117
rect -1981 12117 -1925 12130
rect -1981 12074 -1980 12117
rect -1980 12074 -1926 12117
rect -1926 12074 -1925 12117
rect -1889 11878 -1884 11998
rect -1884 11878 -1838 11998
rect -1838 11878 -1833 11998
rect -2574 11555 -2518 11611
rect -1756 11555 -1700 11611
rect -1403 11438 -1347 11494
rect -6931 11327 -6875 11383
rect -5621 11328 -5565 11384
rect -7601 11220 -7545 11276
rect -7969 10833 -7964 10953
rect -7964 10833 -7918 10953
rect -7918 10833 -7913 10953
rect -7601 10833 -7596 10953
rect -7596 10833 -7550 10953
rect -7550 10833 -7545 10953
rect -7785 10533 -7780 10653
rect -7780 10533 -7734 10653
rect -7734 10533 -7729 10653
rect -7279 10832 -7274 10953
rect -7274 10832 -7228 10953
rect -7228 10832 -7223 10953
rect -7417 10533 -7412 10653
rect -7412 10533 -7366 10653
rect -7366 10533 -7361 10653
rect -7877 10414 -7876 10457
rect -7876 10414 -7822 10457
rect -7822 10414 -7821 10457
rect -7877 10401 -7821 10414
rect -7693 10414 -7692 10457
rect -7692 10414 -7638 10457
rect -7638 10414 -7637 10457
rect -7693 10401 -7637 10414
rect -7509 10414 -7508 10457
rect -7508 10414 -7454 10457
rect -7454 10414 -7453 10457
rect -7509 10401 -7453 10414
rect -7877 10251 -7821 10307
rect -6115 11221 -6059 11277
rect -6483 10834 -6478 10954
rect -6478 10834 -6432 10954
rect -6432 10834 -6427 10954
rect -6115 10834 -6110 10954
rect -6110 10834 -6064 10954
rect -6064 10834 -6059 10954
rect -6299 10534 -6294 10654
rect -6294 10534 -6248 10654
rect -6248 10534 -6243 10654
rect -5793 10833 -5788 10954
rect -5788 10833 -5742 10954
rect -5742 10833 -5737 10954
rect -5931 10534 -5926 10654
rect -5926 10534 -5880 10654
rect -5880 10534 -5875 10654
rect -6391 10415 -6390 10458
rect -6390 10415 -6336 10458
rect -6336 10415 -6335 10458
rect -6391 10402 -6335 10415
rect -6207 10415 -6206 10458
rect -6206 10415 -6152 10458
rect -6152 10415 -6151 10458
rect -6207 10402 -6151 10415
rect -6023 10415 -6022 10458
rect -6022 10415 -5968 10458
rect -5968 10415 -5967 10458
rect -6023 10402 -5967 10415
rect -6391 10252 -6335 10308
rect -7693 10135 -7637 10191
rect -7364 10135 -7308 10191
rect -7107 10135 -7051 10191
rect -6207 10136 -6151 10192
rect -5878 10136 -5822 10192
rect -5445 10136 -5389 10192
rect 2061 12224 2117 12280
rect 207 12117 263 12130
rect 207 12074 208 12117
rect 208 12074 262 12117
rect 262 12074 263 12117
rect 391 12117 447 12130
rect 391 12074 392 12117
rect 392 12074 446 12117
rect 446 12074 447 12117
rect 575 12117 631 12130
rect 575 12074 576 12117
rect 576 12074 630 12117
rect 630 12074 631 12117
rect 667 11878 672 11998
rect 672 11878 718 11998
rect 718 11878 723 11998
rect -18 11555 38 11611
rect 800 11555 856 11611
rect -1039 11438 -983 11494
rect 3441 12340 3497 12396
rect 4433 12340 4489 12396
rect 4762 12340 4818 12396
rect 5195 12340 5251 12396
rect 5919 12340 5975 12396
rect 6248 12340 6304 12396
rect 6505 12340 6561 12396
rect 4617 12224 4673 12280
rect 3275 12152 3331 12208
rect 1693 12117 1749 12130
rect 1693 12074 1694 12117
rect 1694 12074 1748 12117
rect 1748 12074 1749 12117
rect 1877 12117 1933 12130
rect 1877 12074 1878 12117
rect 1878 12074 1932 12117
rect 1932 12074 1933 12117
rect 2061 12117 2117 12130
rect 2061 12074 2062 12117
rect 2062 12074 2116 12117
rect 2116 12074 2117 12117
rect 2153 11878 2158 11998
rect 2158 11878 2204 11998
rect 2204 11878 2209 11998
rect 1468 11555 1524 11611
rect 2286 11555 2342 11611
rect 2639 11438 2695 11494
rect -2889 11327 -2833 11383
rect -1579 11328 -1523 11384
rect -3559 11220 -3503 11276
rect -3927 10833 -3922 10953
rect -3922 10833 -3876 10953
rect -3876 10833 -3871 10953
rect -3559 10833 -3554 10953
rect -3554 10833 -3508 10953
rect -3508 10833 -3503 10953
rect -3743 10533 -3738 10653
rect -3738 10533 -3692 10653
rect -3692 10533 -3687 10653
rect -3237 10832 -3232 10953
rect -3232 10832 -3186 10953
rect -3186 10832 -3181 10953
rect -3375 10533 -3370 10653
rect -3370 10533 -3324 10653
rect -3324 10533 -3319 10653
rect -3835 10414 -3834 10457
rect -3834 10414 -3780 10457
rect -3780 10414 -3779 10457
rect -3835 10401 -3779 10414
rect -3651 10414 -3650 10457
rect -3650 10414 -3596 10457
rect -3596 10414 -3595 10457
rect -3651 10401 -3595 10414
rect -3467 10414 -3466 10457
rect -3466 10414 -3412 10457
rect -3412 10414 -3411 10457
rect -3467 10401 -3411 10414
rect -3835 10251 -3779 10307
rect -2073 11221 -2017 11277
rect -2441 10834 -2436 10954
rect -2436 10834 -2390 10954
rect -2390 10834 -2385 10954
rect -2073 10834 -2068 10954
rect -2068 10834 -2022 10954
rect -2022 10834 -2017 10954
rect -2257 10534 -2252 10654
rect -2252 10534 -2206 10654
rect -2206 10534 -2201 10654
rect -1751 10833 -1746 10954
rect -1746 10833 -1700 10954
rect -1700 10833 -1695 10954
rect -1889 10534 -1884 10654
rect -1884 10534 -1838 10654
rect -1838 10534 -1833 10654
rect -2349 10415 -2348 10458
rect -2348 10415 -2294 10458
rect -2294 10415 -2293 10458
rect -2349 10402 -2293 10415
rect -2165 10415 -2164 10458
rect -2164 10415 -2110 10458
rect -2110 10415 -2109 10458
rect -2165 10402 -2109 10415
rect -1981 10415 -1980 10458
rect -1980 10415 -1926 10458
rect -1926 10415 -1925 10458
rect -1981 10402 -1925 10415
rect -2349 10252 -2293 10308
rect -3651 10135 -3595 10191
rect -3322 10135 -3266 10191
rect -3065 10135 -3009 10191
rect -2165 10136 -2109 10192
rect -1836 10136 -1780 10192
rect -1403 10136 -1347 10192
rect 6103 12224 6159 12280
rect 4249 12117 4305 12130
rect 4249 12074 4250 12117
rect 4250 12074 4304 12117
rect 4304 12074 4305 12117
rect 4433 12117 4489 12130
rect 4433 12074 4434 12117
rect 4434 12074 4488 12117
rect 4488 12074 4489 12117
rect 4617 12117 4673 12130
rect 4617 12074 4618 12117
rect 4618 12074 4672 12117
rect 4672 12074 4673 12117
rect 4709 11878 4714 11998
rect 4714 11878 4760 11998
rect 4760 11878 4765 11998
rect 4024 11555 4080 11611
rect 4842 11555 4898 11611
rect 3003 11438 3059 11494
rect 7483 12340 7539 12396
rect 8475 12340 8531 12396
rect 8804 12340 8860 12396
rect 9237 12340 9293 12396
rect 9961 12340 10017 12396
rect 10290 12340 10346 12396
rect 10547 12340 10603 12396
rect 8659 12224 8715 12280
rect 7317 12152 7373 12208
rect 5735 12117 5791 12130
rect 5735 12074 5736 12117
rect 5736 12074 5790 12117
rect 5790 12074 5791 12117
rect 5919 12117 5975 12130
rect 5919 12074 5920 12117
rect 5920 12074 5974 12117
rect 5974 12074 5975 12117
rect 6103 12117 6159 12130
rect 6103 12074 6104 12117
rect 6104 12074 6158 12117
rect 6158 12074 6159 12117
rect 6195 11878 6200 11998
rect 6200 11878 6246 11998
rect 6246 11878 6251 11998
rect 5510 11555 5566 11611
rect 6328 11555 6384 11611
rect 6681 11438 6737 11494
rect 1153 11327 1209 11383
rect 2463 11328 2519 11384
rect 483 11220 539 11276
rect 115 10833 120 10953
rect 120 10833 166 10953
rect 166 10833 171 10953
rect 483 10833 488 10953
rect 488 10833 534 10953
rect 534 10833 539 10953
rect 299 10533 304 10653
rect 304 10533 350 10653
rect 350 10533 355 10653
rect 805 10832 810 10953
rect 810 10832 856 10953
rect 856 10832 861 10953
rect 667 10533 672 10653
rect 672 10533 718 10653
rect 718 10533 723 10653
rect 207 10414 208 10457
rect 208 10414 262 10457
rect 262 10414 263 10457
rect 207 10401 263 10414
rect 391 10414 392 10457
rect 392 10414 446 10457
rect 446 10414 447 10457
rect 391 10401 447 10414
rect 575 10414 576 10457
rect 576 10414 630 10457
rect 630 10414 631 10457
rect 575 10401 631 10414
rect 207 10251 263 10307
rect 1969 11221 2025 11277
rect 1601 10834 1606 10954
rect 1606 10834 1652 10954
rect 1652 10834 1657 10954
rect 1969 10834 1974 10954
rect 1974 10834 2020 10954
rect 2020 10834 2025 10954
rect 1785 10534 1790 10654
rect 1790 10534 1836 10654
rect 1836 10534 1841 10654
rect 2291 10833 2296 10954
rect 2296 10833 2342 10954
rect 2342 10833 2347 10954
rect 2153 10534 2158 10654
rect 2158 10534 2204 10654
rect 2204 10534 2209 10654
rect 1693 10415 1694 10458
rect 1694 10415 1748 10458
rect 1748 10415 1749 10458
rect 1693 10402 1749 10415
rect 1877 10415 1878 10458
rect 1878 10415 1932 10458
rect 1932 10415 1933 10458
rect 1877 10402 1933 10415
rect 2061 10415 2062 10458
rect 2062 10415 2116 10458
rect 2116 10415 2117 10458
rect 2061 10402 2117 10415
rect 1693 10252 1749 10308
rect 391 10135 447 10191
rect 720 10135 776 10191
rect 977 10135 1033 10191
rect 1877 10136 1933 10192
rect 2206 10136 2262 10192
rect 2639 10136 2695 10192
rect 10145 12224 10201 12280
rect 8291 12117 8347 12130
rect 8291 12074 8292 12117
rect 8292 12074 8346 12117
rect 8346 12074 8347 12117
rect 8475 12117 8531 12130
rect 8475 12074 8476 12117
rect 8476 12074 8530 12117
rect 8530 12074 8531 12117
rect 8659 12117 8715 12130
rect 8659 12074 8660 12117
rect 8660 12074 8714 12117
rect 8714 12074 8715 12117
rect 8751 11878 8756 11998
rect 8756 11878 8802 11998
rect 8802 11878 8807 11998
rect 8066 11555 8122 11611
rect 8884 11555 8940 11611
rect 7045 11438 7101 11494
rect 11525 12340 11581 12396
rect 12517 12340 12573 12396
rect 12846 12340 12902 12396
rect 13279 12340 13335 12396
rect 14003 12340 14059 12396
rect 14332 12340 14388 12396
rect 14589 12340 14645 12396
rect 12701 12224 12757 12280
rect 11359 12152 11415 12208
rect 9777 12117 9833 12130
rect 9777 12074 9778 12117
rect 9778 12074 9832 12117
rect 9832 12074 9833 12117
rect 9961 12117 10017 12130
rect 9961 12074 9962 12117
rect 9962 12074 10016 12117
rect 10016 12074 10017 12117
rect 10145 12117 10201 12130
rect 10145 12074 10146 12117
rect 10146 12074 10200 12117
rect 10200 12074 10201 12117
rect 10237 11878 10242 11998
rect 10242 11878 10288 11998
rect 10288 11878 10293 11998
rect 9552 11555 9608 11611
rect 10370 11555 10426 11611
rect 10723 11438 10779 11494
rect 5195 11327 5251 11383
rect 6505 11328 6561 11384
rect 4525 11220 4581 11276
rect 4157 10833 4162 10953
rect 4162 10833 4208 10953
rect 4208 10833 4213 10953
rect 4525 10833 4530 10953
rect 4530 10833 4576 10953
rect 4576 10833 4581 10953
rect 4341 10533 4346 10653
rect 4346 10533 4392 10653
rect 4392 10533 4397 10653
rect 4847 10832 4852 10953
rect 4852 10832 4898 10953
rect 4898 10832 4903 10953
rect 4709 10533 4714 10653
rect 4714 10533 4760 10653
rect 4760 10533 4765 10653
rect 4249 10414 4250 10457
rect 4250 10414 4304 10457
rect 4304 10414 4305 10457
rect 4249 10401 4305 10414
rect 4433 10414 4434 10457
rect 4434 10414 4488 10457
rect 4488 10414 4489 10457
rect 4433 10401 4489 10414
rect 4617 10414 4618 10457
rect 4618 10414 4672 10457
rect 4672 10414 4673 10457
rect 4617 10401 4673 10414
rect 4249 10251 4305 10307
rect 6011 11221 6067 11277
rect 5643 10834 5648 10954
rect 5648 10834 5694 10954
rect 5694 10834 5699 10954
rect 6011 10834 6016 10954
rect 6016 10834 6062 10954
rect 6062 10834 6067 10954
rect 5827 10534 5832 10654
rect 5832 10534 5878 10654
rect 5878 10534 5883 10654
rect 6333 10833 6338 10954
rect 6338 10833 6384 10954
rect 6384 10833 6389 10954
rect 6195 10534 6200 10654
rect 6200 10534 6246 10654
rect 6246 10534 6251 10654
rect 5735 10415 5736 10458
rect 5736 10415 5790 10458
rect 5790 10415 5791 10458
rect 5735 10402 5791 10415
rect 5919 10415 5920 10458
rect 5920 10415 5974 10458
rect 5974 10415 5975 10458
rect 5919 10402 5975 10415
rect 6103 10415 6104 10458
rect 6104 10415 6158 10458
rect 6158 10415 6159 10458
rect 6103 10402 6159 10415
rect 5735 10252 5791 10308
rect 4433 10135 4489 10191
rect 4762 10135 4818 10191
rect 5019 10135 5075 10191
rect 5919 10136 5975 10192
rect 6248 10136 6304 10192
rect 6681 10136 6737 10192
rect 14187 12224 14243 12280
rect 12333 12117 12389 12130
rect 12333 12074 12334 12117
rect 12334 12074 12388 12117
rect 12388 12074 12389 12117
rect 12517 12117 12573 12130
rect 12517 12074 12518 12117
rect 12518 12074 12572 12117
rect 12572 12074 12573 12117
rect 12701 12117 12757 12130
rect 12701 12074 12702 12117
rect 12702 12074 12756 12117
rect 12756 12074 12757 12117
rect 12793 11878 12798 11998
rect 12798 11878 12844 11998
rect 12844 11878 12849 11998
rect 12108 11555 12164 11611
rect 12926 11555 12982 11611
rect 11087 11438 11143 11494
rect 13819 12117 13875 12130
rect 13819 12074 13820 12117
rect 13820 12074 13874 12117
rect 13874 12074 13875 12117
rect 14003 12117 14059 12130
rect 14003 12074 14004 12117
rect 14004 12074 14058 12117
rect 14058 12074 14059 12117
rect 14187 12117 14243 12130
rect 14187 12074 14188 12117
rect 14188 12074 14242 12117
rect 14242 12074 14243 12117
rect 14279 11878 14284 11998
rect 14284 11878 14330 11998
rect 14330 11878 14335 11998
rect 13594 11555 13650 11611
rect 14412 11555 14468 11611
rect 14765 11438 14821 11494
rect 9237 11327 9293 11383
rect 10547 11328 10603 11384
rect 8567 11220 8623 11276
rect 8199 10833 8204 10953
rect 8204 10833 8250 10953
rect 8250 10833 8255 10953
rect 8567 10833 8572 10953
rect 8572 10833 8618 10953
rect 8618 10833 8623 10953
rect 8383 10533 8388 10653
rect 8388 10533 8434 10653
rect 8434 10533 8439 10653
rect 8889 10832 8894 10953
rect 8894 10832 8940 10953
rect 8940 10832 8945 10953
rect 8751 10533 8756 10653
rect 8756 10533 8802 10653
rect 8802 10533 8807 10653
rect 8291 10414 8292 10457
rect 8292 10414 8346 10457
rect 8346 10414 8347 10457
rect 8291 10401 8347 10414
rect 8475 10414 8476 10457
rect 8476 10414 8530 10457
rect 8530 10414 8531 10457
rect 8475 10401 8531 10414
rect 8659 10414 8660 10457
rect 8660 10414 8714 10457
rect 8714 10414 8715 10457
rect 8659 10401 8715 10414
rect 8291 10251 8347 10307
rect 10053 11221 10109 11277
rect 9685 10834 9690 10954
rect 9690 10834 9736 10954
rect 9736 10834 9741 10954
rect 10053 10834 10058 10954
rect 10058 10834 10104 10954
rect 10104 10834 10109 10954
rect 9869 10534 9874 10654
rect 9874 10534 9920 10654
rect 9920 10534 9925 10654
rect 10375 10833 10380 10954
rect 10380 10833 10426 10954
rect 10426 10833 10431 10954
rect 10237 10534 10242 10654
rect 10242 10534 10288 10654
rect 10288 10534 10293 10654
rect 9777 10415 9778 10458
rect 9778 10415 9832 10458
rect 9832 10415 9833 10458
rect 9777 10402 9833 10415
rect 9961 10415 9962 10458
rect 9962 10415 10016 10458
rect 10016 10415 10017 10458
rect 9961 10402 10017 10415
rect 10145 10415 10146 10458
rect 10146 10415 10200 10458
rect 10200 10415 10201 10458
rect 10145 10402 10201 10415
rect 9777 10252 9833 10308
rect 8475 10135 8531 10191
rect 8804 10135 8860 10191
rect 9061 10135 9117 10191
rect 9961 10136 10017 10192
rect 10290 10136 10346 10192
rect 10723 10136 10779 10192
rect 13279 11327 13335 11383
rect 14589 11328 14645 11384
rect 12609 11220 12665 11276
rect 12241 10833 12246 10953
rect 12246 10833 12292 10953
rect 12292 10833 12297 10953
rect 12609 10833 12614 10953
rect 12614 10833 12660 10953
rect 12660 10833 12665 10953
rect 12425 10533 12430 10653
rect 12430 10533 12476 10653
rect 12476 10533 12481 10653
rect 12931 10832 12936 10953
rect 12936 10832 12982 10953
rect 12982 10832 12987 10953
rect 12793 10533 12798 10653
rect 12798 10533 12844 10653
rect 12844 10533 12849 10653
rect 12333 10414 12334 10457
rect 12334 10414 12388 10457
rect 12388 10414 12389 10457
rect 12333 10401 12389 10414
rect 12517 10414 12518 10457
rect 12518 10414 12572 10457
rect 12572 10414 12573 10457
rect 12517 10401 12573 10414
rect 12701 10414 12702 10457
rect 12702 10414 12756 10457
rect 12756 10414 12757 10457
rect 12701 10401 12757 10414
rect 12333 10251 12389 10307
rect 14095 11221 14151 11277
rect 13727 10834 13732 10954
rect 13732 10834 13778 10954
rect 13778 10834 13783 10954
rect 14095 10834 14100 10954
rect 14100 10834 14146 10954
rect 14146 10834 14151 10954
rect 13911 10534 13916 10654
rect 13916 10534 13962 10654
rect 13962 10534 13967 10654
rect 14417 10833 14422 10954
rect 14422 10833 14468 10954
rect 14468 10833 14473 10954
rect 14279 10534 14284 10654
rect 14284 10534 14330 10654
rect 14330 10534 14335 10654
rect 13819 10415 13820 10458
rect 13820 10415 13874 10458
rect 13874 10415 13875 10458
rect 13819 10402 13875 10415
rect 14003 10415 14004 10458
rect 14004 10415 14058 10458
rect 14058 10415 14059 10458
rect 14003 10402 14059 10415
rect 14187 10415 14188 10458
rect 14188 10415 14242 10458
rect 14242 10415 14243 10458
rect 14187 10402 14243 10415
rect 13819 10252 13875 10308
rect 12517 10135 12573 10191
rect 12846 10135 12902 10191
rect 13103 10135 13159 10191
rect 14003 10136 14059 10192
rect 14332 10136 14388 10192
rect 14765 10136 14821 10192
rect -12561 10019 -12505 10075
rect -11521 10019 -11465 10075
rect -10035 10020 -9979 10076
rect -11889 9912 -11833 9925
rect -11889 9869 -11888 9912
rect -11888 9869 -11834 9912
rect -11834 9869 -11833 9912
rect -11705 9912 -11649 9925
rect -11705 9869 -11704 9912
rect -11704 9869 -11650 9912
rect -11650 9869 -11649 9912
rect -11521 9912 -11465 9925
rect -11521 9869 -11520 9912
rect -11520 9869 -11466 9912
rect -11466 9869 -11465 9912
rect -11429 9673 -11424 9793
rect -11424 9673 -11378 9793
rect -11378 9673 -11373 9793
rect -12114 9350 -12058 9406
rect -11296 9350 -11240 9406
rect -10943 9232 -10887 9288
rect -11119 9124 -11063 9178
rect -11613 9015 -11557 9071
rect -11981 8628 -11976 8748
rect -11976 8628 -11930 8748
rect -11930 8628 -11925 8748
rect -11613 8628 -11608 8748
rect -11608 8628 -11562 8748
rect -11562 8628 -11557 8748
rect -11797 8328 -11792 8448
rect -11792 8328 -11746 8448
rect -11746 8328 -11741 8448
rect -11291 8627 -11286 8748
rect -11286 8627 -11240 8748
rect -11240 8627 -11235 8748
rect -11429 8328 -11424 8448
rect -11424 8328 -11378 8448
rect -11378 8328 -11373 8448
rect -11889 8209 -11888 8252
rect -11888 8209 -11834 8252
rect -11834 8209 -11833 8252
rect -11889 8196 -11833 8209
rect -11705 8209 -11704 8252
rect -11704 8209 -11650 8252
rect -11650 8209 -11649 8252
rect -11705 8196 -11649 8209
rect -11521 8209 -11520 8252
rect -11520 8209 -11466 8252
rect -11466 8209 -11465 8252
rect -11521 8196 -11465 8209
rect -11889 8046 -11833 8102
rect -12697 7930 -12641 7986
rect -11705 7930 -11649 7986
rect -11376 7930 -11320 7986
rect -10943 7930 -10887 7986
rect -12896 7814 -12840 7870
rect -11521 7814 -11465 7870
rect -11889 7707 -11833 7720
rect -11889 7664 -11888 7707
rect -11888 7664 -11834 7707
rect -11834 7664 -11833 7707
rect -11705 7707 -11649 7720
rect -11705 7664 -11704 7707
rect -11704 7664 -11650 7707
rect -11650 7664 -11649 7707
rect -11521 7707 -11465 7720
rect -11521 7664 -11520 7707
rect -11520 7664 -11466 7707
rect -11466 7664 -11465 7707
rect -11429 7468 -11424 7588
rect -11424 7468 -11378 7588
rect -11378 7468 -11373 7588
rect -12114 7145 -12058 7201
rect -11296 7145 -11240 7201
rect -8549 10019 -8493 10075
rect -7509 10019 -7453 10075
rect -10403 9913 -10347 9926
rect -10403 9870 -10402 9913
rect -10402 9870 -10348 9913
rect -10348 9870 -10347 9913
rect -10219 9913 -10163 9926
rect -10219 9870 -10218 9913
rect -10218 9870 -10164 9913
rect -10164 9870 -10163 9913
rect -10035 9913 -9979 9926
rect -10035 9870 -10034 9913
rect -10034 9870 -9980 9913
rect -9980 9870 -9979 9913
rect -9943 9674 -9938 9794
rect -9938 9674 -9892 9794
rect -9892 9674 -9887 9794
rect -10628 9351 -10572 9407
rect -9810 9351 -9754 9407
rect -6023 10020 -5967 10076
rect -7877 9912 -7821 9925
rect -7877 9869 -7876 9912
rect -7876 9869 -7822 9912
rect -7822 9869 -7821 9912
rect -7693 9912 -7637 9925
rect -7693 9869 -7692 9912
rect -7692 9869 -7638 9912
rect -7638 9869 -7637 9912
rect -7509 9912 -7453 9925
rect -7509 9869 -7508 9912
rect -7508 9869 -7454 9912
rect -7454 9869 -7453 9912
rect -7417 9673 -7412 9793
rect -7412 9673 -7366 9793
rect -7366 9673 -7361 9793
rect -8102 9350 -8046 9406
rect -7284 9350 -7228 9406
rect -6931 9232 -6875 9288
rect -7107 9124 -7051 9178
rect -7601 9015 -7545 9071
rect -7969 8628 -7964 8748
rect -7964 8628 -7918 8748
rect -7918 8628 -7913 8748
rect -7601 8628 -7596 8748
rect -7596 8628 -7550 8748
rect -7550 8628 -7545 8748
rect -7785 8328 -7780 8448
rect -7780 8328 -7734 8448
rect -7734 8328 -7729 8448
rect -7279 8627 -7274 8748
rect -7274 8627 -7228 8748
rect -7228 8627 -7223 8748
rect -7417 8328 -7412 8448
rect -7412 8328 -7366 8448
rect -7366 8328 -7361 8448
rect -7877 8209 -7876 8252
rect -7876 8209 -7822 8252
rect -7822 8209 -7821 8252
rect -7877 8196 -7821 8209
rect -7693 8209 -7692 8252
rect -7692 8209 -7638 8252
rect -7638 8209 -7637 8252
rect -7693 8196 -7637 8209
rect -7509 8209 -7508 8252
rect -7508 8209 -7454 8252
rect -7454 8209 -7453 8252
rect -7509 8196 -7453 8209
rect -7877 8046 -7821 8102
rect -8685 7930 -8629 7986
rect -7693 7930 -7637 7986
rect -7364 7930 -7308 7986
rect -6931 7930 -6875 7986
rect -8821 7814 -8765 7870
rect -7509 7814 -7453 7870
rect -7877 7707 -7821 7720
rect -7877 7664 -7876 7707
rect -7876 7664 -7822 7707
rect -7822 7664 -7821 7707
rect -7693 7707 -7637 7720
rect -7693 7664 -7692 7707
rect -7692 7664 -7638 7707
rect -7638 7664 -7637 7707
rect -7509 7707 -7453 7720
rect -7509 7664 -7508 7707
rect -7508 7664 -7454 7707
rect -7454 7664 -7453 7707
rect -7417 7468 -7412 7588
rect -7412 7468 -7366 7588
rect -7366 7468 -7361 7588
rect -8102 7145 -8046 7201
rect -7284 7145 -7228 7201
rect -12896 7027 -12840 7083
rect -12697 7027 -12641 7083
rect -4507 10019 -4451 10075
rect -3467 10019 -3411 10075
rect -6391 9913 -6335 9926
rect -6391 9870 -6390 9913
rect -6390 9870 -6336 9913
rect -6336 9870 -6335 9913
rect -6207 9913 -6151 9926
rect -6207 9870 -6206 9913
rect -6206 9870 -6152 9913
rect -6152 9870 -6151 9913
rect -6023 9913 -5967 9926
rect -6023 9870 -6022 9913
rect -6022 9870 -5968 9913
rect -5968 9870 -5967 9913
rect -5931 9674 -5926 9794
rect -5926 9674 -5880 9794
rect -5880 9674 -5875 9794
rect -6616 9351 -6560 9407
rect -5798 9351 -5742 9407
rect -1981 10020 -1925 10076
rect -3835 9912 -3779 9925
rect -3835 9869 -3834 9912
rect -3834 9869 -3780 9912
rect -3780 9869 -3779 9912
rect -3651 9912 -3595 9925
rect -3651 9869 -3650 9912
rect -3650 9869 -3596 9912
rect -3596 9869 -3595 9912
rect -3467 9912 -3411 9925
rect -3467 9869 -3466 9912
rect -3466 9869 -3412 9912
rect -3412 9869 -3411 9912
rect -3375 9673 -3370 9793
rect -3370 9673 -3324 9793
rect -3324 9673 -3319 9793
rect -4060 9350 -4004 9406
rect -3242 9350 -3186 9406
rect -2889 9232 -2833 9288
rect -3065 9124 -3009 9178
rect -3559 9015 -3503 9071
rect -3927 8628 -3922 8748
rect -3922 8628 -3876 8748
rect -3876 8628 -3871 8748
rect -3559 8628 -3554 8748
rect -3554 8628 -3508 8748
rect -3508 8628 -3503 8748
rect -3743 8328 -3738 8448
rect -3738 8328 -3692 8448
rect -3692 8328 -3687 8448
rect -3237 8627 -3232 8748
rect -3232 8627 -3186 8748
rect -3186 8627 -3181 8748
rect -3375 8328 -3370 8448
rect -3370 8328 -3324 8448
rect -3324 8328 -3319 8448
rect -3835 8209 -3834 8252
rect -3834 8209 -3780 8252
rect -3780 8209 -3779 8252
rect -3835 8196 -3779 8209
rect -3651 8209 -3650 8252
rect -3650 8209 -3596 8252
rect -3596 8209 -3595 8252
rect -3651 8196 -3595 8209
rect -3467 8209 -3466 8252
rect -3466 8209 -3412 8252
rect -3412 8209 -3411 8252
rect -3467 8196 -3411 8209
rect -3835 8046 -3779 8102
rect -4643 7930 -4587 7986
rect -3651 7930 -3595 7986
rect -3322 7930 -3266 7986
rect -2889 7930 -2833 7986
rect -4809 7814 -4753 7870
rect -3467 7814 -3411 7870
rect -3835 7707 -3779 7720
rect -3835 7664 -3834 7707
rect -3834 7664 -3780 7707
rect -3780 7664 -3779 7707
rect -3651 7707 -3595 7720
rect -3651 7664 -3650 7707
rect -3650 7664 -3596 7707
rect -3596 7664 -3595 7707
rect -3467 7707 -3411 7720
rect -3467 7664 -3466 7707
rect -3466 7664 -3412 7707
rect -3412 7664 -3411 7707
rect -3375 7468 -3370 7588
rect -3370 7468 -3324 7588
rect -3324 7468 -3319 7588
rect -4060 7145 -4004 7201
rect -3242 7145 -3186 7201
rect -8957 7027 -8901 7083
rect -8685 7027 -8629 7083
rect -465 10019 -409 10075
rect 575 10019 631 10075
rect -2349 9913 -2293 9926
rect -2349 9870 -2348 9913
rect -2348 9870 -2294 9913
rect -2294 9870 -2293 9913
rect -2165 9913 -2109 9926
rect -2165 9870 -2164 9913
rect -2164 9870 -2110 9913
rect -2110 9870 -2109 9913
rect -1981 9913 -1925 9926
rect -1981 9870 -1980 9913
rect -1980 9870 -1926 9913
rect -1926 9870 -1925 9913
rect -1889 9674 -1884 9794
rect -1884 9674 -1838 9794
rect -1838 9674 -1833 9794
rect -2574 9351 -2518 9407
rect -1756 9351 -1700 9407
rect 2061 10020 2117 10076
rect 207 9912 263 9925
rect 207 9869 208 9912
rect 208 9869 262 9912
rect 262 9869 263 9912
rect 391 9912 447 9925
rect 391 9869 392 9912
rect 392 9869 446 9912
rect 446 9869 447 9912
rect 575 9912 631 9925
rect 575 9869 576 9912
rect 576 9869 630 9912
rect 630 9869 631 9912
rect 667 9673 672 9793
rect 672 9673 718 9793
rect 718 9673 723 9793
rect -18 9350 38 9406
rect 800 9350 856 9406
rect 1153 9232 1209 9288
rect 977 9124 1033 9178
rect 483 9015 539 9071
rect 115 8628 120 8748
rect 120 8628 166 8748
rect 166 8628 171 8748
rect 483 8628 488 8748
rect 488 8628 534 8748
rect 534 8628 539 8748
rect 299 8328 304 8448
rect 304 8328 350 8448
rect 350 8328 355 8448
rect 805 8627 810 8748
rect 810 8627 856 8748
rect 856 8627 861 8748
rect 667 8328 672 8448
rect 672 8328 718 8448
rect 718 8328 723 8448
rect 207 8209 208 8252
rect 208 8209 262 8252
rect 262 8209 263 8252
rect 207 8196 263 8209
rect 391 8209 392 8252
rect 392 8209 446 8252
rect 446 8209 447 8252
rect 391 8196 447 8209
rect 575 8209 576 8252
rect 576 8209 630 8252
rect 630 8209 631 8252
rect 575 8196 631 8209
rect 207 8046 263 8102
rect -601 7930 -545 7986
rect 391 7930 447 7986
rect 720 7930 776 7986
rect 1153 7930 1209 7986
rect -767 7814 -711 7870
rect 575 7814 631 7870
rect 207 7707 263 7720
rect 207 7664 208 7707
rect 208 7664 262 7707
rect 262 7664 263 7707
rect 391 7707 447 7720
rect 391 7664 392 7707
rect 392 7664 446 7707
rect 446 7664 447 7707
rect 575 7707 631 7720
rect 575 7664 576 7707
rect 576 7664 630 7707
rect 630 7664 631 7707
rect 667 7468 672 7588
rect 672 7468 718 7588
rect 718 7468 723 7588
rect -18 7145 38 7201
rect 800 7145 856 7201
rect -4945 7027 -4889 7083
rect -4643 7027 -4587 7083
rect 3577 10019 3633 10075
rect 4617 10019 4673 10075
rect 1693 9913 1749 9926
rect 1693 9870 1694 9913
rect 1694 9870 1748 9913
rect 1748 9870 1749 9913
rect 1877 9913 1933 9926
rect 1877 9870 1878 9913
rect 1878 9870 1932 9913
rect 1932 9870 1933 9913
rect 2061 9913 2117 9926
rect 2061 9870 2062 9913
rect 2062 9870 2116 9913
rect 2116 9870 2117 9913
rect 2153 9674 2158 9794
rect 2158 9674 2204 9794
rect 2204 9674 2209 9794
rect 1468 9351 1524 9407
rect 2286 9351 2342 9407
rect 6103 10020 6159 10076
rect 4249 9912 4305 9925
rect 4249 9869 4250 9912
rect 4250 9869 4304 9912
rect 4304 9869 4305 9912
rect 4433 9912 4489 9925
rect 4433 9869 4434 9912
rect 4434 9869 4488 9912
rect 4488 9869 4489 9912
rect 4617 9912 4673 9925
rect 4617 9869 4618 9912
rect 4618 9869 4672 9912
rect 4672 9869 4673 9912
rect 4709 9673 4714 9793
rect 4714 9673 4760 9793
rect 4760 9673 4765 9793
rect 4024 9350 4080 9406
rect 4842 9350 4898 9406
rect 5195 9232 5251 9288
rect 5019 9124 5075 9178
rect 4525 9015 4581 9071
rect 4157 8628 4162 8748
rect 4162 8628 4208 8748
rect 4208 8628 4213 8748
rect 4525 8628 4530 8748
rect 4530 8628 4576 8748
rect 4576 8628 4581 8748
rect 4341 8328 4346 8448
rect 4346 8328 4392 8448
rect 4392 8328 4397 8448
rect 4847 8627 4852 8748
rect 4852 8627 4898 8748
rect 4898 8627 4903 8748
rect 4709 8328 4714 8448
rect 4714 8328 4760 8448
rect 4760 8328 4765 8448
rect 4249 8209 4250 8252
rect 4250 8209 4304 8252
rect 4304 8209 4305 8252
rect 4249 8196 4305 8209
rect 4433 8209 4434 8252
rect 4434 8209 4488 8252
rect 4488 8209 4489 8252
rect 4433 8196 4489 8209
rect 4617 8209 4618 8252
rect 4618 8209 4672 8252
rect 4672 8209 4673 8252
rect 4617 8196 4673 8209
rect 4249 8046 4305 8102
rect 3441 7930 3497 7986
rect 4433 7930 4489 7986
rect 4762 7930 4818 7986
rect 5195 7930 5251 7986
rect 3275 7814 3331 7870
rect 4617 7814 4673 7870
rect 4249 7707 4305 7720
rect 4249 7664 4250 7707
rect 4250 7664 4304 7707
rect 4304 7664 4305 7707
rect 4433 7707 4489 7720
rect 4433 7664 4434 7707
rect 4434 7664 4488 7707
rect 4488 7664 4489 7707
rect 4617 7707 4673 7720
rect 4617 7664 4618 7707
rect 4618 7664 4672 7707
rect 4672 7664 4673 7707
rect 4709 7468 4714 7588
rect 4714 7468 4760 7588
rect 4760 7468 4765 7588
rect 4024 7145 4080 7201
rect 4842 7145 4898 7201
rect -903 7027 -847 7083
rect -601 7027 -545 7083
rect 7619 10019 7675 10075
rect 8659 10019 8715 10075
rect 5735 9913 5791 9926
rect 5735 9870 5736 9913
rect 5736 9870 5790 9913
rect 5790 9870 5791 9913
rect 5919 9913 5975 9926
rect 5919 9870 5920 9913
rect 5920 9870 5974 9913
rect 5974 9870 5975 9913
rect 6103 9913 6159 9926
rect 6103 9870 6104 9913
rect 6104 9870 6158 9913
rect 6158 9870 6159 9913
rect 6195 9674 6200 9794
rect 6200 9674 6246 9794
rect 6246 9674 6251 9794
rect 5510 9351 5566 9407
rect 6328 9351 6384 9407
rect 10145 10020 10201 10076
rect 8291 9912 8347 9925
rect 8291 9869 8292 9912
rect 8292 9869 8346 9912
rect 8346 9869 8347 9912
rect 8475 9912 8531 9925
rect 8475 9869 8476 9912
rect 8476 9869 8530 9912
rect 8530 9869 8531 9912
rect 8659 9912 8715 9925
rect 8659 9869 8660 9912
rect 8660 9869 8714 9912
rect 8714 9869 8715 9912
rect 8751 9673 8756 9793
rect 8756 9673 8802 9793
rect 8802 9673 8807 9793
rect 8066 9350 8122 9406
rect 8884 9350 8940 9406
rect 9237 9232 9293 9288
rect 9061 9124 9117 9178
rect 8567 9015 8623 9071
rect 8199 8628 8204 8748
rect 8204 8628 8250 8748
rect 8250 8628 8255 8748
rect 8567 8628 8572 8748
rect 8572 8628 8618 8748
rect 8618 8628 8623 8748
rect 8383 8328 8388 8448
rect 8388 8328 8434 8448
rect 8434 8328 8439 8448
rect 8889 8627 8894 8748
rect 8894 8627 8940 8748
rect 8940 8627 8945 8748
rect 8751 8328 8756 8448
rect 8756 8328 8802 8448
rect 8802 8328 8807 8448
rect 8291 8209 8292 8252
rect 8292 8209 8346 8252
rect 8346 8209 8347 8252
rect 8291 8196 8347 8209
rect 8475 8209 8476 8252
rect 8476 8209 8530 8252
rect 8530 8209 8531 8252
rect 8475 8196 8531 8209
rect 8659 8209 8660 8252
rect 8660 8209 8714 8252
rect 8714 8209 8715 8252
rect 8659 8196 8715 8209
rect 8291 8046 8347 8102
rect 7483 7930 7539 7986
rect 8475 7930 8531 7986
rect 8804 7930 8860 7986
rect 9237 7930 9293 7986
rect 7317 7814 7373 7870
rect 8659 7814 8715 7870
rect 8291 7707 8347 7720
rect 8291 7664 8292 7707
rect 8292 7664 8346 7707
rect 8346 7664 8347 7707
rect 8475 7707 8531 7720
rect 8475 7664 8476 7707
rect 8476 7664 8530 7707
rect 8530 7664 8531 7707
rect 8659 7707 8715 7720
rect 8659 7664 8660 7707
rect 8660 7664 8714 7707
rect 8714 7664 8715 7707
rect 8751 7468 8756 7588
rect 8756 7468 8802 7588
rect 8802 7468 8807 7588
rect 8066 7145 8122 7201
rect 8884 7145 8940 7201
rect 3139 7027 3195 7083
rect 3441 7027 3497 7083
rect 11661 10019 11717 10075
rect 12701 10019 12757 10075
rect 9777 9913 9833 9926
rect 9777 9870 9778 9913
rect 9778 9870 9832 9913
rect 9832 9870 9833 9913
rect 9961 9913 10017 9926
rect 9961 9870 9962 9913
rect 9962 9870 10016 9913
rect 10016 9870 10017 9913
rect 10145 9913 10201 9926
rect 10145 9870 10146 9913
rect 10146 9870 10200 9913
rect 10200 9870 10201 9913
rect 10237 9674 10242 9794
rect 10242 9674 10288 9794
rect 10288 9674 10293 9794
rect 9552 9351 9608 9407
rect 10370 9351 10426 9407
rect 14187 10020 14243 10076
rect 12333 9912 12389 9925
rect 12333 9869 12334 9912
rect 12334 9869 12388 9912
rect 12388 9869 12389 9912
rect 12517 9912 12573 9925
rect 12517 9869 12518 9912
rect 12518 9869 12572 9912
rect 12572 9869 12573 9912
rect 12701 9912 12757 9925
rect 12701 9869 12702 9912
rect 12702 9869 12756 9912
rect 12756 9869 12757 9912
rect 12793 9673 12798 9793
rect 12798 9673 12844 9793
rect 12844 9673 12849 9793
rect 12108 9350 12164 9406
rect 12926 9350 12982 9406
rect 13279 9232 13335 9288
rect 13103 9124 13159 9178
rect 12609 9015 12665 9071
rect 12241 8628 12246 8748
rect 12246 8628 12292 8748
rect 12292 8628 12297 8748
rect 12609 8628 12614 8748
rect 12614 8628 12660 8748
rect 12660 8628 12665 8748
rect 12425 8328 12430 8448
rect 12430 8328 12476 8448
rect 12476 8328 12481 8448
rect 12931 8627 12936 8748
rect 12936 8627 12982 8748
rect 12982 8627 12987 8748
rect 12793 8328 12798 8448
rect 12798 8328 12844 8448
rect 12844 8328 12849 8448
rect 12333 8209 12334 8252
rect 12334 8209 12388 8252
rect 12388 8209 12389 8252
rect 12333 8196 12389 8209
rect 12517 8209 12518 8252
rect 12518 8209 12572 8252
rect 12572 8209 12573 8252
rect 12517 8196 12573 8209
rect 12701 8209 12702 8252
rect 12702 8209 12756 8252
rect 12756 8209 12757 8252
rect 12701 8196 12757 8209
rect 12333 8046 12389 8102
rect 11525 7930 11581 7986
rect 12517 7930 12573 7986
rect 12846 7930 12902 7986
rect 13279 7930 13335 7986
rect 11359 7814 11415 7870
rect 12701 7814 12757 7870
rect 12333 7707 12389 7720
rect 12333 7664 12334 7707
rect 12334 7664 12388 7707
rect 12388 7664 12389 7707
rect 12517 7707 12573 7720
rect 12517 7664 12518 7707
rect 12518 7664 12572 7707
rect 12572 7664 12573 7707
rect 12701 7707 12757 7720
rect 12701 7664 12702 7707
rect 12702 7664 12756 7707
rect 12756 7664 12757 7707
rect 12793 7468 12798 7588
rect 12798 7468 12844 7588
rect 12844 7468 12849 7588
rect 12108 7145 12164 7201
rect 12926 7145 12982 7201
rect 7181 7027 7237 7083
rect 7483 7027 7539 7083
rect 13819 9913 13875 9926
rect 13819 9870 13820 9913
rect 13820 9870 13874 9913
rect 13874 9870 13875 9913
rect 14003 9913 14059 9926
rect 14003 9870 14004 9913
rect 14004 9870 14058 9913
rect 14058 9870 14059 9913
rect 14187 9913 14243 9926
rect 14187 9870 14188 9913
rect 14188 9870 14242 9913
rect 14242 9870 14243 9913
rect 14279 9674 14284 9794
rect 14284 9674 14330 9794
rect 14330 9674 14335 9794
rect 13594 9351 13650 9407
rect 14412 9351 14468 9407
rect 11223 7027 11279 7083
rect 11525 7027 11581 7083
rect -4454 6134 -2454 6434
rect -13665 4881 -13607 4939
rect -12366 4880 -12306 4940
rect -10747 4884 -10695 4936
rect -10187 4673 -10135 4676
rect -10187 4627 -10184 4673
rect -10184 4627 -10138 4673
rect -10138 4627 -10135 4673
rect -10187 4624 -10135 4627
rect -8327 4739 -8322 4795
rect -8322 4739 -8276 4795
rect -8276 4739 -8271 4795
rect -8051 4739 -8046 4795
rect -8046 4739 -8000 4795
rect -8000 4739 -7995 4795
rect -8189 4481 -8133 4537
rect -8189 4343 -8133 4399
rect -10519 3300 -10439 3376
rect -8327 3919 -8322 3975
rect -8322 3919 -8276 3975
rect -8276 3919 -8271 3975
rect -8419 3768 -8418 3799
rect -8418 3768 -8364 3799
rect -8364 3768 -8363 3799
rect -8419 3743 -8363 3768
rect -8051 3919 -8046 3975
rect -8046 3919 -8000 3975
rect -8000 3919 -7995 3975
rect -7959 3768 -7958 3799
rect -7958 3768 -7904 3799
rect -7904 3768 -7903 3799
rect -7959 3743 -7903 3768
rect -8419 3300 -8363 3376
rect -12086 2883 -12006 2961
rect -7959 3300 -7903 3376
rect -5883 3300 -5803 3376
rect -5676 2787 -5596 2847
rect -11642 2462 -11551 2551
rect -4764 2542 -4655 2649
rect -11379 2356 -11299 2432
rect -5023 2356 -4943 2432
rect -11029 1530 -11024 1664
rect -11024 1530 -10978 1664
rect -10978 1530 -10973 1664
rect -10845 1530 -10840 1664
rect -10840 1530 -10794 1664
rect -10794 1530 -10789 1664
rect -10707 1530 -10702 1664
rect -10702 1530 -10656 1664
rect -10656 1530 -10651 1664
rect -10169 1530 -10164 1664
rect -10164 1530 -10118 1664
rect -10118 1530 -10113 1664
rect -9985 1530 -9980 1664
rect -9980 1530 -9934 1664
rect -9934 1530 -9929 1664
rect -9847 1530 -9842 1664
rect -9842 1530 -9796 1664
rect -9796 1530 -9791 1664
rect -9405 1533 -9400 1677
rect -9400 1533 -9354 1677
rect -9354 1533 -9349 1677
rect -9101 1520 -9096 1576
rect -9096 1520 -9050 1576
rect -9050 1520 -9045 1576
rect -8797 1533 -8792 1677
rect -8792 1533 -8746 1677
rect -8746 1533 -8741 1677
rect -8493 1520 -8488 1576
rect -8488 1520 -8442 1576
rect -8442 1520 -8437 1576
rect -8189 1533 -8184 1677
rect -8184 1533 -8138 1677
rect -8138 1533 -8133 1677
rect -7885 1520 -7880 1576
rect -7880 1520 -7834 1576
rect -7834 1520 -7829 1576
rect -7581 1533 -7576 1677
rect -7576 1533 -7530 1677
rect -7530 1533 -7525 1677
rect -7277 1520 -7272 1576
rect -7272 1520 -7226 1576
rect -7226 1520 -7221 1576
rect -6973 1533 -6968 1677
rect -6968 1533 -6922 1677
rect -6922 1533 -6917 1677
rect -6531 1530 -6526 1664
rect -6526 1530 -6480 1664
rect -6480 1530 -6475 1664
rect -8298 1464 -8242 1469
rect -8080 1464 -8024 1469
rect -8298 1418 -8242 1464
rect -8080 1418 -8024 1464
rect -6393 1530 -6388 1664
rect -6388 1530 -6342 1664
rect -6342 1530 -6337 1664
rect -6209 1530 -6204 1664
rect -6204 1530 -6158 1664
rect -6158 1530 -6153 1664
rect -8298 1413 -8242 1418
rect -8080 1413 -8024 1418
rect -5671 1530 -5666 1664
rect -5666 1530 -5620 1664
rect -5620 1530 -5615 1664
rect -5533 1530 -5528 1664
rect -5528 1530 -5482 1664
rect -5482 1530 -5477 1664
rect -5349 1530 -5344 1664
rect -5344 1530 -5298 1664
rect -5298 1530 -5293 1664
rect -10519 1077 -10439 1161
rect -9997 1077 -9917 1161
rect -9251 1079 -9171 1159
rect -8643 1079 -8563 1159
rect -8505 1079 -8425 1159
rect -7897 1079 -7817 1159
rect -7759 1079 -7679 1159
rect -7151 1079 -7071 1159
rect -6405 1077 -6325 1161
rect -5883 1077 -5803 1161
rect -8842 820 -8762 865
rect -8842 785 -8762 820
rect -7560 820 -7480 865
rect -9985 271 -9980 415
rect -9980 271 -9934 415
rect -9934 271 -9929 415
rect -9239 577 -9234 721
rect -9234 577 -9188 721
rect -9188 577 -9183 721
rect -9543 361 -9538 505
rect -9538 361 -9492 505
rect -9492 361 -9487 505
rect -8631 577 -8626 721
rect -8626 577 -8580 721
rect -8580 577 -8575 721
rect -8935 361 -8930 505
rect -8930 361 -8884 505
rect -8884 361 -8879 505
rect -7560 785 -7480 820
rect -7747 577 -7742 721
rect -7742 577 -7696 721
rect -7696 577 -7691 721
rect -7139 577 -7134 721
rect -7134 577 -7088 721
rect -7088 577 -7083 721
rect -7443 361 -7438 505
rect -7438 361 -7392 505
rect -7392 361 -7387 505
rect -6835 361 -6830 505
rect -6830 361 -6784 505
rect -6784 361 -6779 505
rect -6393 271 -6388 415
rect -6388 271 -6342 415
rect -6342 271 -6337 415
rect -10857 -85 -10777 -5
rect -9721 -85 -9641 -5
rect -9555 -85 -9475 -5
rect -8947 -85 -8867 -5
rect -7455 -85 -7375 -5
rect -6847 -85 -6767 -5
rect -6681 -85 -6601 -5
rect -5545 -85 -5465 -5
rect -10304 -564 -10204 -403
rect -9709 -974 -9704 -813
rect -9704 -974 -9658 -813
rect -9658 -974 -9653 -813
rect -9405 -1022 -9400 -861
rect -9400 -1022 -9354 -861
rect -9354 -1022 -9349 -861
rect -9101 -994 -9096 -777
rect -9096 -994 -9050 -777
rect -9050 -994 -9045 -777
rect -8493 -833 -8488 -777
rect -8488 -833 -8442 -777
rect -8442 -833 -8437 -777
rect -8797 -1022 -8792 -861
rect -8792 -1022 -8746 -861
rect -8746 -1022 -8741 -861
rect -7885 -833 -7880 -777
rect -7880 -833 -7834 -777
rect -7834 -833 -7829 -777
rect -8189 -1022 -8184 -861
rect -8184 -1022 -8138 -861
rect -8138 -1022 -8133 -861
rect -7581 -1022 -7576 -861
rect -7576 -1022 -7530 -861
rect -7530 -1022 -7525 -861
rect -7277 -1022 -7272 -777
rect -7272 -1022 -7226 -777
rect -7226 -1022 -7221 -777
rect -6973 -1022 -6968 -861
rect -6968 -1022 -6922 -861
rect -6922 -1022 -6917 -861
rect -6669 -974 -6664 -813
rect -6664 -974 -6618 -813
rect -6618 -974 -6613 -813
rect -6118 -564 -6018 -403
rect -9261 -1077 -9191 -1068
rect -8956 -1077 -8886 -1068
rect -8046 -1077 -7976 -1068
rect -7741 -1077 -7671 -1068
rect -6826 -1077 -6756 -1068
rect -9261 -1123 -9191 -1077
rect -8956 -1123 -8886 -1077
rect -8046 -1123 -7976 -1077
rect -7741 -1123 -7671 -1077
rect -6826 -1123 -6756 -1077
rect -9261 -1128 -9191 -1123
rect -8956 -1128 -8886 -1123
rect -8046 -1128 -7976 -1123
rect -7741 -1128 -7671 -1123
rect -6826 -1128 -6756 -1123
rect -13707 -1252 -13634 -1179
rect -9254 -1282 -9198 -1226
rect -8039 -1282 -7983 -1226
rect -6511 -1253 -6451 -1193
rect -13704 -1577 -13631 -1504
rect -8949 -1530 -8893 -1474
rect -7734 -1530 -7678 -1474
rect -6251 -1563 -6191 -1503
rect -9261 -1674 -9191 -1628
rect -8956 -1674 -8886 -1628
rect -8046 -1674 -7976 -1628
rect -7741 -1674 -7671 -1628
rect -6826 -1674 -6756 -1628
rect -9261 -1688 -9191 -1674
rect -8956 -1688 -8886 -1674
rect -8046 -1688 -7976 -1674
rect -7741 -1688 -7671 -1674
rect -6826 -1688 -6756 -1674
rect -10304 -2348 -10204 -2187
rect -9405 -1893 -9400 -1732
rect -9400 -1893 -9354 -1732
rect -9354 -1893 -9349 -1732
rect -9709 -1977 -9704 -1921
rect -9704 -1977 -9658 -1921
rect -9658 -1977 -9653 -1921
rect -9101 -1977 -9096 -1766
rect -9096 -1977 -9050 -1766
rect -9050 -1977 -9045 -1766
rect -8797 -1893 -8792 -1732
rect -8792 -1893 -8746 -1732
rect -8746 -1893 -8741 -1732
rect -8493 -1977 -8488 -1732
rect -8488 -1977 -8442 -1732
rect -8442 -1977 -8437 -1732
rect -8189 -1893 -8184 -1732
rect -8184 -1893 -8138 -1732
rect -8138 -1893 -8133 -1732
rect -7885 -1977 -7880 -1766
rect -7880 -1977 -7834 -1766
rect -7834 -1977 -7829 -1766
rect -7581 -1893 -7576 -1732
rect -7576 -1893 -7530 -1732
rect -7530 -1893 -7525 -1732
rect -7277 -1977 -7272 -1732
rect -7272 -1977 -7226 -1732
rect -7226 -1977 -7221 -1732
rect -6973 -1977 -6968 -1732
rect -6968 -1977 -6922 -1732
rect -6922 -1977 -6917 -1732
rect -6669 -1977 -6664 -1920
rect -6664 -1977 -6618 -1920
rect -6618 -1977 -6613 -1920
rect -6129 -2348 -6118 -2160
rect -6118 -2348 -6024 -2160
rect -6129 -2370 -6024 -2348
rect -8603 -2774 -8598 -2652
rect -8598 -2774 -8552 -2652
rect -8552 -2774 -8547 -2652
rect -8281 -2774 -8276 -2652
rect -8276 -2774 -8230 -2652
rect -8230 -2774 -8225 -2652
rect -8097 -2774 -8092 -2652
rect -8092 -2774 -8046 -2652
rect -8046 -2774 -8041 -2652
rect -13368 -3082 -13290 -3004
rect -11379 -3083 -11299 -3003
rect -5023 -3083 -4943 -3003
rect -11640 -3530 -11555 -3443
rect -10639 -3463 -10550 -3376
rect -10083 -3592 -9728 -3381
rect -6132 -3578 -6018 -3375
rect -5654 -3531 -5550 -3429
rect -4764 -3558 -4655 -3451
rect -4454 -3663 -2454 -3363
<< metal2 >>
rect 40726 39167 40972 39180
rect 40726 39093 40739 39167
rect 40957 39093 40972 39167
rect 40726 39080 40972 39093
rect -8093 33382 -8037 38726
rect 38117 38599 40211 38613
rect 38117 38547 40135 38599
rect 40187 38547 40211 38599
rect 38117 38533 40211 38547
rect 40681 38343 40761 38353
rect 40671 38341 40927 38343
rect 40671 38339 45751 38341
rect 40671 38287 40695 38339
rect 40747 38287 45751 38339
rect 40671 38285 45751 38287
rect 40671 38283 40927 38285
rect 40681 38273 40761 38283
rect 40723 37823 40967 37836
rect 40723 37749 40737 37823
rect 40955 37749 40967 37823
rect 40723 37737 40967 37749
rect -4711 37567 -3965 37579
rect -4711 37511 -4343 37567
rect -4287 37511 -3965 37567
rect -4711 37499 -3965 37511
rect -4711 37246 -4655 37499
rect -4343 37246 -4287 37499
rect -4021 37246 -3965 37499
rect 4761 37567 5507 37579
rect 4761 37511 5129 37567
rect 5185 37511 5507 37567
rect 4761 37499 5507 37511
rect 4761 37246 4817 37499
rect 5129 37246 5185 37499
rect 5451 37246 5507 37499
rect 14233 37568 14979 37580
rect 14233 37512 14601 37568
rect 14657 37512 14979 37568
rect 14233 37500 14979 37512
rect 14233 37247 14289 37500
rect 14601 37247 14657 37500
rect 14923 37247 14979 37500
rect 23705 37568 24451 37580
rect 23705 37512 24073 37568
rect 24129 37512 24451 37568
rect 23705 37500 24451 37512
rect 23705 37247 23761 37500
rect 24073 37247 24129 37500
rect 24395 37247 24451 37500
rect 33177 37568 33923 37580
rect 33177 37512 33545 37568
rect 33601 37512 33923 37568
rect 33177 37500 33923 37512
rect 33177 37247 33233 37500
rect 33545 37247 33601 37500
rect 33867 37247 33923 37500
rect 42649 37568 43395 37580
rect 42649 37512 43017 37568
rect 43073 37512 43395 37568
rect 42649 37500 43395 37512
rect 42649 37247 42705 37500
rect 43017 37247 43073 37500
rect 43339 37247 43395 37500
rect -4723 37244 -4643 37246
rect -4723 37124 -4711 37244
rect -4655 37124 -4643 37244
rect -4723 37122 -4643 37124
rect -4355 37244 -4275 37246
rect -4355 37124 -4343 37244
rect -4287 37124 -4275 37244
rect -4355 37122 -4275 37124
rect -4033 37244 -3953 37246
rect -4033 37123 -4021 37244
rect -3965 37123 -3953 37244
rect -4711 37114 -4655 37122
rect -4343 37114 -4287 37122
rect -4033 37121 -3953 37123
rect 4749 37244 4829 37246
rect 4749 37124 4761 37244
rect 4817 37124 4829 37244
rect 4749 37122 4829 37124
rect 5117 37244 5197 37246
rect 5117 37124 5129 37244
rect 5185 37124 5197 37244
rect 5117 37122 5197 37124
rect 5439 37244 5519 37246
rect 5439 37123 5451 37244
rect 5507 37123 5519 37244
rect 14221 37245 14301 37247
rect 14221 37125 14233 37245
rect 14289 37125 14301 37245
rect 14221 37123 14301 37125
rect 14589 37245 14669 37247
rect 14589 37125 14601 37245
rect 14657 37125 14669 37245
rect 14589 37123 14669 37125
rect 14911 37245 14991 37247
rect 14911 37124 14923 37245
rect 14979 37124 14991 37245
rect -4021 37113 -3965 37121
rect 4761 37114 4817 37122
rect 5129 37114 5185 37122
rect 5439 37121 5519 37123
rect 5451 37113 5507 37121
rect 14233 37115 14289 37123
rect 14601 37115 14657 37123
rect 14911 37122 14991 37124
rect 23693 37245 23773 37247
rect 23693 37125 23705 37245
rect 23761 37125 23773 37245
rect 23693 37123 23773 37125
rect 24061 37245 24141 37247
rect 24061 37125 24073 37245
rect 24129 37125 24141 37245
rect 24061 37123 24141 37125
rect 24383 37245 24463 37247
rect 24383 37124 24395 37245
rect 24451 37124 24463 37245
rect 14923 37114 14979 37122
rect 23705 37115 23761 37123
rect 24073 37115 24129 37123
rect 24383 37122 24463 37124
rect 33165 37245 33245 37247
rect 33165 37125 33177 37245
rect 33233 37125 33245 37245
rect 33165 37123 33245 37125
rect 33533 37245 33613 37247
rect 33533 37125 33545 37245
rect 33601 37125 33613 37245
rect 33533 37123 33613 37125
rect 33855 37245 33935 37247
rect 33855 37124 33867 37245
rect 33923 37124 33935 37245
rect 24395 37114 24451 37122
rect 33177 37115 33233 37123
rect 33545 37115 33601 37123
rect 33855 37122 33935 37124
rect 42637 37245 42717 37247
rect 42637 37125 42649 37245
rect 42705 37125 42717 37245
rect 42637 37123 42717 37125
rect 43005 37245 43085 37247
rect 43005 37125 43017 37245
rect 43073 37125 43085 37245
rect 43005 37123 43085 37125
rect 43327 37245 43407 37247
rect 43327 37124 43339 37245
rect 43395 37124 43407 37245
rect 33867 37114 33923 37122
rect 42649 37115 42705 37123
rect 43017 37115 43073 37123
rect 43327 37122 43407 37124
rect 43339 37114 43395 37122
rect -4527 36946 -4471 36954
rect -4159 36946 -4103 36954
rect 4945 36946 5001 36954
rect 5313 36946 5369 36954
rect 14417 36947 14473 36955
rect 14785 36947 14841 36955
rect 23889 36947 23945 36955
rect 24257 36947 24313 36955
rect 33361 36947 33417 36955
rect 33729 36947 33785 36955
rect 42833 36947 42889 36955
rect 43201 36947 43257 36955
rect -4539 36944 -4050 36946
rect -4539 36824 -4527 36944
rect -4471 36824 -4159 36944
rect -4103 36824 -4050 36944
rect -4539 36822 -4050 36824
rect 4933 36944 5422 36946
rect 4933 36824 4945 36944
rect 5001 36824 5313 36944
rect 5369 36824 5422 36944
rect 4933 36822 5422 36824
rect 14405 36945 14894 36947
rect 14405 36825 14417 36945
rect 14473 36825 14785 36945
rect 14841 36825 14894 36945
rect 14405 36823 14894 36825
rect 23877 36945 24366 36947
rect 23877 36825 23889 36945
rect 23945 36825 24257 36945
rect 24313 36825 24366 36945
rect 23877 36823 24366 36825
rect 33349 36945 33838 36947
rect 33349 36825 33361 36945
rect 33417 36825 33729 36945
rect 33785 36825 33838 36945
rect 33349 36823 33838 36825
rect 42821 36945 43310 36947
rect 42821 36825 42833 36945
rect 42889 36825 43201 36945
rect 43257 36825 43310 36945
rect 42821 36823 43310 36825
rect -4527 36814 -4471 36822
rect -4159 36814 -4050 36822
rect 4945 36814 5001 36822
rect 5313 36814 5422 36822
rect 14417 36815 14473 36823
rect 14785 36815 14894 36823
rect 23889 36815 23945 36823
rect 24257 36815 24366 36823
rect 33361 36815 33417 36823
rect 33729 36815 33838 36823
rect 42833 36815 42889 36823
rect 43201 36815 43310 36823
rect -4631 36748 -4551 36758
rect -4631 36692 -4619 36748
rect -4563 36692 -4551 36748
rect -4631 36682 -4551 36692
rect -4447 36748 -4367 36758
rect -4447 36692 -4435 36748
rect -4379 36692 -4367 36748
rect -4447 36682 -4367 36692
rect -4263 36748 -4183 36758
rect -4263 36692 -4251 36748
rect -4195 36692 -4183 36748
rect -4263 36682 -4183 36692
rect -5521 36598 -5433 36610
rect -4619 36600 -4563 36682
rect -5521 36542 -5507 36598
rect -5451 36542 -5433 36598
rect -5521 36530 -5433 36542
rect -4631 36598 -4551 36600
rect -4631 36542 -4619 36598
rect -4563 36542 -4551 36598
rect -4631 36540 -4551 36542
rect -5303 36482 -5233 36494
rect -5303 36426 -5291 36482
rect -5235 36426 -5233 36482
rect -5303 36414 -5233 36426
rect -5439 34277 -5369 34291
rect -5439 34221 -5427 34277
rect -5371 34221 -5369 34277
rect -5439 34209 -5369 34221
rect -8103 33372 -8027 33382
rect -8103 33316 -8093 33372
rect -8037 33316 -8027 33372
rect -8103 33306 -8027 33316
rect -5721 33375 -5639 33387
rect -5721 33319 -5707 33375
rect -5651 33319 -5639 33375
rect -5721 33307 -5639 33319
rect -6337 31969 -6017 31979
rect -9865 31462 -8693 31472
rect -9865 31222 -9853 31462
rect -9797 31222 -8761 31462
rect -8705 31222 -8693 31462
rect -9865 31212 -8693 31222
rect -10211 31005 -10131 31015
rect -9771 31005 -9693 31017
rect -11141 30949 -10199 31005
rect -10143 30949 -9751 31005
rect -9695 30949 -9693 31005
rect -10211 30939 -10131 30949
rect -9771 30937 -9693 30949
rect -8773 30927 -8693 31212
rect -8293 31462 -8213 31472
rect -8293 31222 -8281 31462
rect -8225 31222 -8213 31462
rect -8471 30927 -8401 30939
rect -8773 30871 -8459 30927
rect -8403 30871 -8401 30927
rect -8951 30849 -8881 30861
rect -11141 30793 -8939 30849
rect -8883 30793 -8881 30849
rect -11029 29507 -10973 30793
rect -8951 30781 -8881 30793
rect -9661 30567 -9581 30577
rect -9661 30511 -9649 30567
rect -9593 30511 -9581 30567
rect -9661 30325 -9581 30511
rect -9181 30567 -9101 30577
rect -9181 30511 -9169 30567
rect -9113 30511 -9101 30567
rect -9181 30501 -9101 30511
rect -8977 30567 -8897 30577
rect -8977 30511 -8965 30567
rect -8909 30511 -8897 30567
rect -8977 30325 -8897 30511
rect -8773 30567 -8693 30871
rect -8471 30859 -8401 30871
rect -8293 30927 -8213 31222
rect -6337 31169 -6327 31969
rect -6027 31169 -6017 31969
rect -6337 31159 -6017 31169
rect -7707 30973 -5915 30985
rect -8293 30871 -7936 30927
rect -8773 30511 -8761 30567
rect -8705 30511 -8693 30567
rect -8773 30501 -8693 30511
rect -8293 30567 -8213 30871
rect -8293 30511 -8281 30567
rect -8225 30511 -8213 30567
rect -8293 30501 -8213 30511
rect -9661 30253 -8897 30325
rect -8767 30199 -8143 30211
rect -9995 30166 -9895 30176
rect -9995 30090 -9985 30166
rect -9905 30090 -9895 30166
rect -9995 30080 -9895 30090
rect -8767 30059 -8755 30199
rect -8155 30059 -8143 30199
rect -10555 30042 -10475 30052
rect -8767 30047 -8143 30059
rect -10555 29802 -10543 30042
rect -10487 29802 -10475 30042
rect -7992 29829 -7936 30871
rect -7707 30833 -7695 30973
rect -5927 30833 -5915 30973
rect -7707 30821 -5915 30833
rect -7433 30570 -6669 30580
rect -7433 30330 -7421 30570
rect -7365 30330 -6737 30570
rect -6681 30330 -6669 30570
rect -7433 30320 -6669 30330
rect -6065 30286 -5985 30296
rect -6953 30236 -6465 30246
rect -6953 29996 -6941 30236
rect -6885 29996 -6533 30236
rect -6477 29996 -6465 30236
rect -6953 29986 -6465 29996
rect -7543 29829 -7447 29841
rect -10733 29507 -10663 29519
rect -11597 29451 -10721 29507
rect -10665 29451 -10663 29507
rect -12268 28112 -12188 28122
rect -12268 27872 -12256 28112
rect -12200 27872 -12188 28112
rect -12446 27577 -12376 27589
rect -13170 27521 -12434 27577
rect -12378 27521 -12376 27577
rect -12446 27509 -12376 27521
rect -12268 27577 -12188 27872
rect -11592 27608 -11536 29451
rect -10733 29439 -10663 29451
rect -10555 29507 -10475 29802
rect -8767 29799 -8143 29811
rect -8767 29659 -8755 29799
rect -8155 29659 -8143 29799
rect -7992 29773 -7523 29829
rect -7467 29773 -7447 29829
rect -7543 29761 -7447 29773
rect -6545 29751 -6465 29986
rect -6065 30046 -6053 30286
rect -5997 30046 -5985 30286
rect -6243 29751 -6173 29763
rect -6545 29695 -6231 29751
rect -6175 29695 -6173 29751
rect -6859 29673 -6763 29683
rect -8767 29647 -8143 29659
rect -7992 29617 -6839 29673
rect -6783 29617 -6763 29673
rect -10555 29451 -10117 29507
rect -10555 29147 -10475 29451
rect -10555 29091 -10543 29147
rect -10487 29091 -10475 29147
rect -10555 29081 -10475 29091
rect -10173 28665 -10117 29451
rect -9865 29122 -8693 29132
rect -9865 28882 -9853 29122
rect -9797 28882 -8761 29122
rect -8705 28882 -8693 29122
rect -9865 28872 -8693 28882
rect -9771 28665 -9693 28677
rect -10173 28609 -9751 28665
rect -9695 28609 -9693 28665
rect -9771 28597 -9693 28609
rect -8773 28587 -8693 28872
rect -8293 29122 -8213 29132
rect -8293 28882 -8281 29122
rect -8225 28882 -8213 29122
rect -8471 28587 -8401 28599
rect -8773 28531 -8459 28587
rect -8403 28531 -8401 28587
rect -8951 28509 -8881 28521
rect -11840 27577 -11764 27587
rect -12268 27521 -11830 27577
rect -11774 27521 -11764 27577
rect -12268 27217 -12188 27521
rect -11840 27511 -11764 27521
rect -11592 27478 -11536 27488
rect -11141 28453 -8939 28509
rect -8883 28453 -8881 28509
rect -12268 27161 -12256 27217
rect -12200 27161 -12188 27217
rect -12268 27151 -12188 27161
rect -11141 26474 -11085 28453
rect -8951 28441 -8881 28453
rect -9661 28227 -9581 28237
rect -9661 28171 -9649 28227
rect -9593 28171 -9581 28227
rect -9661 27985 -9581 28171
rect -9181 28227 -9101 28237
rect -9181 28171 -9169 28227
rect -9113 28171 -9101 28227
rect -9181 28161 -9101 28171
rect -8977 28227 -8897 28237
rect -8977 28171 -8965 28227
rect -8909 28171 -8897 28227
rect -8977 27985 -8897 28171
rect -8773 28227 -8693 28531
rect -8471 28519 -8401 28531
rect -8293 28587 -8213 28882
rect -7992 28587 -7936 29617
rect -6859 29607 -6763 29617
rect -6545 29401 -6465 29695
rect -6243 29683 -6173 29695
rect -6065 29751 -5985 30046
rect -5427 29881 -5371 34209
rect -5291 31968 -5235 36414
rect -4619 36226 -4563 36540
rect -4435 36484 -4379 36682
rect -4447 36482 -4367 36484
rect -4447 36426 -4435 36482
rect -4379 36426 -4367 36482
rect -4447 36424 -4367 36426
rect -4435 36226 -4379 36424
rect -4251 36368 -4195 36682
rect -4118 36484 -4050 36814
rect 4841 36748 4921 36758
rect 4841 36692 4853 36748
rect 4909 36692 4921 36748
rect 4841 36682 4921 36692
rect 5025 36748 5105 36758
rect 5025 36692 5037 36748
rect 5093 36692 5105 36748
rect 5025 36682 5105 36692
rect 5209 36748 5289 36758
rect 5209 36692 5221 36748
rect 5277 36692 5289 36748
rect 5209 36682 5289 36692
rect 3951 36598 4039 36610
rect 4853 36600 4909 36682
rect 3951 36542 3965 36598
rect 4021 36542 4039 36598
rect 3951 36530 4039 36542
rect 4841 36598 4921 36600
rect 4841 36542 4853 36598
rect 4909 36542 4921 36598
rect 4841 36540 4921 36542
rect -4118 36482 -4038 36484
rect -4118 36426 -4106 36482
rect -4050 36426 -4038 36482
rect -4118 36424 -4038 36426
rect -3851 36482 -3781 36494
rect -3851 36426 -3849 36482
rect -3793 36426 -3781 36482
rect -4263 36366 -4183 36368
rect -4263 36310 -4251 36366
rect -4195 36310 -4183 36366
rect -4263 36308 -4183 36310
rect -4251 36226 -4195 36308
rect -4631 36216 -4551 36226
rect -4631 36160 -4619 36216
rect -4563 36160 -4551 36216
rect -4631 36150 -4551 36160
rect -4447 36216 -4367 36226
rect -4447 36160 -4435 36216
rect -4379 36160 -4367 36216
rect -4447 36150 -4367 36160
rect -4263 36216 -4183 36226
rect -4263 36160 -4251 36216
rect -4195 36160 -4183 36216
rect -4263 36150 -4183 36160
rect -4118 36094 -4050 36424
rect -3851 36416 -3781 36426
rect 4169 36482 4239 36494
rect 4169 36426 4181 36482
rect 4237 36426 4239 36482
rect -4159 36086 -4050 36094
rect -4171 36084 -4050 36086
rect -4171 35964 -4159 36084
rect -4103 35964 -4050 36084
rect -4171 35962 -4050 35964
rect -4159 35954 -4103 35962
rect -4856 35697 -3958 35709
rect -4856 35641 -4844 35697
rect -4788 35641 -4026 35697
rect -3970 35641 -3958 35697
rect -4856 35629 -3958 35641
rect -3849 35472 -3793 36416
rect 4169 36414 4239 36426
rect -3685 35579 -3605 35589
rect -3685 35523 -3673 35579
rect -3617 35523 -3605 35579
rect -3685 35521 -3605 35523
rect -3851 35469 -3781 35472
rect -3851 35415 -3849 35469
rect -3793 35415 -3781 35469
rect -3851 35403 -3781 35415
rect -4711 35362 -3965 35374
rect -4711 35306 -4343 35362
rect -4287 35306 -3965 35362
rect -4711 35294 -3965 35306
rect -4711 35041 -4655 35294
rect -4343 35041 -4287 35294
rect -4021 35041 -3965 35294
rect -4723 35039 -4643 35041
rect -4723 34919 -4711 35039
rect -4655 34919 -4643 35039
rect -4723 34917 -4643 34919
rect -4355 35039 -4275 35041
rect -4355 34919 -4343 35039
rect -4287 34919 -4275 35039
rect -4355 34917 -4275 34919
rect -4033 35039 -3953 35041
rect -4033 34918 -4021 35039
rect -3965 34918 -3953 35039
rect -4711 34909 -4655 34917
rect -4343 34909 -4287 34917
rect -4033 34916 -3953 34918
rect -4021 34908 -3965 34916
rect -4527 34741 -4471 34749
rect -4159 34741 -4103 34749
rect -4539 34739 -4050 34741
rect -4539 34619 -4527 34739
rect -4471 34619 -4159 34739
rect -4103 34619 -4050 34739
rect -4539 34617 -4050 34619
rect -4527 34609 -4471 34617
rect -4159 34609 -4050 34617
rect -4631 34543 -4551 34553
rect -4631 34487 -4619 34543
rect -4563 34487 -4551 34543
rect -4631 34477 -4551 34487
rect -4447 34543 -4367 34553
rect -4447 34487 -4435 34543
rect -4379 34487 -4367 34543
rect -4447 34477 -4367 34487
rect -4263 34543 -4183 34553
rect -4263 34487 -4251 34543
rect -4195 34487 -4183 34543
rect -4263 34477 -4183 34487
rect -4619 34395 -4563 34477
rect -4631 34393 -4551 34395
rect -4631 34337 -4619 34393
rect -4563 34337 -4551 34393
rect -4631 34335 -4551 34337
rect -4619 34021 -4563 34335
rect -4435 34279 -4379 34477
rect -4447 34277 -4367 34279
rect -4447 34221 -4435 34277
rect -4379 34221 -4367 34277
rect -4447 34219 -4367 34221
rect -4435 34021 -4379 34219
rect -4251 34163 -4195 34477
rect -4118 34279 -4050 34609
rect -3673 34287 -3617 35521
rect -3225 35362 -2479 35374
rect -3225 35306 -2857 35362
rect -2801 35306 -2479 35362
rect -3225 35294 -2479 35306
rect -3225 35041 -3169 35294
rect -2857 35041 -2801 35294
rect -2535 35041 -2479 35294
rect -3237 35039 -3157 35041
rect -3237 34919 -3225 35039
rect -3169 34919 -3157 35039
rect -3237 34917 -3157 34919
rect -2869 35039 -2789 35041
rect -2869 34919 -2857 35039
rect -2801 34919 -2789 35039
rect -2869 34917 -2789 34919
rect -2547 35039 -2467 35041
rect -2547 34918 -2535 35039
rect -2479 34918 -2467 35039
rect -3225 34909 -3169 34917
rect -2857 34909 -2801 34917
rect -2547 34916 -2467 34918
rect -2535 34908 -2479 34916
rect -3041 34741 -2985 34749
rect -2673 34741 -2617 34749
rect -3053 34739 -2564 34741
rect -3053 34619 -3041 34739
rect -2985 34619 -2673 34739
rect -2617 34619 -2564 34739
rect -3053 34617 -2564 34619
rect -3041 34609 -2985 34617
rect -2673 34609 -2564 34617
rect -3145 34543 -3065 34553
rect -3145 34487 -3133 34543
rect -3077 34487 -3065 34543
rect -3145 34477 -3065 34487
rect -2961 34543 -2881 34553
rect -2961 34487 -2949 34543
rect -2893 34487 -2881 34543
rect -2961 34477 -2881 34487
rect -2777 34543 -2697 34553
rect -2777 34487 -2765 34543
rect -2709 34487 -2697 34543
rect -2777 34477 -2697 34487
rect -3133 34395 -3077 34477
rect -3145 34393 -3065 34395
rect -3145 34337 -3133 34393
rect -3077 34337 -3065 34393
rect -3145 34335 -3065 34337
rect -4118 34277 -4038 34279
rect -4118 34221 -4106 34277
rect -4050 34221 -4038 34277
rect -4118 34219 -4038 34221
rect -3675 34277 -3615 34287
rect -3675 34221 -3673 34277
rect -3617 34221 -3615 34277
rect -4263 34161 -4183 34163
rect -4263 34105 -4251 34161
rect -4195 34105 -4183 34161
rect -4263 34103 -4183 34105
rect -4251 34021 -4195 34103
rect -4631 34011 -4551 34021
rect -4631 33955 -4619 34011
rect -4563 33955 -4551 34011
rect -4631 33945 -4551 33955
rect -4447 34011 -4367 34021
rect -4447 33955 -4435 34011
rect -4379 33955 -4367 34011
rect -4447 33945 -4367 33955
rect -4263 34011 -4183 34021
rect -4263 33955 -4251 34011
rect -4195 33955 -4183 34011
rect -4263 33945 -4183 33955
rect -4118 33889 -4050 34219
rect -3675 34209 -3615 34221
rect -4159 33881 -4050 33889
rect -4171 33879 -4050 33881
rect -4171 33759 -4159 33879
rect -4103 33759 -4050 33879
rect -4171 33757 -4050 33759
rect -4159 33749 -4103 33757
rect -4856 33492 -3960 33504
rect -4856 33436 -4844 33492
rect -4788 33436 -4026 33492
rect -3970 33436 -3960 33492
rect -4856 33424 -3960 33436
rect -3673 33266 -3617 34209
rect -3133 34021 -3077 34335
rect -2949 34279 -2893 34477
rect -2961 34277 -2881 34279
rect -2961 34221 -2949 34277
rect -2893 34221 -2881 34277
rect -2961 34219 -2881 34221
rect -2949 34021 -2893 34219
rect -2765 34163 -2709 34477
rect -2632 34279 -2564 34609
rect -2632 34277 -2552 34279
rect -2632 34221 -2620 34277
rect -2564 34221 -2552 34277
rect -2632 34219 -2552 34221
rect -2365 34277 -2295 34289
rect 4033 34277 4103 34291
rect -2365 34221 -2363 34277
rect -2307 34221 -1609 34277
rect -2777 34161 -2697 34163
rect -2777 34105 -2765 34161
rect -2709 34105 -2697 34161
rect -2777 34103 -2697 34105
rect -2765 34021 -2709 34103
rect -3145 34011 -3065 34021
rect -3145 33955 -3133 34011
rect -3077 33955 -3065 34011
rect -3145 33945 -3065 33955
rect -2961 34011 -2881 34021
rect -2961 33955 -2949 34011
rect -2893 33955 -2881 34011
rect -2961 33945 -2881 33955
rect -2777 34011 -2697 34021
rect -2777 33955 -2765 34011
rect -2709 33955 -2697 34011
rect -2777 33945 -2697 33955
rect -2632 33889 -2564 34219
rect -2365 34211 -2295 34221
rect -2673 33881 -2564 33889
rect -2685 33879 -2564 33881
rect -2685 33759 -2673 33879
rect -2617 33759 -2564 33879
rect -2685 33757 -2564 33759
rect -2673 33749 -2617 33757
rect -3370 33492 -2474 33504
rect -3370 33436 -3358 33492
rect -3302 33436 -2540 33492
rect -2484 33436 -2474 33492
rect -3370 33424 -2474 33436
rect -2363 33267 -2307 34211
rect -2199 33375 -2119 33385
rect -2199 33319 -2187 33375
rect -2131 33319 -2119 33375
rect -2199 33317 -2119 33319
rect -3675 33264 -3605 33266
rect -3675 33208 -3673 33264
rect -3617 33208 -3605 33264
rect -3675 33196 -3605 33208
rect -2375 33265 -2295 33267
rect -2375 33209 -2363 33265
rect -2307 33209 -2295 33265
rect -2375 33197 -2295 33209
rect -4711 33157 -3965 33169
rect -4711 33101 -4343 33157
rect -4287 33101 -3965 33157
rect -4711 33089 -3965 33101
rect -4711 32836 -4655 33089
rect -4343 32836 -4287 33089
rect -4021 32836 -3965 33089
rect -3225 33158 -2479 33170
rect -3225 33102 -2857 33158
rect -2801 33102 -2479 33158
rect -3225 33090 -2479 33102
rect -3225 32837 -3169 33090
rect -2857 32837 -2801 33090
rect -2535 32837 -2479 33090
rect -4723 32834 -4643 32836
rect -4723 32714 -4711 32834
rect -4655 32714 -4643 32834
rect -4723 32712 -4643 32714
rect -4355 32834 -4275 32836
rect -4355 32714 -4343 32834
rect -4287 32714 -4275 32834
rect -4355 32712 -4275 32714
rect -4033 32834 -3953 32836
rect -4033 32713 -4021 32834
rect -3965 32713 -3953 32834
rect -3237 32835 -3157 32837
rect -3237 32715 -3225 32835
rect -3169 32715 -3157 32835
rect -3237 32713 -3157 32715
rect -2869 32835 -2789 32837
rect -2869 32715 -2857 32835
rect -2801 32715 -2789 32835
rect -2869 32713 -2789 32715
rect -2547 32835 -2467 32837
rect -2547 32714 -2535 32835
rect -2479 32714 -2467 32835
rect -4711 32704 -4655 32712
rect -4343 32704 -4287 32712
rect -4033 32711 -3953 32713
rect -4021 32703 -3965 32711
rect -3225 32705 -3169 32713
rect -2857 32705 -2801 32713
rect -2547 32712 -2467 32714
rect -2535 32704 -2479 32712
rect -4527 32536 -4471 32544
rect -4159 32536 -4103 32544
rect -3041 32537 -2985 32545
rect -2673 32537 -2617 32545
rect -4539 32534 -4050 32536
rect -4539 32414 -4527 32534
rect -4471 32414 -4159 32534
rect -4103 32414 -4050 32534
rect -4539 32412 -4050 32414
rect -3053 32535 -2564 32537
rect -3053 32415 -3041 32535
rect -2985 32415 -2673 32535
rect -2617 32415 -2564 32535
rect -3053 32413 -2564 32415
rect -4527 32404 -4471 32412
rect -4159 32404 -4050 32412
rect -3041 32405 -2985 32413
rect -2673 32405 -2564 32413
rect -4631 32338 -4551 32348
rect -4631 32282 -4619 32338
rect -4563 32282 -4551 32338
rect -4631 32272 -4551 32282
rect -4447 32338 -4367 32348
rect -4447 32282 -4435 32338
rect -4379 32282 -4367 32338
rect -4447 32272 -4367 32282
rect -4263 32338 -4183 32348
rect -4263 32282 -4251 32338
rect -4195 32282 -4183 32338
rect -4263 32272 -4183 32282
rect -4619 32190 -4563 32272
rect -4631 32188 -4551 32190
rect -4631 32132 -4619 32188
rect -4563 32132 -4551 32188
rect -4631 32130 -4551 32132
rect -5303 31956 -5233 31968
rect -5303 31900 -5291 31956
rect -5235 31900 -5233 31956
rect -5303 31888 -5233 31900
rect -4619 31816 -4563 32130
rect -4435 32074 -4379 32272
rect -4447 32072 -4367 32074
rect -4447 32016 -4435 32072
rect -4379 32016 -4367 32072
rect -4447 32014 -4367 32016
rect -4435 31816 -4379 32014
rect -4251 31958 -4195 32272
rect -4118 32074 -4050 32404
rect -3145 32339 -3065 32349
rect -3145 32283 -3133 32339
rect -3077 32283 -3065 32339
rect -3145 32273 -3065 32283
rect -2961 32339 -2881 32349
rect -2961 32283 -2949 32339
rect -2893 32283 -2881 32339
rect -2961 32273 -2881 32283
rect -2777 32339 -2697 32349
rect -2777 32283 -2765 32339
rect -2709 32283 -2697 32339
rect -2777 32273 -2697 32283
rect -3133 32191 -3077 32273
rect -3145 32189 -3065 32191
rect -3145 32133 -3133 32189
rect -3077 32133 -3065 32189
rect -3145 32131 -3065 32133
rect -4118 32072 -4038 32074
rect -4118 32016 -4106 32072
rect -4050 32016 -4038 32072
rect -4118 32014 -4038 32016
rect -3851 32072 -3781 32084
rect -3851 32016 -3849 32072
rect -3793 32016 -3781 32072
rect -4263 31956 -4183 31958
rect -4263 31900 -4251 31956
rect -4195 31900 -4183 31956
rect -4263 31898 -4183 31900
rect -4251 31816 -4195 31898
rect -4631 31806 -4551 31816
rect -4631 31750 -4619 31806
rect -4563 31750 -4551 31806
rect -4631 31740 -4551 31750
rect -4447 31806 -4367 31816
rect -4447 31750 -4435 31806
rect -4379 31750 -4367 31806
rect -4447 31740 -4367 31750
rect -4263 31806 -4183 31816
rect -4263 31750 -4251 31806
rect -4195 31750 -4183 31806
rect -4263 31740 -4183 31750
rect -4118 31684 -4050 32014
rect -3851 32006 -3781 32016
rect -4159 31676 -4050 31684
rect -4171 31674 -4050 31676
rect -4171 31554 -4159 31674
rect -4103 31554 -4050 31674
rect -4171 31552 -4050 31554
rect -4159 31544 -4103 31552
rect -4856 31287 -3960 31299
rect -4856 31231 -4844 31287
rect -4788 31231 -4026 31287
rect -3970 31231 -3960 31287
rect -4856 31219 -3960 31231
rect -3849 31062 -3793 32006
rect -3133 31817 -3077 32131
rect -2949 32075 -2893 32273
rect -2961 32073 -2881 32075
rect -2961 32017 -2949 32073
rect -2893 32017 -2881 32073
rect -2961 32015 -2881 32017
rect -2949 31817 -2893 32015
rect -2765 31959 -2709 32273
rect -2632 32075 -2564 32405
rect -2187 32083 -2131 33317
rect -2632 32073 -2552 32075
rect -2632 32017 -2620 32073
rect -2564 32017 -2552 32073
rect -2632 32015 -2552 32017
rect -2189 32073 -2119 32083
rect -2189 32017 -2187 32073
rect -2131 32017 -2039 32073
rect -2777 31957 -2697 31959
rect -2777 31901 -2765 31957
rect -2709 31901 -2697 31957
rect -2777 31899 -2697 31901
rect -2765 31817 -2709 31899
rect -3145 31807 -3065 31817
rect -3145 31751 -3133 31807
rect -3077 31751 -3065 31807
rect -3145 31741 -3065 31751
rect -2961 31807 -2881 31817
rect -2961 31751 -2949 31807
rect -2893 31751 -2881 31807
rect -2961 31741 -2881 31751
rect -2777 31807 -2697 31817
rect -2777 31751 -2765 31807
rect -2709 31751 -2697 31807
rect -2777 31741 -2697 31751
rect -2632 31685 -2564 32015
rect -2189 32005 -2119 32017
rect -2673 31677 -2564 31685
rect -2685 31675 -2564 31677
rect -2685 31555 -2673 31675
rect -2617 31555 -2564 31675
rect -2685 31553 -2564 31555
rect -2673 31545 -2617 31553
rect -3370 31288 -2474 31300
rect -3370 31232 -3358 31288
rect -3302 31232 -2540 31288
rect -2484 31232 -2474 31288
rect -3370 31220 -2474 31232
rect -3685 31169 -3605 31179
rect -3685 31113 -3673 31169
rect -3617 31113 -3605 31169
rect -3685 31111 -3605 31113
rect -3851 31059 -3781 31062
rect -3851 31005 -3849 31059
rect -3793 31005 -3781 31059
rect -3851 30993 -3781 31005
rect -4711 30952 -3965 30964
rect -4711 30896 -4343 30952
rect -4287 30896 -3965 30952
rect -4711 30884 -3965 30896
rect -4711 30631 -4655 30884
rect -4343 30631 -4287 30884
rect -4021 30631 -3965 30884
rect -4723 30629 -4643 30631
rect -4723 30509 -4711 30629
rect -4655 30509 -4643 30629
rect -4723 30507 -4643 30509
rect -4355 30629 -4275 30631
rect -4355 30509 -4343 30629
rect -4287 30509 -4275 30629
rect -4355 30507 -4275 30509
rect -4033 30629 -3953 30631
rect -4033 30508 -4021 30629
rect -3965 30508 -3953 30629
rect -4711 30499 -4655 30507
rect -4343 30499 -4287 30507
rect -4033 30506 -3953 30508
rect -4021 30498 -3965 30506
rect -4527 30331 -4471 30339
rect -4159 30331 -4103 30339
rect -4539 30329 -4050 30331
rect -4539 30209 -4527 30329
rect -4471 30209 -4159 30329
rect -4103 30209 -4050 30329
rect -4539 30207 -4050 30209
rect -4527 30199 -4471 30207
rect -4159 30199 -4050 30207
rect -4631 30133 -4551 30143
rect -4631 30077 -4619 30133
rect -4563 30077 -4551 30133
rect -4631 30067 -4551 30077
rect -4447 30133 -4367 30143
rect -4447 30077 -4435 30133
rect -4379 30077 -4367 30133
rect -4447 30067 -4367 30077
rect -4263 30133 -4183 30143
rect -4263 30077 -4251 30133
rect -4195 30077 -4183 30133
rect -4263 30067 -4183 30077
rect -4619 29985 -4563 30067
rect -4631 29983 -4551 29985
rect -4631 29927 -4619 29983
rect -4563 29927 -4551 29983
rect -4631 29925 -4551 29927
rect -5439 29867 -5369 29881
rect -5439 29811 -5427 29867
rect -5371 29811 -5369 29867
rect -5439 29799 -5369 29811
rect -5673 29751 -5595 29762
rect -6065 29750 -5595 29751
rect -6065 29696 -5661 29750
rect -5607 29696 -5595 29750
rect -6065 29695 -5595 29696
rect -7637 29391 -6465 29401
rect -7637 29335 -7625 29391
rect -7569 29335 -6737 29391
rect -6681 29335 -6465 29391
rect -7637 29325 -6465 29335
rect -6065 29391 -5985 29695
rect -5673 29684 -5595 29695
rect -6065 29335 -6053 29391
rect -5997 29335 -5985 29391
rect -6065 29325 -5985 29335
rect -7707 29013 -5915 29025
rect -7707 28873 -7695 29013
rect -5927 28873 -5915 29013
rect -5622 28964 -5536 28976
rect -5427 28968 -5371 29799
rect -4619 29611 -4563 29925
rect -4435 29869 -4379 30067
rect -4447 29867 -4367 29869
rect -4447 29811 -4435 29867
rect -4379 29811 -4367 29867
rect -4447 29809 -4367 29811
rect -4435 29611 -4379 29809
rect -4251 29753 -4195 30067
rect -4118 29869 -4050 30199
rect -3673 29879 -3617 31111
rect -1665 31005 -1609 34221
rect 4033 34221 4045 34277
rect 4101 34221 4103 34277
rect 4033 34209 4103 34221
rect 3751 33375 3833 33387
rect 3751 33319 3765 33375
rect 3821 33319 3833 33375
rect 3751 33307 3833 33319
rect -1255 31969 -1035 31979
rect -1255 31169 -1245 31969
rect -1045 31169 -1035 31969
rect 3135 31969 3455 31979
rect -393 31462 779 31472
rect -393 31222 -381 31462
rect -325 31222 711 31462
rect 767 31222 779 31462
rect -393 31212 779 31222
rect -1255 31159 -1035 31169
rect -299 31005 -221 31017
rect -1669 30949 -279 31005
rect -223 30949 -221 31005
rect -299 30937 -221 30949
rect 699 30927 779 31212
rect 1179 31462 1259 31472
rect 1179 31222 1191 31462
rect 1247 31222 1259 31462
rect 1001 30927 1071 30939
rect 699 30871 1013 30927
rect 1069 30871 1071 30927
rect 521 30849 591 30861
rect -1669 30793 533 30849
rect 589 30793 591 30849
rect -4118 29867 -4038 29869
rect -4118 29811 -4106 29867
rect -4050 29811 -4038 29867
rect -4118 29809 -4038 29811
rect -3675 29867 -3615 29879
rect -3675 29811 -3673 29867
rect -3617 29811 -3615 29867
rect -4263 29751 -4183 29753
rect -4263 29695 -4251 29751
rect -4195 29695 -4183 29751
rect -4263 29693 -4183 29695
rect -4251 29611 -4195 29693
rect -4631 29601 -4551 29611
rect -4631 29545 -4619 29601
rect -4563 29545 -4551 29601
rect -4631 29535 -4551 29545
rect -4447 29601 -4367 29611
rect -4447 29545 -4435 29601
rect -4379 29545 -4367 29601
rect -4447 29535 -4367 29545
rect -4263 29601 -4183 29611
rect -4263 29545 -4251 29601
rect -4195 29545 -4183 29601
rect -4263 29535 -4183 29545
rect -4118 29479 -4050 29809
rect -3675 29799 -3615 29811
rect -1557 29508 -1501 30793
rect 521 30781 591 30793
rect -189 30567 -109 30577
rect -189 30511 -177 30567
rect -121 30511 -109 30567
rect -189 30325 -109 30511
rect 291 30567 371 30577
rect 291 30511 303 30567
rect 359 30511 371 30567
rect 291 30501 371 30511
rect 495 30567 575 30577
rect 495 30511 507 30567
rect 563 30511 575 30567
rect 495 30325 575 30511
rect 699 30567 779 30871
rect 1001 30859 1071 30871
rect 1179 30927 1259 31222
rect 3135 31169 3145 31969
rect 3445 31169 3455 31969
rect 3135 31159 3455 31169
rect 1765 30973 3557 30985
rect 1179 30871 1536 30927
rect 699 30511 711 30567
rect 767 30511 779 30567
rect 699 30501 779 30511
rect 1179 30567 1259 30871
rect 1179 30511 1191 30567
rect 1247 30511 1259 30567
rect 1179 30501 1259 30511
rect -189 30253 575 30325
rect 705 30199 1329 30211
rect 705 30059 717 30199
rect 1317 30059 1329 30199
rect -1083 30042 -1003 30052
rect 705 30047 1329 30059
rect -1083 29802 -1071 30042
rect -1015 29802 -1003 30042
rect 1480 29829 1536 30871
rect 1765 30833 1777 30973
rect 3545 30833 3557 30973
rect 1765 30821 3557 30833
rect 2039 30570 2803 30580
rect 2039 30330 2051 30570
rect 2107 30330 2735 30570
rect 2791 30330 2803 30570
rect 2039 30320 2803 30330
rect 3407 30286 3487 30296
rect 2519 30236 3007 30246
rect 2519 29996 2531 30236
rect 2587 29996 2939 30236
rect 2995 29996 3007 30236
rect 2519 29986 3007 29996
rect 1929 29829 2025 29841
rect -4159 29471 -4050 29479
rect -4171 29469 -4050 29471
rect -4171 29349 -4159 29469
rect -4103 29349 -4050 29469
rect -2069 29507 -1501 29508
rect -1261 29507 -1191 29519
rect -2069 29452 -1249 29507
rect -4171 29347 -4050 29349
rect -4159 29339 -4103 29347
rect -4856 29082 -3958 29094
rect -4856 29026 -4844 29082
rect -4788 29026 -4026 29082
rect -3970 29026 -3958 29082
rect -4856 29014 -3958 29026
rect -5622 28908 -5610 28964
rect -5554 28908 -5536 28964
rect -5622 28896 -5536 28908
rect -5429 28964 -5369 28968
rect -5429 28908 -5427 28964
rect -5371 28908 -5369 28964
rect -5429 28896 -5369 28908
rect -7707 28861 -5915 28873
rect -8293 28531 -7936 28587
rect -6337 28689 -6017 28699
rect -8773 28171 -8761 28227
rect -8705 28171 -8693 28227
rect -8773 28161 -8693 28171
rect -8293 28227 -8213 28531
rect -8293 28171 -8281 28227
rect -8225 28171 -8213 28227
rect -8293 28161 -8213 28171
rect -9661 27913 -8897 27985
rect -6337 27889 -6327 28689
rect -6027 27889 -6017 28689
rect -6337 27879 -6017 27889
rect -2064 27609 -2008 29452
rect -1557 29451 -1249 29452
rect -1193 29451 -1191 29507
rect -1261 29439 -1191 29451
rect -1083 29507 -1003 29802
rect 705 29799 1329 29811
rect 705 29659 717 29799
rect 1317 29659 1329 29799
rect 1480 29773 1949 29829
rect 2005 29773 2025 29829
rect 1929 29761 2025 29773
rect 2927 29751 3007 29986
rect 3407 30046 3419 30286
rect 3475 30046 3487 30286
rect 3229 29751 3299 29763
rect 2927 29695 3241 29751
rect 3297 29695 3299 29751
rect 2613 29673 2709 29683
rect 705 29647 1329 29659
rect 1480 29617 2633 29673
rect 2689 29617 2709 29673
rect -1083 29451 -645 29507
rect -1083 29147 -1003 29451
rect -1083 29091 -1071 29147
rect -1015 29091 -1003 29147
rect -1083 29081 -1003 29091
rect -701 28665 -645 29451
rect -393 29122 779 29132
rect -393 28882 -381 29122
rect -325 28882 711 29122
rect 767 28882 779 29122
rect -393 28872 779 28882
rect -299 28665 -221 28677
rect -701 28609 -279 28665
rect -223 28609 -221 28665
rect -299 28597 -221 28609
rect 699 28587 779 28872
rect 1179 29122 1259 29132
rect 1179 28882 1191 29122
rect 1247 28882 1259 29122
rect 1001 28587 1071 28599
rect 699 28531 1013 28587
rect 1069 28531 1071 28587
rect 521 28509 591 28521
rect -2064 27479 -2008 27489
rect -1669 28453 533 28509
rect 589 28453 591 28509
rect -5081 26474 -5025 26489
rect -11141 26418 -5025 26474
rect -1669 26484 -1613 28453
rect 521 28441 591 28453
rect -189 28227 -109 28237
rect -189 28171 -177 28227
rect -121 28171 -109 28227
rect -189 27985 -109 28171
rect 291 28227 371 28237
rect 291 28171 303 28227
rect 359 28171 371 28227
rect 291 28161 371 28171
rect 495 28227 575 28237
rect 495 28171 507 28227
rect 563 28171 575 28227
rect 495 27985 575 28171
rect 699 28227 779 28531
rect 1001 28519 1071 28531
rect 1179 28587 1259 28882
rect 1480 28587 1536 29617
rect 2613 29607 2709 29617
rect 2927 29401 3007 29695
rect 3229 29683 3299 29695
rect 3407 29751 3487 30046
rect 4045 29881 4101 34209
rect 4181 31968 4237 36414
rect 4853 36226 4909 36540
rect 5037 36484 5093 36682
rect 5025 36482 5105 36484
rect 5025 36426 5037 36482
rect 5093 36426 5105 36482
rect 5025 36424 5105 36426
rect 5037 36226 5093 36424
rect 5221 36368 5277 36682
rect 5354 36484 5422 36814
rect 14313 36749 14393 36759
rect 14313 36693 14325 36749
rect 14381 36693 14393 36749
rect 14313 36683 14393 36693
rect 14497 36749 14577 36759
rect 14497 36693 14509 36749
rect 14565 36693 14577 36749
rect 14497 36683 14577 36693
rect 14681 36749 14761 36759
rect 14681 36693 14693 36749
rect 14749 36693 14761 36749
rect 14681 36683 14761 36693
rect 13423 36599 13511 36611
rect 14325 36601 14381 36683
rect 13423 36543 13437 36599
rect 13493 36543 13511 36599
rect 13423 36531 13511 36543
rect 14313 36599 14393 36601
rect 14313 36543 14325 36599
rect 14381 36543 14393 36599
rect 14313 36541 14393 36543
rect 5354 36482 5434 36484
rect 5354 36426 5366 36482
rect 5422 36426 5434 36482
rect 5354 36424 5434 36426
rect 5621 36482 5691 36494
rect 5621 36426 5623 36482
rect 5679 36426 5691 36482
rect 5209 36366 5289 36368
rect 5209 36310 5221 36366
rect 5277 36310 5289 36366
rect 5209 36308 5289 36310
rect 5221 36226 5277 36308
rect 4841 36216 4921 36226
rect 4841 36160 4853 36216
rect 4909 36160 4921 36216
rect 4841 36150 4921 36160
rect 5025 36216 5105 36226
rect 5025 36160 5037 36216
rect 5093 36160 5105 36216
rect 5025 36150 5105 36160
rect 5209 36216 5289 36226
rect 5209 36160 5221 36216
rect 5277 36160 5289 36216
rect 5209 36150 5289 36160
rect 5354 36094 5422 36424
rect 5621 36416 5691 36426
rect 13641 36483 13711 36495
rect 13641 36427 13653 36483
rect 13709 36427 13711 36483
rect 5313 36086 5422 36094
rect 5301 36084 5422 36086
rect 5301 35964 5313 36084
rect 5369 35964 5422 36084
rect 5301 35962 5422 35964
rect 5313 35954 5369 35962
rect 4616 35697 5514 35709
rect 4616 35641 4628 35697
rect 4684 35641 5446 35697
rect 5502 35641 5514 35697
rect 4616 35629 5514 35641
rect 5623 35472 5679 36416
rect 13641 36415 13711 36427
rect 5787 35579 5867 35589
rect 5787 35523 5799 35579
rect 5855 35523 5867 35579
rect 5787 35521 5867 35523
rect 5621 35469 5691 35472
rect 5621 35415 5623 35469
rect 5679 35415 5691 35469
rect 5621 35403 5691 35415
rect 4761 35362 5507 35374
rect 4761 35306 5129 35362
rect 5185 35306 5507 35362
rect 4761 35294 5507 35306
rect 4761 35041 4817 35294
rect 5129 35041 5185 35294
rect 5451 35041 5507 35294
rect 4749 35039 4829 35041
rect 4749 34919 4761 35039
rect 4817 34919 4829 35039
rect 4749 34917 4829 34919
rect 5117 35039 5197 35041
rect 5117 34919 5129 35039
rect 5185 34919 5197 35039
rect 5117 34917 5197 34919
rect 5439 35039 5519 35041
rect 5439 34918 5451 35039
rect 5507 34918 5519 35039
rect 4761 34909 4817 34917
rect 5129 34909 5185 34917
rect 5439 34916 5519 34918
rect 5451 34908 5507 34916
rect 4945 34741 5001 34749
rect 5313 34741 5369 34749
rect 4933 34739 5422 34741
rect 4933 34619 4945 34739
rect 5001 34619 5313 34739
rect 5369 34619 5422 34739
rect 4933 34617 5422 34619
rect 4945 34609 5001 34617
rect 5313 34609 5422 34617
rect 4841 34543 4921 34553
rect 4841 34487 4853 34543
rect 4909 34487 4921 34543
rect 4841 34477 4921 34487
rect 5025 34543 5105 34553
rect 5025 34487 5037 34543
rect 5093 34487 5105 34543
rect 5025 34477 5105 34487
rect 5209 34543 5289 34553
rect 5209 34487 5221 34543
rect 5277 34487 5289 34543
rect 5209 34477 5289 34487
rect 4853 34395 4909 34477
rect 4841 34393 4921 34395
rect 4841 34337 4853 34393
rect 4909 34337 4921 34393
rect 4841 34335 4921 34337
rect 4853 34021 4909 34335
rect 5037 34279 5093 34477
rect 5025 34277 5105 34279
rect 5025 34221 5037 34277
rect 5093 34221 5105 34277
rect 5025 34219 5105 34221
rect 5037 34021 5093 34219
rect 5221 34163 5277 34477
rect 5354 34279 5422 34609
rect 5799 34287 5855 35521
rect 6247 35362 6993 35374
rect 6247 35306 6615 35362
rect 6671 35306 6993 35362
rect 6247 35294 6993 35306
rect 6247 35041 6303 35294
rect 6615 35041 6671 35294
rect 6937 35041 6993 35294
rect 6235 35039 6315 35041
rect 6235 34919 6247 35039
rect 6303 34919 6315 35039
rect 6235 34917 6315 34919
rect 6603 35039 6683 35041
rect 6603 34919 6615 35039
rect 6671 34919 6683 35039
rect 6603 34917 6683 34919
rect 6925 35039 7005 35041
rect 6925 34918 6937 35039
rect 6993 34918 7005 35039
rect 6247 34909 6303 34917
rect 6615 34909 6671 34917
rect 6925 34916 7005 34918
rect 6937 34908 6993 34916
rect 6431 34741 6487 34749
rect 6799 34741 6855 34749
rect 6419 34739 6908 34741
rect 6419 34619 6431 34739
rect 6487 34619 6799 34739
rect 6855 34619 6908 34739
rect 6419 34617 6908 34619
rect 6431 34609 6487 34617
rect 6799 34609 6908 34617
rect 6327 34543 6407 34553
rect 6327 34487 6339 34543
rect 6395 34487 6407 34543
rect 6327 34477 6407 34487
rect 6511 34543 6591 34553
rect 6511 34487 6523 34543
rect 6579 34487 6591 34543
rect 6511 34477 6591 34487
rect 6695 34543 6775 34553
rect 6695 34487 6707 34543
rect 6763 34487 6775 34543
rect 6695 34477 6775 34487
rect 6339 34395 6395 34477
rect 6327 34393 6407 34395
rect 6327 34337 6339 34393
rect 6395 34337 6407 34393
rect 6327 34335 6407 34337
rect 5354 34277 5434 34279
rect 5354 34221 5366 34277
rect 5422 34221 5434 34277
rect 5354 34219 5434 34221
rect 5797 34277 5857 34287
rect 5797 34221 5799 34277
rect 5855 34221 5857 34277
rect 5209 34161 5289 34163
rect 5209 34105 5221 34161
rect 5277 34105 5289 34161
rect 5209 34103 5289 34105
rect 5221 34021 5277 34103
rect 4841 34011 4921 34021
rect 4841 33955 4853 34011
rect 4909 33955 4921 34011
rect 4841 33945 4921 33955
rect 5025 34011 5105 34021
rect 5025 33955 5037 34011
rect 5093 33955 5105 34011
rect 5025 33945 5105 33955
rect 5209 34011 5289 34021
rect 5209 33955 5221 34011
rect 5277 33955 5289 34011
rect 5209 33945 5289 33955
rect 5354 33889 5422 34219
rect 5797 34209 5857 34221
rect 5313 33881 5422 33889
rect 5301 33879 5422 33881
rect 5301 33759 5313 33879
rect 5369 33759 5422 33879
rect 5301 33757 5422 33759
rect 5313 33749 5369 33757
rect 4616 33492 5512 33504
rect 4616 33436 4628 33492
rect 4684 33436 5446 33492
rect 5502 33436 5512 33492
rect 4616 33424 5512 33436
rect 5799 33266 5855 34209
rect 6339 34021 6395 34335
rect 6523 34279 6579 34477
rect 6511 34277 6591 34279
rect 6511 34221 6523 34277
rect 6579 34221 6591 34277
rect 6511 34219 6591 34221
rect 6523 34021 6579 34219
rect 6707 34163 6763 34477
rect 6840 34279 6908 34609
rect 6840 34277 6920 34279
rect 6840 34221 6852 34277
rect 6908 34221 6920 34277
rect 6840 34219 6920 34221
rect 7107 34277 7177 34289
rect 13505 34278 13575 34292
rect 7107 34221 7109 34277
rect 7165 34221 7863 34277
rect 6695 34161 6775 34163
rect 6695 34105 6707 34161
rect 6763 34105 6775 34161
rect 6695 34103 6775 34105
rect 6707 34021 6763 34103
rect 6327 34011 6407 34021
rect 6327 33955 6339 34011
rect 6395 33955 6407 34011
rect 6327 33945 6407 33955
rect 6511 34011 6591 34021
rect 6511 33955 6523 34011
rect 6579 33955 6591 34011
rect 6511 33945 6591 33955
rect 6695 34011 6775 34021
rect 6695 33955 6707 34011
rect 6763 33955 6775 34011
rect 6695 33945 6775 33955
rect 6840 33889 6908 34219
rect 7107 34211 7177 34221
rect 6799 33881 6908 33889
rect 6787 33879 6908 33881
rect 6787 33759 6799 33879
rect 6855 33759 6908 33879
rect 6787 33757 6908 33759
rect 6799 33749 6855 33757
rect 6102 33492 6998 33504
rect 6102 33436 6114 33492
rect 6170 33436 6932 33492
rect 6988 33436 6998 33492
rect 6102 33424 6998 33436
rect 7109 33267 7165 34211
rect 7273 33375 7353 33385
rect 7273 33319 7285 33375
rect 7341 33319 7353 33375
rect 7273 33317 7353 33319
rect 5797 33264 5867 33266
rect 5797 33208 5799 33264
rect 5855 33208 5867 33264
rect 5797 33196 5867 33208
rect 7097 33265 7177 33267
rect 7097 33209 7109 33265
rect 7165 33209 7177 33265
rect 7097 33197 7177 33209
rect 4761 33157 5507 33169
rect 4761 33101 5129 33157
rect 5185 33101 5507 33157
rect 4761 33089 5507 33101
rect 4761 32836 4817 33089
rect 5129 32836 5185 33089
rect 5451 32836 5507 33089
rect 6247 33158 6993 33170
rect 6247 33102 6615 33158
rect 6671 33102 6993 33158
rect 6247 33090 6993 33102
rect 6247 32837 6303 33090
rect 6615 32837 6671 33090
rect 6937 32837 6993 33090
rect 4749 32834 4829 32836
rect 4749 32714 4761 32834
rect 4817 32714 4829 32834
rect 4749 32712 4829 32714
rect 5117 32834 5197 32836
rect 5117 32714 5129 32834
rect 5185 32714 5197 32834
rect 5117 32712 5197 32714
rect 5439 32834 5519 32836
rect 5439 32713 5451 32834
rect 5507 32713 5519 32834
rect 6235 32835 6315 32837
rect 6235 32715 6247 32835
rect 6303 32715 6315 32835
rect 6235 32713 6315 32715
rect 6603 32835 6683 32837
rect 6603 32715 6615 32835
rect 6671 32715 6683 32835
rect 6603 32713 6683 32715
rect 6925 32835 7005 32837
rect 6925 32714 6937 32835
rect 6993 32714 7005 32835
rect 4761 32704 4817 32712
rect 5129 32704 5185 32712
rect 5439 32711 5519 32713
rect 5451 32703 5507 32711
rect 6247 32705 6303 32713
rect 6615 32705 6671 32713
rect 6925 32712 7005 32714
rect 6937 32704 6993 32712
rect 4945 32536 5001 32544
rect 5313 32536 5369 32544
rect 6431 32537 6487 32545
rect 6799 32537 6855 32545
rect 4933 32534 5422 32536
rect 4933 32414 4945 32534
rect 5001 32414 5313 32534
rect 5369 32414 5422 32534
rect 4933 32412 5422 32414
rect 6419 32535 6908 32537
rect 6419 32415 6431 32535
rect 6487 32415 6799 32535
rect 6855 32415 6908 32535
rect 6419 32413 6908 32415
rect 4945 32404 5001 32412
rect 5313 32404 5422 32412
rect 6431 32405 6487 32413
rect 6799 32405 6908 32413
rect 4841 32338 4921 32348
rect 4841 32282 4853 32338
rect 4909 32282 4921 32338
rect 4841 32272 4921 32282
rect 5025 32338 5105 32348
rect 5025 32282 5037 32338
rect 5093 32282 5105 32338
rect 5025 32272 5105 32282
rect 5209 32338 5289 32348
rect 5209 32282 5221 32338
rect 5277 32282 5289 32338
rect 5209 32272 5289 32282
rect 4853 32190 4909 32272
rect 4841 32188 4921 32190
rect 4841 32132 4853 32188
rect 4909 32132 4921 32188
rect 4841 32130 4921 32132
rect 4169 31956 4239 31968
rect 4169 31900 4181 31956
rect 4237 31900 4239 31956
rect 4169 31888 4239 31900
rect 4853 31816 4909 32130
rect 5037 32074 5093 32272
rect 5025 32072 5105 32074
rect 5025 32016 5037 32072
rect 5093 32016 5105 32072
rect 5025 32014 5105 32016
rect 5037 31816 5093 32014
rect 5221 31958 5277 32272
rect 5354 32074 5422 32404
rect 6327 32339 6407 32349
rect 6327 32283 6339 32339
rect 6395 32283 6407 32339
rect 6327 32273 6407 32283
rect 6511 32339 6591 32349
rect 6511 32283 6523 32339
rect 6579 32283 6591 32339
rect 6511 32273 6591 32283
rect 6695 32339 6775 32349
rect 6695 32283 6707 32339
rect 6763 32283 6775 32339
rect 6695 32273 6775 32283
rect 6339 32191 6395 32273
rect 6327 32189 6407 32191
rect 6327 32133 6339 32189
rect 6395 32133 6407 32189
rect 6327 32131 6407 32133
rect 5354 32072 5434 32074
rect 5354 32016 5366 32072
rect 5422 32016 5434 32072
rect 5354 32014 5434 32016
rect 5621 32072 5691 32084
rect 5621 32016 5623 32072
rect 5679 32016 5691 32072
rect 5209 31956 5289 31958
rect 5209 31900 5221 31956
rect 5277 31900 5289 31956
rect 5209 31898 5289 31900
rect 5221 31816 5277 31898
rect 4841 31806 4921 31816
rect 4841 31750 4853 31806
rect 4909 31750 4921 31806
rect 4841 31740 4921 31750
rect 5025 31806 5105 31816
rect 5025 31750 5037 31806
rect 5093 31750 5105 31806
rect 5025 31740 5105 31750
rect 5209 31806 5289 31816
rect 5209 31750 5221 31806
rect 5277 31750 5289 31806
rect 5209 31740 5289 31750
rect 5354 31684 5422 32014
rect 5621 32006 5691 32016
rect 5313 31676 5422 31684
rect 5301 31674 5422 31676
rect 5301 31554 5313 31674
rect 5369 31554 5422 31674
rect 5301 31552 5422 31554
rect 5313 31544 5369 31552
rect 4616 31287 5512 31299
rect 4616 31231 4628 31287
rect 4684 31231 5446 31287
rect 5502 31231 5512 31287
rect 4616 31219 5512 31231
rect 5623 31062 5679 32006
rect 6339 31817 6395 32131
rect 6523 32075 6579 32273
rect 6511 32073 6591 32075
rect 6511 32017 6523 32073
rect 6579 32017 6591 32073
rect 6511 32015 6591 32017
rect 6523 31817 6579 32015
rect 6707 31959 6763 32273
rect 6840 32075 6908 32405
rect 7285 32083 7341 33317
rect 6840 32073 6920 32075
rect 6840 32017 6852 32073
rect 6908 32017 6920 32073
rect 6840 32015 6920 32017
rect 7283 32073 7353 32083
rect 7283 32017 7285 32073
rect 7341 32017 7433 32073
rect 6695 31957 6775 31959
rect 6695 31901 6707 31957
rect 6763 31901 6775 31957
rect 6695 31899 6775 31901
rect 6707 31817 6763 31899
rect 6327 31807 6407 31817
rect 6327 31751 6339 31807
rect 6395 31751 6407 31807
rect 6327 31741 6407 31751
rect 6511 31807 6591 31817
rect 6511 31751 6523 31807
rect 6579 31751 6591 31807
rect 6511 31741 6591 31751
rect 6695 31807 6775 31817
rect 6695 31751 6707 31807
rect 6763 31751 6775 31807
rect 6695 31741 6775 31751
rect 6840 31685 6908 32015
rect 7283 32005 7353 32017
rect 6799 31677 6908 31685
rect 6787 31675 6908 31677
rect 6787 31555 6799 31675
rect 6855 31555 6908 31675
rect 6787 31553 6908 31555
rect 6799 31545 6855 31553
rect 6102 31288 6998 31300
rect 6102 31232 6114 31288
rect 6170 31232 6932 31288
rect 6988 31232 6998 31288
rect 6102 31220 6998 31232
rect 5787 31169 5867 31179
rect 5787 31113 5799 31169
rect 5855 31113 5867 31169
rect 5787 31111 5867 31113
rect 5621 31059 5691 31062
rect 5621 31005 5623 31059
rect 5679 31005 5691 31059
rect 5621 30993 5691 31005
rect 4761 30952 5507 30964
rect 4761 30896 5129 30952
rect 5185 30896 5507 30952
rect 4761 30884 5507 30896
rect 4761 30631 4817 30884
rect 5129 30631 5185 30884
rect 5451 30631 5507 30884
rect 4749 30629 4829 30631
rect 4749 30509 4761 30629
rect 4817 30509 4829 30629
rect 4749 30507 4829 30509
rect 5117 30629 5197 30631
rect 5117 30509 5129 30629
rect 5185 30509 5197 30629
rect 5117 30507 5197 30509
rect 5439 30629 5519 30631
rect 5439 30508 5451 30629
rect 5507 30508 5519 30629
rect 4761 30499 4817 30507
rect 5129 30499 5185 30507
rect 5439 30506 5519 30508
rect 5451 30498 5507 30506
rect 4945 30331 5001 30339
rect 5313 30331 5369 30339
rect 4933 30329 5422 30331
rect 4933 30209 4945 30329
rect 5001 30209 5313 30329
rect 5369 30209 5422 30329
rect 4933 30207 5422 30209
rect 4945 30199 5001 30207
rect 5313 30199 5422 30207
rect 4841 30133 4921 30143
rect 4841 30077 4853 30133
rect 4909 30077 4921 30133
rect 4841 30067 4921 30077
rect 5025 30133 5105 30143
rect 5025 30077 5037 30133
rect 5093 30077 5105 30133
rect 5025 30067 5105 30077
rect 5209 30133 5289 30143
rect 5209 30077 5221 30133
rect 5277 30077 5289 30133
rect 5209 30067 5289 30077
rect 4853 29985 4909 30067
rect 4841 29983 4921 29985
rect 4841 29927 4853 29983
rect 4909 29927 4921 29983
rect 4841 29925 4921 29927
rect 4033 29867 4103 29881
rect 4033 29811 4045 29867
rect 4101 29811 4103 29867
rect 4033 29799 4103 29811
rect 3799 29751 3877 29762
rect 3407 29750 3877 29751
rect 3407 29696 3811 29750
rect 3865 29696 3877 29750
rect 3407 29695 3877 29696
rect 1835 29391 3007 29401
rect 1835 29335 1847 29391
rect 1903 29335 2735 29391
rect 2791 29335 3007 29391
rect 1835 29325 3007 29335
rect 3407 29391 3487 29695
rect 3799 29684 3877 29695
rect 3407 29335 3419 29391
rect 3475 29335 3487 29391
rect 3407 29325 3487 29335
rect 1765 29013 3557 29025
rect 1765 28873 1777 29013
rect 3545 28873 3557 29013
rect 3850 28964 3936 28976
rect 4045 28968 4101 29799
rect 4853 29611 4909 29925
rect 5037 29869 5093 30067
rect 5025 29867 5105 29869
rect 5025 29811 5037 29867
rect 5093 29811 5105 29867
rect 5025 29809 5105 29811
rect 5037 29611 5093 29809
rect 5221 29753 5277 30067
rect 5354 29869 5422 30199
rect 5799 29879 5855 31111
rect 7807 31006 7863 34221
rect 13505 34222 13517 34278
rect 13573 34222 13575 34278
rect 13505 34210 13575 34222
rect 13223 33376 13305 33388
rect 13223 33320 13237 33376
rect 13293 33320 13305 33376
rect 13223 33308 13305 33320
rect 8217 31970 8437 31980
rect 8217 31170 8227 31970
rect 8427 31170 8437 31970
rect 12607 31970 12927 31980
rect 9079 31463 10251 31473
rect 9079 31223 9091 31463
rect 9147 31223 10183 31463
rect 10239 31223 10251 31463
rect 9079 31213 10251 31223
rect 8217 31160 8437 31170
rect 9173 31006 9251 31018
rect 7803 30950 9193 31006
rect 9249 30950 9251 31006
rect 7807 30949 7863 30950
rect 9173 30938 9251 30950
rect 10171 30928 10251 31213
rect 10651 31463 10731 31473
rect 10651 31223 10663 31463
rect 10719 31223 10731 31463
rect 10473 30928 10543 30940
rect 10171 30872 10485 30928
rect 10541 30872 10543 30928
rect 9993 30850 10063 30862
rect 7803 30794 10005 30850
rect 10061 30794 10063 30850
rect 5354 29867 5434 29869
rect 5354 29811 5366 29867
rect 5422 29811 5434 29867
rect 5354 29809 5434 29811
rect 5797 29867 5857 29879
rect 5797 29811 5799 29867
rect 5855 29811 5857 29867
rect 5209 29751 5289 29753
rect 5209 29695 5221 29751
rect 5277 29695 5289 29751
rect 5209 29693 5289 29695
rect 5221 29611 5277 29693
rect 4841 29601 4921 29611
rect 4841 29545 4853 29601
rect 4909 29545 4921 29601
rect 4841 29535 4921 29545
rect 5025 29601 5105 29611
rect 5025 29545 5037 29601
rect 5093 29545 5105 29601
rect 5025 29535 5105 29545
rect 5209 29601 5289 29611
rect 5209 29545 5221 29601
rect 5277 29545 5289 29601
rect 5209 29535 5289 29545
rect 5354 29479 5422 29809
rect 5797 29799 5857 29811
rect 7915 29508 7971 30794
rect 9993 30782 10063 30794
rect 9283 30568 9363 30578
rect 9283 30512 9295 30568
rect 9351 30512 9363 30568
rect 9283 30326 9363 30512
rect 9763 30568 9843 30578
rect 9763 30512 9775 30568
rect 9831 30512 9843 30568
rect 9763 30502 9843 30512
rect 9967 30568 10047 30578
rect 9967 30512 9979 30568
rect 10035 30512 10047 30568
rect 9967 30326 10047 30512
rect 10171 30568 10251 30872
rect 10473 30860 10543 30872
rect 10651 30928 10731 31223
rect 12607 31170 12617 31970
rect 12917 31170 12927 31970
rect 12607 31160 12927 31170
rect 11237 30974 13029 30986
rect 10651 30872 11008 30928
rect 10171 30512 10183 30568
rect 10239 30512 10251 30568
rect 10171 30502 10251 30512
rect 10651 30568 10731 30872
rect 10651 30512 10663 30568
rect 10719 30512 10731 30568
rect 10651 30502 10731 30512
rect 9283 30254 10047 30326
rect 10177 30200 10801 30212
rect 10177 30060 10189 30200
rect 10789 30060 10801 30200
rect 8389 30043 8469 30053
rect 10177 30048 10801 30060
rect 8389 29803 8401 30043
rect 8457 29803 8469 30043
rect 10952 29830 11008 30872
rect 11237 30834 11249 30974
rect 13017 30834 13029 30974
rect 11237 30822 13029 30834
rect 11511 30571 12275 30581
rect 11511 30331 11523 30571
rect 11579 30331 12207 30571
rect 12263 30331 12275 30571
rect 11511 30321 12275 30331
rect 12879 30287 12959 30297
rect 11991 30237 12479 30247
rect 11991 29997 12003 30237
rect 12059 29997 12411 30237
rect 12467 29997 12479 30237
rect 11991 29987 12479 29997
rect 11401 29830 11497 29842
rect 8211 29508 8281 29520
rect 5313 29471 5422 29479
rect 5301 29469 5422 29471
rect 5301 29349 5313 29469
rect 5369 29349 5422 29469
rect 7403 29452 8223 29508
rect 8279 29452 8281 29508
rect 5301 29347 5422 29349
rect 5313 29339 5369 29347
rect 4616 29082 5514 29094
rect 4616 29026 4628 29082
rect 4684 29026 5446 29082
rect 5502 29026 5514 29082
rect 4616 29014 5514 29026
rect 3850 28908 3862 28964
rect 3918 28908 3936 28964
rect 3850 28896 3936 28908
rect 4043 28964 4103 28968
rect 4043 28908 4045 28964
rect 4101 28908 4103 28964
rect 4043 28896 4103 28908
rect 1765 28861 3557 28873
rect 1179 28531 1536 28587
rect 3135 28689 3455 28699
rect 699 28171 711 28227
rect 767 28171 779 28227
rect 699 28161 779 28171
rect 1179 28227 1259 28531
rect 1179 28171 1191 28227
rect 1247 28171 1259 28227
rect 1179 28161 1259 28171
rect -189 27913 575 27985
rect 3135 27889 3145 28689
rect 3445 27889 3455 28689
rect 3135 27879 3455 27889
rect 7408 27609 7464 29452
rect 8211 29440 8281 29452
rect 8389 29508 8469 29803
rect 10177 29800 10801 29812
rect 10177 29660 10189 29800
rect 10789 29660 10801 29800
rect 10952 29774 11421 29830
rect 11477 29774 11497 29830
rect 11401 29762 11497 29774
rect 12399 29752 12479 29987
rect 12879 30047 12891 30287
rect 12947 30047 12959 30287
rect 12701 29752 12771 29764
rect 12399 29696 12713 29752
rect 12769 29696 12771 29752
rect 12085 29674 12181 29684
rect 10177 29648 10801 29660
rect 10952 29618 12105 29674
rect 12161 29618 12181 29674
rect 8389 29452 8827 29508
rect 8389 29148 8469 29452
rect 8389 29092 8401 29148
rect 8457 29092 8469 29148
rect 8389 29082 8469 29092
rect 8771 28666 8827 29452
rect 9079 29123 10251 29133
rect 9079 28883 9091 29123
rect 9147 28883 10183 29123
rect 10239 28883 10251 29123
rect 9079 28873 10251 28883
rect 9173 28666 9251 28678
rect 8771 28610 9193 28666
rect 9249 28610 9251 28666
rect 9173 28598 9251 28610
rect 10171 28588 10251 28873
rect 10651 29123 10731 29133
rect 10651 28883 10663 29123
rect 10719 28883 10731 29123
rect 10473 28588 10543 28600
rect 10171 28532 10485 28588
rect 10541 28532 10543 28588
rect 9993 28510 10063 28522
rect 7408 27479 7464 27489
rect 7803 28454 10005 28510
rect 10061 28454 10063 28510
rect 7803 27345 7859 28454
rect 9993 28442 10063 28454
rect 9283 28228 9363 28238
rect 9283 28172 9295 28228
rect 9351 28172 9363 28228
rect 9283 27986 9363 28172
rect 9763 28228 9843 28238
rect 9763 28172 9775 28228
rect 9831 28172 9843 28228
rect 9763 28162 9843 28172
rect 9967 28228 10047 28238
rect 9967 28172 9979 28228
rect 10035 28172 10047 28228
rect 9967 27986 10047 28172
rect 10171 28228 10251 28532
rect 10473 28520 10543 28532
rect 10651 28588 10731 28883
rect 10952 28588 11008 29618
rect 12085 29608 12181 29618
rect 12399 29402 12479 29696
rect 12701 29684 12771 29696
rect 12879 29752 12959 30047
rect 13517 29882 13573 34210
rect 13653 31969 13709 36415
rect 14325 36227 14381 36541
rect 14509 36485 14565 36683
rect 14497 36483 14577 36485
rect 14497 36427 14509 36483
rect 14565 36427 14577 36483
rect 14497 36425 14577 36427
rect 14509 36227 14565 36425
rect 14693 36369 14749 36683
rect 14826 36485 14894 36815
rect 23785 36749 23865 36759
rect 23785 36693 23797 36749
rect 23853 36693 23865 36749
rect 23785 36683 23865 36693
rect 23969 36749 24049 36759
rect 23969 36693 23981 36749
rect 24037 36693 24049 36749
rect 23969 36683 24049 36693
rect 24153 36749 24233 36759
rect 24153 36693 24165 36749
rect 24221 36693 24233 36749
rect 24153 36683 24233 36693
rect 22895 36599 22983 36611
rect 23797 36601 23853 36683
rect 22895 36543 22909 36599
rect 22965 36543 22983 36599
rect 22895 36531 22983 36543
rect 23785 36599 23865 36601
rect 23785 36543 23797 36599
rect 23853 36543 23865 36599
rect 23785 36541 23865 36543
rect 14826 36483 14906 36485
rect 14826 36427 14838 36483
rect 14894 36427 14906 36483
rect 14826 36425 14906 36427
rect 15093 36483 15163 36495
rect 15093 36427 15095 36483
rect 15151 36427 15163 36483
rect 14681 36367 14761 36369
rect 14681 36311 14693 36367
rect 14749 36311 14761 36367
rect 14681 36309 14761 36311
rect 14693 36227 14749 36309
rect 14313 36217 14393 36227
rect 14313 36161 14325 36217
rect 14381 36161 14393 36217
rect 14313 36151 14393 36161
rect 14497 36217 14577 36227
rect 14497 36161 14509 36217
rect 14565 36161 14577 36217
rect 14497 36151 14577 36161
rect 14681 36217 14761 36227
rect 14681 36161 14693 36217
rect 14749 36161 14761 36217
rect 14681 36151 14761 36161
rect 14826 36095 14894 36425
rect 15093 36417 15163 36427
rect 23113 36483 23183 36495
rect 23113 36427 23125 36483
rect 23181 36427 23183 36483
rect 14785 36087 14894 36095
rect 14773 36085 14894 36087
rect 14773 35965 14785 36085
rect 14841 35965 14894 36085
rect 14773 35963 14894 35965
rect 14785 35955 14841 35963
rect 14088 35698 14986 35710
rect 14088 35642 14100 35698
rect 14156 35642 14918 35698
rect 14974 35642 14986 35698
rect 14088 35630 14986 35642
rect 15095 35473 15151 36417
rect 23113 36415 23183 36427
rect 15259 35580 15339 35590
rect 15259 35524 15271 35580
rect 15327 35524 15339 35580
rect 15259 35522 15339 35524
rect 15093 35470 15163 35473
rect 15093 35416 15095 35470
rect 15151 35416 15163 35470
rect 15093 35404 15163 35416
rect 14233 35363 14979 35375
rect 14233 35307 14601 35363
rect 14657 35307 14979 35363
rect 14233 35295 14979 35307
rect 14233 35042 14289 35295
rect 14601 35042 14657 35295
rect 14923 35042 14979 35295
rect 14221 35040 14301 35042
rect 14221 34920 14233 35040
rect 14289 34920 14301 35040
rect 14221 34918 14301 34920
rect 14589 35040 14669 35042
rect 14589 34920 14601 35040
rect 14657 34920 14669 35040
rect 14589 34918 14669 34920
rect 14911 35040 14991 35042
rect 14911 34919 14923 35040
rect 14979 34919 14991 35040
rect 14233 34910 14289 34918
rect 14601 34910 14657 34918
rect 14911 34917 14991 34919
rect 14923 34909 14979 34917
rect 14417 34742 14473 34750
rect 14785 34742 14841 34750
rect 14405 34740 14894 34742
rect 14405 34620 14417 34740
rect 14473 34620 14785 34740
rect 14841 34620 14894 34740
rect 14405 34618 14894 34620
rect 14417 34610 14473 34618
rect 14785 34610 14894 34618
rect 14313 34544 14393 34554
rect 14313 34488 14325 34544
rect 14381 34488 14393 34544
rect 14313 34478 14393 34488
rect 14497 34544 14577 34554
rect 14497 34488 14509 34544
rect 14565 34488 14577 34544
rect 14497 34478 14577 34488
rect 14681 34544 14761 34554
rect 14681 34488 14693 34544
rect 14749 34488 14761 34544
rect 14681 34478 14761 34488
rect 14325 34396 14381 34478
rect 14313 34394 14393 34396
rect 14313 34338 14325 34394
rect 14381 34338 14393 34394
rect 14313 34336 14393 34338
rect 14325 34022 14381 34336
rect 14509 34280 14565 34478
rect 14497 34278 14577 34280
rect 14497 34222 14509 34278
rect 14565 34222 14577 34278
rect 14497 34220 14577 34222
rect 14509 34022 14565 34220
rect 14693 34164 14749 34478
rect 14826 34280 14894 34610
rect 15271 34288 15327 35522
rect 15719 35363 16465 35375
rect 15719 35307 16087 35363
rect 16143 35307 16465 35363
rect 15719 35295 16465 35307
rect 15719 35042 15775 35295
rect 16087 35042 16143 35295
rect 16409 35042 16465 35295
rect 15707 35040 15787 35042
rect 15707 34920 15719 35040
rect 15775 34920 15787 35040
rect 15707 34918 15787 34920
rect 16075 35040 16155 35042
rect 16075 34920 16087 35040
rect 16143 34920 16155 35040
rect 16075 34918 16155 34920
rect 16397 35040 16477 35042
rect 16397 34919 16409 35040
rect 16465 34919 16477 35040
rect 15719 34910 15775 34918
rect 16087 34910 16143 34918
rect 16397 34917 16477 34919
rect 16409 34909 16465 34917
rect 15903 34742 15959 34750
rect 16271 34742 16327 34750
rect 15891 34740 16380 34742
rect 15891 34620 15903 34740
rect 15959 34620 16271 34740
rect 16327 34620 16380 34740
rect 15891 34618 16380 34620
rect 15903 34610 15959 34618
rect 16271 34610 16380 34618
rect 15799 34544 15879 34554
rect 15799 34488 15811 34544
rect 15867 34488 15879 34544
rect 15799 34478 15879 34488
rect 15983 34544 16063 34554
rect 15983 34488 15995 34544
rect 16051 34488 16063 34544
rect 15983 34478 16063 34488
rect 16167 34544 16247 34554
rect 16167 34488 16179 34544
rect 16235 34488 16247 34544
rect 16167 34478 16247 34488
rect 15811 34396 15867 34478
rect 15799 34394 15879 34396
rect 15799 34338 15811 34394
rect 15867 34338 15879 34394
rect 15799 34336 15879 34338
rect 14826 34278 14906 34280
rect 14826 34222 14838 34278
rect 14894 34222 14906 34278
rect 14826 34220 14906 34222
rect 15269 34278 15329 34288
rect 15269 34222 15271 34278
rect 15327 34222 15329 34278
rect 14681 34162 14761 34164
rect 14681 34106 14693 34162
rect 14749 34106 14761 34162
rect 14681 34104 14761 34106
rect 14693 34022 14749 34104
rect 14313 34012 14393 34022
rect 14313 33956 14325 34012
rect 14381 33956 14393 34012
rect 14313 33946 14393 33956
rect 14497 34012 14577 34022
rect 14497 33956 14509 34012
rect 14565 33956 14577 34012
rect 14497 33946 14577 33956
rect 14681 34012 14761 34022
rect 14681 33956 14693 34012
rect 14749 33956 14761 34012
rect 14681 33946 14761 33956
rect 14826 33890 14894 34220
rect 15269 34210 15329 34222
rect 14785 33882 14894 33890
rect 14773 33880 14894 33882
rect 14773 33760 14785 33880
rect 14841 33760 14894 33880
rect 14773 33758 14894 33760
rect 14785 33750 14841 33758
rect 14088 33493 14984 33505
rect 14088 33437 14100 33493
rect 14156 33437 14918 33493
rect 14974 33437 14984 33493
rect 14088 33425 14984 33437
rect 15271 33267 15327 34210
rect 15811 34022 15867 34336
rect 15995 34280 16051 34478
rect 15983 34278 16063 34280
rect 15983 34222 15995 34278
rect 16051 34222 16063 34278
rect 15983 34220 16063 34222
rect 15995 34022 16051 34220
rect 16179 34164 16235 34478
rect 16312 34280 16380 34610
rect 16312 34278 16392 34280
rect 16312 34222 16324 34278
rect 16380 34222 16392 34278
rect 16312 34220 16392 34222
rect 16579 34278 16649 34290
rect 22977 34278 23047 34292
rect 16579 34222 16581 34278
rect 16637 34222 17335 34278
rect 16167 34162 16247 34164
rect 16167 34106 16179 34162
rect 16235 34106 16247 34162
rect 16167 34104 16247 34106
rect 16179 34022 16235 34104
rect 15799 34012 15879 34022
rect 15799 33956 15811 34012
rect 15867 33956 15879 34012
rect 15799 33946 15879 33956
rect 15983 34012 16063 34022
rect 15983 33956 15995 34012
rect 16051 33956 16063 34012
rect 15983 33946 16063 33956
rect 16167 34012 16247 34022
rect 16167 33956 16179 34012
rect 16235 33956 16247 34012
rect 16167 33946 16247 33956
rect 16312 33890 16380 34220
rect 16579 34212 16649 34222
rect 16271 33882 16380 33890
rect 16259 33880 16380 33882
rect 16259 33760 16271 33880
rect 16327 33760 16380 33880
rect 16259 33758 16380 33760
rect 16271 33750 16327 33758
rect 15574 33493 16470 33505
rect 15574 33437 15586 33493
rect 15642 33437 16404 33493
rect 16460 33437 16470 33493
rect 15574 33425 16470 33437
rect 16581 33268 16637 34212
rect 16745 33376 16825 33386
rect 16745 33320 16757 33376
rect 16813 33320 16825 33376
rect 16745 33318 16825 33320
rect 15269 33265 15339 33267
rect 15269 33209 15271 33265
rect 15327 33209 15339 33265
rect 15269 33197 15339 33209
rect 16569 33266 16649 33268
rect 16569 33210 16581 33266
rect 16637 33210 16649 33266
rect 16569 33198 16649 33210
rect 14233 33158 14979 33170
rect 14233 33102 14601 33158
rect 14657 33102 14979 33158
rect 14233 33090 14979 33102
rect 14233 32837 14289 33090
rect 14601 32837 14657 33090
rect 14923 32837 14979 33090
rect 15719 33159 16465 33171
rect 15719 33103 16087 33159
rect 16143 33103 16465 33159
rect 15719 33091 16465 33103
rect 15719 32838 15775 33091
rect 16087 32838 16143 33091
rect 16409 32838 16465 33091
rect 14221 32835 14301 32837
rect 14221 32715 14233 32835
rect 14289 32715 14301 32835
rect 14221 32713 14301 32715
rect 14589 32835 14669 32837
rect 14589 32715 14601 32835
rect 14657 32715 14669 32835
rect 14589 32713 14669 32715
rect 14911 32835 14991 32837
rect 14911 32714 14923 32835
rect 14979 32714 14991 32835
rect 15707 32836 15787 32838
rect 15707 32716 15719 32836
rect 15775 32716 15787 32836
rect 15707 32714 15787 32716
rect 16075 32836 16155 32838
rect 16075 32716 16087 32836
rect 16143 32716 16155 32836
rect 16075 32714 16155 32716
rect 16397 32836 16477 32838
rect 16397 32715 16409 32836
rect 16465 32715 16477 32836
rect 14233 32705 14289 32713
rect 14601 32705 14657 32713
rect 14911 32712 14991 32714
rect 14923 32704 14979 32712
rect 15719 32706 15775 32714
rect 16087 32706 16143 32714
rect 16397 32713 16477 32715
rect 16409 32705 16465 32713
rect 14417 32537 14473 32545
rect 14785 32537 14841 32545
rect 15903 32538 15959 32546
rect 16271 32538 16327 32546
rect 14405 32535 14894 32537
rect 14405 32415 14417 32535
rect 14473 32415 14785 32535
rect 14841 32415 14894 32535
rect 14405 32413 14894 32415
rect 15891 32536 16380 32538
rect 15891 32416 15903 32536
rect 15959 32416 16271 32536
rect 16327 32416 16380 32536
rect 15891 32414 16380 32416
rect 14417 32405 14473 32413
rect 14785 32405 14894 32413
rect 15903 32406 15959 32414
rect 16271 32406 16380 32414
rect 14313 32339 14393 32349
rect 14313 32283 14325 32339
rect 14381 32283 14393 32339
rect 14313 32273 14393 32283
rect 14497 32339 14577 32349
rect 14497 32283 14509 32339
rect 14565 32283 14577 32339
rect 14497 32273 14577 32283
rect 14681 32339 14761 32349
rect 14681 32283 14693 32339
rect 14749 32283 14761 32339
rect 14681 32273 14761 32283
rect 14325 32191 14381 32273
rect 14313 32189 14393 32191
rect 14313 32133 14325 32189
rect 14381 32133 14393 32189
rect 14313 32131 14393 32133
rect 13641 31957 13711 31969
rect 13641 31901 13653 31957
rect 13709 31901 13711 31957
rect 13641 31889 13711 31901
rect 14325 31817 14381 32131
rect 14509 32075 14565 32273
rect 14497 32073 14577 32075
rect 14497 32017 14509 32073
rect 14565 32017 14577 32073
rect 14497 32015 14577 32017
rect 14509 31817 14565 32015
rect 14693 31959 14749 32273
rect 14826 32075 14894 32405
rect 15799 32340 15879 32350
rect 15799 32284 15811 32340
rect 15867 32284 15879 32340
rect 15799 32274 15879 32284
rect 15983 32340 16063 32350
rect 15983 32284 15995 32340
rect 16051 32284 16063 32340
rect 15983 32274 16063 32284
rect 16167 32340 16247 32350
rect 16167 32284 16179 32340
rect 16235 32284 16247 32340
rect 16167 32274 16247 32284
rect 15811 32192 15867 32274
rect 15799 32190 15879 32192
rect 15799 32134 15811 32190
rect 15867 32134 15879 32190
rect 15799 32132 15879 32134
rect 14826 32073 14906 32075
rect 14826 32017 14838 32073
rect 14894 32017 14906 32073
rect 14826 32015 14906 32017
rect 15093 32073 15163 32085
rect 15093 32017 15095 32073
rect 15151 32017 15163 32073
rect 14681 31957 14761 31959
rect 14681 31901 14693 31957
rect 14749 31901 14761 31957
rect 14681 31899 14761 31901
rect 14693 31817 14749 31899
rect 14313 31807 14393 31817
rect 14313 31751 14325 31807
rect 14381 31751 14393 31807
rect 14313 31741 14393 31751
rect 14497 31807 14577 31817
rect 14497 31751 14509 31807
rect 14565 31751 14577 31807
rect 14497 31741 14577 31751
rect 14681 31807 14761 31817
rect 14681 31751 14693 31807
rect 14749 31751 14761 31807
rect 14681 31741 14761 31751
rect 14826 31685 14894 32015
rect 15093 32007 15163 32017
rect 14785 31677 14894 31685
rect 14773 31675 14894 31677
rect 14773 31555 14785 31675
rect 14841 31555 14894 31675
rect 14773 31553 14894 31555
rect 14785 31545 14841 31553
rect 14088 31288 14984 31300
rect 14088 31232 14100 31288
rect 14156 31232 14918 31288
rect 14974 31232 14984 31288
rect 14088 31220 14984 31232
rect 15095 31063 15151 32007
rect 15811 31818 15867 32132
rect 15995 32076 16051 32274
rect 15983 32074 16063 32076
rect 15983 32018 15995 32074
rect 16051 32018 16063 32074
rect 15983 32016 16063 32018
rect 15995 31818 16051 32016
rect 16179 31960 16235 32274
rect 16312 32076 16380 32406
rect 16757 32084 16813 33318
rect 16312 32074 16392 32076
rect 16312 32018 16324 32074
rect 16380 32018 16392 32074
rect 16312 32016 16392 32018
rect 16755 32074 16825 32084
rect 16755 32018 16757 32074
rect 16813 32018 16905 32074
rect 16167 31958 16247 31960
rect 16167 31902 16179 31958
rect 16235 31902 16247 31958
rect 16167 31900 16247 31902
rect 16179 31818 16235 31900
rect 15799 31808 15879 31818
rect 15799 31752 15811 31808
rect 15867 31752 15879 31808
rect 15799 31742 15879 31752
rect 15983 31808 16063 31818
rect 15983 31752 15995 31808
rect 16051 31752 16063 31808
rect 15983 31742 16063 31752
rect 16167 31808 16247 31818
rect 16167 31752 16179 31808
rect 16235 31752 16247 31808
rect 16167 31742 16247 31752
rect 16312 31686 16380 32016
rect 16755 32006 16825 32018
rect 16271 31678 16380 31686
rect 16259 31676 16380 31678
rect 16259 31556 16271 31676
rect 16327 31556 16380 31676
rect 16259 31554 16380 31556
rect 16271 31546 16327 31554
rect 15574 31289 16470 31301
rect 15574 31233 15586 31289
rect 15642 31233 16404 31289
rect 16460 31233 16470 31289
rect 15574 31221 16470 31233
rect 15259 31170 15339 31180
rect 15259 31114 15271 31170
rect 15327 31114 15339 31170
rect 15259 31112 15339 31114
rect 15093 31060 15163 31063
rect 15093 31006 15095 31060
rect 15151 31006 15163 31060
rect 15093 30994 15163 31006
rect 14233 30953 14979 30965
rect 14233 30897 14601 30953
rect 14657 30897 14979 30953
rect 14233 30885 14979 30897
rect 14233 30632 14289 30885
rect 14601 30632 14657 30885
rect 14923 30632 14979 30885
rect 14221 30630 14301 30632
rect 14221 30510 14233 30630
rect 14289 30510 14301 30630
rect 14221 30508 14301 30510
rect 14589 30630 14669 30632
rect 14589 30510 14601 30630
rect 14657 30510 14669 30630
rect 14589 30508 14669 30510
rect 14911 30630 14991 30632
rect 14911 30509 14923 30630
rect 14979 30509 14991 30630
rect 14233 30500 14289 30508
rect 14601 30500 14657 30508
rect 14911 30507 14991 30509
rect 14923 30499 14979 30507
rect 14417 30332 14473 30340
rect 14785 30332 14841 30340
rect 14405 30330 14894 30332
rect 14405 30210 14417 30330
rect 14473 30210 14785 30330
rect 14841 30210 14894 30330
rect 14405 30208 14894 30210
rect 14417 30200 14473 30208
rect 14785 30200 14894 30208
rect 14313 30134 14393 30144
rect 14313 30078 14325 30134
rect 14381 30078 14393 30134
rect 14313 30068 14393 30078
rect 14497 30134 14577 30144
rect 14497 30078 14509 30134
rect 14565 30078 14577 30134
rect 14497 30068 14577 30078
rect 14681 30134 14761 30144
rect 14681 30078 14693 30134
rect 14749 30078 14761 30134
rect 14681 30068 14761 30078
rect 14325 29986 14381 30068
rect 14313 29984 14393 29986
rect 14313 29928 14325 29984
rect 14381 29928 14393 29984
rect 14313 29926 14393 29928
rect 13505 29868 13575 29882
rect 13505 29812 13517 29868
rect 13573 29812 13575 29868
rect 13505 29800 13575 29812
rect 13271 29752 13349 29763
rect 12879 29751 13349 29752
rect 12879 29697 13283 29751
rect 13337 29697 13349 29751
rect 12879 29696 13349 29697
rect 11307 29392 12479 29402
rect 11307 29336 11319 29392
rect 11375 29336 12207 29392
rect 12263 29336 12479 29392
rect 11307 29326 12479 29336
rect 12879 29392 12959 29696
rect 13271 29685 13349 29696
rect 12879 29336 12891 29392
rect 12947 29336 12959 29392
rect 12879 29326 12959 29336
rect 11237 29014 13029 29026
rect 11237 28874 11249 29014
rect 13017 28874 13029 29014
rect 13322 28965 13408 28977
rect 13517 28969 13573 29800
rect 14325 29612 14381 29926
rect 14509 29870 14565 30068
rect 14497 29868 14577 29870
rect 14497 29812 14509 29868
rect 14565 29812 14577 29868
rect 14497 29810 14577 29812
rect 14509 29612 14565 29810
rect 14693 29754 14749 30068
rect 14826 29870 14894 30200
rect 15271 29880 15327 31112
rect 17279 31006 17335 34222
rect 22977 34222 22989 34278
rect 23045 34222 23047 34278
rect 22977 34210 23047 34222
rect 22695 33376 22777 33388
rect 22695 33320 22709 33376
rect 22765 33320 22777 33376
rect 22695 33308 22777 33320
rect 17689 31970 17909 31980
rect 17689 31170 17699 31970
rect 17899 31170 17909 31970
rect 22079 31970 22399 31980
rect 18551 31463 19723 31473
rect 18551 31223 18563 31463
rect 18619 31223 19655 31463
rect 19711 31223 19723 31463
rect 18551 31213 19723 31223
rect 17689 31160 17909 31170
rect 18645 31006 18723 31018
rect 17275 30950 18665 31006
rect 18721 30950 18723 31006
rect 18645 30938 18723 30950
rect 19643 30928 19723 31213
rect 20123 31463 20203 31473
rect 20123 31223 20135 31463
rect 20191 31223 20203 31463
rect 19945 30928 20015 30940
rect 19643 30872 19957 30928
rect 20013 30872 20015 30928
rect 19465 30850 19535 30862
rect 17275 30794 19477 30850
rect 19533 30794 19535 30850
rect 14826 29868 14906 29870
rect 14826 29812 14838 29868
rect 14894 29812 14906 29868
rect 14826 29810 14906 29812
rect 15269 29868 15329 29880
rect 15269 29812 15271 29868
rect 15327 29812 15329 29868
rect 14681 29752 14761 29754
rect 14681 29696 14693 29752
rect 14749 29696 14761 29752
rect 14681 29694 14761 29696
rect 14693 29612 14749 29694
rect 14313 29602 14393 29612
rect 14313 29546 14325 29602
rect 14381 29546 14393 29602
rect 14313 29536 14393 29546
rect 14497 29602 14577 29612
rect 14497 29546 14509 29602
rect 14565 29546 14577 29602
rect 14497 29536 14577 29546
rect 14681 29602 14761 29612
rect 14681 29546 14693 29602
rect 14749 29546 14761 29602
rect 14681 29536 14761 29546
rect 14826 29480 14894 29810
rect 15269 29800 15329 29812
rect 17387 29509 17443 30794
rect 19465 30782 19535 30794
rect 18755 30568 18835 30578
rect 18755 30512 18767 30568
rect 18823 30512 18835 30568
rect 18755 30326 18835 30512
rect 19235 30568 19315 30578
rect 19235 30512 19247 30568
rect 19303 30512 19315 30568
rect 19235 30502 19315 30512
rect 19439 30568 19519 30578
rect 19439 30512 19451 30568
rect 19507 30512 19519 30568
rect 19439 30326 19519 30512
rect 19643 30568 19723 30872
rect 19945 30860 20015 30872
rect 20123 30928 20203 31223
rect 22079 31170 22089 31970
rect 22389 31170 22399 31970
rect 22079 31160 22399 31170
rect 20709 30974 22501 30986
rect 20123 30872 20480 30928
rect 19643 30512 19655 30568
rect 19711 30512 19723 30568
rect 19643 30502 19723 30512
rect 20123 30568 20203 30872
rect 20123 30512 20135 30568
rect 20191 30512 20203 30568
rect 20123 30502 20203 30512
rect 18755 30254 19519 30326
rect 19649 30200 20273 30212
rect 19649 30060 19661 30200
rect 20261 30060 20273 30200
rect 17861 30043 17941 30053
rect 19649 30048 20273 30060
rect 17861 29803 17873 30043
rect 17929 29803 17941 30043
rect 20424 29830 20480 30872
rect 20709 30834 20721 30974
rect 22489 30834 22501 30974
rect 20709 30822 22501 30834
rect 20983 30571 21747 30581
rect 20983 30331 20995 30571
rect 21051 30331 21679 30571
rect 21735 30331 21747 30571
rect 20983 30321 21747 30331
rect 22351 30287 22431 30297
rect 21463 30237 21951 30247
rect 21463 29997 21475 30237
rect 21531 29997 21883 30237
rect 21939 29997 21951 30237
rect 21463 29987 21951 29997
rect 20873 29830 20969 29842
rect 14785 29472 14894 29480
rect 14773 29470 14894 29472
rect 14773 29350 14785 29470
rect 14841 29350 14894 29470
rect 16875 29508 17443 29509
rect 17683 29508 17753 29520
rect 16875 29453 17695 29508
rect 14773 29348 14894 29350
rect 14785 29340 14841 29348
rect 14088 29083 14986 29095
rect 14088 29027 14100 29083
rect 14156 29027 14918 29083
rect 14974 29027 14986 29083
rect 14088 29015 14986 29027
rect 13322 28909 13334 28965
rect 13390 28909 13408 28965
rect 13322 28897 13408 28909
rect 13515 28965 13575 28969
rect 13515 28909 13517 28965
rect 13573 28909 13575 28965
rect 13515 28897 13575 28909
rect 11237 28862 13029 28874
rect 10651 28532 11008 28588
rect 12607 28690 12927 28700
rect 10171 28172 10183 28228
rect 10239 28172 10251 28228
rect 10171 28162 10251 28172
rect 10651 28228 10731 28532
rect 10651 28172 10663 28228
rect 10719 28172 10731 28228
rect 10651 28162 10731 28172
rect 9283 27914 10047 27986
rect 12607 27890 12617 28690
rect 12917 27890 12927 28690
rect 12607 27880 12927 27890
rect 16880 27610 16936 29453
rect 17387 29452 17695 29453
rect 17751 29452 17753 29508
rect 17683 29440 17753 29452
rect 17861 29508 17941 29803
rect 19649 29800 20273 29812
rect 19649 29660 19661 29800
rect 20261 29660 20273 29800
rect 20424 29774 20893 29830
rect 20949 29774 20969 29830
rect 20873 29762 20969 29774
rect 21871 29752 21951 29987
rect 22351 30047 22363 30287
rect 22419 30047 22431 30287
rect 22173 29752 22243 29764
rect 21871 29696 22185 29752
rect 22241 29696 22243 29752
rect 21557 29674 21653 29684
rect 19649 29648 20273 29660
rect 20424 29618 21577 29674
rect 21633 29618 21653 29674
rect 17861 29452 18299 29508
rect 17861 29148 17941 29452
rect 17861 29092 17873 29148
rect 17929 29092 17941 29148
rect 17861 29082 17941 29092
rect 18243 28666 18299 29452
rect 18551 29123 19723 29133
rect 18551 28883 18563 29123
rect 18619 28883 19655 29123
rect 19711 28883 19723 29123
rect 18551 28873 19723 28883
rect 18645 28666 18723 28678
rect 18243 28610 18665 28666
rect 18721 28610 18723 28666
rect 18645 28598 18723 28610
rect 19643 28588 19723 28873
rect 20123 29123 20203 29133
rect 20123 28883 20135 29123
rect 20191 28883 20203 29123
rect 19945 28588 20015 28600
rect 19643 28532 19957 28588
rect 20013 28532 20015 28588
rect 19465 28510 19535 28522
rect 16880 27480 16936 27490
rect 17275 28454 19477 28510
rect 19533 28454 19535 28510
rect 3069 27289 7859 27345
rect -1027 26484 -971 26486
rect -1669 26428 -971 26484
rect -8887 25722 -8817 25734
rect -8887 25666 -8875 25722
rect -8819 25666 -8817 25722
rect -8887 25664 -8817 25666
rect -9241 24296 -9171 24308
rect -9241 24240 -9229 24296
rect -9173 24240 -9171 24296
rect -9241 24238 -9171 24240
rect -9513 17449 -9443 17461
rect -9513 17393 -9501 17449
rect -9445 17393 -9443 17449
rect -9513 17381 -9443 17393
rect -13224 16499 -12777 16509
rect -13224 16399 -12833 16499
rect -13224 16389 -12777 16399
rect -9501 16499 -9445 17381
rect -9501 16389 -9445 16399
rect -13233 15989 -12777 15999
rect -13233 15889 -12833 15989
rect -13233 15879 -12777 15889
rect -12833 14729 -12777 15879
rect -11981 15686 -11235 15698
rect -11981 15630 -11613 15686
rect -11557 15630 -11235 15686
rect -11981 15618 -11235 15630
rect -11981 15365 -11925 15618
rect -11613 15365 -11557 15618
rect -11291 15365 -11235 15618
rect -11993 15363 -11913 15365
rect -11993 15243 -11981 15363
rect -11925 15243 -11913 15363
rect -11993 15241 -11913 15243
rect -11625 15363 -11545 15365
rect -11625 15243 -11613 15363
rect -11557 15243 -11545 15363
rect -11625 15241 -11545 15243
rect -11303 15363 -11223 15365
rect -11303 15242 -11291 15363
rect -11235 15242 -11223 15363
rect -11981 15233 -11925 15241
rect -11613 15233 -11557 15241
rect -11303 15240 -11223 15242
rect -11291 15232 -11235 15240
rect -11797 15065 -11741 15073
rect -11429 15065 -11373 15073
rect -11809 15063 -11320 15065
rect -11809 14943 -11797 15063
rect -11741 14943 -11429 15063
rect -11373 14943 -11320 15063
rect -11809 14941 -11320 14943
rect -11797 14933 -11741 14941
rect -11429 14933 -11320 14941
rect -11901 14867 -11821 14877
rect -11901 14811 -11889 14867
rect -11833 14811 -11821 14867
rect -11901 14801 -11821 14811
rect -11717 14867 -11637 14877
rect -11717 14811 -11705 14867
rect -11649 14811 -11637 14867
rect -11717 14801 -11637 14811
rect -11533 14867 -11453 14877
rect -11533 14811 -11521 14867
rect -11465 14811 -11453 14867
rect -11533 14801 -11453 14811
rect -12845 14717 -12775 14729
rect -11889 14719 -11833 14801
rect -12845 14661 -12833 14717
rect -12777 14661 -12775 14717
rect -12845 14649 -12775 14661
rect -11901 14717 -11821 14719
rect -11901 14661 -11889 14717
rect -11833 14661 -11821 14717
rect -11901 14659 -11821 14661
rect -12573 14601 -12503 14613
rect -12573 14545 -12561 14601
rect -12505 14545 -12503 14601
rect -12573 14533 -12503 14545
rect -12709 12396 -12639 12410
rect -12709 12340 -12697 12396
rect -12641 12340 -12639 12396
rect -12709 12328 -12639 12340
rect -13117 11494 -13047 11506
rect -13117 11438 -13105 11494
rect -13049 11438 -13047 11494
rect -13117 11426 -13047 11438
rect -13105 6930 -13049 11426
rect -12697 8000 -12641 12328
rect -12561 10087 -12505 14533
rect -11889 14345 -11833 14659
rect -11705 14603 -11649 14801
rect -11717 14601 -11637 14603
rect -11717 14545 -11705 14601
rect -11649 14545 -11637 14601
rect -11717 14543 -11637 14545
rect -11705 14345 -11649 14543
rect -11521 14487 -11465 14801
rect -11388 14603 -11320 14933
rect -11388 14601 -11308 14603
rect -11388 14545 -11376 14601
rect -11320 14545 -11308 14601
rect -11388 14543 -11308 14545
rect -11121 14601 -11051 14613
rect -11121 14545 -11119 14601
rect -11063 14545 -11051 14601
rect -11533 14485 -11453 14487
rect -11533 14429 -11521 14485
rect -11465 14429 -11453 14485
rect -11533 14427 -11453 14429
rect -11521 14345 -11465 14427
rect -11901 14335 -11821 14345
rect -11901 14279 -11889 14335
rect -11833 14279 -11821 14335
rect -11901 14269 -11821 14279
rect -11717 14335 -11637 14345
rect -11717 14279 -11705 14335
rect -11649 14279 -11637 14335
rect -11717 14269 -11637 14279
rect -11533 14335 -11453 14345
rect -11533 14279 -11521 14335
rect -11465 14279 -11453 14335
rect -11533 14269 -11453 14279
rect -11388 14213 -11320 14543
rect -11121 14535 -11051 14545
rect -11429 14205 -11320 14213
rect -11441 14203 -11320 14205
rect -11441 14083 -11429 14203
rect -11373 14083 -11320 14203
rect -11441 14081 -11320 14083
rect -11429 14073 -11373 14081
rect -12126 13816 -11228 13828
rect -12126 13760 -12114 13816
rect -12058 13760 -11296 13816
rect -11240 13760 -11228 13816
rect -12126 13748 -11228 13760
rect -11119 13591 -11063 14535
rect -10955 13698 -10875 13708
rect -10955 13642 -10943 13698
rect -10887 13642 -10875 13698
rect -10955 13640 -10875 13642
rect -11121 13588 -11051 13591
rect -11121 13534 -11119 13588
rect -11063 13534 -11051 13588
rect -11121 13522 -11051 13534
rect -11981 13481 -11235 13493
rect -11981 13425 -11613 13481
rect -11557 13425 -11235 13481
rect -11981 13413 -11235 13425
rect -11981 13160 -11925 13413
rect -11613 13160 -11557 13413
rect -11291 13160 -11235 13413
rect -11993 13158 -11913 13160
rect -11993 13038 -11981 13158
rect -11925 13038 -11913 13158
rect -11993 13036 -11913 13038
rect -11625 13158 -11545 13160
rect -11625 13038 -11613 13158
rect -11557 13038 -11545 13158
rect -11625 13036 -11545 13038
rect -11303 13158 -11223 13160
rect -11303 13037 -11291 13158
rect -11235 13037 -11223 13158
rect -11981 13028 -11925 13036
rect -11613 13028 -11557 13036
rect -11303 13035 -11223 13037
rect -11291 13027 -11235 13035
rect -11797 12860 -11741 12868
rect -11429 12860 -11373 12868
rect -11809 12858 -11320 12860
rect -11809 12738 -11797 12858
rect -11741 12738 -11429 12858
rect -11373 12738 -11320 12858
rect -11809 12736 -11320 12738
rect -11797 12728 -11741 12736
rect -11429 12728 -11320 12736
rect -11901 12662 -11821 12672
rect -11901 12606 -11889 12662
rect -11833 12606 -11821 12662
rect -11901 12596 -11821 12606
rect -11717 12662 -11637 12672
rect -11717 12606 -11705 12662
rect -11649 12606 -11637 12662
rect -11717 12596 -11637 12606
rect -11533 12662 -11453 12672
rect -11533 12606 -11521 12662
rect -11465 12606 -11453 12662
rect -11533 12596 -11453 12606
rect -11889 12514 -11833 12596
rect -11901 12512 -11821 12514
rect -11901 12456 -11889 12512
rect -11833 12456 -11821 12512
rect -11901 12454 -11821 12456
rect -11889 12140 -11833 12454
rect -11705 12398 -11649 12596
rect -11717 12396 -11637 12398
rect -11717 12340 -11705 12396
rect -11649 12340 -11637 12396
rect -11717 12338 -11637 12340
rect -11705 12140 -11649 12338
rect -11521 12282 -11465 12596
rect -11388 12398 -11320 12728
rect -10943 12406 -10887 13640
rect -10495 13481 -9749 13493
rect -10495 13425 -10127 13481
rect -10071 13425 -9749 13481
rect -10495 13413 -9749 13425
rect -10495 13160 -10439 13413
rect -10127 13160 -10071 13413
rect -9805 13160 -9749 13413
rect -10507 13158 -10427 13160
rect -10507 13038 -10495 13158
rect -10439 13038 -10427 13158
rect -10507 13036 -10427 13038
rect -10139 13158 -10059 13160
rect -10139 13038 -10127 13158
rect -10071 13038 -10059 13158
rect -10139 13036 -10059 13038
rect -9817 13158 -9737 13160
rect -9817 13037 -9805 13158
rect -9749 13037 -9737 13158
rect -10495 13028 -10439 13036
rect -10127 13028 -10071 13036
rect -9817 13035 -9737 13037
rect -9805 13027 -9749 13035
rect -10311 12860 -10255 12868
rect -9943 12860 -9887 12868
rect -10323 12858 -9834 12860
rect -10323 12738 -10311 12858
rect -10255 12738 -9943 12858
rect -9887 12738 -9834 12858
rect -10323 12736 -9834 12738
rect -10311 12728 -10255 12736
rect -9943 12728 -9834 12736
rect -10415 12662 -10335 12672
rect -10415 12606 -10403 12662
rect -10347 12606 -10335 12662
rect -10415 12596 -10335 12606
rect -10231 12662 -10151 12672
rect -10231 12606 -10219 12662
rect -10163 12606 -10151 12662
rect -10231 12596 -10151 12606
rect -10047 12662 -9967 12672
rect -10047 12606 -10035 12662
rect -9979 12606 -9967 12662
rect -10047 12596 -9967 12606
rect -10403 12514 -10347 12596
rect -10415 12512 -10335 12514
rect -10415 12456 -10403 12512
rect -10347 12456 -10335 12512
rect -10415 12454 -10335 12456
rect -11388 12396 -11308 12398
rect -11388 12340 -11376 12396
rect -11320 12340 -11308 12396
rect -11388 12338 -11308 12340
rect -10945 12396 -10885 12406
rect -10945 12340 -10943 12396
rect -10887 12340 -10885 12396
rect -11533 12280 -11453 12282
rect -11533 12224 -11521 12280
rect -11465 12224 -11453 12280
rect -11533 12222 -11453 12224
rect -11521 12140 -11465 12222
rect -11901 12130 -11821 12140
rect -11901 12074 -11889 12130
rect -11833 12074 -11821 12130
rect -11901 12064 -11821 12074
rect -11717 12130 -11637 12140
rect -11717 12074 -11705 12130
rect -11649 12074 -11637 12130
rect -11717 12064 -11637 12074
rect -11533 12130 -11453 12140
rect -11533 12074 -11521 12130
rect -11465 12074 -11453 12130
rect -11533 12064 -11453 12074
rect -11388 12008 -11320 12338
rect -10945 12328 -10885 12340
rect -11429 12000 -11320 12008
rect -11441 11998 -11320 12000
rect -11441 11878 -11429 11998
rect -11373 11878 -11320 11998
rect -11441 11876 -11320 11878
rect -11429 11868 -11373 11876
rect -12126 11611 -11230 11623
rect -12126 11555 -12114 11611
rect -12058 11555 -11296 11611
rect -11240 11555 -11230 11611
rect -12126 11543 -11230 11555
rect -10943 11385 -10887 12328
rect -10403 12140 -10347 12454
rect -10219 12398 -10163 12596
rect -10231 12396 -10151 12398
rect -10231 12340 -10219 12396
rect -10163 12340 -10151 12396
rect -10231 12338 -10151 12340
rect -10219 12140 -10163 12338
rect -10035 12282 -9979 12596
rect -9902 12398 -9834 12728
rect -9902 12396 -9822 12398
rect -9902 12340 -9890 12396
rect -9834 12340 -9822 12396
rect -9902 12338 -9822 12340
rect -9635 12396 -9565 12408
rect -9635 12340 -9633 12396
rect -9577 12340 -9309 12396
rect -10047 12280 -9967 12282
rect -10047 12224 -10035 12280
rect -9979 12224 -9967 12280
rect -10047 12222 -9967 12224
rect -10035 12140 -9979 12222
rect -10415 12130 -10335 12140
rect -10415 12074 -10403 12130
rect -10347 12074 -10335 12130
rect -10415 12064 -10335 12074
rect -10231 12130 -10151 12140
rect -10231 12074 -10219 12130
rect -10163 12074 -10151 12130
rect -10231 12064 -10151 12074
rect -10047 12130 -9967 12140
rect -10047 12074 -10035 12130
rect -9979 12074 -9967 12130
rect -10047 12064 -9967 12074
rect -9902 12008 -9834 12338
rect -9635 12330 -9565 12340
rect -9943 12000 -9834 12008
rect -9955 11998 -9834 12000
rect -9955 11878 -9943 11998
rect -9887 11878 -9834 11998
rect -9955 11876 -9834 11878
rect -9943 11868 -9887 11876
rect -10640 11611 -9744 11623
rect -10640 11555 -10628 11611
rect -10572 11555 -9810 11611
rect -9754 11555 -9744 11611
rect -10640 11543 -9744 11555
rect -9633 11386 -9577 12330
rect -9469 11494 -9389 11504
rect -9469 11438 -9457 11494
rect -9401 11438 -9389 11494
rect -9469 11436 -9389 11438
rect -10945 11383 -10875 11385
rect -10945 11327 -10943 11383
rect -10887 11327 -10875 11383
rect -10945 11315 -10875 11327
rect -9645 11384 -9565 11386
rect -9645 11328 -9633 11384
rect -9577 11328 -9565 11384
rect -9645 11316 -9565 11328
rect -11981 11276 -11235 11288
rect -11981 11220 -11613 11276
rect -11557 11220 -11235 11276
rect -11981 11208 -11235 11220
rect -11981 10955 -11925 11208
rect -11613 10955 -11557 11208
rect -11291 10955 -11235 11208
rect -10495 11277 -9749 11289
rect -10495 11221 -10127 11277
rect -10071 11221 -9749 11277
rect -10495 11209 -9749 11221
rect -10495 10956 -10439 11209
rect -10127 10956 -10071 11209
rect -9805 10956 -9749 11209
rect -11993 10953 -11913 10955
rect -11993 10833 -11981 10953
rect -11925 10833 -11913 10953
rect -11993 10831 -11913 10833
rect -11625 10953 -11545 10955
rect -11625 10833 -11613 10953
rect -11557 10833 -11545 10953
rect -11625 10831 -11545 10833
rect -11303 10953 -11223 10955
rect -11303 10832 -11291 10953
rect -11235 10832 -11223 10953
rect -10507 10954 -10427 10956
rect -10507 10834 -10495 10954
rect -10439 10834 -10427 10954
rect -10507 10832 -10427 10834
rect -10139 10954 -10059 10956
rect -10139 10834 -10127 10954
rect -10071 10834 -10059 10954
rect -10139 10832 -10059 10834
rect -9817 10954 -9737 10956
rect -9817 10833 -9805 10954
rect -9749 10833 -9737 10954
rect -11981 10823 -11925 10831
rect -11613 10823 -11557 10831
rect -11303 10830 -11223 10832
rect -11291 10822 -11235 10830
rect -10495 10824 -10439 10832
rect -10127 10824 -10071 10832
rect -9817 10831 -9737 10833
rect -9805 10823 -9749 10831
rect -11797 10655 -11741 10663
rect -11429 10655 -11373 10663
rect -10311 10656 -10255 10664
rect -9943 10656 -9887 10664
rect -11809 10653 -11320 10655
rect -11809 10533 -11797 10653
rect -11741 10533 -11429 10653
rect -11373 10533 -11320 10653
rect -11809 10531 -11320 10533
rect -10323 10654 -9834 10656
rect -10323 10534 -10311 10654
rect -10255 10534 -9943 10654
rect -9887 10534 -9834 10654
rect -10323 10532 -9834 10534
rect -11797 10523 -11741 10531
rect -11429 10523 -11320 10531
rect -10311 10524 -10255 10532
rect -9943 10524 -9834 10532
rect -11901 10457 -11821 10467
rect -11901 10401 -11889 10457
rect -11833 10401 -11821 10457
rect -11901 10391 -11821 10401
rect -11717 10457 -11637 10467
rect -11717 10401 -11705 10457
rect -11649 10401 -11637 10457
rect -11717 10391 -11637 10401
rect -11533 10457 -11453 10467
rect -11533 10401 -11521 10457
rect -11465 10401 -11453 10457
rect -11533 10391 -11453 10401
rect -11889 10309 -11833 10391
rect -11901 10307 -11821 10309
rect -11901 10251 -11889 10307
rect -11833 10251 -11821 10307
rect -11901 10249 -11821 10251
rect -12573 10075 -12503 10087
rect -12573 10019 -12561 10075
rect -12505 10019 -12503 10075
rect -12573 10007 -12503 10019
rect -11889 9935 -11833 10249
rect -11705 10193 -11649 10391
rect -11717 10191 -11637 10193
rect -11717 10135 -11705 10191
rect -11649 10135 -11637 10191
rect -11717 10133 -11637 10135
rect -11705 9935 -11649 10133
rect -11521 10077 -11465 10391
rect -11388 10193 -11320 10523
rect -10415 10458 -10335 10468
rect -10415 10402 -10403 10458
rect -10347 10402 -10335 10458
rect -10415 10392 -10335 10402
rect -10231 10458 -10151 10468
rect -10231 10402 -10219 10458
rect -10163 10402 -10151 10458
rect -10231 10392 -10151 10402
rect -10047 10458 -9967 10468
rect -10047 10402 -10035 10458
rect -9979 10402 -9967 10458
rect -10047 10392 -9967 10402
rect -10403 10310 -10347 10392
rect -10415 10308 -10335 10310
rect -10415 10252 -10403 10308
rect -10347 10252 -10335 10308
rect -10415 10250 -10335 10252
rect -11388 10191 -11308 10193
rect -11388 10135 -11376 10191
rect -11320 10135 -11308 10191
rect -11388 10133 -11308 10135
rect -11121 10191 -11051 10203
rect -11121 10135 -11119 10191
rect -11063 10135 -11051 10191
rect -11533 10075 -11453 10077
rect -11533 10019 -11521 10075
rect -11465 10019 -11453 10075
rect -11533 10017 -11453 10019
rect -11521 9935 -11465 10017
rect -11901 9925 -11821 9935
rect -11901 9869 -11889 9925
rect -11833 9869 -11821 9925
rect -11901 9859 -11821 9869
rect -11717 9925 -11637 9935
rect -11717 9869 -11705 9925
rect -11649 9869 -11637 9925
rect -11717 9859 -11637 9869
rect -11533 9925 -11453 9935
rect -11533 9869 -11521 9925
rect -11465 9869 -11453 9925
rect -11533 9859 -11453 9869
rect -11388 9803 -11320 10133
rect -11121 10125 -11051 10135
rect -11429 9795 -11320 9803
rect -11441 9793 -11320 9795
rect -11441 9673 -11429 9793
rect -11373 9673 -11320 9793
rect -11441 9671 -11320 9673
rect -11429 9663 -11373 9671
rect -12126 9406 -11230 9418
rect -12126 9350 -12114 9406
rect -12058 9350 -11296 9406
rect -11240 9350 -11230 9406
rect -12126 9338 -11230 9350
rect -11119 9181 -11063 10125
rect -10403 9936 -10347 10250
rect -10219 10194 -10163 10392
rect -10231 10192 -10151 10194
rect -10231 10136 -10219 10192
rect -10163 10136 -10151 10192
rect -10231 10134 -10151 10136
rect -10219 9936 -10163 10134
rect -10035 10078 -9979 10392
rect -9902 10194 -9834 10524
rect -9457 10202 -9401 11436
rect -9902 10192 -9822 10194
rect -9902 10136 -9890 10192
rect -9834 10136 -9822 10192
rect -9902 10134 -9822 10136
rect -9459 10192 -9389 10202
rect -9229 10192 -9173 24238
rect -8875 21075 -8819 25664
rect -7969 25265 -7223 25277
rect -7969 25209 -7601 25265
rect -7545 25209 -7223 25265
rect -7969 25197 -7223 25209
rect -7969 24944 -7913 25197
rect -7601 24944 -7545 25197
rect -7279 24944 -7223 25197
rect -7981 24942 -7901 24944
rect -7981 24822 -7969 24942
rect -7913 24822 -7901 24942
rect -7981 24820 -7901 24822
rect -7613 24942 -7533 24944
rect -7613 24822 -7601 24942
rect -7545 24822 -7533 24942
rect -7613 24820 -7533 24822
rect -7291 24942 -7211 24944
rect -7291 24821 -7279 24942
rect -7223 24821 -7211 24942
rect -7969 24812 -7913 24820
rect -7601 24812 -7545 24820
rect -7291 24819 -7211 24821
rect -7279 24811 -7223 24819
rect -7785 24644 -7729 24652
rect -7417 24644 -7361 24652
rect -7797 24642 -7308 24644
rect -7797 24522 -7785 24642
rect -7729 24522 -7417 24642
rect -7361 24522 -7308 24642
rect -7797 24520 -7308 24522
rect -7785 24512 -7729 24520
rect -7417 24512 -7308 24520
rect -7889 24446 -7809 24456
rect -7889 24390 -7877 24446
rect -7821 24390 -7809 24446
rect -7889 24380 -7809 24390
rect -7705 24446 -7625 24456
rect -7705 24390 -7693 24446
rect -7637 24390 -7625 24446
rect -7705 24380 -7625 24390
rect -7521 24446 -7441 24456
rect -7521 24390 -7509 24446
rect -7453 24390 -7441 24446
rect -7521 24380 -7441 24390
rect -7877 24298 -7821 24380
rect -7889 24296 -7809 24298
rect -7889 24240 -7877 24296
rect -7821 24240 -7809 24296
rect -7889 24238 -7809 24240
rect -8561 24180 -8491 24192
rect -8561 24124 -8549 24180
rect -8493 24124 -8491 24180
rect -8561 24112 -8491 24124
rect -8697 21975 -8627 21989
rect -8697 21919 -8685 21975
rect -8629 21919 -8627 21975
rect -8697 21907 -8627 21919
rect -8887 21073 -8817 21075
rect -8887 21017 -8875 21073
rect -8819 21017 -8817 21073
rect -8887 21005 -8817 21017
rect -8685 17579 -8629 21907
rect -8549 19666 -8493 24112
rect -7877 23924 -7821 24238
rect -7693 24182 -7637 24380
rect -7705 24180 -7625 24182
rect -7705 24124 -7693 24180
rect -7637 24124 -7625 24180
rect -7705 24122 -7625 24124
rect -7693 23924 -7637 24122
rect -7509 24066 -7453 24380
rect -7376 24182 -7308 24512
rect -5229 24293 -5159 24305
rect -5229 24237 -5217 24293
rect -5161 24237 -5159 24293
rect -5229 24235 -5159 24237
rect -7376 24180 -7296 24182
rect -7376 24124 -7364 24180
rect -7308 24124 -7296 24180
rect -7376 24122 -7296 24124
rect -7109 24180 -7039 24192
rect -7109 24124 -7107 24180
rect -7051 24124 -7039 24180
rect -7521 24064 -7441 24066
rect -7521 24008 -7509 24064
rect -7453 24008 -7441 24064
rect -7521 24006 -7441 24008
rect -7509 23924 -7453 24006
rect -7889 23914 -7809 23924
rect -7889 23858 -7877 23914
rect -7821 23858 -7809 23914
rect -7889 23848 -7809 23858
rect -7705 23914 -7625 23924
rect -7705 23858 -7693 23914
rect -7637 23858 -7625 23914
rect -7705 23848 -7625 23858
rect -7521 23914 -7441 23924
rect -7521 23858 -7509 23914
rect -7453 23858 -7441 23914
rect -7521 23848 -7441 23858
rect -7376 23792 -7308 24122
rect -7109 24114 -7039 24124
rect -7417 23784 -7308 23792
rect -7429 23782 -7308 23784
rect -7429 23662 -7417 23782
rect -7361 23662 -7308 23782
rect -7429 23660 -7308 23662
rect -7417 23652 -7361 23660
rect -8114 23395 -7216 23407
rect -8114 23339 -8102 23395
rect -8046 23339 -7284 23395
rect -7228 23339 -7216 23395
rect -8114 23327 -7216 23339
rect -7107 23170 -7051 24114
rect -6943 23277 -6863 23287
rect -6943 23221 -6931 23277
rect -6875 23221 -6863 23277
rect -6943 23219 -6863 23221
rect -7109 23167 -7039 23170
rect -7109 23113 -7107 23167
rect -7051 23113 -7039 23167
rect -7109 23101 -7039 23113
rect -7969 23060 -7223 23072
rect -7969 23004 -7601 23060
rect -7545 23004 -7223 23060
rect -7969 22992 -7223 23004
rect -7969 22739 -7913 22992
rect -7601 22739 -7545 22992
rect -7279 22739 -7223 22992
rect -7981 22737 -7901 22739
rect -7981 22617 -7969 22737
rect -7913 22617 -7901 22737
rect -7981 22615 -7901 22617
rect -7613 22737 -7533 22739
rect -7613 22617 -7601 22737
rect -7545 22617 -7533 22737
rect -7613 22615 -7533 22617
rect -7291 22737 -7211 22739
rect -7291 22616 -7279 22737
rect -7223 22616 -7211 22737
rect -7969 22607 -7913 22615
rect -7601 22607 -7545 22615
rect -7291 22614 -7211 22616
rect -7279 22606 -7223 22614
rect -7785 22439 -7729 22447
rect -7417 22439 -7361 22447
rect -7797 22437 -7308 22439
rect -7797 22317 -7785 22437
rect -7729 22317 -7417 22437
rect -7361 22317 -7308 22437
rect -7797 22315 -7308 22317
rect -7785 22307 -7729 22315
rect -7417 22307 -7308 22315
rect -7889 22241 -7809 22251
rect -7889 22185 -7877 22241
rect -7821 22185 -7809 22241
rect -7889 22175 -7809 22185
rect -7705 22241 -7625 22251
rect -7705 22185 -7693 22241
rect -7637 22185 -7625 22241
rect -7705 22175 -7625 22185
rect -7521 22241 -7441 22251
rect -7521 22185 -7509 22241
rect -7453 22185 -7441 22241
rect -7521 22175 -7441 22185
rect -7877 22093 -7821 22175
rect -7889 22091 -7809 22093
rect -7889 22035 -7877 22091
rect -7821 22035 -7809 22091
rect -7889 22033 -7809 22035
rect -7877 21719 -7821 22033
rect -7693 21977 -7637 22175
rect -7705 21975 -7625 21977
rect -7705 21919 -7693 21975
rect -7637 21919 -7625 21975
rect -7705 21917 -7625 21919
rect -7693 21719 -7637 21917
rect -7509 21861 -7453 22175
rect -7376 21977 -7308 22307
rect -6931 21985 -6875 23219
rect -6483 23060 -5737 23072
rect -6483 23004 -6115 23060
rect -6059 23004 -5737 23060
rect -6483 22992 -5737 23004
rect -6483 22739 -6427 22992
rect -6115 22739 -6059 22992
rect -5793 22739 -5737 22992
rect -6495 22737 -6415 22739
rect -6495 22617 -6483 22737
rect -6427 22617 -6415 22737
rect -6495 22615 -6415 22617
rect -6127 22737 -6047 22739
rect -6127 22617 -6115 22737
rect -6059 22617 -6047 22737
rect -6127 22615 -6047 22617
rect -5805 22737 -5725 22739
rect -5805 22616 -5793 22737
rect -5737 22616 -5725 22737
rect -6483 22607 -6427 22615
rect -6115 22607 -6059 22615
rect -5805 22614 -5725 22616
rect -5793 22606 -5737 22614
rect -6299 22439 -6243 22447
rect -5931 22439 -5875 22447
rect -6311 22437 -5822 22439
rect -6311 22317 -6299 22437
rect -6243 22317 -5931 22437
rect -5875 22317 -5822 22437
rect -6311 22315 -5822 22317
rect -6299 22307 -6243 22315
rect -5931 22307 -5822 22315
rect -6403 22241 -6323 22251
rect -6403 22185 -6391 22241
rect -6335 22185 -6323 22241
rect -6403 22175 -6323 22185
rect -6219 22241 -6139 22251
rect -6219 22185 -6207 22241
rect -6151 22185 -6139 22241
rect -6219 22175 -6139 22185
rect -6035 22241 -5955 22251
rect -6035 22185 -6023 22241
rect -5967 22185 -5955 22241
rect -6035 22175 -5955 22185
rect -6391 22093 -6335 22175
rect -6403 22091 -6323 22093
rect -6403 22035 -6391 22091
rect -6335 22035 -6323 22091
rect -6403 22033 -6323 22035
rect -7376 21975 -7296 21977
rect -7376 21919 -7364 21975
rect -7308 21919 -7296 21975
rect -7376 21917 -7296 21919
rect -6933 21975 -6873 21985
rect -6933 21919 -6931 21975
rect -6875 21919 -6873 21975
rect -7521 21859 -7441 21861
rect -7521 21803 -7509 21859
rect -7453 21803 -7441 21859
rect -7521 21801 -7441 21803
rect -7509 21719 -7453 21801
rect -7889 21709 -7809 21719
rect -7889 21653 -7877 21709
rect -7821 21653 -7809 21709
rect -7889 21643 -7809 21653
rect -7705 21709 -7625 21719
rect -7705 21653 -7693 21709
rect -7637 21653 -7625 21709
rect -7705 21643 -7625 21653
rect -7521 21709 -7441 21719
rect -7521 21653 -7509 21709
rect -7453 21653 -7441 21709
rect -7521 21643 -7441 21653
rect -7376 21587 -7308 21917
rect -6933 21907 -6873 21919
rect -7417 21579 -7308 21587
rect -7429 21577 -7308 21579
rect -7429 21457 -7417 21577
rect -7361 21457 -7308 21577
rect -7429 21455 -7308 21457
rect -7417 21447 -7361 21455
rect -8114 21190 -7218 21202
rect -8114 21134 -8102 21190
rect -8046 21134 -7284 21190
rect -7228 21134 -7218 21190
rect -8114 21122 -7218 21134
rect -6931 20964 -6875 21907
rect -6391 21719 -6335 22033
rect -6207 21977 -6151 22175
rect -6219 21975 -6139 21977
rect -6219 21919 -6207 21975
rect -6151 21919 -6139 21975
rect -6219 21917 -6139 21919
rect -6207 21719 -6151 21917
rect -6023 21861 -5967 22175
rect -5890 21977 -5822 22307
rect -5890 21975 -5810 21977
rect -5890 21919 -5878 21975
rect -5822 21919 -5810 21975
rect -5890 21917 -5810 21919
rect -5623 21975 -5553 21987
rect -5623 21919 -5621 21975
rect -5565 21919 -5297 21975
rect -6035 21859 -5955 21861
rect -6035 21803 -6023 21859
rect -5967 21803 -5955 21859
rect -6035 21801 -5955 21803
rect -6023 21719 -5967 21801
rect -6403 21709 -6323 21719
rect -6403 21653 -6391 21709
rect -6335 21653 -6323 21709
rect -6403 21643 -6323 21653
rect -6219 21709 -6139 21719
rect -6219 21653 -6207 21709
rect -6151 21653 -6139 21709
rect -6219 21643 -6139 21653
rect -6035 21709 -5955 21719
rect -6035 21653 -6023 21709
rect -5967 21653 -5955 21709
rect -6035 21643 -5955 21653
rect -5890 21587 -5822 21917
rect -5623 21909 -5553 21919
rect -5931 21579 -5822 21587
rect -5943 21577 -5822 21579
rect -5943 21457 -5931 21577
rect -5875 21457 -5822 21577
rect -5943 21455 -5822 21457
rect -5931 21447 -5875 21455
rect -6628 21190 -5732 21202
rect -6628 21134 -6616 21190
rect -6560 21134 -5798 21190
rect -5742 21134 -5732 21190
rect -6628 21122 -5732 21134
rect -5621 20965 -5565 21909
rect -5457 21073 -5377 21083
rect -5457 21017 -5445 21073
rect -5389 21017 -5377 21073
rect -5457 21015 -5377 21017
rect -6933 20962 -6863 20964
rect -6933 20906 -6931 20962
rect -6875 20906 -6863 20962
rect -6933 20894 -6863 20906
rect -5633 20963 -5553 20965
rect -5633 20907 -5621 20963
rect -5565 20907 -5553 20963
rect -5633 20895 -5553 20907
rect -7969 20855 -7223 20867
rect -7969 20799 -7601 20855
rect -7545 20799 -7223 20855
rect -7969 20787 -7223 20799
rect -7969 20534 -7913 20787
rect -7601 20534 -7545 20787
rect -7279 20534 -7223 20787
rect -6483 20856 -5737 20868
rect -6483 20800 -6115 20856
rect -6059 20800 -5737 20856
rect -6483 20788 -5737 20800
rect -6483 20535 -6427 20788
rect -6115 20535 -6059 20788
rect -5793 20535 -5737 20788
rect -7981 20532 -7901 20534
rect -7981 20412 -7969 20532
rect -7913 20412 -7901 20532
rect -7981 20410 -7901 20412
rect -7613 20532 -7533 20534
rect -7613 20412 -7601 20532
rect -7545 20412 -7533 20532
rect -7613 20410 -7533 20412
rect -7291 20532 -7211 20534
rect -7291 20411 -7279 20532
rect -7223 20411 -7211 20532
rect -6495 20533 -6415 20535
rect -6495 20413 -6483 20533
rect -6427 20413 -6415 20533
rect -6495 20411 -6415 20413
rect -6127 20533 -6047 20535
rect -6127 20413 -6115 20533
rect -6059 20413 -6047 20533
rect -6127 20411 -6047 20413
rect -5805 20533 -5725 20535
rect -5805 20412 -5793 20533
rect -5737 20412 -5725 20533
rect -7969 20402 -7913 20410
rect -7601 20402 -7545 20410
rect -7291 20409 -7211 20411
rect -7279 20401 -7223 20409
rect -6483 20403 -6427 20411
rect -6115 20403 -6059 20411
rect -5805 20410 -5725 20412
rect -5793 20402 -5737 20410
rect -7785 20234 -7729 20242
rect -7417 20234 -7361 20242
rect -6299 20235 -6243 20243
rect -5931 20235 -5875 20243
rect -7797 20232 -7308 20234
rect -7797 20112 -7785 20232
rect -7729 20112 -7417 20232
rect -7361 20112 -7308 20232
rect -7797 20110 -7308 20112
rect -6311 20233 -5822 20235
rect -6311 20113 -6299 20233
rect -6243 20113 -5931 20233
rect -5875 20113 -5822 20233
rect -6311 20111 -5822 20113
rect -7785 20102 -7729 20110
rect -7417 20102 -7308 20110
rect -6299 20103 -6243 20111
rect -5931 20103 -5822 20111
rect -7889 20036 -7809 20046
rect -7889 19980 -7877 20036
rect -7821 19980 -7809 20036
rect -7889 19970 -7809 19980
rect -7705 20036 -7625 20046
rect -7705 19980 -7693 20036
rect -7637 19980 -7625 20036
rect -7705 19970 -7625 19980
rect -7521 20036 -7441 20046
rect -7521 19980 -7509 20036
rect -7453 19980 -7441 20036
rect -7521 19970 -7441 19980
rect -7877 19888 -7821 19970
rect -7889 19886 -7809 19888
rect -7889 19830 -7877 19886
rect -7821 19830 -7809 19886
rect -7889 19828 -7809 19830
rect -8561 19654 -8491 19666
rect -8561 19598 -8549 19654
rect -8493 19598 -8491 19654
rect -8561 19586 -8491 19598
rect -7877 19514 -7821 19828
rect -7693 19772 -7637 19970
rect -7705 19770 -7625 19772
rect -7705 19714 -7693 19770
rect -7637 19714 -7625 19770
rect -7705 19712 -7625 19714
rect -7693 19514 -7637 19712
rect -7509 19656 -7453 19970
rect -7376 19772 -7308 20102
rect -6403 20037 -6323 20047
rect -6403 19981 -6391 20037
rect -6335 19981 -6323 20037
rect -6403 19971 -6323 19981
rect -6219 20037 -6139 20047
rect -6219 19981 -6207 20037
rect -6151 19981 -6139 20037
rect -6219 19971 -6139 19981
rect -6035 20037 -5955 20047
rect -6035 19981 -6023 20037
rect -5967 19981 -5955 20037
rect -6035 19971 -5955 19981
rect -6391 19889 -6335 19971
rect -6403 19887 -6323 19889
rect -6403 19831 -6391 19887
rect -6335 19831 -6323 19887
rect -6403 19829 -6323 19831
rect -7376 19770 -7296 19772
rect -7376 19714 -7364 19770
rect -7308 19714 -7296 19770
rect -7376 19712 -7296 19714
rect -7109 19770 -7039 19782
rect -7109 19714 -7107 19770
rect -7051 19714 -7039 19770
rect -7521 19654 -7441 19656
rect -7521 19598 -7509 19654
rect -7453 19598 -7441 19654
rect -7521 19596 -7441 19598
rect -7509 19514 -7453 19596
rect -7889 19504 -7809 19514
rect -7889 19448 -7877 19504
rect -7821 19448 -7809 19504
rect -7889 19438 -7809 19448
rect -7705 19504 -7625 19514
rect -7705 19448 -7693 19504
rect -7637 19448 -7625 19504
rect -7705 19438 -7625 19448
rect -7521 19504 -7441 19514
rect -7521 19448 -7509 19504
rect -7453 19448 -7441 19504
rect -7521 19438 -7441 19448
rect -7376 19382 -7308 19712
rect -7109 19704 -7039 19714
rect -7417 19374 -7308 19382
rect -7429 19372 -7308 19374
rect -7429 19252 -7417 19372
rect -7361 19252 -7308 19372
rect -7429 19250 -7308 19252
rect -7417 19242 -7361 19250
rect -8114 18985 -7218 18997
rect -8114 18929 -8102 18985
rect -8046 18929 -7284 18985
rect -7228 18929 -7218 18985
rect -8114 18917 -7218 18929
rect -7107 18760 -7051 19704
rect -6391 19515 -6335 19829
rect -6207 19773 -6151 19971
rect -6219 19771 -6139 19773
rect -6219 19715 -6207 19771
rect -6151 19715 -6139 19771
rect -6219 19713 -6139 19715
rect -6207 19515 -6151 19713
rect -6023 19657 -5967 19971
rect -5890 19773 -5822 20103
rect -5445 19781 -5389 21015
rect -5890 19771 -5810 19773
rect -5890 19715 -5878 19771
rect -5822 19715 -5810 19771
rect -5890 19713 -5810 19715
rect -5447 19771 -5377 19781
rect -5447 19715 -5445 19771
rect -5389 19715 -5297 19771
rect -6035 19655 -5955 19657
rect -6035 19599 -6023 19655
rect -5967 19599 -5955 19655
rect -6035 19597 -5955 19599
rect -6023 19515 -5967 19597
rect -6403 19505 -6323 19515
rect -6403 19449 -6391 19505
rect -6335 19449 -6323 19505
rect -6403 19439 -6323 19449
rect -6219 19505 -6139 19515
rect -6219 19449 -6207 19505
rect -6151 19449 -6139 19505
rect -6219 19439 -6139 19449
rect -6035 19505 -5955 19515
rect -6035 19449 -6023 19505
rect -5967 19449 -5955 19505
rect -6035 19439 -5955 19449
rect -5890 19383 -5822 19713
rect -5447 19703 -5377 19715
rect -5931 19375 -5822 19383
rect -5943 19373 -5822 19375
rect -5943 19253 -5931 19373
rect -5875 19253 -5822 19373
rect -5943 19251 -5822 19253
rect -5931 19243 -5875 19251
rect -6628 18986 -5732 18998
rect -6628 18930 -6616 18986
rect -6560 18930 -5798 18986
rect -5742 18930 -5732 18986
rect -6628 18918 -5732 18930
rect -6943 18867 -6863 18877
rect -6943 18811 -6931 18867
rect -6875 18811 -6863 18867
rect -6943 18809 -6863 18811
rect -7109 18757 -7039 18760
rect -7109 18703 -7107 18757
rect -7051 18703 -7039 18757
rect -7109 18691 -7039 18703
rect -7969 18650 -7223 18662
rect -7969 18594 -7601 18650
rect -7545 18594 -7223 18650
rect -7969 18582 -7223 18594
rect -7969 18329 -7913 18582
rect -7601 18329 -7545 18582
rect -7279 18329 -7223 18582
rect -7981 18327 -7901 18329
rect -7981 18207 -7969 18327
rect -7913 18207 -7901 18327
rect -7981 18205 -7901 18207
rect -7613 18327 -7533 18329
rect -7613 18207 -7601 18327
rect -7545 18207 -7533 18327
rect -7613 18205 -7533 18207
rect -7291 18327 -7211 18329
rect -7291 18206 -7279 18327
rect -7223 18206 -7211 18327
rect -7969 18197 -7913 18205
rect -7601 18197 -7545 18205
rect -7291 18204 -7211 18206
rect -7279 18196 -7223 18204
rect -7785 18029 -7729 18037
rect -7417 18029 -7361 18037
rect -7797 18027 -7308 18029
rect -7797 17907 -7785 18027
rect -7729 17907 -7417 18027
rect -7361 17907 -7308 18027
rect -7797 17905 -7308 17907
rect -7785 17897 -7729 17905
rect -7417 17897 -7308 17905
rect -7889 17831 -7809 17841
rect -7889 17775 -7877 17831
rect -7821 17775 -7809 17831
rect -7889 17765 -7809 17775
rect -7705 17831 -7625 17841
rect -7705 17775 -7693 17831
rect -7637 17775 -7625 17831
rect -7705 17765 -7625 17775
rect -7521 17831 -7441 17841
rect -7521 17775 -7509 17831
rect -7453 17775 -7441 17831
rect -7521 17765 -7441 17775
rect -7877 17683 -7821 17765
rect -7889 17681 -7809 17683
rect -7889 17625 -7877 17681
rect -7821 17625 -7809 17681
rect -7889 17623 -7809 17625
rect -8697 17565 -8627 17579
rect -8697 17509 -8685 17565
rect -8629 17509 -8627 17565
rect -8697 17497 -8627 17509
rect -8969 16662 -8899 16674
rect -8685 16666 -8629 17497
rect -7877 17309 -7821 17623
rect -7693 17567 -7637 17765
rect -7705 17565 -7625 17567
rect -7705 17509 -7693 17565
rect -7637 17509 -7625 17565
rect -7705 17507 -7625 17509
rect -7693 17309 -7637 17507
rect -7509 17451 -7453 17765
rect -7376 17567 -7308 17897
rect -6931 17577 -6875 18809
rect -7376 17565 -7296 17567
rect -7376 17509 -7364 17565
rect -7308 17509 -7296 17565
rect -7376 17507 -7296 17509
rect -6933 17565 -6873 17577
rect -6933 17509 -6931 17565
rect -6875 17509 -6873 17565
rect -7521 17449 -7441 17451
rect -7521 17393 -7509 17449
rect -7453 17393 -7441 17449
rect -7521 17391 -7441 17393
rect -7509 17309 -7453 17391
rect -7889 17299 -7809 17309
rect -7889 17243 -7877 17299
rect -7821 17243 -7809 17299
rect -7889 17233 -7809 17243
rect -7705 17299 -7625 17309
rect -7705 17243 -7693 17299
rect -7637 17243 -7625 17299
rect -7705 17233 -7625 17243
rect -7521 17299 -7441 17309
rect -7521 17243 -7509 17299
rect -7453 17243 -7441 17299
rect -7521 17233 -7441 17243
rect -7376 17177 -7308 17507
rect -6933 17497 -6873 17509
rect -5501 17446 -5431 17458
rect -5501 17390 -5489 17446
rect -5433 17390 -5431 17446
rect -5501 17378 -5431 17390
rect -7417 17169 -7308 17177
rect -7429 17167 -7308 17169
rect -7429 17047 -7417 17167
rect -7361 17047 -7308 17167
rect -7429 17045 -7308 17047
rect -7417 17037 -7361 17045
rect -8114 16780 -7216 16792
rect -8114 16724 -8102 16780
rect -8046 16724 -7284 16780
rect -7228 16724 -7216 16780
rect -8114 16712 -7216 16724
rect -8969 16606 -8957 16662
rect -8901 16606 -8899 16662
rect -8969 16604 -8899 16606
rect -8687 16662 -8627 16666
rect -8687 16606 -8685 16662
rect -8629 16606 -8627 16662
rect -8957 15992 -8901 16604
rect -8687 16594 -8627 16606
rect -5489 16499 -5433 17378
rect -5489 16389 -5433 16399
rect -9105 11494 -9035 11506
rect -9105 11438 -9093 11494
rect -9037 11438 -9035 11494
rect -9105 11426 -9035 11438
rect -9459 10136 -9457 10192
rect -9401 10136 -9173 10192
rect -10047 10076 -9967 10078
rect -10047 10020 -10035 10076
rect -9979 10020 -9967 10076
rect -10047 10018 -9967 10020
rect -10035 9936 -9979 10018
rect -10415 9926 -10335 9936
rect -10415 9870 -10403 9926
rect -10347 9870 -10335 9926
rect -10415 9860 -10335 9870
rect -10231 9926 -10151 9936
rect -10231 9870 -10219 9926
rect -10163 9870 -10151 9926
rect -10231 9860 -10151 9870
rect -10047 9926 -9967 9936
rect -10047 9870 -10035 9926
rect -9979 9870 -9967 9926
rect -10047 9860 -9967 9870
rect -9902 9804 -9834 10134
rect -9459 10124 -9389 10136
rect -9943 9796 -9834 9804
rect -9955 9794 -9834 9796
rect -9955 9674 -9943 9794
rect -9887 9674 -9834 9794
rect -9955 9672 -9834 9674
rect -9943 9664 -9887 9672
rect -10640 9407 -9744 9419
rect -10640 9351 -10628 9407
rect -10572 9351 -9810 9407
rect -9754 9351 -9744 9407
rect -10640 9339 -9744 9351
rect -10955 9288 -10875 9298
rect -10955 9232 -10943 9288
rect -10887 9232 -10875 9288
rect -10955 9230 -10875 9232
rect -11121 9178 -11051 9181
rect -11121 9124 -11119 9178
rect -11063 9124 -11051 9178
rect -11121 9112 -11051 9124
rect -11981 9071 -11235 9083
rect -11981 9015 -11613 9071
rect -11557 9015 -11235 9071
rect -11981 9003 -11235 9015
rect -11981 8750 -11925 9003
rect -11613 8750 -11557 9003
rect -11291 8750 -11235 9003
rect -11993 8748 -11913 8750
rect -11993 8628 -11981 8748
rect -11925 8628 -11913 8748
rect -11993 8626 -11913 8628
rect -11625 8748 -11545 8750
rect -11625 8628 -11613 8748
rect -11557 8628 -11545 8748
rect -11625 8626 -11545 8628
rect -11303 8748 -11223 8750
rect -11303 8627 -11291 8748
rect -11235 8627 -11223 8748
rect -11981 8618 -11925 8626
rect -11613 8618 -11557 8626
rect -11303 8625 -11223 8627
rect -11291 8617 -11235 8625
rect -11797 8450 -11741 8458
rect -11429 8450 -11373 8458
rect -11809 8448 -11320 8450
rect -11809 8328 -11797 8448
rect -11741 8328 -11429 8448
rect -11373 8328 -11320 8448
rect -11809 8326 -11320 8328
rect -11797 8318 -11741 8326
rect -11429 8318 -11320 8326
rect -11901 8252 -11821 8262
rect -11901 8196 -11889 8252
rect -11833 8196 -11821 8252
rect -11901 8186 -11821 8196
rect -11717 8252 -11637 8262
rect -11717 8196 -11705 8252
rect -11649 8196 -11637 8252
rect -11717 8186 -11637 8196
rect -11533 8252 -11453 8262
rect -11533 8196 -11521 8252
rect -11465 8196 -11453 8252
rect -11533 8186 -11453 8196
rect -11889 8104 -11833 8186
rect -11901 8102 -11821 8104
rect -11901 8046 -11889 8102
rect -11833 8046 -11821 8102
rect -11901 8044 -11821 8046
rect -12709 7986 -12639 8000
rect -12709 7930 -12697 7986
rect -12641 7930 -12639 7986
rect -12709 7918 -12639 7930
rect -12908 7870 -12828 7882
rect -12908 7814 -12896 7870
rect -12840 7814 -12828 7870
rect -12908 7802 -12828 7814
rect -12908 7083 -12822 7095
rect -12697 7087 -12641 7918
rect -11889 7730 -11833 8044
rect -11705 7988 -11649 8186
rect -11717 7986 -11637 7988
rect -11717 7930 -11705 7986
rect -11649 7930 -11637 7986
rect -11717 7928 -11637 7930
rect -11705 7730 -11649 7928
rect -11521 7872 -11465 8186
rect -11388 7988 -11320 8318
rect -10943 7998 -10887 9230
rect -11388 7986 -11308 7988
rect -11388 7930 -11376 7986
rect -11320 7930 -11308 7986
rect -11388 7928 -11308 7930
rect -10945 7986 -10885 7998
rect -10945 7930 -10943 7986
rect -10887 7930 -10885 7986
rect -11533 7870 -11453 7872
rect -11533 7814 -11521 7870
rect -11465 7814 -11453 7870
rect -11533 7812 -11453 7814
rect -11521 7730 -11465 7812
rect -11901 7720 -11821 7730
rect -11901 7664 -11889 7720
rect -11833 7664 -11821 7720
rect -11901 7654 -11821 7664
rect -11717 7720 -11637 7730
rect -11717 7664 -11705 7720
rect -11649 7664 -11637 7720
rect -11717 7654 -11637 7664
rect -11533 7720 -11453 7730
rect -11533 7664 -11521 7720
rect -11465 7664 -11453 7720
rect -11533 7654 -11453 7664
rect -11388 7598 -11320 7928
rect -10945 7918 -10885 7930
rect -11429 7590 -11320 7598
rect -11441 7588 -11320 7590
rect -11441 7468 -11429 7588
rect -11373 7468 -11320 7588
rect -11441 7466 -11320 7468
rect -11429 7458 -11373 7466
rect -12126 7201 -11228 7213
rect -12126 7145 -12114 7201
rect -12058 7145 -11296 7201
rect -11240 7145 -11228 7201
rect -12126 7133 -11228 7145
rect -12908 7027 -12896 7083
rect -12840 7027 -12822 7083
rect -12908 7015 -12822 7027
rect -12699 7083 -12639 7087
rect -12699 7027 -12697 7083
rect -12641 7027 -12639 7083
rect -12699 7015 -12639 7027
rect -13369 6920 -13049 6930
rect -13369 6820 -13105 6920
rect -13369 6810 -13049 6820
rect -9093 6920 -9037 11426
rect -8957 7095 -8901 15892
rect -7969 15686 -7223 15698
rect -7969 15630 -7601 15686
rect -7545 15630 -7223 15686
rect -7969 15618 -7223 15630
rect -7969 15365 -7913 15618
rect -7601 15365 -7545 15618
rect -7279 15365 -7223 15618
rect -7981 15363 -7901 15365
rect -7981 15243 -7969 15363
rect -7913 15243 -7901 15363
rect -7981 15241 -7901 15243
rect -7613 15363 -7533 15365
rect -7613 15243 -7601 15363
rect -7545 15243 -7533 15363
rect -7613 15241 -7533 15243
rect -7291 15363 -7211 15365
rect -7291 15242 -7279 15363
rect -7223 15242 -7211 15363
rect -7969 15233 -7913 15241
rect -7601 15233 -7545 15241
rect -7291 15240 -7211 15242
rect -7279 15232 -7223 15240
rect -7785 15065 -7729 15073
rect -7417 15065 -7361 15073
rect -7797 15063 -7308 15065
rect -7797 14943 -7785 15063
rect -7729 14943 -7417 15063
rect -7361 14943 -7308 15063
rect -7797 14941 -7308 14943
rect -7785 14933 -7729 14941
rect -7417 14933 -7308 14941
rect -7889 14867 -7809 14877
rect -7889 14811 -7877 14867
rect -7821 14811 -7809 14867
rect -7889 14801 -7809 14811
rect -7705 14867 -7625 14877
rect -7705 14811 -7693 14867
rect -7637 14811 -7625 14867
rect -7705 14801 -7625 14811
rect -7521 14867 -7441 14877
rect -7521 14811 -7509 14867
rect -7453 14811 -7441 14867
rect -7521 14801 -7441 14811
rect -8777 14717 -8691 14729
rect -7877 14719 -7821 14801
rect -8777 14661 -8765 14717
rect -8709 14661 -8691 14717
rect -8777 14649 -8691 14661
rect -7889 14717 -7809 14719
rect -7889 14661 -7877 14717
rect -7821 14661 -7809 14717
rect -7889 14659 -7809 14661
rect -8561 14601 -8491 14613
rect -8561 14545 -8549 14601
rect -8493 14545 -8491 14601
rect -8561 14533 -8491 14545
rect -8697 12396 -8627 12410
rect -8697 12340 -8685 12396
rect -8629 12340 -8627 12396
rect -8697 12328 -8627 12340
rect -8833 12208 -8753 12218
rect -8833 12152 -8821 12208
rect -8765 12152 -8753 12208
rect -8833 12150 -8753 12152
rect -8821 7882 -8765 12150
rect -8685 8000 -8629 12328
rect -8549 10087 -8493 14533
rect -7877 14345 -7821 14659
rect -7693 14603 -7637 14801
rect -7705 14601 -7625 14603
rect -7705 14545 -7693 14601
rect -7637 14545 -7625 14601
rect -7705 14543 -7625 14545
rect -7693 14345 -7637 14543
rect -7509 14487 -7453 14801
rect -7376 14603 -7308 14933
rect -7376 14601 -7296 14603
rect -7376 14545 -7364 14601
rect -7308 14545 -7296 14601
rect -7376 14543 -7296 14545
rect -7109 14601 -7039 14613
rect -7109 14545 -7107 14601
rect -7051 14545 -7039 14601
rect -7521 14485 -7441 14487
rect -7521 14429 -7509 14485
rect -7453 14429 -7441 14485
rect -7521 14427 -7441 14429
rect -7509 14345 -7453 14427
rect -7889 14335 -7809 14345
rect -7889 14279 -7877 14335
rect -7821 14279 -7809 14335
rect -7889 14269 -7809 14279
rect -7705 14335 -7625 14345
rect -7705 14279 -7693 14335
rect -7637 14279 -7625 14335
rect -7705 14269 -7625 14279
rect -7521 14335 -7441 14345
rect -7521 14279 -7509 14335
rect -7453 14279 -7441 14335
rect -7521 14269 -7441 14279
rect -7376 14213 -7308 14543
rect -7109 14535 -7039 14545
rect -7417 14205 -7308 14213
rect -7429 14203 -7308 14205
rect -7429 14083 -7417 14203
rect -7361 14083 -7308 14203
rect -7429 14081 -7308 14083
rect -7417 14073 -7361 14081
rect -8114 13816 -7216 13828
rect -8114 13760 -8102 13816
rect -8046 13760 -7284 13816
rect -7228 13760 -7216 13816
rect -8114 13748 -7216 13760
rect -7107 13591 -7051 14535
rect -6943 13698 -6863 13708
rect -6943 13642 -6931 13698
rect -6875 13642 -6863 13698
rect -6943 13640 -6863 13642
rect -7109 13588 -7039 13591
rect -7109 13534 -7107 13588
rect -7051 13534 -7039 13588
rect -7109 13522 -7039 13534
rect -7969 13481 -7223 13493
rect -7969 13425 -7601 13481
rect -7545 13425 -7223 13481
rect -7969 13413 -7223 13425
rect -7969 13160 -7913 13413
rect -7601 13160 -7545 13413
rect -7279 13160 -7223 13413
rect -7981 13158 -7901 13160
rect -7981 13038 -7969 13158
rect -7913 13038 -7901 13158
rect -7981 13036 -7901 13038
rect -7613 13158 -7533 13160
rect -7613 13038 -7601 13158
rect -7545 13038 -7533 13158
rect -7613 13036 -7533 13038
rect -7291 13158 -7211 13160
rect -7291 13037 -7279 13158
rect -7223 13037 -7211 13158
rect -7969 13028 -7913 13036
rect -7601 13028 -7545 13036
rect -7291 13035 -7211 13037
rect -7279 13027 -7223 13035
rect -7785 12860 -7729 12868
rect -7417 12860 -7361 12868
rect -7797 12858 -7308 12860
rect -7797 12738 -7785 12858
rect -7729 12738 -7417 12858
rect -7361 12738 -7308 12858
rect -7797 12736 -7308 12738
rect -7785 12728 -7729 12736
rect -7417 12728 -7308 12736
rect -7889 12662 -7809 12672
rect -7889 12606 -7877 12662
rect -7821 12606 -7809 12662
rect -7889 12596 -7809 12606
rect -7705 12662 -7625 12672
rect -7705 12606 -7693 12662
rect -7637 12606 -7625 12662
rect -7705 12596 -7625 12606
rect -7521 12662 -7441 12672
rect -7521 12606 -7509 12662
rect -7453 12606 -7441 12662
rect -7521 12596 -7441 12606
rect -7877 12514 -7821 12596
rect -7889 12512 -7809 12514
rect -7889 12456 -7877 12512
rect -7821 12456 -7809 12512
rect -7889 12454 -7809 12456
rect -7877 12140 -7821 12454
rect -7693 12398 -7637 12596
rect -7705 12396 -7625 12398
rect -7705 12340 -7693 12396
rect -7637 12340 -7625 12396
rect -7705 12338 -7625 12340
rect -7693 12140 -7637 12338
rect -7509 12282 -7453 12596
rect -7376 12398 -7308 12728
rect -6931 12406 -6875 13640
rect -6483 13481 -5737 13493
rect -6483 13425 -6115 13481
rect -6059 13425 -5737 13481
rect -6483 13413 -5737 13425
rect -6483 13160 -6427 13413
rect -6115 13160 -6059 13413
rect -5793 13160 -5737 13413
rect -6495 13158 -6415 13160
rect -6495 13038 -6483 13158
rect -6427 13038 -6415 13158
rect -6495 13036 -6415 13038
rect -6127 13158 -6047 13160
rect -6127 13038 -6115 13158
rect -6059 13038 -6047 13158
rect -6127 13036 -6047 13038
rect -5805 13158 -5725 13160
rect -5805 13037 -5793 13158
rect -5737 13037 -5725 13158
rect -6483 13028 -6427 13036
rect -6115 13028 -6059 13036
rect -5805 13035 -5725 13037
rect -5793 13027 -5737 13035
rect -6299 12860 -6243 12868
rect -5931 12860 -5875 12868
rect -6311 12858 -5822 12860
rect -6311 12738 -6299 12858
rect -6243 12738 -5931 12858
rect -5875 12738 -5822 12858
rect -6311 12736 -5822 12738
rect -6299 12728 -6243 12736
rect -5931 12728 -5822 12736
rect -6403 12662 -6323 12672
rect -6403 12606 -6391 12662
rect -6335 12606 -6323 12662
rect -6403 12596 -6323 12606
rect -6219 12662 -6139 12672
rect -6219 12606 -6207 12662
rect -6151 12606 -6139 12662
rect -6219 12596 -6139 12606
rect -6035 12662 -5955 12672
rect -6035 12606 -6023 12662
rect -5967 12606 -5955 12662
rect -6035 12596 -5955 12606
rect -6391 12514 -6335 12596
rect -6403 12512 -6323 12514
rect -6403 12456 -6391 12512
rect -6335 12456 -6323 12512
rect -6403 12454 -6323 12456
rect -7376 12396 -7296 12398
rect -7376 12340 -7364 12396
rect -7308 12340 -7296 12396
rect -7376 12338 -7296 12340
rect -6933 12396 -6873 12406
rect -6933 12340 -6931 12396
rect -6875 12340 -6873 12396
rect -7521 12280 -7441 12282
rect -7521 12224 -7509 12280
rect -7453 12224 -7441 12280
rect -7521 12222 -7441 12224
rect -7509 12140 -7453 12222
rect -7889 12130 -7809 12140
rect -7889 12074 -7877 12130
rect -7821 12074 -7809 12130
rect -7889 12064 -7809 12074
rect -7705 12130 -7625 12140
rect -7705 12074 -7693 12130
rect -7637 12074 -7625 12130
rect -7705 12064 -7625 12074
rect -7521 12130 -7441 12140
rect -7521 12074 -7509 12130
rect -7453 12074 -7441 12130
rect -7521 12064 -7441 12074
rect -7376 12008 -7308 12338
rect -6933 12328 -6873 12340
rect -7417 12000 -7308 12008
rect -7429 11998 -7308 12000
rect -7429 11878 -7417 11998
rect -7361 11878 -7308 11998
rect -7429 11876 -7308 11878
rect -7417 11868 -7361 11876
rect -8114 11611 -7218 11623
rect -8114 11555 -8102 11611
rect -8046 11555 -7284 11611
rect -7228 11555 -7218 11611
rect -8114 11543 -7218 11555
rect -6931 11385 -6875 12328
rect -6391 12140 -6335 12454
rect -6207 12398 -6151 12596
rect -6219 12396 -6139 12398
rect -6219 12340 -6207 12396
rect -6151 12340 -6139 12396
rect -6219 12338 -6139 12340
rect -6207 12140 -6151 12338
rect -6023 12282 -5967 12596
rect -5890 12398 -5822 12728
rect -5890 12396 -5810 12398
rect -5890 12340 -5878 12396
rect -5822 12340 -5810 12396
rect -5890 12338 -5810 12340
rect -5623 12396 -5553 12408
rect -5623 12340 -5621 12396
rect -5565 12340 -5297 12396
rect -6035 12280 -5955 12282
rect -6035 12224 -6023 12280
rect -5967 12224 -5955 12280
rect -6035 12222 -5955 12224
rect -6023 12140 -5967 12222
rect -6403 12130 -6323 12140
rect -6403 12074 -6391 12130
rect -6335 12074 -6323 12130
rect -6403 12064 -6323 12074
rect -6219 12130 -6139 12140
rect -6219 12074 -6207 12130
rect -6151 12074 -6139 12130
rect -6219 12064 -6139 12074
rect -6035 12130 -5955 12140
rect -6035 12074 -6023 12130
rect -5967 12074 -5955 12130
rect -6035 12064 -5955 12074
rect -5890 12008 -5822 12338
rect -5623 12330 -5553 12340
rect -5931 12000 -5822 12008
rect -5943 11998 -5822 12000
rect -5943 11878 -5931 11998
rect -5875 11878 -5822 11998
rect -5943 11876 -5822 11878
rect -5931 11868 -5875 11876
rect -6628 11611 -5732 11623
rect -6628 11555 -6616 11611
rect -6560 11555 -5798 11611
rect -5742 11555 -5732 11611
rect -6628 11543 -5732 11555
rect -5621 11386 -5565 12330
rect -5457 11494 -5377 11504
rect -5457 11438 -5445 11494
rect -5389 11438 -5377 11494
rect -5457 11436 -5377 11438
rect -6933 11383 -6863 11385
rect -6933 11327 -6931 11383
rect -6875 11327 -6863 11383
rect -6933 11315 -6863 11327
rect -5633 11384 -5553 11386
rect -5633 11328 -5621 11384
rect -5565 11328 -5553 11384
rect -5633 11316 -5553 11328
rect -7969 11276 -7223 11288
rect -7969 11220 -7601 11276
rect -7545 11220 -7223 11276
rect -7969 11208 -7223 11220
rect -7969 10955 -7913 11208
rect -7601 10955 -7545 11208
rect -7279 10955 -7223 11208
rect -6483 11277 -5737 11289
rect -6483 11221 -6115 11277
rect -6059 11221 -5737 11277
rect -6483 11209 -5737 11221
rect -6483 10956 -6427 11209
rect -6115 10956 -6059 11209
rect -5793 10956 -5737 11209
rect -7981 10953 -7901 10955
rect -7981 10833 -7969 10953
rect -7913 10833 -7901 10953
rect -7981 10831 -7901 10833
rect -7613 10953 -7533 10955
rect -7613 10833 -7601 10953
rect -7545 10833 -7533 10953
rect -7613 10831 -7533 10833
rect -7291 10953 -7211 10955
rect -7291 10832 -7279 10953
rect -7223 10832 -7211 10953
rect -6495 10954 -6415 10956
rect -6495 10834 -6483 10954
rect -6427 10834 -6415 10954
rect -6495 10832 -6415 10834
rect -6127 10954 -6047 10956
rect -6127 10834 -6115 10954
rect -6059 10834 -6047 10954
rect -6127 10832 -6047 10834
rect -5805 10954 -5725 10956
rect -5805 10833 -5793 10954
rect -5737 10833 -5725 10954
rect -7969 10823 -7913 10831
rect -7601 10823 -7545 10831
rect -7291 10830 -7211 10832
rect -7279 10822 -7223 10830
rect -6483 10824 -6427 10832
rect -6115 10824 -6059 10832
rect -5805 10831 -5725 10833
rect -5793 10823 -5737 10831
rect -7785 10655 -7729 10663
rect -7417 10655 -7361 10663
rect -6299 10656 -6243 10664
rect -5931 10656 -5875 10664
rect -7797 10653 -7308 10655
rect -7797 10533 -7785 10653
rect -7729 10533 -7417 10653
rect -7361 10533 -7308 10653
rect -7797 10531 -7308 10533
rect -6311 10654 -5822 10656
rect -6311 10534 -6299 10654
rect -6243 10534 -5931 10654
rect -5875 10534 -5822 10654
rect -6311 10532 -5822 10534
rect -7785 10523 -7729 10531
rect -7417 10523 -7308 10531
rect -6299 10524 -6243 10532
rect -5931 10524 -5822 10532
rect -7889 10457 -7809 10467
rect -7889 10401 -7877 10457
rect -7821 10401 -7809 10457
rect -7889 10391 -7809 10401
rect -7705 10457 -7625 10467
rect -7705 10401 -7693 10457
rect -7637 10401 -7625 10457
rect -7705 10391 -7625 10401
rect -7521 10457 -7441 10467
rect -7521 10401 -7509 10457
rect -7453 10401 -7441 10457
rect -7521 10391 -7441 10401
rect -7877 10309 -7821 10391
rect -7889 10307 -7809 10309
rect -7889 10251 -7877 10307
rect -7821 10251 -7809 10307
rect -7889 10249 -7809 10251
rect -8561 10075 -8491 10087
rect -8561 10019 -8549 10075
rect -8493 10019 -8491 10075
rect -8561 10007 -8491 10019
rect -7877 9935 -7821 10249
rect -7693 10193 -7637 10391
rect -7705 10191 -7625 10193
rect -7705 10135 -7693 10191
rect -7637 10135 -7625 10191
rect -7705 10133 -7625 10135
rect -7693 9935 -7637 10133
rect -7509 10077 -7453 10391
rect -7376 10193 -7308 10523
rect -6403 10458 -6323 10468
rect -6403 10402 -6391 10458
rect -6335 10402 -6323 10458
rect -6403 10392 -6323 10402
rect -6219 10458 -6139 10468
rect -6219 10402 -6207 10458
rect -6151 10402 -6139 10458
rect -6219 10392 -6139 10402
rect -6035 10458 -5955 10468
rect -6035 10402 -6023 10458
rect -5967 10402 -5955 10458
rect -6035 10392 -5955 10402
rect -6391 10310 -6335 10392
rect -6403 10308 -6323 10310
rect -6403 10252 -6391 10308
rect -6335 10252 -6323 10308
rect -6403 10250 -6323 10252
rect -7376 10191 -7296 10193
rect -7376 10135 -7364 10191
rect -7308 10135 -7296 10191
rect -7376 10133 -7296 10135
rect -7109 10191 -7039 10203
rect -7109 10135 -7107 10191
rect -7051 10135 -7039 10191
rect -7521 10075 -7441 10077
rect -7521 10019 -7509 10075
rect -7453 10019 -7441 10075
rect -7521 10017 -7441 10019
rect -7509 9935 -7453 10017
rect -7889 9925 -7809 9935
rect -7889 9869 -7877 9925
rect -7821 9869 -7809 9925
rect -7889 9859 -7809 9869
rect -7705 9925 -7625 9935
rect -7705 9869 -7693 9925
rect -7637 9869 -7625 9925
rect -7705 9859 -7625 9869
rect -7521 9925 -7441 9935
rect -7521 9869 -7509 9925
rect -7453 9869 -7441 9925
rect -7521 9859 -7441 9869
rect -7376 9803 -7308 10133
rect -7109 10125 -7039 10135
rect -7417 9795 -7308 9803
rect -7429 9793 -7308 9795
rect -7429 9673 -7417 9793
rect -7361 9673 -7308 9793
rect -7429 9671 -7308 9673
rect -7417 9663 -7361 9671
rect -8114 9406 -7218 9418
rect -8114 9350 -8102 9406
rect -8046 9350 -7284 9406
rect -7228 9350 -7218 9406
rect -8114 9338 -7218 9350
rect -7107 9181 -7051 10125
rect -6391 9936 -6335 10250
rect -6207 10194 -6151 10392
rect -6219 10192 -6139 10194
rect -6219 10136 -6207 10192
rect -6151 10136 -6139 10192
rect -6219 10134 -6139 10136
rect -6207 9936 -6151 10134
rect -6023 10078 -5967 10392
rect -5890 10194 -5822 10524
rect -5445 10202 -5389 11436
rect -5890 10192 -5810 10194
rect -5890 10136 -5878 10192
rect -5822 10136 -5810 10192
rect -5890 10134 -5810 10136
rect -5447 10192 -5377 10202
rect -5217 10192 -5161 24235
rect -5081 21977 -5025 26418
rect -1027 25724 -971 26428
rect -749 26074 -679 26086
rect -749 26018 -737 26074
rect -681 26018 -679 26074
rect -749 26016 -679 26018
rect -1029 25722 -959 25724
rect -1029 25666 -1027 25722
rect -971 25666 -959 25722
rect -1029 25664 -959 25666
rect -4791 25546 -4721 25558
rect -4791 25490 -4779 25546
rect -4723 25490 -4721 25546
rect -4791 25488 -4721 25490
rect -5083 21975 -5013 21977
rect -5083 21919 -5081 21975
rect -5025 21919 -5013 21975
rect -5083 21907 -5013 21919
rect -4779 21072 -4723 25488
rect -3927 25262 -3181 25274
rect -3927 25206 -3559 25262
rect -3503 25206 -3181 25262
rect -3927 25194 -3181 25206
rect -3927 24941 -3871 25194
rect -3559 24941 -3503 25194
rect -3237 24941 -3181 25194
rect -3939 24939 -3859 24941
rect -3939 24819 -3927 24939
rect -3871 24819 -3859 24939
rect -3939 24817 -3859 24819
rect -3571 24939 -3491 24941
rect -3571 24819 -3559 24939
rect -3503 24819 -3491 24939
rect -3571 24817 -3491 24819
rect -3249 24939 -3169 24941
rect -3249 24818 -3237 24939
rect -3181 24818 -3169 24939
rect -3927 24809 -3871 24817
rect -3559 24809 -3503 24817
rect -3249 24816 -3169 24818
rect -3237 24808 -3181 24816
rect -3743 24641 -3687 24649
rect -3375 24641 -3319 24649
rect -3755 24639 -3266 24641
rect -3755 24519 -3743 24639
rect -3687 24519 -3375 24639
rect -3319 24519 -3266 24639
rect -3755 24517 -3266 24519
rect -3743 24509 -3687 24517
rect -3375 24509 -3266 24517
rect -3847 24443 -3767 24453
rect -3847 24387 -3835 24443
rect -3779 24387 -3767 24443
rect -3847 24377 -3767 24387
rect -3663 24443 -3583 24453
rect -3663 24387 -3651 24443
rect -3595 24387 -3583 24443
rect -3663 24377 -3583 24387
rect -3479 24443 -3399 24453
rect -3479 24387 -3467 24443
rect -3411 24387 -3399 24443
rect -3479 24377 -3399 24387
rect -3835 24295 -3779 24377
rect -3847 24293 -3767 24295
rect -3847 24237 -3835 24293
rect -3779 24237 -3767 24293
rect -3847 24235 -3767 24237
rect -4519 24177 -4449 24189
rect -4519 24121 -4507 24177
rect -4451 24121 -4449 24177
rect -4519 24109 -4449 24121
rect -4655 21972 -4585 21986
rect -4655 21916 -4643 21972
rect -4587 21916 -4585 21972
rect -4655 21904 -4585 21916
rect -4791 21070 -4721 21072
rect -4791 21014 -4779 21070
rect -4723 21014 -4721 21070
rect -4791 21002 -4721 21014
rect -4643 17576 -4587 21904
rect -4507 19663 -4451 24109
rect -3835 23921 -3779 24235
rect -3651 24179 -3595 24377
rect -3663 24177 -3583 24179
rect -3663 24121 -3651 24177
rect -3595 24121 -3583 24177
rect -3663 24119 -3583 24121
rect -3651 23921 -3595 24119
rect -3467 24063 -3411 24377
rect -3334 24179 -3266 24509
rect -1187 24293 -1117 24305
rect -1187 24237 -1175 24293
rect -1119 24237 -1117 24293
rect -1187 24235 -1117 24237
rect -3334 24177 -3254 24179
rect -3334 24121 -3322 24177
rect -3266 24121 -3254 24177
rect -3334 24119 -3254 24121
rect -3067 24177 -2997 24189
rect -3067 24121 -3065 24177
rect -3009 24121 -2997 24177
rect -3479 24061 -3399 24063
rect -3479 24005 -3467 24061
rect -3411 24005 -3399 24061
rect -3479 24003 -3399 24005
rect -3467 23921 -3411 24003
rect -3847 23911 -3767 23921
rect -3847 23855 -3835 23911
rect -3779 23855 -3767 23911
rect -3847 23845 -3767 23855
rect -3663 23911 -3583 23921
rect -3663 23855 -3651 23911
rect -3595 23855 -3583 23911
rect -3663 23845 -3583 23855
rect -3479 23911 -3399 23921
rect -3479 23855 -3467 23911
rect -3411 23855 -3399 23911
rect -3479 23845 -3399 23855
rect -3334 23789 -3266 24119
rect -3067 24111 -2997 24121
rect -3375 23781 -3266 23789
rect -3387 23779 -3266 23781
rect -3387 23659 -3375 23779
rect -3319 23659 -3266 23779
rect -3387 23657 -3266 23659
rect -3375 23649 -3319 23657
rect -4072 23392 -3174 23404
rect -4072 23336 -4060 23392
rect -4004 23336 -3242 23392
rect -3186 23336 -3174 23392
rect -4072 23324 -3174 23336
rect -3065 23167 -3009 24111
rect -2901 23274 -2821 23284
rect -2901 23218 -2889 23274
rect -2833 23218 -2821 23274
rect -2901 23216 -2821 23218
rect -3067 23164 -2997 23167
rect -3067 23110 -3065 23164
rect -3009 23110 -2997 23164
rect -3067 23098 -2997 23110
rect -3927 23057 -3181 23069
rect -3927 23001 -3559 23057
rect -3503 23001 -3181 23057
rect -3927 22989 -3181 23001
rect -3927 22736 -3871 22989
rect -3559 22736 -3503 22989
rect -3237 22736 -3181 22989
rect -3939 22734 -3859 22736
rect -3939 22614 -3927 22734
rect -3871 22614 -3859 22734
rect -3939 22612 -3859 22614
rect -3571 22734 -3491 22736
rect -3571 22614 -3559 22734
rect -3503 22614 -3491 22734
rect -3571 22612 -3491 22614
rect -3249 22734 -3169 22736
rect -3249 22613 -3237 22734
rect -3181 22613 -3169 22734
rect -3927 22604 -3871 22612
rect -3559 22604 -3503 22612
rect -3249 22611 -3169 22613
rect -3237 22603 -3181 22611
rect -3743 22436 -3687 22444
rect -3375 22436 -3319 22444
rect -3755 22434 -3266 22436
rect -3755 22314 -3743 22434
rect -3687 22314 -3375 22434
rect -3319 22314 -3266 22434
rect -3755 22312 -3266 22314
rect -3743 22304 -3687 22312
rect -3375 22304 -3266 22312
rect -3847 22238 -3767 22248
rect -3847 22182 -3835 22238
rect -3779 22182 -3767 22238
rect -3847 22172 -3767 22182
rect -3663 22238 -3583 22248
rect -3663 22182 -3651 22238
rect -3595 22182 -3583 22238
rect -3663 22172 -3583 22182
rect -3479 22238 -3399 22248
rect -3479 22182 -3467 22238
rect -3411 22182 -3399 22238
rect -3479 22172 -3399 22182
rect -3835 22090 -3779 22172
rect -3847 22088 -3767 22090
rect -3847 22032 -3835 22088
rect -3779 22032 -3767 22088
rect -3847 22030 -3767 22032
rect -3835 21716 -3779 22030
rect -3651 21974 -3595 22172
rect -3663 21972 -3583 21974
rect -3663 21916 -3651 21972
rect -3595 21916 -3583 21972
rect -3663 21914 -3583 21916
rect -3651 21716 -3595 21914
rect -3467 21858 -3411 22172
rect -3334 21974 -3266 22304
rect -2889 21982 -2833 23216
rect -2441 23057 -1695 23069
rect -2441 23001 -2073 23057
rect -2017 23001 -1695 23057
rect -2441 22989 -1695 23001
rect -2441 22736 -2385 22989
rect -2073 22736 -2017 22989
rect -1751 22736 -1695 22989
rect -2453 22734 -2373 22736
rect -2453 22614 -2441 22734
rect -2385 22614 -2373 22734
rect -2453 22612 -2373 22614
rect -2085 22734 -2005 22736
rect -2085 22614 -2073 22734
rect -2017 22614 -2005 22734
rect -2085 22612 -2005 22614
rect -1763 22734 -1683 22736
rect -1763 22613 -1751 22734
rect -1695 22613 -1683 22734
rect -2441 22604 -2385 22612
rect -2073 22604 -2017 22612
rect -1763 22611 -1683 22613
rect -1751 22603 -1695 22611
rect -2257 22436 -2201 22444
rect -1889 22436 -1833 22444
rect -2269 22434 -1780 22436
rect -2269 22314 -2257 22434
rect -2201 22314 -1889 22434
rect -1833 22314 -1780 22434
rect -2269 22312 -1780 22314
rect -2257 22304 -2201 22312
rect -1889 22304 -1780 22312
rect -2361 22238 -2281 22248
rect -2361 22182 -2349 22238
rect -2293 22182 -2281 22238
rect -2361 22172 -2281 22182
rect -2177 22238 -2097 22248
rect -2177 22182 -2165 22238
rect -2109 22182 -2097 22238
rect -2177 22172 -2097 22182
rect -1993 22238 -1913 22248
rect -1993 22182 -1981 22238
rect -1925 22182 -1913 22238
rect -1993 22172 -1913 22182
rect -2349 22090 -2293 22172
rect -2361 22088 -2281 22090
rect -2361 22032 -2349 22088
rect -2293 22032 -2281 22088
rect -2361 22030 -2281 22032
rect -3334 21972 -3254 21974
rect -3334 21916 -3322 21972
rect -3266 21916 -3254 21972
rect -3334 21914 -3254 21916
rect -2891 21972 -2831 21982
rect -2891 21916 -2889 21972
rect -2833 21916 -2831 21972
rect -3479 21856 -3399 21858
rect -3479 21800 -3467 21856
rect -3411 21800 -3399 21856
rect -3479 21798 -3399 21800
rect -3467 21716 -3411 21798
rect -3847 21706 -3767 21716
rect -3847 21650 -3835 21706
rect -3779 21650 -3767 21706
rect -3847 21640 -3767 21650
rect -3663 21706 -3583 21716
rect -3663 21650 -3651 21706
rect -3595 21650 -3583 21706
rect -3663 21640 -3583 21650
rect -3479 21706 -3399 21716
rect -3479 21650 -3467 21706
rect -3411 21650 -3399 21706
rect -3479 21640 -3399 21650
rect -3334 21584 -3266 21914
rect -2891 21904 -2831 21916
rect -3375 21576 -3266 21584
rect -3387 21574 -3266 21576
rect -3387 21454 -3375 21574
rect -3319 21454 -3266 21574
rect -3387 21452 -3266 21454
rect -3375 21444 -3319 21452
rect -4072 21187 -3176 21199
rect -4072 21131 -4060 21187
rect -4004 21131 -3242 21187
rect -3186 21131 -3176 21187
rect -4072 21119 -3176 21131
rect -2889 20961 -2833 21904
rect -2349 21716 -2293 22030
rect -2165 21974 -2109 22172
rect -2177 21972 -2097 21974
rect -2177 21916 -2165 21972
rect -2109 21916 -2097 21972
rect -2177 21914 -2097 21916
rect -2165 21716 -2109 21914
rect -1981 21858 -1925 22172
rect -1848 21974 -1780 22304
rect -1848 21972 -1768 21974
rect -1848 21916 -1836 21972
rect -1780 21916 -1768 21972
rect -1848 21914 -1768 21916
rect -1581 21972 -1511 21984
rect -1581 21916 -1579 21972
rect -1523 21916 -1255 21972
rect -1993 21856 -1913 21858
rect -1993 21800 -1981 21856
rect -1925 21800 -1913 21856
rect -1993 21798 -1913 21800
rect -1981 21716 -1925 21798
rect -2361 21706 -2281 21716
rect -2361 21650 -2349 21706
rect -2293 21650 -2281 21706
rect -2361 21640 -2281 21650
rect -2177 21706 -2097 21716
rect -2177 21650 -2165 21706
rect -2109 21650 -2097 21706
rect -2177 21640 -2097 21650
rect -1993 21706 -1913 21716
rect -1993 21650 -1981 21706
rect -1925 21650 -1913 21706
rect -1993 21640 -1913 21650
rect -1848 21584 -1780 21914
rect -1581 21906 -1511 21916
rect -1889 21576 -1780 21584
rect -1901 21574 -1780 21576
rect -1901 21454 -1889 21574
rect -1833 21454 -1780 21574
rect -1901 21452 -1780 21454
rect -1889 21444 -1833 21452
rect -2586 21187 -1690 21199
rect -2586 21131 -2574 21187
rect -2518 21131 -1756 21187
rect -1700 21131 -1690 21187
rect -2586 21119 -1690 21131
rect -1579 20962 -1523 21906
rect -1415 21070 -1335 21080
rect -1415 21014 -1403 21070
rect -1347 21014 -1335 21070
rect -1415 21012 -1335 21014
rect -2891 20959 -2821 20961
rect -2891 20903 -2889 20959
rect -2833 20903 -2821 20959
rect -2891 20891 -2821 20903
rect -1591 20960 -1511 20962
rect -1591 20904 -1579 20960
rect -1523 20904 -1511 20960
rect -1591 20892 -1511 20904
rect -3927 20852 -3181 20864
rect -3927 20796 -3559 20852
rect -3503 20796 -3181 20852
rect -3927 20784 -3181 20796
rect -3927 20531 -3871 20784
rect -3559 20531 -3503 20784
rect -3237 20531 -3181 20784
rect -2441 20853 -1695 20865
rect -2441 20797 -2073 20853
rect -2017 20797 -1695 20853
rect -2441 20785 -1695 20797
rect -2441 20532 -2385 20785
rect -2073 20532 -2017 20785
rect -1751 20532 -1695 20785
rect -3939 20529 -3859 20531
rect -3939 20409 -3927 20529
rect -3871 20409 -3859 20529
rect -3939 20407 -3859 20409
rect -3571 20529 -3491 20531
rect -3571 20409 -3559 20529
rect -3503 20409 -3491 20529
rect -3571 20407 -3491 20409
rect -3249 20529 -3169 20531
rect -3249 20408 -3237 20529
rect -3181 20408 -3169 20529
rect -2453 20530 -2373 20532
rect -2453 20410 -2441 20530
rect -2385 20410 -2373 20530
rect -2453 20408 -2373 20410
rect -2085 20530 -2005 20532
rect -2085 20410 -2073 20530
rect -2017 20410 -2005 20530
rect -2085 20408 -2005 20410
rect -1763 20530 -1683 20532
rect -1763 20409 -1751 20530
rect -1695 20409 -1683 20530
rect -3927 20399 -3871 20407
rect -3559 20399 -3503 20407
rect -3249 20406 -3169 20408
rect -3237 20398 -3181 20406
rect -2441 20400 -2385 20408
rect -2073 20400 -2017 20408
rect -1763 20407 -1683 20409
rect -1751 20399 -1695 20407
rect -3743 20231 -3687 20239
rect -3375 20231 -3319 20239
rect -2257 20232 -2201 20240
rect -1889 20232 -1833 20240
rect -3755 20229 -3266 20231
rect -3755 20109 -3743 20229
rect -3687 20109 -3375 20229
rect -3319 20109 -3266 20229
rect -3755 20107 -3266 20109
rect -2269 20230 -1780 20232
rect -2269 20110 -2257 20230
rect -2201 20110 -1889 20230
rect -1833 20110 -1780 20230
rect -2269 20108 -1780 20110
rect -3743 20099 -3687 20107
rect -3375 20099 -3266 20107
rect -2257 20100 -2201 20108
rect -1889 20100 -1780 20108
rect -3847 20033 -3767 20043
rect -3847 19977 -3835 20033
rect -3779 19977 -3767 20033
rect -3847 19967 -3767 19977
rect -3663 20033 -3583 20043
rect -3663 19977 -3651 20033
rect -3595 19977 -3583 20033
rect -3663 19967 -3583 19977
rect -3479 20033 -3399 20043
rect -3479 19977 -3467 20033
rect -3411 19977 -3399 20033
rect -3479 19967 -3399 19977
rect -3835 19885 -3779 19967
rect -3847 19883 -3767 19885
rect -3847 19827 -3835 19883
rect -3779 19827 -3767 19883
rect -3847 19825 -3767 19827
rect -4519 19651 -4449 19663
rect -4519 19595 -4507 19651
rect -4451 19595 -4449 19651
rect -4519 19583 -4449 19595
rect -3835 19511 -3779 19825
rect -3651 19769 -3595 19967
rect -3663 19767 -3583 19769
rect -3663 19711 -3651 19767
rect -3595 19711 -3583 19767
rect -3663 19709 -3583 19711
rect -3651 19511 -3595 19709
rect -3467 19653 -3411 19967
rect -3334 19769 -3266 20099
rect -2361 20034 -2281 20044
rect -2361 19978 -2349 20034
rect -2293 19978 -2281 20034
rect -2361 19968 -2281 19978
rect -2177 20034 -2097 20044
rect -2177 19978 -2165 20034
rect -2109 19978 -2097 20034
rect -2177 19968 -2097 19978
rect -1993 20034 -1913 20044
rect -1993 19978 -1981 20034
rect -1925 19978 -1913 20034
rect -1993 19968 -1913 19978
rect -2349 19886 -2293 19968
rect -2361 19884 -2281 19886
rect -2361 19828 -2349 19884
rect -2293 19828 -2281 19884
rect -2361 19826 -2281 19828
rect -3334 19767 -3254 19769
rect -3334 19711 -3322 19767
rect -3266 19711 -3254 19767
rect -3334 19709 -3254 19711
rect -3067 19767 -2997 19779
rect -3067 19711 -3065 19767
rect -3009 19711 -2997 19767
rect -3479 19651 -3399 19653
rect -3479 19595 -3467 19651
rect -3411 19595 -3399 19651
rect -3479 19593 -3399 19595
rect -3467 19511 -3411 19593
rect -3847 19501 -3767 19511
rect -3847 19445 -3835 19501
rect -3779 19445 -3767 19501
rect -3847 19435 -3767 19445
rect -3663 19501 -3583 19511
rect -3663 19445 -3651 19501
rect -3595 19445 -3583 19501
rect -3663 19435 -3583 19445
rect -3479 19501 -3399 19511
rect -3479 19445 -3467 19501
rect -3411 19445 -3399 19501
rect -3479 19435 -3399 19445
rect -3334 19379 -3266 19709
rect -3067 19701 -2997 19711
rect -3375 19371 -3266 19379
rect -3387 19369 -3266 19371
rect -3387 19249 -3375 19369
rect -3319 19249 -3266 19369
rect -3387 19247 -3266 19249
rect -3375 19239 -3319 19247
rect -4072 18982 -3176 18994
rect -4072 18926 -4060 18982
rect -4004 18926 -3242 18982
rect -3186 18926 -3176 18982
rect -4072 18914 -3176 18926
rect -3065 18757 -3009 19701
rect -2349 19512 -2293 19826
rect -2165 19770 -2109 19968
rect -2177 19768 -2097 19770
rect -2177 19712 -2165 19768
rect -2109 19712 -2097 19768
rect -2177 19710 -2097 19712
rect -2165 19512 -2109 19710
rect -1981 19654 -1925 19968
rect -1848 19770 -1780 20100
rect -1403 19778 -1347 21012
rect -1848 19768 -1768 19770
rect -1848 19712 -1836 19768
rect -1780 19712 -1768 19768
rect -1848 19710 -1768 19712
rect -1405 19768 -1335 19778
rect -1405 19712 -1403 19768
rect -1347 19712 -1255 19768
rect -1993 19652 -1913 19654
rect -1993 19596 -1981 19652
rect -1925 19596 -1913 19652
rect -1993 19594 -1913 19596
rect -1981 19512 -1925 19594
rect -2361 19502 -2281 19512
rect -2361 19446 -2349 19502
rect -2293 19446 -2281 19502
rect -2361 19436 -2281 19446
rect -2177 19502 -2097 19512
rect -2177 19446 -2165 19502
rect -2109 19446 -2097 19502
rect -2177 19436 -2097 19446
rect -1993 19502 -1913 19512
rect -1993 19446 -1981 19502
rect -1925 19446 -1913 19502
rect -1993 19436 -1913 19446
rect -1848 19380 -1780 19710
rect -1405 19700 -1335 19712
rect -1889 19372 -1780 19380
rect -1901 19370 -1780 19372
rect -1901 19250 -1889 19370
rect -1833 19250 -1780 19370
rect -1901 19248 -1780 19250
rect -1889 19240 -1833 19248
rect -2586 18983 -1690 18995
rect -2586 18927 -2574 18983
rect -2518 18927 -1756 18983
rect -1700 18927 -1690 18983
rect -2586 18915 -1690 18927
rect -2901 18864 -2821 18874
rect -2901 18808 -2889 18864
rect -2833 18808 -2821 18864
rect -2901 18806 -2821 18808
rect -3067 18754 -2997 18757
rect -3067 18700 -3065 18754
rect -3009 18700 -2997 18754
rect -3067 18688 -2997 18700
rect -3927 18647 -3181 18659
rect -3927 18591 -3559 18647
rect -3503 18591 -3181 18647
rect -3927 18579 -3181 18591
rect -3927 18326 -3871 18579
rect -3559 18326 -3503 18579
rect -3237 18326 -3181 18579
rect -3939 18324 -3859 18326
rect -3939 18204 -3927 18324
rect -3871 18204 -3859 18324
rect -3939 18202 -3859 18204
rect -3571 18324 -3491 18326
rect -3571 18204 -3559 18324
rect -3503 18204 -3491 18324
rect -3571 18202 -3491 18204
rect -3249 18324 -3169 18326
rect -3249 18203 -3237 18324
rect -3181 18203 -3169 18324
rect -3927 18194 -3871 18202
rect -3559 18194 -3503 18202
rect -3249 18201 -3169 18203
rect -3237 18193 -3181 18201
rect -3743 18026 -3687 18034
rect -3375 18026 -3319 18034
rect -3755 18024 -3266 18026
rect -3755 17904 -3743 18024
rect -3687 17904 -3375 18024
rect -3319 17904 -3266 18024
rect -3755 17902 -3266 17904
rect -3743 17894 -3687 17902
rect -3375 17894 -3266 17902
rect -3847 17828 -3767 17838
rect -3847 17772 -3835 17828
rect -3779 17772 -3767 17828
rect -3847 17762 -3767 17772
rect -3663 17828 -3583 17838
rect -3663 17772 -3651 17828
rect -3595 17772 -3583 17828
rect -3663 17762 -3583 17772
rect -3479 17828 -3399 17838
rect -3479 17772 -3467 17828
rect -3411 17772 -3399 17828
rect -3479 17762 -3399 17772
rect -3835 17680 -3779 17762
rect -3847 17678 -3767 17680
rect -3847 17622 -3835 17678
rect -3779 17622 -3767 17678
rect -3847 17620 -3767 17622
rect -4655 17562 -4585 17576
rect -4655 17506 -4643 17562
rect -4587 17506 -4585 17562
rect -4655 17494 -4585 17506
rect -4957 16659 -4887 16671
rect -4643 16663 -4587 17494
rect -3835 17306 -3779 17620
rect -3651 17564 -3595 17762
rect -3663 17562 -3583 17564
rect -3663 17506 -3651 17562
rect -3595 17506 -3583 17562
rect -3663 17504 -3583 17506
rect -3651 17306 -3595 17504
rect -3467 17448 -3411 17762
rect -3334 17564 -3266 17894
rect -2889 17574 -2833 18806
rect -3334 17562 -3254 17564
rect -3334 17506 -3322 17562
rect -3266 17506 -3254 17562
rect -3334 17504 -3254 17506
rect -2891 17562 -2831 17574
rect -2891 17506 -2889 17562
rect -2833 17506 -2831 17562
rect -3479 17446 -3399 17448
rect -3479 17390 -3467 17446
rect -3411 17390 -3399 17446
rect -3479 17388 -3399 17390
rect -3467 17306 -3411 17388
rect -3847 17296 -3767 17306
rect -3847 17240 -3835 17296
rect -3779 17240 -3767 17296
rect -3847 17230 -3767 17240
rect -3663 17296 -3583 17306
rect -3663 17240 -3651 17296
rect -3595 17240 -3583 17296
rect -3663 17230 -3583 17240
rect -3479 17296 -3399 17306
rect -3479 17240 -3467 17296
rect -3411 17240 -3399 17296
rect -3479 17230 -3399 17240
rect -3334 17174 -3266 17504
rect -2891 17494 -2831 17506
rect -1459 17446 -1389 17458
rect -1459 17390 -1447 17446
rect -1391 17390 -1389 17446
rect -1459 17378 -1389 17390
rect -3375 17166 -3266 17174
rect -3387 17164 -3266 17166
rect -3387 17044 -3375 17164
rect -3319 17044 -3266 17164
rect -3387 17042 -3266 17044
rect -3375 17034 -3319 17042
rect -4072 16777 -3174 16789
rect -4072 16721 -4060 16777
rect -4004 16721 -3242 16777
rect -3186 16721 -3174 16777
rect -4072 16709 -3174 16721
rect -4957 16603 -4945 16659
rect -4889 16603 -4887 16659
rect -4957 16601 -4887 16603
rect -4645 16659 -4585 16663
rect -4645 16603 -4643 16659
rect -4587 16603 -4585 16659
rect -4945 15989 -4889 16601
rect -4645 16591 -4585 16603
rect -1447 16499 -1391 17378
rect -1447 16389 -1391 16399
rect -5093 11494 -5023 11506
rect -5093 11438 -5081 11494
rect -5025 11438 -5023 11494
rect -5093 11426 -5023 11438
rect -5447 10136 -5445 10192
rect -5389 10136 -5161 10192
rect -6035 10076 -5955 10078
rect -6035 10020 -6023 10076
rect -5967 10020 -5955 10076
rect -6035 10018 -5955 10020
rect -6023 9936 -5967 10018
rect -6403 9926 -6323 9936
rect -6403 9870 -6391 9926
rect -6335 9870 -6323 9926
rect -6403 9860 -6323 9870
rect -6219 9926 -6139 9936
rect -6219 9870 -6207 9926
rect -6151 9870 -6139 9926
rect -6219 9860 -6139 9870
rect -6035 9926 -5955 9936
rect -6035 9870 -6023 9926
rect -5967 9870 -5955 9926
rect -6035 9860 -5955 9870
rect -5890 9804 -5822 10134
rect -5447 10124 -5377 10136
rect -5931 9796 -5822 9804
rect -5943 9794 -5822 9796
rect -5943 9674 -5931 9794
rect -5875 9674 -5822 9794
rect -5943 9672 -5822 9674
rect -5931 9664 -5875 9672
rect -6628 9407 -5732 9419
rect -6628 9351 -6616 9407
rect -6560 9351 -5798 9407
rect -5742 9351 -5732 9407
rect -6628 9339 -5732 9351
rect -6943 9288 -6863 9298
rect -6943 9232 -6931 9288
rect -6875 9232 -6863 9288
rect -6943 9230 -6863 9232
rect -7109 9178 -7039 9181
rect -7109 9124 -7107 9178
rect -7051 9124 -7039 9178
rect -7109 9112 -7039 9124
rect -7969 9071 -7223 9083
rect -7969 9015 -7601 9071
rect -7545 9015 -7223 9071
rect -7969 9003 -7223 9015
rect -7969 8750 -7913 9003
rect -7601 8750 -7545 9003
rect -7279 8750 -7223 9003
rect -7981 8748 -7901 8750
rect -7981 8628 -7969 8748
rect -7913 8628 -7901 8748
rect -7981 8626 -7901 8628
rect -7613 8748 -7533 8750
rect -7613 8628 -7601 8748
rect -7545 8628 -7533 8748
rect -7613 8626 -7533 8628
rect -7291 8748 -7211 8750
rect -7291 8627 -7279 8748
rect -7223 8627 -7211 8748
rect -7969 8618 -7913 8626
rect -7601 8618 -7545 8626
rect -7291 8625 -7211 8627
rect -7279 8617 -7223 8625
rect -7785 8450 -7729 8458
rect -7417 8450 -7361 8458
rect -7797 8448 -7308 8450
rect -7797 8328 -7785 8448
rect -7729 8328 -7417 8448
rect -7361 8328 -7308 8448
rect -7797 8326 -7308 8328
rect -7785 8318 -7729 8326
rect -7417 8318 -7308 8326
rect -7889 8252 -7809 8262
rect -7889 8196 -7877 8252
rect -7821 8196 -7809 8252
rect -7889 8186 -7809 8196
rect -7705 8252 -7625 8262
rect -7705 8196 -7693 8252
rect -7637 8196 -7625 8252
rect -7705 8186 -7625 8196
rect -7521 8252 -7441 8262
rect -7521 8196 -7509 8252
rect -7453 8196 -7441 8252
rect -7521 8186 -7441 8196
rect -7877 8104 -7821 8186
rect -7889 8102 -7809 8104
rect -7889 8046 -7877 8102
rect -7821 8046 -7809 8102
rect -7889 8044 -7809 8046
rect -8697 7986 -8627 8000
rect -8697 7930 -8685 7986
rect -8629 7930 -8627 7986
rect -8697 7918 -8627 7930
rect -8833 7870 -8763 7882
rect -8833 7814 -8821 7870
rect -8765 7814 -8763 7870
rect -8833 7802 -8763 7814
rect -8969 7083 -8899 7095
rect -8685 7087 -8629 7918
rect -7877 7730 -7821 8044
rect -7693 7988 -7637 8186
rect -7705 7986 -7625 7988
rect -7705 7930 -7693 7986
rect -7637 7930 -7625 7986
rect -7705 7928 -7625 7930
rect -7693 7730 -7637 7928
rect -7509 7872 -7453 8186
rect -7376 7988 -7308 8318
rect -6931 7998 -6875 9230
rect -7376 7986 -7296 7988
rect -7376 7930 -7364 7986
rect -7308 7930 -7296 7986
rect -7376 7928 -7296 7930
rect -6933 7986 -6873 7998
rect -6933 7930 -6931 7986
rect -6875 7930 -6873 7986
rect -7521 7870 -7441 7872
rect -7521 7814 -7509 7870
rect -7453 7814 -7441 7870
rect -7521 7812 -7441 7814
rect -7509 7730 -7453 7812
rect -7889 7720 -7809 7730
rect -7889 7664 -7877 7720
rect -7821 7664 -7809 7720
rect -7889 7654 -7809 7664
rect -7705 7720 -7625 7730
rect -7705 7664 -7693 7720
rect -7637 7664 -7625 7720
rect -7705 7654 -7625 7664
rect -7521 7720 -7441 7730
rect -7521 7664 -7509 7720
rect -7453 7664 -7441 7720
rect -7521 7654 -7441 7664
rect -7376 7598 -7308 7928
rect -6933 7918 -6873 7930
rect -7417 7590 -7308 7598
rect -7429 7588 -7308 7590
rect -7429 7468 -7417 7588
rect -7361 7468 -7308 7588
rect -7429 7466 -7308 7468
rect -7417 7458 -7361 7466
rect -8114 7201 -7216 7213
rect -8114 7145 -8102 7201
rect -8046 7145 -7284 7201
rect -7228 7145 -7216 7201
rect -8114 7133 -7216 7145
rect -8969 7027 -8957 7083
rect -8901 7027 -8899 7083
rect -8969 7015 -8899 7027
rect -8687 7083 -8627 7087
rect -8687 7027 -8685 7083
rect -8629 7027 -8627 7083
rect -8687 7015 -8627 7027
rect -9093 6810 -9037 6820
rect -5081 6920 -5025 11426
rect -4945 7095 -4889 15889
rect -3927 15686 -3181 15698
rect -3927 15630 -3559 15686
rect -3503 15630 -3181 15686
rect -3927 15618 -3181 15630
rect -3927 15365 -3871 15618
rect -3559 15365 -3503 15618
rect -3237 15365 -3181 15618
rect -3939 15363 -3859 15365
rect -3939 15243 -3927 15363
rect -3871 15243 -3859 15363
rect -3939 15241 -3859 15243
rect -3571 15363 -3491 15365
rect -3571 15243 -3559 15363
rect -3503 15243 -3491 15363
rect -3571 15241 -3491 15243
rect -3249 15363 -3169 15365
rect -3249 15242 -3237 15363
rect -3181 15242 -3169 15363
rect -3927 15233 -3871 15241
rect -3559 15233 -3503 15241
rect -3249 15240 -3169 15242
rect -3237 15232 -3181 15240
rect -3743 15065 -3687 15073
rect -3375 15065 -3319 15073
rect -3755 15063 -3266 15065
rect -3755 14943 -3743 15063
rect -3687 14943 -3375 15063
rect -3319 14943 -3266 15063
rect -3755 14941 -3266 14943
rect -3743 14933 -3687 14941
rect -3375 14933 -3266 14941
rect -3847 14867 -3767 14877
rect -3847 14811 -3835 14867
rect -3779 14811 -3767 14867
rect -3847 14801 -3767 14811
rect -3663 14867 -3583 14877
rect -3663 14811 -3651 14867
rect -3595 14811 -3583 14867
rect -3663 14801 -3583 14811
rect -3479 14867 -3399 14877
rect -3479 14811 -3467 14867
rect -3411 14811 -3399 14867
rect -3479 14801 -3399 14811
rect -4735 14717 -4649 14729
rect -3835 14719 -3779 14801
rect -4735 14661 -4723 14717
rect -4667 14661 -4649 14717
rect -4735 14649 -4649 14661
rect -3847 14717 -3767 14719
rect -3847 14661 -3835 14717
rect -3779 14661 -3767 14717
rect -3847 14659 -3767 14661
rect -4519 14601 -4449 14613
rect -4519 14545 -4507 14601
rect -4451 14545 -4449 14601
rect -4519 14533 -4449 14545
rect -4655 12396 -4585 12410
rect -4655 12340 -4643 12396
rect -4587 12340 -4585 12396
rect -4655 12328 -4585 12340
rect -4821 12208 -4741 12218
rect -4821 12152 -4809 12208
rect -4753 12152 -4741 12208
rect -4821 12150 -4741 12152
rect -4809 7882 -4753 12150
rect -4643 8000 -4587 12328
rect -4507 10087 -4451 14533
rect -3835 14345 -3779 14659
rect -3651 14603 -3595 14801
rect -3663 14601 -3583 14603
rect -3663 14545 -3651 14601
rect -3595 14545 -3583 14601
rect -3663 14543 -3583 14545
rect -3651 14345 -3595 14543
rect -3467 14487 -3411 14801
rect -3334 14603 -3266 14933
rect -3334 14601 -3254 14603
rect -3334 14545 -3322 14601
rect -3266 14545 -3254 14601
rect -3334 14543 -3254 14545
rect -3067 14601 -2997 14613
rect -3067 14545 -3065 14601
rect -3009 14545 -2997 14601
rect -3479 14485 -3399 14487
rect -3479 14429 -3467 14485
rect -3411 14429 -3399 14485
rect -3479 14427 -3399 14429
rect -3467 14345 -3411 14427
rect -3847 14335 -3767 14345
rect -3847 14279 -3835 14335
rect -3779 14279 -3767 14335
rect -3847 14269 -3767 14279
rect -3663 14335 -3583 14345
rect -3663 14279 -3651 14335
rect -3595 14279 -3583 14335
rect -3663 14269 -3583 14279
rect -3479 14335 -3399 14345
rect -3479 14279 -3467 14335
rect -3411 14279 -3399 14335
rect -3479 14269 -3399 14279
rect -3334 14213 -3266 14543
rect -3067 14535 -2997 14545
rect -3375 14205 -3266 14213
rect -3387 14203 -3266 14205
rect -3387 14083 -3375 14203
rect -3319 14083 -3266 14203
rect -3387 14081 -3266 14083
rect -3375 14073 -3319 14081
rect -4072 13816 -3174 13828
rect -4072 13760 -4060 13816
rect -4004 13760 -3242 13816
rect -3186 13760 -3174 13816
rect -4072 13748 -3174 13760
rect -3065 13591 -3009 14535
rect -2901 13698 -2821 13708
rect -2901 13642 -2889 13698
rect -2833 13642 -2821 13698
rect -2901 13640 -2821 13642
rect -3067 13588 -2997 13591
rect -3067 13534 -3065 13588
rect -3009 13534 -2997 13588
rect -3067 13522 -2997 13534
rect -3927 13481 -3181 13493
rect -3927 13425 -3559 13481
rect -3503 13425 -3181 13481
rect -3927 13413 -3181 13425
rect -3927 13160 -3871 13413
rect -3559 13160 -3503 13413
rect -3237 13160 -3181 13413
rect -3939 13158 -3859 13160
rect -3939 13038 -3927 13158
rect -3871 13038 -3859 13158
rect -3939 13036 -3859 13038
rect -3571 13158 -3491 13160
rect -3571 13038 -3559 13158
rect -3503 13038 -3491 13158
rect -3571 13036 -3491 13038
rect -3249 13158 -3169 13160
rect -3249 13037 -3237 13158
rect -3181 13037 -3169 13158
rect -3927 13028 -3871 13036
rect -3559 13028 -3503 13036
rect -3249 13035 -3169 13037
rect -3237 13027 -3181 13035
rect -3743 12860 -3687 12868
rect -3375 12860 -3319 12868
rect -3755 12858 -3266 12860
rect -3755 12738 -3743 12858
rect -3687 12738 -3375 12858
rect -3319 12738 -3266 12858
rect -3755 12736 -3266 12738
rect -3743 12728 -3687 12736
rect -3375 12728 -3266 12736
rect -3847 12662 -3767 12672
rect -3847 12606 -3835 12662
rect -3779 12606 -3767 12662
rect -3847 12596 -3767 12606
rect -3663 12662 -3583 12672
rect -3663 12606 -3651 12662
rect -3595 12606 -3583 12662
rect -3663 12596 -3583 12606
rect -3479 12662 -3399 12672
rect -3479 12606 -3467 12662
rect -3411 12606 -3399 12662
rect -3479 12596 -3399 12606
rect -3835 12514 -3779 12596
rect -3847 12512 -3767 12514
rect -3847 12456 -3835 12512
rect -3779 12456 -3767 12512
rect -3847 12454 -3767 12456
rect -3835 12140 -3779 12454
rect -3651 12398 -3595 12596
rect -3663 12396 -3583 12398
rect -3663 12340 -3651 12396
rect -3595 12340 -3583 12396
rect -3663 12338 -3583 12340
rect -3651 12140 -3595 12338
rect -3467 12282 -3411 12596
rect -3334 12398 -3266 12728
rect -2889 12406 -2833 13640
rect -2441 13481 -1695 13493
rect -2441 13425 -2073 13481
rect -2017 13425 -1695 13481
rect -2441 13413 -1695 13425
rect -2441 13160 -2385 13413
rect -2073 13160 -2017 13413
rect -1751 13160 -1695 13413
rect -2453 13158 -2373 13160
rect -2453 13038 -2441 13158
rect -2385 13038 -2373 13158
rect -2453 13036 -2373 13038
rect -2085 13158 -2005 13160
rect -2085 13038 -2073 13158
rect -2017 13038 -2005 13158
rect -2085 13036 -2005 13038
rect -1763 13158 -1683 13160
rect -1763 13037 -1751 13158
rect -1695 13037 -1683 13158
rect -2441 13028 -2385 13036
rect -2073 13028 -2017 13036
rect -1763 13035 -1683 13037
rect -1751 13027 -1695 13035
rect -2257 12860 -2201 12868
rect -1889 12860 -1833 12868
rect -2269 12858 -1780 12860
rect -2269 12738 -2257 12858
rect -2201 12738 -1889 12858
rect -1833 12738 -1780 12858
rect -2269 12736 -1780 12738
rect -2257 12728 -2201 12736
rect -1889 12728 -1780 12736
rect -2361 12662 -2281 12672
rect -2361 12606 -2349 12662
rect -2293 12606 -2281 12662
rect -2361 12596 -2281 12606
rect -2177 12662 -2097 12672
rect -2177 12606 -2165 12662
rect -2109 12606 -2097 12662
rect -2177 12596 -2097 12606
rect -1993 12662 -1913 12672
rect -1993 12606 -1981 12662
rect -1925 12606 -1913 12662
rect -1993 12596 -1913 12606
rect -2349 12514 -2293 12596
rect -2361 12512 -2281 12514
rect -2361 12456 -2349 12512
rect -2293 12456 -2281 12512
rect -2361 12454 -2281 12456
rect -3334 12396 -3254 12398
rect -3334 12340 -3322 12396
rect -3266 12340 -3254 12396
rect -3334 12338 -3254 12340
rect -2891 12396 -2831 12406
rect -2891 12340 -2889 12396
rect -2833 12340 -2831 12396
rect -3479 12280 -3399 12282
rect -3479 12224 -3467 12280
rect -3411 12224 -3399 12280
rect -3479 12222 -3399 12224
rect -3467 12140 -3411 12222
rect -3847 12130 -3767 12140
rect -3847 12074 -3835 12130
rect -3779 12074 -3767 12130
rect -3847 12064 -3767 12074
rect -3663 12130 -3583 12140
rect -3663 12074 -3651 12130
rect -3595 12074 -3583 12130
rect -3663 12064 -3583 12074
rect -3479 12130 -3399 12140
rect -3479 12074 -3467 12130
rect -3411 12074 -3399 12130
rect -3479 12064 -3399 12074
rect -3334 12008 -3266 12338
rect -2891 12328 -2831 12340
rect -3375 12000 -3266 12008
rect -3387 11998 -3266 12000
rect -3387 11878 -3375 11998
rect -3319 11878 -3266 11998
rect -3387 11876 -3266 11878
rect -3375 11868 -3319 11876
rect -4072 11611 -3176 11623
rect -4072 11555 -4060 11611
rect -4004 11555 -3242 11611
rect -3186 11555 -3176 11611
rect -4072 11543 -3176 11555
rect -2889 11385 -2833 12328
rect -2349 12140 -2293 12454
rect -2165 12398 -2109 12596
rect -2177 12396 -2097 12398
rect -2177 12340 -2165 12396
rect -2109 12340 -2097 12396
rect -2177 12338 -2097 12340
rect -2165 12140 -2109 12338
rect -1981 12282 -1925 12596
rect -1848 12398 -1780 12728
rect -1848 12396 -1768 12398
rect -1848 12340 -1836 12396
rect -1780 12340 -1768 12396
rect -1848 12338 -1768 12340
rect -1581 12396 -1511 12408
rect -1581 12340 -1579 12396
rect -1523 12340 -1255 12396
rect -1993 12280 -1913 12282
rect -1993 12224 -1981 12280
rect -1925 12224 -1913 12280
rect -1993 12222 -1913 12224
rect -1981 12140 -1925 12222
rect -2361 12130 -2281 12140
rect -2361 12074 -2349 12130
rect -2293 12074 -2281 12130
rect -2361 12064 -2281 12074
rect -2177 12130 -2097 12140
rect -2177 12074 -2165 12130
rect -2109 12074 -2097 12130
rect -2177 12064 -2097 12074
rect -1993 12130 -1913 12140
rect -1993 12074 -1981 12130
rect -1925 12074 -1913 12130
rect -1993 12064 -1913 12074
rect -1848 12008 -1780 12338
rect -1581 12330 -1511 12340
rect -1889 12000 -1780 12008
rect -1901 11998 -1780 12000
rect -1901 11878 -1889 11998
rect -1833 11878 -1780 11998
rect -1901 11876 -1780 11878
rect -1889 11868 -1833 11876
rect -2586 11611 -1690 11623
rect -2586 11555 -2574 11611
rect -2518 11555 -1756 11611
rect -1700 11555 -1690 11611
rect -2586 11543 -1690 11555
rect -1579 11386 -1523 12330
rect -1415 11494 -1335 11504
rect -1415 11438 -1403 11494
rect -1347 11438 -1335 11494
rect -1415 11436 -1335 11438
rect -2891 11383 -2821 11385
rect -2891 11327 -2889 11383
rect -2833 11327 -2821 11383
rect -2891 11315 -2821 11327
rect -1591 11384 -1511 11386
rect -1591 11328 -1579 11384
rect -1523 11328 -1511 11384
rect -1591 11316 -1511 11328
rect -3927 11276 -3181 11288
rect -3927 11220 -3559 11276
rect -3503 11220 -3181 11276
rect -3927 11208 -3181 11220
rect -3927 10955 -3871 11208
rect -3559 10955 -3503 11208
rect -3237 10955 -3181 11208
rect -2441 11277 -1695 11289
rect -2441 11221 -2073 11277
rect -2017 11221 -1695 11277
rect -2441 11209 -1695 11221
rect -2441 10956 -2385 11209
rect -2073 10956 -2017 11209
rect -1751 10956 -1695 11209
rect -3939 10953 -3859 10955
rect -3939 10833 -3927 10953
rect -3871 10833 -3859 10953
rect -3939 10831 -3859 10833
rect -3571 10953 -3491 10955
rect -3571 10833 -3559 10953
rect -3503 10833 -3491 10953
rect -3571 10831 -3491 10833
rect -3249 10953 -3169 10955
rect -3249 10832 -3237 10953
rect -3181 10832 -3169 10953
rect -2453 10954 -2373 10956
rect -2453 10834 -2441 10954
rect -2385 10834 -2373 10954
rect -2453 10832 -2373 10834
rect -2085 10954 -2005 10956
rect -2085 10834 -2073 10954
rect -2017 10834 -2005 10954
rect -2085 10832 -2005 10834
rect -1763 10954 -1683 10956
rect -1763 10833 -1751 10954
rect -1695 10833 -1683 10954
rect -3927 10823 -3871 10831
rect -3559 10823 -3503 10831
rect -3249 10830 -3169 10832
rect -3237 10822 -3181 10830
rect -2441 10824 -2385 10832
rect -2073 10824 -2017 10832
rect -1763 10831 -1683 10833
rect -1751 10823 -1695 10831
rect -3743 10655 -3687 10663
rect -3375 10655 -3319 10663
rect -2257 10656 -2201 10664
rect -1889 10656 -1833 10664
rect -3755 10653 -3266 10655
rect -3755 10533 -3743 10653
rect -3687 10533 -3375 10653
rect -3319 10533 -3266 10653
rect -3755 10531 -3266 10533
rect -2269 10654 -1780 10656
rect -2269 10534 -2257 10654
rect -2201 10534 -1889 10654
rect -1833 10534 -1780 10654
rect -2269 10532 -1780 10534
rect -3743 10523 -3687 10531
rect -3375 10523 -3266 10531
rect -2257 10524 -2201 10532
rect -1889 10524 -1780 10532
rect -3847 10457 -3767 10467
rect -3847 10401 -3835 10457
rect -3779 10401 -3767 10457
rect -3847 10391 -3767 10401
rect -3663 10457 -3583 10467
rect -3663 10401 -3651 10457
rect -3595 10401 -3583 10457
rect -3663 10391 -3583 10401
rect -3479 10457 -3399 10467
rect -3479 10401 -3467 10457
rect -3411 10401 -3399 10457
rect -3479 10391 -3399 10401
rect -3835 10309 -3779 10391
rect -3847 10307 -3767 10309
rect -3847 10251 -3835 10307
rect -3779 10251 -3767 10307
rect -3847 10249 -3767 10251
rect -4519 10075 -4449 10087
rect -4519 10019 -4507 10075
rect -4451 10019 -4449 10075
rect -4519 10007 -4449 10019
rect -3835 9935 -3779 10249
rect -3651 10193 -3595 10391
rect -3663 10191 -3583 10193
rect -3663 10135 -3651 10191
rect -3595 10135 -3583 10191
rect -3663 10133 -3583 10135
rect -3651 9935 -3595 10133
rect -3467 10077 -3411 10391
rect -3334 10193 -3266 10523
rect -2361 10458 -2281 10468
rect -2361 10402 -2349 10458
rect -2293 10402 -2281 10458
rect -2361 10392 -2281 10402
rect -2177 10458 -2097 10468
rect -2177 10402 -2165 10458
rect -2109 10402 -2097 10458
rect -2177 10392 -2097 10402
rect -1993 10458 -1913 10468
rect -1993 10402 -1981 10458
rect -1925 10402 -1913 10458
rect -1993 10392 -1913 10402
rect -2349 10310 -2293 10392
rect -2361 10308 -2281 10310
rect -2361 10252 -2349 10308
rect -2293 10252 -2281 10308
rect -2361 10250 -2281 10252
rect -3334 10191 -3254 10193
rect -3334 10135 -3322 10191
rect -3266 10135 -3254 10191
rect -3334 10133 -3254 10135
rect -3067 10191 -2997 10203
rect -3067 10135 -3065 10191
rect -3009 10135 -2997 10191
rect -3479 10075 -3399 10077
rect -3479 10019 -3467 10075
rect -3411 10019 -3399 10075
rect -3479 10017 -3399 10019
rect -3467 9935 -3411 10017
rect -3847 9925 -3767 9935
rect -3847 9869 -3835 9925
rect -3779 9869 -3767 9925
rect -3847 9859 -3767 9869
rect -3663 9925 -3583 9935
rect -3663 9869 -3651 9925
rect -3595 9869 -3583 9925
rect -3663 9859 -3583 9869
rect -3479 9925 -3399 9935
rect -3479 9869 -3467 9925
rect -3411 9869 -3399 9925
rect -3479 9859 -3399 9869
rect -3334 9803 -3266 10133
rect -3067 10125 -2997 10135
rect -3375 9795 -3266 9803
rect -3387 9793 -3266 9795
rect -3387 9673 -3375 9793
rect -3319 9673 -3266 9793
rect -3387 9671 -3266 9673
rect -3375 9663 -3319 9671
rect -4072 9406 -3176 9418
rect -4072 9350 -4060 9406
rect -4004 9350 -3242 9406
rect -3186 9350 -3176 9406
rect -4072 9338 -3176 9350
rect -3065 9181 -3009 10125
rect -2349 9936 -2293 10250
rect -2165 10194 -2109 10392
rect -2177 10192 -2097 10194
rect -2177 10136 -2165 10192
rect -2109 10136 -2097 10192
rect -2177 10134 -2097 10136
rect -2165 9936 -2109 10134
rect -1981 10078 -1925 10392
rect -1848 10194 -1780 10524
rect -1403 10202 -1347 11436
rect -1848 10192 -1768 10194
rect -1848 10136 -1836 10192
rect -1780 10136 -1768 10192
rect -1848 10134 -1768 10136
rect -1405 10192 -1335 10202
rect -1175 10192 -1119 24235
rect -1027 21984 -971 25664
rect -1029 21972 -959 21984
rect -1029 21916 -1027 21972
rect -971 21916 -959 21972
rect -1029 21904 -959 21916
rect -737 21072 -681 26016
rect 3069 25548 3125 27289
rect 17275 27078 17331 28454
rect 19465 28442 19535 28454
rect 18755 28228 18835 28238
rect 18755 28172 18767 28228
rect 18823 28172 18835 28228
rect 18755 27986 18835 28172
rect 19235 28228 19315 28238
rect 19235 28172 19247 28228
rect 19303 28172 19315 28228
rect 19235 28162 19315 28172
rect 19439 28228 19519 28238
rect 19439 28172 19451 28228
rect 19507 28172 19519 28228
rect 19439 27986 19519 28172
rect 19643 28228 19723 28532
rect 19945 28520 20015 28532
rect 20123 28588 20203 28883
rect 20424 28588 20480 29618
rect 21557 29608 21653 29618
rect 21871 29402 21951 29696
rect 22173 29684 22243 29696
rect 22351 29752 22431 30047
rect 22989 29882 23045 34210
rect 23125 31969 23181 36415
rect 23797 36227 23853 36541
rect 23981 36485 24037 36683
rect 23969 36483 24049 36485
rect 23969 36427 23981 36483
rect 24037 36427 24049 36483
rect 23969 36425 24049 36427
rect 23981 36227 24037 36425
rect 24165 36369 24221 36683
rect 24298 36485 24366 36815
rect 33257 36749 33337 36759
rect 33257 36693 33269 36749
rect 33325 36693 33337 36749
rect 33257 36683 33337 36693
rect 33441 36749 33521 36759
rect 33441 36693 33453 36749
rect 33509 36693 33521 36749
rect 33441 36683 33521 36693
rect 33625 36749 33705 36759
rect 33625 36693 33637 36749
rect 33693 36693 33705 36749
rect 33625 36683 33705 36693
rect 32367 36599 32455 36611
rect 33269 36601 33325 36683
rect 32367 36543 32381 36599
rect 32437 36543 32455 36599
rect 32367 36531 32455 36543
rect 33257 36599 33337 36601
rect 33257 36543 33269 36599
rect 33325 36543 33337 36599
rect 33257 36541 33337 36543
rect 24298 36483 24378 36485
rect 24298 36427 24310 36483
rect 24366 36427 24378 36483
rect 24298 36425 24378 36427
rect 24565 36483 24635 36495
rect 24565 36427 24567 36483
rect 24623 36427 24635 36483
rect 24153 36367 24233 36369
rect 24153 36311 24165 36367
rect 24221 36311 24233 36367
rect 24153 36309 24233 36311
rect 24165 36227 24221 36309
rect 23785 36217 23865 36227
rect 23785 36161 23797 36217
rect 23853 36161 23865 36217
rect 23785 36151 23865 36161
rect 23969 36217 24049 36227
rect 23969 36161 23981 36217
rect 24037 36161 24049 36217
rect 23969 36151 24049 36161
rect 24153 36217 24233 36227
rect 24153 36161 24165 36217
rect 24221 36161 24233 36217
rect 24153 36151 24233 36161
rect 24298 36095 24366 36425
rect 24565 36417 24635 36427
rect 32585 36483 32655 36495
rect 32585 36427 32597 36483
rect 32653 36427 32655 36483
rect 24257 36087 24366 36095
rect 24245 36085 24366 36087
rect 24245 35965 24257 36085
rect 24313 35965 24366 36085
rect 24245 35963 24366 35965
rect 24257 35955 24313 35963
rect 23560 35698 24458 35710
rect 23560 35642 23572 35698
rect 23628 35642 24390 35698
rect 24446 35642 24458 35698
rect 23560 35630 24458 35642
rect 24567 35473 24623 36417
rect 32585 36415 32655 36427
rect 24731 35580 24811 35590
rect 24731 35524 24743 35580
rect 24799 35524 24811 35580
rect 24731 35522 24811 35524
rect 24565 35470 24635 35473
rect 24565 35416 24567 35470
rect 24623 35416 24635 35470
rect 24565 35404 24635 35416
rect 23705 35363 24451 35375
rect 23705 35307 24073 35363
rect 24129 35307 24451 35363
rect 23705 35295 24451 35307
rect 23705 35042 23761 35295
rect 24073 35042 24129 35295
rect 24395 35042 24451 35295
rect 23693 35040 23773 35042
rect 23693 34920 23705 35040
rect 23761 34920 23773 35040
rect 23693 34918 23773 34920
rect 24061 35040 24141 35042
rect 24061 34920 24073 35040
rect 24129 34920 24141 35040
rect 24061 34918 24141 34920
rect 24383 35040 24463 35042
rect 24383 34919 24395 35040
rect 24451 34919 24463 35040
rect 23705 34910 23761 34918
rect 24073 34910 24129 34918
rect 24383 34917 24463 34919
rect 24395 34909 24451 34917
rect 23889 34742 23945 34750
rect 24257 34742 24313 34750
rect 23877 34740 24366 34742
rect 23877 34620 23889 34740
rect 23945 34620 24257 34740
rect 24313 34620 24366 34740
rect 23877 34618 24366 34620
rect 23889 34610 23945 34618
rect 24257 34610 24366 34618
rect 23785 34544 23865 34554
rect 23785 34488 23797 34544
rect 23853 34488 23865 34544
rect 23785 34478 23865 34488
rect 23969 34544 24049 34554
rect 23969 34488 23981 34544
rect 24037 34488 24049 34544
rect 23969 34478 24049 34488
rect 24153 34544 24233 34554
rect 24153 34488 24165 34544
rect 24221 34488 24233 34544
rect 24153 34478 24233 34488
rect 23797 34396 23853 34478
rect 23785 34394 23865 34396
rect 23785 34338 23797 34394
rect 23853 34338 23865 34394
rect 23785 34336 23865 34338
rect 23797 34022 23853 34336
rect 23981 34280 24037 34478
rect 23969 34278 24049 34280
rect 23969 34222 23981 34278
rect 24037 34222 24049 34278
rect 23969 34220 24049 34222
rect 23981 34022 24037 34220
rect 24165 34164 24221 34478
rect 24298 34280 24366 34610
rect 24743 34288 24799 35522
rect 25191 35363 25937 35375
rect 25191 35307 25559 35363
rect 25615 35307 25937 35363
rect 25191 35295 25937 35307
rect 25191 35042 25247 35295
rect 25559 35042 25615 35295
rect 25881 35042 25937 35295
rect 25179 35040 25259 35042
rect 25179 34920 25191 35040
rect 25247 34920 25259 35040
rect 25179 34918 25259 34920
rect 25547 35040 25627 35042
rect 25547 34920 25559 35040
rect 25615 34920 25627 35040
rect 25547 34918 25627 34920
rect 25869 35040 25949 35042
rect 25869 34919 25881 35040
rect 25937 34919 25949 35040
rect 25191 34910 25247 34918
rect 25559 34910 25615 34918
rect 25869 34917 25949 34919
rect 25881 34909 25937 34917
rect 25375 34742 25431 34750
rect 25743 34742 25799 34750
rect 25363 34740 25852 34742
rect 25363 34620 25375 34740
rect 25431 34620 25743 34740
rect 25799 34620 25852 34740
rect 25363 34618 25852 34620
rect 25375 34610 25431 34618
rect 25743 34610 25852 34618
rect 25271 34544 25351 34554
rect 25271 34488 25283 34544
rect 25339 34488 25351 34544
rect 25271 34478 25351 34488
rect 25455 34544 25535 34554
rect 25455 34488 25467 34544
rect 25523 34488 25535 34544
rect 25455 34478 25535 34488
rect 25639 34544 25719 34554
rect 25639 34488 25651 34544
rect 25707 34488 25719 34544
rect 25639 34478 25719 34488
rect 25283 34396 25339 34478
rect 25271 34394 25351 34396
rect 25271 34338 25283 34394
rect 25339 34338 25351 34394
rect 25271 34336 25351 34338
rect 24298 34278 24378 34280
rect 24298 34222 24310 34278
rect 24366 34222 24378 34278
rect 24298 34220 24378 34222
rect 24741 34278 24801 34288
rect 24741 34222 24743 34278
rect 24799 34222 24801 34278
rect 24153 34162 24233 34164
rect 24153 34106 24165 34162
rect 24221 34106 24233 34162
rect 24153 34104 24233 34106
rect 24165 34022 24221 34104
rect 23785 34012 23865 34022
rect 23785 33956 23797 34012
rect 23853 33956 23865 34012
rect 23785 33946 23865 33956
rect 23969 34012 24049 34022
rect 23969 33956 23981 34012
rect 24037 33956 24049 34012
rect 23969 33946 24049 33956
rect 24153 34012 24233 34022
rect 24153 33956 24165 34012
rect 24221 33956 24233 34012
rect 24153 33946 24233 33956
rect 24298 33890 24366 34220
rect 24741 34210 24801 34222
rect 24257 33882 24366 33890
rect 24245 33880 24366 33882
rect 24245 33760 24257 33880
rect 24313 33760 24366 33880
rect 24245 33758 24366 33760
rect 24257 33750 24313 33758
rect 23560 33493 24456 33505
rect 23560 33437 23572 33493
rect 23628 33437 24390 33493
rect 24446 33437 24456 33493
rect 23560 33425 24456 33437
rect 24743 33267 24799 34210
rect 25283 34022 25339 34336
rect 25467 34280 25523 34478
rect 25455 34278 25535 34280
rect 25455 34222 25467 34278
rect 25523 34222 25535 34278
rect 25455 34220 25535 34222
rect 25467 34022 25523 34220
rect 25651 34164 25707 34478
rect 25784 34280 25852 34610
rect 25784 34278 25864 34280
rect 25784 34222 25796 34278
rect 25852 34222 25864 34278
rect 25784 34220 25864 34222
rect 26051 34278 26121 34290
rect 32449 34278 32519 34292
rect 26051 34222 26053 34278
rect 26109 34222 26807 34278
rect 25639 34162 25719 34164
rect 25639 34106 25651 34162
rect 25707 34106 25719 34162
rect 25639 34104 25719 34106
rect 25651 34022 25707 34104
rect 25271 34012 25351 34022
rect 25271 33956 25283 34012
rect 25339 33956 25351 34012
rect 25271 33946 25351 33956
rect 25455 34012 25535 34022
rect 25455 33956 25467 34012
rect 25523 33956 25535 34012
rect 25455 33946 25535 33956
rect 25639 34012 25719 34022
rect 25639 33956 25651 34012
rect 25707 33956 25719 34012
rect 25639 33946 25719 33956
rect 25784 33890 25852 34220
rect 26051 34212 26121 34222
rect 25743 33882 25852 33890
rect 25731 33880 25852 33882
rect 25731 33760 25743 33880
rect 25799 33760 25852 33880
rect 25731 33758 25852 33760
rect 25743 33750 25799 33758
rect 25046 33493 25942 33505
rect 25046 33437 25058 33493
rect 25114 33437 25876 33493
rect 25932 33437 25942 33493
rect 25046 33425 25942 33437
rect 26053 33268 26109 34212
rect 26217 33376 26297 33386
rect 26217 33320 26229 33376
rect 26285 33320 26297 33376
rect 26217 33318 26297 33320
rect 24741 33265 24811 33267
rect 24741 33209 24743 33265
rect 24799 33209 24811 33265
rect 24741 33197 24811 33209
rect 26041 33266 26121 33268
rect 26041 33210 26053 33266
rect 26109 33210 26121 33266
rect 26041 33198 26121 33210
rect 23705 33158 24451 33170
rect 23705 33102 24073 33158
rect 24129 33102 24451 33158
rect 23705 33090 24451 33102
rect 23705 32837 23761 33090
rect 24073 32837 24129 33090
rect 24395 32837 24451 33090
rect 25191 33159 25937 33171
rect 25191 33103 25559 33159
rect 25615 33103 25937 33159
rect 25191 33091 25937 33103
rect 25191 32838 25247 33091
rect 25559 32838 25615 33091
rect 25881 32838 25937 33091
rect 23693 32835 23773 32837
rect 23693 32715 23705 32835
rect 23761 32715 23773 32835
rect 23693 32713 23773 32715
rect 24061 32835 24141 32837
rect 24061 32715 24073 32835
rect 24129 32715 24141 32835
rect 24061 32713 24141 32715
rect 24383 32835 24463 32837
rect 24383 32714 24395 32835
rect 24451 32714 24463 32835
rect 25179 32836 25259 32838
rect 25179 32716 25191 32836
rect 25247 32716 25259 32836
rect 25179 32714 25259 32716
rect 25547 32836 25627 32838
rect 25547 32716 25559 32836
rect 25615 32716 25627 32836
rect 25547 32714 25627 32716
rect 25869 32836 25949 32838
rect 25869 32715 25881 32836
rect 25937 32715 25949 32836
rect 23705 32705 23761 32713
rect 24073 32705 24129 32713
rect 24383 32712 24463 32714
rect 24395 32704 24451 32712
rect 25191 32706 25247 32714
rect 25559 32706 25615 32714
rect 25869 32713 25949 32715
rect 25881 32705 25937 32713
rect 23889 32537 23945 32545
rect 24257 32537 24313 32545
rect 25375 32538 25431 32546
rect 25743 32538 25799 32546
rect 23877 32535 24366 32537
rect 23877 32415 23889 32535
rect 23945 32415 24257 32535
rect 24313 32415 24366 32535
rect 23877 32413 24366 32415
rect 25363 32536 25852 32538
rect 25363 32416 25375 32536
rect 25431 32416 25743 32536
rect 25799 32416 25852 32536
rect 25363 32414 25852 32416
rect 23889 32405 23945 32413
rect 24257 32405 24366 32413
rect 25375 32406 25431 32414
rect 25743 32406 25852 32414
rect 23785 32339 23865 32349
rect 23785 32283 23797 32339
rect 23853 32283 23865 32339
rect 23785 32273 23865 32283
rect 23969 32339 24049 32349
rect 23969 32283 23981 32339
rect 24037 32283 24049 32339
rect 23969 32273 24049 32283
rect 24153 32339 24233 32349
rect 24153 32283 24165 32339
rect 24221 32283 24233 32339
rect 24153 32273 24233 32283
rect 23797 32191 23853 32273
rect 23785 32189 23865 32191
rect 23785 32133 23797 32189
rect 23853 32133 23865 32189
rect 23785 32131 23865 32133
rect 23113 31957 23183 31969
rect 23113 31901 23125 31957
rect 23181 31901 23183 31957
rect 23113 31889 23183 31901
rect 23797 31817 23853 32131
rect 23981 32075 24037 32273
rect 23969 32073 24049 32075
rect 23969 32017 23981 32073
rect 24037 32017 24049 32073
rect 23969 32015 24049 32017
rect 23981 31817 24037 32015
rect 24165 31959 24221 32273
rect 24298 32075 24366 32405
rect 25271 32340 25351 32350
rect 25271 32284 25283 32340
rect 25339 32284 25351 32340
rect 25271 32274 25351 32284
rect 25455 32340 25535 32350
rect 25455 32284 25467 32340
rect 25523 32284 25535 32340
rect 25455 32274 25535 32284
rect 25639 32340 25719 32350
rect 25639 32284 25651 32340
rect 25707 32284 25719 32340
rect 25639 32274 25719 32284
rect 25283 32192 25339 32274
rect 25271 32190 25351 32192
rect 25271 32134 25283 32190
rect 25339 32134 25351 32190
rect 25271 32132 25351 32134
rect 24298 32073 24378 32075
rect 24298 32017 24310 32073
rect 24366 32017 24378 32073
rect 24298 32015 24378 32017
rect 24565 32073 24635 32085
rect 24565 32017 24567 32073
rect 24623 32017 24635 32073
rect 24153 31957 24233 31959
rect 24153 31901 24165 31957
rect 24221 31901 24233 31957
rect 24153 31899 24233 31901
rect 24165 31817 24221 31899
rect 23785 31807 23865 31817
rect 23785 31751 23797 31807
rect 23853 31751 23865 31807
rect 23785 31741 23865 31751
rect 23969 31807 24049 31817
rect 23969 31751 23981 31807
rect 24037 31751 24049 31807
rect 23969 31741 24049 31751
rect 24153 31807 24233 31817
rect 24153 31751 24165 31807
rect 24221 31751 24233 31807
rect 24153 31741 24233 31751
rect 24298 31685 24366 32015
rect 24565 32007 24635 32017
rect 24257 31677 24366 31685
rect 24245 31675 24366 31677
rect 24245 31555 24257 31675
rect 24313 31555 24366 31675
rect 24245 31553 24366 31555
rect 24257 31545 24313 31553
rect 23560 31288 24456 31300
rect 23560 31232 23572 31288
rect 23628 31232 24390 31288
rect 24446 31232 24456 31288
rect 23560 31220 24456 31232
rect 24567 31063 24623 32007
rect 25283 31818 25339 32132
rect 25467 32076 25523 32274
rect 25455 32074 25535 32076
rect 25455 32018 25467 32074
rect 25523 32018 25535 32074
rect 25455 32016 25535 32018
rect 25467 31818 25523 32016
rect 25651 31960 25707 32274
rect 25784 32076 25852 32406
rect 26229 32084 26285 33318
rect 25784 32074 25864 32076
rect 25784 32018 25796 32074
rect 25852 32018 25864 32074
rect 25784 32016 25864 32018
rect 26227 32074 26297 32084
rect 26227 32018 26229 32074
rect 26285 32018 26377 32074
rect 25639 31958 25719 31960
rect 25639 31902 25651 31958
rect 25707 31902 25719 31958
rect 25639 31900 25719 31902
rect 25651 31818 25707 31900
rect 25271 31808 25351 31818
rect 25271 31752 25283 31808
rect 25339 31752 25351 31808
rect 25271 31742 25351 31752
rect 25455 31808 25535 31818
rect 25455 31752 25467 31808
rect 25523 31752 25535 31808
rect 25455 31742 25535 31752
rect 25639 31808 25719 31818
rect 25639 31752 25651 31808
rect 25707 31752 25719 31808
rect 25639 31742 25719 31752
rect 25784 31686 25852 32016
rect 26227 32006 26297 32018
rect 25743 31678 25852 31686
rect 25731 31676 25852 31678
rect 25731 31556 25743 31676
rect 25799 31556 25852 31676
rect 25731 31554 25852 31556
rect 25743 31546 25799 31554
rect 25046 31289 25942 31301
rect 25046 31233 25058 31289
rect 25114 31233 25876 31289
rect 25932 31233 25942 31289
rect 25046 31221 25942 31233
rect 24731 31170 24811 31180
rect 24731 31114 24743 31170
rect 24799 31114 24811 31170
rect 24731 31112 24811 31114
rect 24565 31060 24635 31063
rect 24565 31006 24567 31060
rect 24623 31006 24635 31060
rect 24565 30994 24635 31006
rect 23705 30953 24451 30965
rect 23705 30897 24073 30953
rect 24129 30897 24451 30953
rect 23705 30885 24451 30897
rect 23705 30632 23761 30885
rect 24073 30632 24129 30885
rect 24395 30632 24451 30885
rect 23693 30630 23773 30632
rect 23693 30510 23705 30630
rect 23761 30510 23773 30630
rect 23693 30508 23773 30510
rect 24061 30630 24141 30632
rect 24061 30510 24073 30630
rect 24129 30510 24141 30630
rect 24061 30508 24141 30510
rect 24383 30630 24463 30632
rect 24383 30509 24395 30630
rect 24451 30509 24463 30630
rect 23705 30500 23761 30508
rect 24073 30500 24129 30508
rect 24383 30507 24463 30509
rect 24395 30499 24451 30507
rect 23889 30332 23945 30340
rect 24257 30332 24313 30340
rect 23877 30330 24366 30332
rect 23877 30210 23889 30330
rect 23945 30210 24257 30330
rect 24313 30210 24366 30330
rect 23877 30208 24366 30210
rect 23889 30200 23945 30208
rect 24257 30200 24366 30208
rect 23785 30134 23865 30144
rect 23785 30078 23797 30134
rect 23853 30078 23865 30134
rect 23785 30068 23865 30078
rect 23969 30134 24049 30144
rect 23969 30078 23981 30134
rect 24037 30078 24049 30134
rect 23969 30068 24049 30078
rect 24153 30134 24233 30144
rect 24153 30078 24165 30134
rect 24221 30078 24233 30134
rect 24153 30068 24233 30078
rect 23797 29986 23853 30068
rect 23785 29984 23865 29986
rect 23785 29928 23797 29984
rect 23853 29928 23865 29984
rect 23785 29926 23865 29928
rect 22977 29868 23047 29882
rect 22977 29812 22989 29868
rect 23045 29812 23047 29868
rect 22977 29800 23047 29812
rect 22743 29752 22821 29763
rect 22351 29751 22821 29752
rect 22351 29697 22755 29751
rect 22809 29697 22821 29751
rect 22351 29696 22821 29697
rect 20779 29392 21951 29402
rect 20779 29336 20791 29392
rect 20847 29336 21679 29392
rect 21735 29336 21951 29392
rect 20779 29326 21951 29336
rect 22351 29392 22431 29696
rect 22743 29685 22821 29696
rect 22351 29336 22363 29392
rect 22419 29336 22431 29392
rect 22351 29326 22431 29336
rect 20709 29014 22501 29026
rect 20709 28874 20721 29014
rect 22489 28874 22501 29014
rect 22794 28965 22880 28977
rect 22989 28969 23045 29800
rect 23797 29612 23853 29926
rect 23981 29870 24037 30068
rect 23969 29868 24049 29870
rect 23969 29812 23981 29868
rect 24037 29812 24049 29868
rect 23969 29810 24049 29812
rect 23981 29612 24037 29810
rect 24165 29754 24221 30068
rect 24298 29870 24366 30200
rect 24743 29880 24799 31112
rect 26751 31006 26807 34222
rect 32449 34222 32461 34278
rect 32517 34222 32519 34278
rect 32449 34210 32519 34222
rect 32167 33376 32249 33388
rect 32167 33320 32181 33376
rect 32237 33320 32249 33376
rect 32167 33308 32249 33320
rect 27161 31970 27381 31980
rect 27161 31170 27171 31970
rect 27371 31170 27381 31970
rect 31551 31970 31871 31980
rect 28023 31463 29195 31473
rect 28023 31223 28035 31463
rect 28091 31223 29127 31463
rect 29183 31223 29195 31463
rect 28023 31213 29195 31223
rect 27161 31160 27381 31170
rect 28117 31006 28195 31018
rect 26747 30950 28137 31006
rect 28193 30950 28195 31006
rect 28117 30938 28195 30950
rect 29115 30928 29195 31213
rect 29595 31463 29675 31473
rect 29595 31223 29607 31463
rect 29663 31223 29675 31463
rect 29417 30928 29487 30940
rect 29115 30872 29429 30928
rect 29485 30872 29487 30928
rect 28937 30850 29007 30862
rect 26747 30794 28949 30850
rect 29005 30794 29007 30850
rect 24298 29868 24378 29870
rect 24298 29812 24310 29868
rect 24366 29812 24378 29868
rect 24298 29810 24378 29812
rect 24741 29868 24801 29880
rect 24741 29812 24743 29868
rect 24799 29812 24801 29868
rect 24153 29752 24233 29754
rect 24153 29696 24165 29752
rect 24221 29696 24233 29752
rect 24153 29694 24233 29696
rect 24165 29612 24221 29694
rect 23785 29602 23865 29612
rect 23785 29546 23797 29602
rect 23853 29546 23865 29602
rect 23785 29536 23865 29546
rect 23969 29602 24049 29612
rect 23969 29546 23981 29602
rect 24037 29546 24049 29602
rect 23969 29536 24049 29546
rect 24153 29602 24233 29612
rect 24153 29546 24165 29602
rect 24221 29546 24233 29602
rect 24153 29536 24233 29546
rect 24298 29480 24366 29810
rect 24741 29800 24801 29812
rect 26859 29509 26915 30794
rect 28937 30782 29007 30794
rect 28227 30568 28307 30578
rect 28227 30512 28239 30568
rect 28295 30512 28307 30568
rect 28227 30326 28307 30512
rect 28707 30568 28787 30578
rect 28707 30512 28719 30568
rect 28775 30512 28787 30568
rect 28707 30502 28787 30512
rect 28911 30568 28991 30578
rect 28911 30512 28923 30568
rect 28979 30512 28991 30568
rect 28911 30326 28991 30512
rect 29115 30568 29195 30872
rect 29417 30860 29487 30872
rect 29595 30928 29675 31223
rect 31551 31170 31561 31970
rect 31861 31170 31871 31970
rect 31551 31160 31871 31170
rect 30181 30974 31973 30986
rect 29595 30872 29952 30928
rect 29115 30512 29127 30568
rect 29183 30512 29195 30568
rect 29115 30502 29195 30512
rect 29595 30568 29675 30872
rect 29595 30512 29607 30568
rect 29663 30512 29675 30568
rect 29595 30502 29675 30512
rect 28227 30254 28991 30326
rect 29121 30200 29745 30212
rect 29121 30060 29133 30200
rect 29733 30060 29745 30200
rect 27333 30043 27413 30053
rect 29121 30048 29745 30060
rect 27333 29803 27345 30043
rect 27401 29803 27413 30043
rect 29896 29830 29952 30872
rect 30181 30834 30193 30974
rect 31961 30834 31973 30974
rect 30181 30822 31973 30834
rect 30455 30571 31219 30581
rect 30455 30331 30467 30571
rect 30523 30331 31151 30571
rect 31207 30331 31219 30571
rect 30455 30321 31219 30331
rect 31823 30287 31903 30297
rect 30935 30237 31423 30247
rect 30935 29997 30947 30237
rect 31003 29997 31355 30237
rect 31411 29997 31423 30237
rect 30935 29987 31423 29997
rect 30345 29830 30441 29842
rect 24257 29472 24366 29480
rect 24245 29470 24366 29472
rect 24245 29350 24257 29470
rect 24313 29350 24366 29470
rect 26347 29508 26915 29509
rect 27155 29508 27225 29520
rect 26347 29453 27167 29508
rect 24245 29348 24366 29350
rect 24257 29340 24313 29348
rect 23560 29083 24458 29095
rect 23560 29027 23572 29083
rect 23628 29027 24390 29083
rect 24446 29027 24458 29083
rect 23560 29015 24458 29027
rect 22794 28909 22806 28965
rect 22862 28909 22880 28965
rect 22794 28897 22880 28909
rect 22987 28965 23047 28969
rect 22987 28909 22989 28965
rect 23045 28909 23047 28965
rect 22987 28897 23047 28909
rect 20709 28862 22501 28874
rect 20123 28532 20480 28588
rect 22079 28690 22399 28700
rect 19643 28172 19655 28228
rect 19711 28172 19723 28228
rect 19643 28162 19723 28172
rect 20123 28228 20203 28532
rect 20123 28172 20135 28228
rect 20191 28172 20203 28228
rect 20123 28162 20203 28172
rect 18755 27914 19519 27986
rect 22079 27890 22089 28690
rect 22389 27890 22399 28690
rect 22079 27880 22399 27890
rect 26352 27610 26408 29453
rect 26859 29452 27167 29453
rect 27223 29452 27225 29508
rect 27155 29440 27225 29452
rect 27333 29508 27413 29803
rect 29121 29800 29745 29812
rect 29121 29660 29133 29800
rect 29733 29660 29745 29800
rect 29896 29774 30365 29830
rect 30421 29774 30441 29830
rect 30345 29762 30441 29774
rect 31343 29752 31423 29987
rect 31823 30047 31835 30287
rect 31891 30047 31903 30287
rect 31645 29752 31715 29764
rect 31343 29696 31657 29752
rect 31713 29696 31715 29752
rect 31029 29674 31125 29684
rect 29121 29648 29745 29660
rect 29896 29618 31049 29674
rect 31105 29618 31125 29674
rect 27333 29452 27771 29508
rect 27333 29148 27413 29452
rect 27333 29092 27345 29148
rect 27401 29092 27413 29148
rect 27333 29082 27413 29092
rect 27715 28666 27771 29452
rect 28023 29123 29195 29133
rect 28023 28883 28035 29123
rect 28091 28883 29127 29123
rect 29183 28883 29195 29123
rect 28023 28873 29195 28883
rect 28117 28666 28195 28678
rect 27715 28610 28137 28666
rect 28193 28610 28195 28666
rect 28117 28598 28195 28610
rect 29115 28588 29195 28873
rect 29595 29123 29675 29133
rect 29595 28883 29607 29123
rect 29663 28883 29675 29123
rect 29417 28588 29487 28600
rect 29115 28532 29429 28588
rect 29485 28532 29487 28588
rect 28937 28510 29007 28522
rect 26352 27480 26408 27490
rect 26747 28454 28949 28510
rect 29005 28454 29007 28510
rect 7111 27022 17331 27078
rect 7111 26076 7167 27022
rect 26747 26814 26803 28454
rect 28937 28442 29007 28454
rect 28227 28228 28307 28238
rect 28227 28172 28239 28228
rect 28295 28172 28307 28228
rect 28227 27986 28307 28172
rect 28707 28228 28787 28238
rect 28707 28172 28719 28228
rect 28775 28172 28787 28228
rect 28707 28162 28787 28172
rect 28911 28228 28991 28238
rect 28911 28172 28923 28228
rect 28979 28172 28991 28228
rect 28911 27986 28991 28172
rect 29115 28228 29195 28532
rect 29417 28520 29487 28532
rect 29595 28588 29675 28883
rect 29896 28588 29952 29618
rect 31029 29608 31125 29618
rect 31343 29402 31423 29696
rect 31645 29684 31715 29696
rect 31823 29752 31903 30047
rect 32461 29882 32517 34210
rect 32597 31969 32653 36415
rect 33269 36227 33325 36541
rect 33453 36485 33509 36683
rect 33441 36483 33521 36485
rect 33441 36427 33453 36483
rect 33509 36427 33521 36483
rect 33441 36425 33521 36427
rect 33453 36227 33509 36425
rect 33637 36369 33693 36683
rect 33770 36485 33838 36815
rect 42729 36749 42809 36759
rect 42729 36693 42741 36749
rect 42797 36693 42809 36749
rect 42729 36683 42809 36693
rect 42913 36749 42993 36759
rect 42913 36693 42925 36749
rect 42981 36693 42993 36749
rect 42913 36683 42993 36693
rect 43097 36749 43177 36759
rect 43097 36693 43109 36749
rect 43165 36693 43177 36749
rect 43097 36683 43177 36693
rect 41839 36599 41927 36611
rect 42741 36601 42797 36683
rect 41839 36543 41853 36599
rect 41909 36543 41927 36599
rect 41839 36531 41927 36543
rect 42729 36599 42809 36601
rect 42729 36543 42741 36599
rect 42797 36543 42809 36599
rect 42729 36541 42809 36543
rect 33770 36483 33850 36485
rect 33770 36427 33782 36483
rect 33838 36427 33850 36483
rect 33770 36425 33850 36427
rect 34037 36483 34107 36495
rect 34037 36427 34039 36483
rect 34095 36427 34107 36483
rect 33625 36367 33705 36369
rect 33625 36311 33637 36367
rect 33693 36311 33705 36367
rect 33625 36309 33705 36311
rect 33637 36227 33693 36309
rect 33257 36217 33337 36227
rect 33257 36161 33269 36217
rect 33325 36161 33337 36217
rect 33257 36151 33337 36161
rect 33441 36217 33521 36227
rect 33441 36161 33453 36217
rect 33509 36161 33521 36217
rect 33441 36151 33521 36161
rect 33625 36217 33705 36227
rect 33625 36161 33637 36217
rect 33693 36161 33705 36217
rect 33625 36151 33705 36161
rect 33770 36095 33838 36425
rect 34037 36417 34107 36427
rect 42057 36483 42127 36495
rect 42057 36427 42069 36483
rect 42125 36427 42127 36483
rect 33729 36087 33838 36095
rect 33717 36085 33838 36087
rect 33717 35965 33729 36085
rect 33785 35965 33838 36085
rect 33717 35963 33838 35965
rect 33729 35955 33785 35963
rect 33032 35698 33930 35710
rect 33032 35642 33044 35698
rect 33100 35642 33862 35698
rect 33918 35642 33930 35698
rect 33032 35630 33930 35642
rect 34039 35473 34095 36417
rect 42057 36415 42127 36427
rect 34203 35580 34283 35590
rect 34203 35524 34215 35580
rect 34271 35524 34283 35580
rect 34203 35522 34283 35524
rect 34037 35470 34107 35473
rect 34037 35416 34039 35470
rect 34095 35416 34107 35470
rect 34037 35404 34107 35416
rect 33177 35363 33923 35375
rect 33177 35307 33545 35363
rect 33601 35307 33923 35363
rect 33177 35295 33923 35307
rect 33177 35042 33233 35295
rect 33545 35042 33601 35295
rect 33867 35042 33923 35295
rect 33165 35040 33245 35042
rect 33165 34920 33177 35040
rect 33233 34920 33245 35040
rect 33165 34918 33245 34920
rect 33533 35040 33613 35042
rect 33533 34920 33545 35040
rect 33601 34920 33613 35040
rect 33533 34918 33613 34920
rect 33855 35040 33935 35042
rect 33855 34919 33867 35040
rect 33923 34919 33935 35040
rect 33177 34910 33233 34918
rect 33545 34910 33601 34918
rect 33855 34917 33935 34919
rect 33867 34909 33923 34917
rect 33361 34742 33417 34750
rect 33729 34742 33785 34750
rect 33349 34740 33838 34742
rect 33349 34620 33361 34740
rect 33417 34620 33729 34740
rect 33785 34620 33838 34740
rect 33349 34618 33838 34620
rect 33361 34610 33417 34618
rect 33729 34610 33838 34618
rect 33257 34544 33337 34554
rect 33257 34488 33269 34544
rect 33325 34488 33337 34544
rect 33257 34478 33337 34488
rect 33441 34544 33521 34554
rect 33441 34488 33453 34544
rect 33509 34488 33521 34544
rect 33441 34478 33521 34488
rect 33625 34544 33705 34554
rect 33625 34488 33637 34544
rect 33693 34488 33705 34544
rect 33625 34478 33705 34488
rect 33269 34396 33325 34478
rect 33257 34394 33337 34396
rect 33257 34338 33269 34394
rect 33325 34338 33337 34394
rect 33257 34336 33337 34338
rect 33269 34022 33325 34336
rect 33453 34280 33509 34478
rect 33441 34278 33521 34280
rect 33441 34222 33453 34278
rect 33509 34222 33521 34278
rect 33441 34220 33521 34222
rect 33453 34022 33509 34220
rect 33637 34164 33693 34478
rect 33770 34280 33838 34610
rect 34215 34288 34271 35522
rect 34663 35363 35409 35375
rect 34663 35307 35031 35363
rect 35087 35307 35409 35363
rect 34663 35295 35409 35307
rect 34663 35042 34719 35295
rect 35031 35042 35087 35295
rect 35353 35042 35409 35295
rect 34651 35040 34731 35042
rect 34651 34920 34663 35040
rect 34719 34920 34731 35040
rect 34651 34918 34731 34920
rect 35019 35040 35099 35042
rect 35019 34920 35031 35040
rect 35087 34920 35099 35040
rect 35019 34918 35099 34920
rect 35341 35040 35421 35042
rect 35341 34919 35353 35040
rect 35409 34919 35421 35040
rect 34663 34910 34719 34918
rect 35031 34910 35087 34918
rect 35341 34917 35421 34919
rect 35353 34909 35409 34917
rect 34847 34742 34903 34750
rect 35215 34742 35271 34750
rect 34835 34740 35324 34742
rect 34835 34620 34847 34740
rect 34903 34620 35215 34740
rect 35271 34620 35324 34740
rect 34835 34618 35324 34620
rect 34847 34610 34903 34618
rect 35215 34610 35324 34618
rect 34743 34544 34823 34554
rect 34743 34488 34755 34544
rect 34811 34488 34823 34544
rect 34743 34478 34823 34488
rect 34927 34544 35007 34554
rect 34927 34488 34939 34544
rect 34995 34488 35007 34544
rect 34927 34478 35007 34488
rect 35111 34544 35191 34554
rect 35111 34488 35123 34544
rect 35179 34488 35191 34544
rect 35111 34478 35191 34488
rect 34755 34396 34811 34478
rect 34743 34394 34823 34396
rect 34743 34338 34755 34394
rect 34811 34338 34823 34394
rect 34743 34336 34823 34338
rect 33770 34278 33850 34280
rect 33770 34222 33782 34278
rect 33838 34222 33850 34278
rect 33770 34220 33850 34222
rect 34213 34278 34273 34288
rect 34213 34222 34215 34278
rect 34271 34222 34273 34278
rect 33625 34162 33705 34164
rect 33625 34106 33637 34162
rect 33693 34106 33705 34162
rect 33625 34104 33705 34106
rect 33637 34022 33693 34104
rect 33257 34012 33337 34022
rect 33257 33956 33269 34012
rect 33325 33956 33337 34012
rect 33257 33946 33337 33956
rect 33441 34012 33521 34022
rect 33441 33956 33453 34012
rect 33509 33956 33521 34012
rect 33441 33946 33521 33956
rect 33625 34012 33705 34022
rect 33625 33956 33637 34012
rect 33693 33956 33705 34012
rect 33625 33946 33705 33956
rect 33770 33890 33838 34220
rect 34213 34210 34273 34222
rect 33729 33882 33838 33890
rect 33717 33880 33838 33882
rect 33717 33760 33729 33880
rect 33785 33760 33838 33880
rect 33717 33758 33838 33760
rect 33729 33750 33785 33758
rect 33032 33493 33928 33505
rect 33032 33437 33044 33493
rect 33100 33437 33862 33493
rect 33918 33437 33928 33493
rect 33032 33425 33928 33437
rect 34215 33267 34271 34210
rect 34755 34022 34811 34336
rect 34939 34280 34995 34478
rect 34927 34278 35007 34280
rect 34927 34222 34939 34278
rect 34995 34222 35007 34278
rect 34927 34220 35007 34222
rect 34939 34022 34995 34220
rect 35123 34164 35179 34478
rect 35256 34280 35324 34610
rect 35256 34278 35336 34280
rect 35256 34222 35268 34278
rect 35324 34222 35336 34278
rect 35256 34220 35336 34222
rect 35523 34278 35593 34290
rect 41921 34278 41991 34292
rect 35523 34222 35525 34278
rect 35581 34222 36279 34278
rect 35111 34162 35191 34164
rect 35111 34106 35123 34162
rect 35179 34106 35191 34162
rect 35111 34104 35191 34106
rect 35123 34022 35179 34104
rect 34743 34012 34823 34022
rect 34743 33956 34755 34012
rect 34811 33956 34823 34012
rect 34743 33946 34823 33956
rect 34927 34012 35007 34022
rect 34927 33956 34939 34012
rect 34995 33956 35007 34012
rect 34927 33946 35007 33956
rect 35111 34012 35191 34022
rect 35111 33956 35123 34012
rect 35179 33956 35191 34012
rect 35111 33946 35191 33956
rect 35256 33890 35324 34220
rect 35523 34212 35593 34222
rect 35215 33882 35324 33890
rect 35203 33880 35324 33882
rect 35203 33760 35215 33880
rect 35271 33760 35324 33880
rect 35203 33758 35324 33760
rect 35215 33750 35271 33758
rect 34518 33493 35414 33505
rect 34518 33437 34530 33493
rect 34586 33437 35348 33493
rect 35404 33437 35414 33493
rect 34518 33425 35414 33437
rect 35525 33268 35581 34212
rect 35689 33376 35769 33386
rect 35689 33320 35701 33376
rect 35757 33320 35769 33376
rect 35689 33318 35769 33320
rect 34213 33265 34283 33267
rect 34213 33209 34215 33265
rect 34271 33209 34283 33265
rect 34213 33197 34283 33209
rect 35513 33266 35593 33268
rect 35513 33210 35525 33266
rect 35581 33210 35593 33266
rect 35513 33198 35593 33210
rect 33177 33158 33923 33170
rect 33177 33102 33545 33158
rect 33601 33102 33923 33158
rect 33177 33090 33923 33102
rect 33177 32837 33233 33090
rect 33545 32837 33601 33090
rect 33867 32837 33923 33090
rect 34663 33159 35409 33171
rect 34663 33103 35031 33159
rect 35087 33103 35409 33159
rect 34663 33091 35409 33103
rect 34663 32838 34719 33091
rect 35031 32838 35087 33091
rect 35353 32838 35409 33091
rect 33165 32835 33245 32837
rect 33165 32715 33177 32835
rect 33233 32715 33245 32835
rect 33165 32713 33245 32715
rect 33533 32835 33613 32837
rect 33533 32715 33545 32835
rect 33601 32715 33613 32835
rect 33533 32713 33613 32715
rect 33855 32835 33935 32837
rect 33855 32714 33867 32835
rect 33923 32714 33935 32835
rect 34651 32836 34731 32838
rect 34651 32716 34663 32836
rect 34719 32716 34731 32836
rect 34651 32714 34731 32716
rect 35019 32836 35099 32838
rect 35019 32716 35031 32836
rect 35087 32716 35099 32836
rect 35019 32714 35099 32716
rect 35341 32836 35421 32838
rect 35341 32715 35353 32836
rect 35409 32715 35421 32836
rect 33177 32705 33233 32713
rect 33545 32705 33601 32713
rect 33855 32712 33935 32714
rect 33867 32704 33923 32712
rect 34663 32706 34719 32714
rect 35031 32706 35087 32714
rect 35341 32713 35421 32715
rect 35353 32705 35409 32713
rect 33361 32537 33417 32545
rect 33729 32537 33785 32545
rect 34847 32538 34903 32546
rect 35215 32538 35271 32546
rect 33349 32535 33838 32537
rect 33349 32415 33361 32535
rect 33417 32415 33729 32535
rect 33785 32415 33838 32535
rect 33349 32413 33838 32415
rect 34835 32536 35324 32538
rect 34835 32416 34847 32536
rect 34903 32416 35215 32536
rect 35271 32416 35324 32536
rect 34835 32414 35324 32416
rect 33361 32405 33417 32413
rect 33729 32405 33838 32413
rect 34847 32406 34903 32414
rect 35215 32406 35324 32414
rect 33257 32339 33337 32349
rect 33257 32283 33269 32339
rect 33325 32283 33337 32339
rect 33257 32273 33337 32283
rect 33441 32339 33521 32349
rect 33441 32283 33453 32339
rect 33509 32283 33521 32339
rect 33441 32273 33521 32283
rect 33625 32339 33705 32349
rect 33625 32283 33637 32339
rect 33693 32283 33705 32339
rect 33625 32273 33705 32283
rect 33269 32191 33325 32273
rect 33257 32189 33337 32191
rect 33257 32133 33269 32189
rect 33325 32133 33337 32189
rect 33257 32131 33337 32133
rect 32585 31957 32655 31969
rect 32585 31901 32597 31957
rect 32653 31901 32655 31957
rect 32585 31889 32655 31901
rect 33269 31817 33325 32131
rect 33453 32075 33509 32273
rect 33441 32073 33521 32075
rect 33441 32017 33453 32073
rect 33509 32017 33521 32073
rect 33441 32015 33521 32017
rect 33453 31817 33509 32015
rect 33637 31959 33693 32273
rect 33770 32075 33838 32405
rect 34743 32340 34823 32350
rect 34743 32284 34755 32340
rect 34811 32284 34823 32340
rect 34743 32274 34823 32284
rect 34927 32340 35007 32350
rect 34927 32284 34939 32340
rect 34995 32284 35007 32340
rect 34927 32274 35007 32284
rect 35111 32340 35191 32350
rect 35111 32284 35123 32340
rect 35179 32284 35191 32340
rect 35111 32274 35191 32284
rect 34755 32192 34811 32274
rect 34743 32190 34823 32192
rect 34743 32134 34755 32190
rect 34811 32134 34823 32190
rect 34743 32132 34823 32134
rect 33770 32073 33850 32075
rect 33770 32017 33782 32073
rect 33838 32017 33850 32073
rect 33770 32015 33850 32017
rect 34037 32073 34107 32085
rect 34037 32017 34039 32073
rect 34095 32017 34107 32073
rect 33625 31957 33705 31959
rect 33625 31901 33637 31957
rect 33693 31901 33705 31957
rect 33625 31899 33705 31901
rect 33637 31817 33693 31899
rect 33257 31807 33337 31817
rect 33257 31751 33269 31807
rect 33325 31751 33337 31807
rect 33257 31741 33337 31751
rect 33441 31807 33521 31817
rect 33441 31751 33453 31807
rect 33509 31751 33521 31807
rect 33441 31741 33521 31751
rect 33625 31807 33705 31817
rect 33625 31751 33637 31807
rect 33693 31751 33705 31807
rect 33625 31741 33705 31751
rect 33770 31685 33838 32015
rect 34037 32007 34107 32017
rect 33729 31677 33838 31685
rect 33717 31675 33838 31677
rect 33717 31555 33729 31675
rect 33785 31555 33838 31675
rect 33717 31553 33838 31555
rect 33729 31545 33785 31553
rect 33032 31288 33928 31300
rect 33032 31232 33044 31288
rect 33100 31232 33862 31288
rect 33918 31232 33928 31288
rect 33032 31220 33928 31232
rect 34039 31063 34095 32007
rect 34755 31818 34811 32132
rect 34939 32076 34995 32274
rect 34927 32074 35007 32076
rect 34927 32018 34939 32074
rect 34995 32018 35007 32074
rect 34927 32016 35007 32018
rect 34939 31818 34995 32016
rect 35123 31960 35179 32274
rect 35256 32076 35324 32406
rect 35701 32084 35757 33318
rect 35256 32074 35336 32076
rect 35256 32018 35268 32074
rect 35324 32018 35336 32074
rect 35256 32016 35336 32018
rect 35699 32074 35769 32084
rect 35699 32018 35701 32074
rect 35757 32018 35849 32074
rect 35111 31958 35191 31960
rect 35111 31902 35123 31958
rect 35179 31902 35191 31958
rect 35111 31900 35191 31902
rect 35123 31818 35179 31900
rect 34743 31808 34823 31818
rect 34743 31752 34755 31808
rect 34811 31752 34823 31808
rect 34743 31742 34823 31752
rect 34927 31808 35007 31818
rect 34927 31752 34939 31808
rect 34995 31752 35007 31808
rect 34927 31742 35007 31752
rect 35111 31808 35191 31818
rect 35111 31752 35123 31808
rect 35179 31752 35191 31808
rect 35111 31742 35191 31752
rect 35256 31686 35324 32016
rect 35699 32006 35769 32018
rect 35215 31678 35324 31686
rect 35203 31676 35324 31678
rect 35203 31556 35215 31676
rect 35271 31556 35324 31676
rect 35203 31554 35324 31556
rect 35215 31546 35271 31554
rect 34518 31289 35414 31301
rect 34518 31233 34530 31289
rect 34586 31233 35348 31289
rect 35404 31233 35414 31289
rect 34518 31221 35414 31233
rect 34203 31170 34283 31180
rect 34203 31114 34215 31170
rect 34271 31114 34283 31170
rect 34203 31112 34283 31114
rect 34037 31060 34107 31063
rect 34037 31006 34039 31060
rect 34095 31006 34107 31060
rect 34037 30994 34107 31006
rect 33177 30953 33923 30965
rect 33177 30897 33545 30953
rect 33601 30897 33923 30953
rect 33177 30885 33923 30897
rect 33177 30632 33233 30885
rect 33545 30632 33601 30885
rect 33867 30632 33923 30885
rect 33165 30630 33245 30632
rect 33165 30510 33177 30630
rect 33233 30510 33245 30630
rect 33165 30508 33245 30510
rect 33533 30630 33613 30632
rect 33533 30510 33545 30630
rect 33601 30510 33613 30630
rect 33533 30508 33613 30510
rect 33855 30630 33935 30632
rect 33855 30509 33867 30630
rect 33923 30509 33935 30630
rect 33177 30500 33233 30508
rect 33545 30500 33601 30508
rect 33855 30507 33935 30509
rect 33867 30499 33923 30507
rect 33361 30332 33417 30340
rect 33729 30332 33785 30340
rect 33349 30330 33838 30332
rect 33349 30210 33361 30330
rect 33417 30210 33729 30330
rect 33785 30210 33838 30330
rect 33349 30208 33838 30210
rect 33361 30200 33417 30208
rect 33729 30200 33838 30208
rect 33257 30134 33337 30144
rect 33257 30078 33269 30134
rect 33325 30078 33337 30134
rect 33257 30068 33337 30078
rect 33441 30134 33521 30144
rect 33441 30078 33453 30134
rect 33509 30078 33521 30134
rect 33441 30068 33521 30078
rect 33625 30134 33705 30144
rect 33625 30078 33637 30134
rect 33693 30078 33705 30134
rect 33625 30068 33705 30078
rect 33269 29986 33325 30068
rect 33257 29984 33337 29986
rect 33257 29928 33269 29984
rect 33325 29928 33337 29984
rect 33257 29926 33337 29928
rect 32449 29868 32519 29882
rect 32449 29812 32461 29868
rect 32517 29812 32519 29868
rect 32449 29800 32519 29812
rect 32215 29752 32293 29763
rect 31823 29751 32293 29752
rect 31823 29697 32227 29751
rect 32281 29697 32293 29751
rect 31823 29696 32293 29697
rect 30251 29392 31423 29402
rect 30251 29336 30263 29392
rect 30319 29336 31151 29392
rect 31207 29336 31423 29392
rect 30251 29326 31423 29336
rect 31823 29392 31903 29696
rect 32215 29685 32293 29696
rect 31823 29336 31835 29392
rect 31891 29336 31903 29392
rect 31823 29326 31903 29336
rect 30181 29014 31973 29026
rect 30181 28874 30193 29014
rect 31961 28874 31973 29014
rect 32266 28965 32352 28977
rect 32461 28969 32517 29800
rect 33269 29612 33325 29926
rect 33453 29870 33509 30068
rect 33441 29868 33521 29870
rect 33441 29812 33453 29868
rect 33509 29812 33521 29868
rect 33441 29810 33521 29812
rect 33453 29612 33509 29810
rect 33637 29754 33693 30068
rect 33770 29870 33838 30200
rect 34215 29880 34271 31112
rect 36223 31006 36279 34222
rect 41921 34222 41933 34278
rect 41989 34222 41991 34278
rect 41921 34210 41991 34222
rect 41639 33376 41721 33388
rect 41639 33320 41653 33376
rect 41709 33320 41721 33376
rect 41639 33308 41721 33320
rect 36633 31970 36853 31980
rect 36633 31170 36643 31970
rect 36843 31170 36853 31970
rect 41023 31970 41343 31980
rect 37495 31463 38667 31473
rect 37495 31223 37507 31463
rect 37563 31223 38599 31463
rect 38655 31223 38667 31463
rect 37495 31213 38667 31223
rect 36633 31160 36853 31170
rect 37589 31006 37667 31018
rect 36219 30950 37609 31006
rect 37665 30950 37667 31006
rect 37589 30938 37667 30950
rect 38587 30928 38667 31213
rect 39067 31463 39147 31473
rect 39067 31223 39079 31463
rect 39135 31223 39147 31463
rect 38889 30928 38959 30940
rect 38587 30872 38901 30928
rect 38957 30872 38959 30928
rect 38409 30850 38479 30862
rect 36219 30794 38421 30850
rect 38477 30794 38479 30850
rect 33770 29868 33850 29870
rect 33770 29812 33782 29868
rect 33838 29812 33850 29868
rect 33770 29810 33850 29812
rect 34213 29868 34273 29880
rect 34213 29812 34215 29868
rect 34271 29812 34273 29868
rect 33625 29752 33705 29754
rect 33625 29696 33637 29752
rect 33693 29696 33705 29752
rect 33625 29694 33705 29696
rect 33637 29612 33693 29694
rect 33257 29602 33337 29612
rect 33257 29546 33269 29602
rect 33325 29546 33337 29602
rect 33257 29536 33337 29546
rect 33441 29602 33521 29612
rect 33441 29546 33453 29602
rect 33509 29546 33521 29602
rect 33441 29536 33521 29546
rect 33625 29602 33705 29612
rect 33625 29546 33637 29602
rect 33693 29546 33705 29602
rect 33625 29536 33705 29546
rect 33770 29480 33838 29810
rect 34213 29800 34273 29812
rect 36331 29509 36387 30794
rect 38409 30782 38479 30794
rect 37699 30568 37779 30578
rect 37699 30512 37711 30568
rect 37767 30512 37779 30568
rect 37699 30326 37779 30512
rect 38179 30568 38259 30578
rect 38179 30512 38191 30568
rect 38247 30512 38259 30568
rect 38179 30502 38259 30512
rect 38383 30568 38463 30578
rect 38383 30512 38395 30568
rect 38451 30512 38463 30568
rect 38383 30326 38463 30512
rect 38587 30568 38667 30872
rect 38889 30860 38959 30872
rect 39067 30928 39147 31223
rect 41023 31170 41033 31970
rect 41333 31170 41343 31970
rect 41023 31160 41343 31170
rect 39653 30974 41445 30986
rect 39067 30872 39424 30928
rect 38587 30512 38599 30568
rect 38655 30512 38667 30568
rect 38587 30502 38667 30512
rect 39067 30568 39147 30872
rect 39067 30512 39079 30568
rect 39135 30512 39147 30568
rect 39067 30502 39147 30512
rect 37699 30254 38463 30326
rect 38593 30200 39217 30212
rect 38593 30060 38605 30200
rect 39205 30060 39217 30200
rect 36805 30043 36885 30053
rect 38593 30048 39217 30060
rect 36805 29803 36817 30043
rect 36873 29803 36885 30043
rect 39368 29830 39424 30872
rect 39653 30834 39665 30974
rect 41433 30834 41445 30974
rect 39653 30822 41445 30834
rect 39927 30571 40691 30581
rect 39927 30331 39939 30571
rect 39995 30331 40623 30571
rect 40679 30331 40691 30571
rect 39927 30321 40691 30331
rect 41295 30287 41375 30297
rect 40407 30237 40895 30247
rect 40407 29997 40419 30237
rect 40475 29997 40827 30237
rect 40883 29997 40895 30237
rect 40407 29987 40895 29997
rect 39817 29830 39913 29842
rect 33729 29472 33838 29480
rect 33717 29470 33838 29472
rect 33717 29350 33729 29470
rect 33785 29350 33838 29470
rect 35819 29508 36387 29509
rect 36627 29508 36697 29520
rect 35819 29453 36639 29508
rect 33717 29348 33838 29350
rect 33729 29340 33785 29348
rect 33032 29083 33930 29095
rect 33032 29027 33044 29083
rect 33100 29027 33862 29083
rect 33918 29027 33930 29083
rect 33032 29015 33930 29027
rect 32266 28909 32278 28965
rect 32334 28909 32352 28965
rect 32266 28897 32352 28909
rect 32459 28965 32519 28969
rect 32459 28909 32461 28965
rect 32517 28909 32519 28965
rect 32459 28897 32519 28909
rect 30181 28862 31973 28874
rect 29595 28532 29952 28588
rect 31551 28690 31871 28700
rect 29115 28172 29127 28228
rect 29183 28172 29195 28228
rect 29115 28162 29195 28172
rect 29595 28228 29675 28532
rect 29595 28172 29607 28228
rect 29663 28172 29675 28228
rect 29595 28162 29675 28172
rect 28227 27914 28991 27986
rect 31551 27890 31561 28690
rect 31861 27890 31871 28690
rect 31551 27880 31871 27890
rect 35824 27610 35880 29453
rect 36331 29452 36639 29453
rect 36695 29452 36697 29508
rect 36627 29440 36697 29452
rect 36805 29508 36885 29803
rect 38593 29800 39217 29812
rect 38593 29660 38605 29800
rect 39205 29660 39217 29800
rect 39368 29774 39837 29830
rect 39893 29774 39913 29830
rect 39817 29762 39913 29774
rect 40815 29752 40895 29987
rect 41295 30047 41307 30287
rect 41363 30047 41375 30287
rect 41117 29752 41187 29764
rect 40815 29696 41129 29752
rect 41185 29696 41187 29752
rect 40501 29674 40597 29684
rect 38593 29648 39217 29660
rect 39368 29618 40521 29674
rect 40577 29618 40597 29674
rect 36805 29452 37243 29508
rect 36805 29148 36885 29452
rect 36805 29092 36817 29148
rect 36873 29092 36885 29148
rect 36805 29082 36885 29092
rect 37187 28666 37243 29452
rect 37495 29123 38667 29133
rect 37495 28883 37507 29123
rect 37563 28883 38599 29123
rect 38655 28883 38667 29123
rect 37495 28873 38667 28883
rect 37589 28666 37667 28678
rect 37187 28610 37609 28666
rect 37665 28610 37667 28666
rect 37589 28598 37667 28610
rect 38587 28588 38667 28873
rect 39067 29123 39147 29133
rect 39067 28883 39079 29123
rect 39135 28883 39147 29123
rect 38889 28588 38959 28600
rect 38587 28532 38901 28588
rect 38957 28532 38959 28588
rect 38409 28510 38479 28522
rect 35824 27480 35880 27490
rect 36219 28454 38421 28510
rect 38477 28454 38479 28510
rect 11153 26758 26803 26814
rect 7109 26074 7179 26076
rect 7109 26018 7111 26074
rect 7167 26018 7179 26074
rect 7109 26016 7179 26018
rect 3293 25898 3363 25910
rect 3293 25842 3305 25898
rect 3361 25842 3363 25898
rect 3293 25840 3363 25842
rect 3067 25546 3137 25548
rect 3067 25490 3069 25546
rect 3125 25490 3137 25546
rect 3067 25488 3137 25490
rect 115 25262 861 25274
rect 115 25206 483 25262
rect 539 25206 861 25262
rect 115 25194 861 25206
rect 115 24941 171 25194
rect 483 24941 539 25194
rect 805 24941 861 25194
rect 103 24939 183 24941
rect 103 24819 115 24939
rect 171 24819 183 24939
rect 103 24817 183 24819
rect 471 24939 551 24941
rect 471 24819 483 24939
rect 539 24819 551 24939
rect 471 24817 551 24819
rect 793 24939 873 24941
rect 793 24818 805 24939
rect 861 24818 873 24939
rect 115 24809 171 24817
rect 483 24809 539 24817
rect 793 24816 873 24818
rect 805 24808 861 24816
rect 299 24641 355 24649
rect 667 24641 723 24649
rect 287 24639 776 24641
rect 287 24519 299 24639
rect 355 24519 667 24639
rect 723 24519 776 24639
rect 287 24517 776 24519
rect 299 24509 355 24517
rect 667 24509 776 24517
rect 195 24443 275 24453
rect 195 24387 207 24443
rect 263 24387 275 24443
rect 195 24377 275 24387
rect 379 24443 459 24453
rect 379 24387 391 24443
rect 447 24387 459 24443
rect 379 24377 459 24387
rect 563 24443 643 24453
rect 563 24387 575 24443
rect 631 24387 643 24443
rect 563 24377 643 24387
rect 207 24295 263 24377
rect 195 24293 275 24295
rect 195 24237 207 24293
rect 263 24237 275 24293
rect 195 24235 275 24237
rect -477 24177 -407 24189
rect -477 24121 -465 24177
rect -409 24121 -407 24177
rect -477 24109 -407 24121
rect -613 21972 -543 21986
rect -613 21916 -601 21972
rect -545 21916 -543 21972
rect -613 21904 -543 21916
rect -749 21070 -679 21072
rect -749 21014 -737 21070
rect -681 21014 -679 21070
rect -749 21002 -679 21014
rect -601 17576 -545 21904
rect -465 19663 -409 24109
rect 207 23921 263 24235
rect 391 24179 447 24377
rect 379 24177 459 24179
rect 379 24121 391 24177
rect 447 24121 459 24177
rect 379 24119 459 24121
rect 391 23921 447 24119
rect 575 24063 631 24377
rect 708 24179 776 24509
rect 2855 24293 2925 24305
rect 2855 24237 2867 24293
rect 2923 24237 2925 24293
rect 2855 24235 2925 24237
rect 708 24177 788 24179
rect 708 24121 720 24177
rect 776 24121 788 24177
rect 708 24119 788 24121
rect 975 24177 1045 24189
rect 975 24121 977 24177
rect 1033 24121 1045 24177
rect 563 24061 643 24063
rect 563 24005 575 24061
rect 631 24005 643 24061
rect 563 24003 643 24005
rect 575 23921 631 24003
rect 195 23911 275 23921
rect 195 23855 207 23911
rect 263 23855 275 23911
rect 195 23845 275 23855
rect 379 23911 459 23921
rect 379 23855 391 23911
rect 447 23855 459 23911
rect 379 23845 459 23855
rect 563 23911 643 23921
rect 563 23855 575 23911
rect 631 23855 643 23911
rect 563 23845 643 23855
rect 708 23789 776 24119
rect 975 24111 1045 24121
rect 667 23781 776 23789
rect 655 23779 776 23781
rect 655 23659 667 23779
rect 723 23659 776 23779
rect 655 23657 776 23659
rect 667 23649 723 23657
rect -30 23392 868 23404
rect -30 23336 -18 23392
rect 38 23336 800 23392
rect 856 23336 868 23392
rect -30 23324 868 23336
rect 977 23167 1033 24111
rect 1141 23274 1221 23284
rect 1141 23218 1153 23274
rect 1209 23218 1221 23274
rect 1141 23216 1221 23218
rect 975 23164 1045 23167
rect 975 23110 977 23164
rect 1033 23110 1045 23164
rect 975 23098 1045 23110
rect 115 23057 861 23069
rect 115 23001 483 23057
rect 539 23001 861 23057
rect 115 22989 861 23001
rect 115 22736 171 22989
rect 483 22736 539 22989
rect 805 22736 861 22989
rect 103 22734 183 22736
rect 103 22614 115 22734
rect 171 22614 183 22734
rect 103 22612 183 22614
rect 471 22734 551 22736
rect 471 22614 483 22734
rect 539 22614 551 22734
rect 471 22612 551 22614
rect 793 22734 873 22736
rect 793 22613 805 22734
rect 861 22613 873 22734
rect 115 22604 171 22612
rect 483 22604 539 22612
rect 793 22611 873 22613
rect 805 22603 861 22611
rect 299 22436 355 22444
rect 667 22436 723 22444
rect 287 22434 776 22436
rect 287 22314 299 22434
rect 355 22314 667 22434
rect 723 22314 776 22434
rect 287 22312 776 22314
rect 299 22304 355 22312
rect 667 22304 776 22312
rect 195 22238 275 22248
rect 195 22182 207 22238
rect 263 22182 275 22238
rect 195 22172 275 22182
rect 379 22238 459 22248
rect 379 22182 391 22238
rect 447 22182 459 22238
rect 379 22172 459 22182
rect 563 22238 643 22248
rect 563 22182 575 22238
rect 631 22182 643 22238
rect 563 22172 643 22182
rect 207 22090 263 22172
rect 195 22088 275 22090
rect 195 22032 207 22088
rect 263 22032 275 22088
rect 195 22030 275 22032
rect 207 21716 263 22030
rect 391 21974 447 22172
rect 379 21972 459 21974
rect 379 21916 391 21972
rect 447 21916 459 21972
rect 379 21914 459 21916
rect 391 21716 447 21914
rect 575 21858 631 22172
rect 708 21974 776 22304
rect 1153 21982 1209 23216
rect 1601 23057 2347 23069
rect 1601 23001 1969 23057
rect 2025 23001 2347 23057
rect 1601 22989 2347 23001
rect 1601 22736 1657 22989
rect 1969 22736 2025 22989
rect 2291 22736 2347 22989
rect 1589 22734 1669 22736
rect 1589 22614 1601 22734
rect 1657 22614 1669 22734
rect 1589 22612 1669 22614
rect 1957 22734 2037 22736
rect 1957 22614 1969 22734
rect 2025 22614 2037 22734
rect 1957 22612 2037 22614
rect 2279 22734 2359 22736
rect 2279 22613 2291 22734
rect 2347 22613 2359 22734
rect 1601 22604 1657 22612
rect 1969 22604 2025 22612
rect 2279 22611 2359 22613
rect 2291 22603 2347 22611
rect 1785 22436 1841 22444
rect 2153 22436 2209 22444
rect 1773 22434 2262 22436
rect 1773 22314 1785 22434
rect 1841 22314 2153 22434
rect 2209 22314 2262 22434
rect 1773 22312 2262 22314
rect 1785 22304 1841 22312
rect 2153 22304 2262 22312
rect 1681 22238 1761 22248
rect 1681 22182 1693 22238
rect 1749 22182 1761 22238
rect 1681 22172 1761 22182
rect 1865 22238 1945 22248
rect 1865 22182 1877 22238
rect 1933 22182 1945 22238
rect 1865 22172 1945 22182
rect 2049 22238 2129 22248
rect 2049 22182 2061 22238
rect 2117 22182 2129 22238
rect 2049 22172 2129 22182
rect 1693 22090 1749 22172
rect 1681 22088 1761 22090
rect 1681 22032 1693 22088
rect 1749 22032 1761 22088
rect 1681 22030 1761 22032
rect 708 21972 788 21974
rect 708 21916 720 21972
rect 776 21916 788 21972
rect 708 21914 788 21916
rect 1151 21972 1211 21982
rect 1151 21916 1153 21972
rect 1209 21916 1211 21972
rect 563 21856 643 21858
rect 563 21800 575 21856
rect 631 21800 643 21856
rect 563 21798 643 21800
rect 575 21716 631 21798
rect 195 21706 275 21716
rect 195 21650 207 21706
rect 263 21650 275 21706
rect 195 21640 275 21650
rect 379 21706 459 21716
rect 379 21650 391 21706
rect 447 21650 459 21706
rect 379 21640 459 21650
rect 563 21706 643 21716
rect 563 21650 575 21706
rect 631 21650 643 21706
rect 563 21640 643 21650
rect 708 21584 776 21914
rect 1151 21904 1211 21916
rect 667 21576 776 21584
rect 655 21574 776 21576
rect 655 21454 667 21574
rect 723 21454 776 21574
rect 655 21452 776 21454
rect 667 21444 723 21452
rect -30 21187 866 21199
rect -30 21131 -18 21187
rect 38 21131 800 21187
rect 856 21131 866 21187
rect -30 21119 866 21131
rect 1153 20961 1209 21904
rect 1693 21716 1749 22030
rect 1877 21974 1933 22172
rect 1865 21972 1945 21974
rect 1865 21916 1877 21972
rect 1933 21916 1945 21972
rect 1865 21914 1945 21916
rect 1877 21716 1933 21914
rect 2061 21858 2117 22172
rect 2194 21974 2262 22304
rect 2194 21972 2274 21974
rect 2194 21916 2206 21972
rect 2262 21916 2274 21972
rect 2194 21914 2274 21916
rect 2461 21972 2531 21984
rect 2461 21916 2463 21972
rect 2519 21916 2787 21972
rect 2049 21856 2129 21858
rect 2049 21800 2061 21856
rect 2117 21800 2129 21856
rect 2049 21798 2129 21800
rect 2061 21716 2117 21798
rect 1681 21706 1761 21716
rect 1681 21650 1693 21706
rect 1749 21650 1761 21706
rect 1681 21640 1761 21650
rect 1865 21706 1945 21716
rect 1865 21650 1877 21706
rect 1933 21650 1945 21706
rect 1865 21640 1945 21650
rect 2049 21706 2129 21716
rect 2049 21650 2061 21706
rect 2117 21650 2129 21706
rect 2049 21640 2129 21650
rect 2194 21584 2262 21914
rect 2461 21906 2531 21916
rect 2153 21576 2262 21584
rect 2141 21574 2262 21576
rect 2141 21454 2153 21574
rect 2209 21454 2262 21574
rect 2141 21452 2262 21454
rect 2153 21444 2209 21452
rect 1456 21187 2352 21199
rect 1456 21131 1468 21187
rect 1524 21131 2286 21187
rect 2342 21131 2352 21187
rect 1456 21119 2352 21131
rect 2463 20962 2519 21906
rect 2627 21070 2707 21080
rect 2627 21014 2639 21070
rect 2695 21014 2707 21070
rect 2627 21012 2707 21014
rect 1151 20959 1221 20961
rect 1151 20903 1153 20959
rect 1209 20903 1221 20959
rect 1151 20891 1221 20903
rect 2451 20960 2531 20962
rect 2451 20904 2463 20960
rect 2519 20904 2531 20960
rect 2451 20892 2531 20904
rect 115 20852 861 20864
rect 115 20796 483 20852
rect 539 20796 861 20852
rect 115 20784 861 20796
rect 115 20531 171 20784
rect 483 20531 539 20784
rect 805 20531 861 20784
rect 1601 20853 2347 20865
rect 1601 20797 1969 20853
rect 2025 20797 2347 20853
rect 1601 20785 2347 20797
rect 1601 20532 1657 20785
rect 1969 20532 2025 20785
rect 2291 20532 2347 20785
rect 103 20529 183 20531
rect 103 20409 115 20529
rect 171 20409 183 20529
rect 103 20407 183 20409
rect 471 20529 551 20531
rect 471 20409 483 20529
rect 539 20409 551 20529
rect 471 20407 551 20409
rect 793 20529 873 20531
rect 793 20408 805 20529
rect 861 20408 873 20529
rect 1589 20530 1669 20532
rect 1589 20410 1601 20530
rect 1657 20410 1669 20530
rect 1589 20408 1669 20410
rect 1957 20530 2037 20532
rect 1957 20410 1969 20530
rect 2025 20410 2037 20530
rect 1957 20408 2037 20410
rect 2279 20530 2359 20532
rect 2279 20409 2291 20530
rect 2347 20409 2359 20530
rect 115 20399 171 20407
rect 483 20399 539 20407
rect 793 20406 873 20408
rect 805 20398 861 20406
rect 1601 20400 1657 20408
rect 1969 20400 2025 20408
rect 2279 20407 2359 20409
rect 2291 20399 2347 20407
rect 299 20231 355 20239
rect 667 20231 723 20239
rect 1785 20232 1841 20240
rect 2153 20232 2209 20240
rect 287 20229 776 20231
rect 287 20109 299 20229
rect 355 20109 667 20229
rect 723 20109 776 20229
rect 287 20107 776 20109
rect 1773 20230 2262 20232
rect 1773 20110 1785 20230
rect 1841 20110 2153 20230
rect 2209 20110 2262 20230
rect 1773 20108 2262 20110
rect 299 20099 355 20107
rect 667 20099 776 20107
rect 1785 20100 1841 20108
rect 2153 20100 2262 20108
rect 195 20033 275 20043
rect 195 19977 207 20033
rect 263 19977 275 20033
rect 195 19967 275 19977
rect 379 20033 459 20043
rect 379 19977 391 20033
rect 447 19977 459 20033
rect 379 19967 459 19977
rect 563 20033 643 20043
rect 563 19977 575 20033
rect 631 19977 643 20033
rect 563 19967 643 19977
rect 207 19885 263 19967
rect 195 19883 275 19885
rect 195 19827 207 19883
rect 263 19827 275 19883
rect 195 19825 275 19827
rect -477 19651 -407 19663
rect -477 19595 -465 19651
rect -409 19595 -407 19651
rect -477 19583 -407 19595
rect 207 19511 263 19825
rect 391 19769 447 19967
rect 379 19767 459 19769
rect 379 19711 391 19767
rect 447 19711 459 19767
rect 379 19709 459 19711
rect 391 19511 447 19709
rect 575 19653 631 19967
rect 708 19769 776 20099
rect 1681 20034 1761 20044
rect 1681 19978 1693 20034
rect 1749 19978 1761 20034
rect 1681 19968 1761 19978
rect 1865 20034 1945 20044
rect 1865 19978 1877 20034
rect 1933 19978 1945 20034
rect 1865 19968 1945 19978
rect 2049 20034 2129 20044
rect 2049 19978 2061 20034
rect 2117 19978 2129 20034
rect 2049 19968 2129 19978
rect 1693 19886 1749 19968
rect 1681 19884 1761 19886
rect 1681 19828 1693 19884
rect 1749 19828 1761 19884
rect 1681 19826 1761 19828
rect 708 19767 788 19769
rect 708 19711 720 19767
rect 776 19711 788 19767
rect 708 19709 788 19711
rect 975 19767 1045 19779
rect 975 19711 977 19767
rect 1033 19711 1045 19767
rect 563 19651 643 19653
rect 563 19595 575 19651
rect 631 19595 643 19651
rect 563 19593 643 19595
rect 575 19511 631 19593
rect 195 19501 275 19511
rect 195 19445 207 19501
rect 263 19445 275 19501
rect 195 19435 275 19445
rect 379 19501 459 19511
rect 379 19445 391 19501
rect 447 19445 459 19501
rect 379 19435 459 19445
rect 563 19501 643 19511
rect 563 19445 575 19501
rect 631 19445 643 19501
rect 563 19435 643 19445
rect 708 19379 776 19709
rect 975 19701 1045 19711
rect 667 19371 776 19379
rect 655 19369 776 19371
rect 655 19249 667 19369
rect 723 19249 776 19369
rect 655 19247 776 19249
rect 667 19239 723 19247
rect -30 18982 866 18994
rect -30 18926 -18 18982
rect 38 18926 800 18982
rect 856 18926 866 18982
rect -30 18914 866 18926
rect 977 18757 1033 19701
rect 1693 19512 1749 19826
rect 1877 19770 1933 19968
rect 1865 19768 1945 19770
rect 1865 19712 1877 19768
rect 1933 19712 1945 19768
rect 1865 19710 1945 19712
rect 1877 19512 1933 19710
rect 2061 19654 2117 19968
rect 2194 19770 2262 20100
rect 2639 19778 2695 21012
rect 2194 19768 2274 19770
rect 2194 19712 2206 19768
rect 2262 19712 2274 19768
rect 2194 19710 2274 19712
rect 2637 19768 2707 19778
rect 2637 19712 2639 19768
rect 2695 19712 2787 19768
rect 2049 19652 2129 19654
rect 2049 19596 2061 19652
rect 2117 19596 2129 19652
rect 2049 19594 2129 19596
rect 2061 19512 2117 19594
rect 1681 19502 1761 19512
rect 1681 19446 1693 19502
rect 1749 19446 1761 19502
rect 1681 19436 1761 19446
rect 1865 19502 1945 19512
rect 1865 19446 1877 19502
rect 1933 19446 1945 19502
rect 1865 19436 1945 19446
rect 2049 19502 2129 19512
rect 2049 19446 2061 19502
rect 2117 19446 2129 19502
rect 2049 19436 2129 19446
rect 2194 19380 2262 19710
rect 2637 19700 2707 19712
rect 2153 19372 2262 19380
rect 2141 19370 2262 19372
rect 2141 19250 2153 19370
rect 2209 19250 2262 19370
rect 2141 19248 2262 19250
rect 2153 19240 2209 19248
rect 1456 18983 2352 18995
rect 1456 18927 1468 18983
rect 1524 18927 2286 18983
rect 2342 18927 2352 18983
rect 1456 18915 2352 18927
rect 1141 18864 1221 18874
rect 1141 18808 1153 18864
rect 1209 18808 1221 18864
rect 1141 18806 1221 18808
rect 975 18754 1045 18757
rect 975 18700 977 18754
rect 1033 18700 1045 18754
rect 975 18688 1045 18700
rect 115 18647 861 18659
rect 115 18591 483 18647
rect 539 18591 861 18647
rect 115 18579 861 18591
rect 115 18326 171 18579
rect 483 18326 539 18579
rect 805 18326 861 18579
rect 103 18324 183 18326
rect 103 18204 115 18324
rect 171 18204 183 18324
rect 103 18202 183 18204
rect 471 18324 551 18326
rect 471 18204 483 18324
rect 539 18204 551 18324
rect 471 18202 551 18204
rect 793 18324 873 18326
rect 793 18203 805 18324
rect 861 18203 873 18324
rect 115 18194 171 18202
rect 483 18194 539 18202
rect 793 18201 873 18203
rect 805 18193 861 18201
rect 299 18026 355 18034
rect 667 18026 723 18034
rect 287 18024 776 18026
rect 287 17904 299 18024
rect 355 17904 667 18024
rect 723 17904 776 18024
rect 287 17902 776 17904
rect 299 17894 355 17902
rect 667 17894 776 17902
rect 195 17828 275 17838
rect 195 17772 207 17828
rect 263 17772 275 17828
rect 195 17762 275 17772
rect 379 17828 459 17838
rect 379 17772 391 17828
rect 447 17772 459 17828
rect 379 17762 459 17772
rect 563 17828 643 17838
rect 563 17772 575 17828
rect 631 17772 643 17828
rect 563 17762 643 17772
rect 207 17680 263 17762
rect 195 17678 275 17680
rect 195 17622 207 17678
rect 263 17622 275 17678
rect 195 17620 275 17622
rect -613 17562 -543 17576
rect -613 17506 -601 17562
rect -545 17506 -543 17562
rect -613 17494 -543 17506
rect -915 16659 -845 16671
rect -601 16663 -545 17494
rect 207 17306 263 17620
rect 391 17564 447 17762
rect 379 17562 459 17564
rect 379 17506 391 17562
rect 447 17506 459 17562
rect 379 17504 459 17506
rect 391 17306 447 17504
rect 575 17448 631 17762
rect 708 17564 776 17894
rect 1153 17574 1209 18806
rect 708 17562 788 17564
rect 708 17506 720 17562
rect 776 17506 788 17562
rect 708 17504 788 17506
rect 1151 17562 1211 17574
rect 1151 17506 1153 17562
rect 1209 17506 1211 17562
rect 563 17446 643 17448
rect 563 17390 575 17446
rect 631 17390 643 17446
rect 563 17388 643 17390
rect 575 17306 631 17388
rect 195 17296 275 17306
rect 195 17240 207 17296
rect 263 17240 275 17296
rect 195 17230 275 17240
rect 379 17296 459 17306
rect 379 17240 391 17296
rect 447 17240 459 17296
rect 379 17230 459 17240
rect 563 17296 643 17306
rect 563 17240 575 17296
rect 631 17240 643 17296
rect 563 17230 643 17240
rect 708 17174 776 17504
rect 1151 17494 1211 17506
rect 2583 17446 2653 17458
rect 2583 17390 2595 17446
rect 2651 17390 2653 17446
rect 2583 17378 2653 17390
rect 667 17166 776 17174
rect 655 17164 776 17166
rect 655 17044 667 17164
rect 723 17044 776 17164
rect 655 17042 776 17044
rect 667 17034 723 17042
rect -30 16777 868 16789
rect -30 16721 -18 16777
rect 38 16721 800 16777
rect 856 16721 868 16777
rect -30 16709 868 16721
rect -915 16603 -903 16659
rect -847 16603 -845 16659
rect -915 16601 -845 16603
rect -603 16659 -543 16663
rect -603 16603 -601 16659
rect -545 16603 -543 16659
rect -903 15989 -847 16601
rect -603 16591 -543 16603
rect 2595 16499 2651 17378
rect 2595 16389 2651 16399
rect -1051 11494 -981 11506
rect -1051 11438 -1039 11494
rect -983 11438 -981 11494
rect -1051 11426 -981 11438
rect -1405 10136 -1403 10192
rect -1347 10136 -1119 10192
rect -1993 10076 -1913 10078
rect -1993 10020 -1981 10076
rect -1925 10020 -1913 10076
rect -1993 10018 -1913 10020
rect -1981 9936 -1925 10018
rect -2361 9926 -2281 9936
rect -2361 9870 -2349 9926
rect -2293 9870 -2281 9926
rect -2361 9860 -2281 9870
rect -2177 9926 -2097 9936
rect -2177 9870 -2165 9926
rect -2109 9870 -2097 9926
rect -2177 9860 -2097 9870
rect -1993 9926 -1913 9936
rect -1993 9870 -1981 9926
rect -1925 9870 -1913 9926
rect -1993 9860 -1913 9870
rect -1848 9804 -1780 10134
rect -1405 10124 -1335 10136
rect -1889 9796 -1780 9804
rect -1901 9794 -1780 9796
rect -1901 9674 -1889 9794
rect -1833 9674 -1780 9794
rect -1901 9672 -1780 9674
rect -1889 9664 -1833 9672
rect -2586 9407 -1690 9419
rect -2586 9351 -2574 9407
rect -2518 9351 -1756 9407
rect -1700 9351 -1690 9407
rect -2586 9339 -1690 9351
rect -2901 9288 -2821 9298
rect -2901 9232 -2889 9288
rect -2833 9232 -2821 9288
rect -2901 9230 -2821 9232
rect -3067 9178 -2997 9181
rect -3067 9124 -3065 9178
rect -3009 9124 -2997 9178
rect -3067 9112 -2997 9124
rect -3927 9071 -3181 9083
rect -3927 9015 -3559 9071
rect -3503 9015 -3181 9071
rect -3927 9003 -3181 9015
rect -3927 8750 -3871 9003
rect -3559 8750 -3503 9003
rect -3237 8750 -3181 9003
rect -3939 8748 -3859 8750
rect -3939 8628 -3927 8748
rect -3871 8628 -3859 8748
rect -3939 8626 -3859 8628
rect -3571 8748 -3491 8750
rect -3571 8628 -3559 8748
rect -3503 8628 -3491 8748
rect -3571 8626 -3491 8628
rect -3249 8748 -3169 8750
rect -3249 8627 -3237 8748
rect -3181 8627 -3169 8748
rect -3927 8618 -3871 8626
rect -3559 8618 -3503 8626
rect -3249 8625 -3169 8627
rect -3237 8617 -3181 8625
rect -3743 8450 -3687 8458
rect -3375 8450 -3319 8458
rect -3755 8448 -3266 8450
rect -3755 8328 -3743 8448
rect -3687 8328 -3375 8448
rect -3319 8328 -3266 8448
rect -3755 8326 -3266 8328
rect -3743 8318 -3687 8326
rect -3375 8318 -3266 8326
rect -3847 8252 -3767 8262
rect -3847 8196 -3835 8252
rect -3779 8196 -3767 8252
rect -3847 8186 -3767 8196
rect -3663 8252 -3583 8262
rect -3663 8196 -3651 8252
rect -3595 8196 -3583 8252
rect -3663 8186 -3583 8196
rect -3479 8252 -3399 8262
rect -3479 8196 -3467 8252
rect -3411 8196 -3399 8252
rect -3479 8186 -3399 8196
rect -3835 8104 -3779 8186
rect -3847 8102 -3767 8104
rect -3847 8046 -3835 8102
rect -3779 8046 -3767 8102
rect -3847 8044 -3767 8046
rect -4655 7986 -4585 8000
rect -4655 7930 -4643 7986
rect -4587 7930 -4585 7986
rect -4655 7918 -4585 7930
rect -4821 7870 -4741 7882
rect -4821 7814 -4809 7870
rect -4753 7814 -4741 7870
rect -4821 7802 -4741 7814
rect -4957 7083 -4887 7095
rect -4643 7087 -4587 7918
rect -3835 7730 -3779 8044
rect -3651 7988 -3595 8186
rect -3663 7986 -3583 7988
rect -3663 7930 -3651 7986
rect -3595 7930 -3583 7986
rect -3663 7928 -3583 7930
rect -3651 7730 -3595 7928
rect -3467 7872 -3411 8186
rect -3334 7988 -3266 8318
rect -2889 7998 -2833 9230
rect -3334 7986 -3254 7988
rect -3334 7930 -3322 7986
rect -3266 7930 -3254 7986
rect -3334 7928 -3254 7930
rect -2891 7986 -2831 7998
rect -2891 7930 -2889 7986
rect -2833 7930 -2831 7986
rect -3479 7870 -3399 7872
rect -3479 7814 -3467 7870
rect -3411 7814 -3399 7870
rect -3479 7812 -3399 7814
rect -3467 7730 -3411 7812
rect -3847 7720 -3767 7730
rect -3847 7664 -3835 7720
rect -3779 7664 -3767 7720
rect -3847 7654 -3767 7664
rect -3663 7720 -3583 7730
rect -3663 7664 -3651 7720
rect -3595 7664 -3583 7720
rect -3663 7654 -3583 7664
rect -3479 7720 -3399 7730
rect -3479 7664 -3467 7720
rect -3411 7664 -3399 7720
rect -3479 7654 -3399 7664
rect -3334 7598 -3266 7928
rect -2891 7918 -2831 7930
rect -3375 7590 -3266 7598
rect -3387 7588 -3266 7590
rect -3387 7468 -3375 7588
rect -3319 7468 -3266 7588
rect -3387 7466 -3266 7468
rect -3375 7458 -3319 7466
rect -4072 7201 -3174 7213
rect -4072 7145 -4060 7201
rect -4004 7145 -3242 7201
rect -3186 7145 -3174 7201
rect -4072 7133 -3174 7145
rect -4957 7027 -4945 7083
rect -4889 7027 -4887 7083
rect -4957 7015 -4887 7027
rect -4645 7083 -4585 7087
rect -4645 7027 -4643 7083
rect -4587 7027 -4585 7083
rect -4645 7015 -4585 7027
rect -5081 6810 -5025 6820
rect -1039 6920 -983 11426
rect -903 7095 -847 15889
rect 115 15686 861 15698
rect 115 15630 483 15686
rect 539 15630 861 15686
rect 115 15618 861 15630
rect 115 15365 171 15618
rect 483 15365 539 15618
rect 805 15365 861 15618
rect 103 15363 183 15365
rect 103 15243 115 15363
rect 171 15243 183 15363
rect 103 15241 183 15243
rect 471 15363 551 15365
rect 471 15243 483 15363
rect 539 15243 551 15363
rect 471 15241 551 15243
rect 793 15363 873 15365
rect 793 15242 805 15363
rect 861 15242 873 15363
rect 115 15233 171 15241
rect 483 15233 539 15241
rect 793 15240 873 15242
rect 805 15232 861 15240
rect 299 15065 355 15073
rect 667 15065 723 15073
rect 287 15063 776 15065
rect 287 14943 299 15063
rect 355 14943 667 15063
rect 723 14943 776 15063
rect 287 14941 776 14943
rect 299 14933 355 14941
rect 667 14933 776 14941
rect 195 14867 275 14877
rect 195 14811 207 14867
rect 263 14811 275 14867
rect 195 14801 275 14811
rect 379 14867 459 14877
rect 379 14811 391 14867
rect 447 14811 459 14867
rect 379 14801 459 14811
rect 563 14867 643 14877
rect 563 14811 575 14867
rect 631 14811 643 14867
rect 563 14801 643 14811
rect -693 14717 -607 14729
rect 207 14719 263 14801
rect -693 14661 -681 14717
rect -625 14661 -607 14717
rect -693 14649 -607 14661
rect 195 14717 275 14719
rect 195 14661 207 14717
rect 263 14661 275 14717
rect 195 14659 275 14661
rect -477 14601 -407 14613
rect -477 14545 -465 14601
rect -409 14545 -407 14601
rect -477 14533 -407 14545
rect -613 12396 -543 12410
rect -613 12340 -601 12396
rect -545 12340 -543 12396
rect -613 12328 -543 12340
rect -779 12208 -699 12218
rect -779 12152 -767 12208
rect -711 12152 -699 12208
rect -779 12150 -699 12152
rect -767 7882 -711 12150
rect -601 8000 -545 12328
rect -465 10087 -409 14533
rect 207 14345 263 14659
rect 391 14603 447 14801
rect 379 14601 459 14603
rect 379 14545 391 14601
rect 447 14545 459 14601
rect 379 14543 459 14545
rect 391 14345 447 14543
rect 575 14487 631 14801
rect 708 14603 776 14933
rect 708 14601 788 14603
rect 708 14545 720 14601
rect 776 14545 788 14601
rect 708 14543 788 14545
rect 975 14601 1045 14613
rect 975 14545 977 14601
rect 1033 14545 1045 14601
rect 563 14485 643 14487
rect 563 14429 575 14485
rect 631 14429 643 14485
rect 563 14427 643 14429
rect 575 14345 631 14427
rect 195 14335 275 14345
rect 195 14279 207 14335
rect 263 14279 275 14335
rect 195 14269 275 14279
rect 379 14335 459 14345
rect 379 14279 391 14335
rect 447 14279 459 14335
rect 379 14269 459 14279
rect 563 14335 643 14345
rect 563 14279 575 14335
rect 631 14279 643 14335
rect 563 14269 643 14279
rect 708 14213 776 14543
rect 975 14535 1045 14545
rect 667 14205 776 14213
rect 655 14203 776 14205
rect 655 14083 667 14203
rect 723 14083 776 14203
rect 655 14081 776 14083
rect 667 14073 723 14081
rect -30 13816 868 13828
rect -30 13760 -18 13816
rect 38 13760 800 13816
rect 856 13760 868 13816
rect -30 13748 868 13760
rect 977 13591 1033 14535
rect 1141 13698 1221 13708
rect 1141 13642 1153 13698
rect 1209 13642 1221 13698
rect 1141 13640 1221 13642
rect 975 13588 1045 13591
rect 975 13534 977 13588
rect 1033 13534 1045 13588
rect 975 13522 1045 13534
rect 115 13481 861 13493
rect 115 13425 483 13481
rect 539 13425 861 13481
rect 115 13413 861 13425
rect 115 13160 171 13413
rect 483 13160 539 13413
rect 805 13160 861 13413
rect 103 13158 183 13160
rect 103 13038 115 13158
rect 171 13038 183 13158
rect 103 13036 183 13038
rect 471 13158 551 13160
rect 471 13038 483 13158
rect 539 13038 551 13158
rect 471 13036 551 13038
rect 793 13158 873 13160
rect 793 13037 805 13158
rect 861 13037 873 13158
rect 115 13028 171 13036
rect 483 13028 539 13036
rect 793 13035 873 13037
rect 805 13027 861 13035
rect 299 12860 355 12868
rect 667 12860 723 12868
rect 287 12858 776 12860
rect 287 12738 299 12858
rect 355 12738 667 12858
rect 723 12738 776 12858
rect 287 12736 776 12738
rect 299 12728 355 12736
rect 667 12728 776 12736
rect 195 12662 275 12672
rect 195 12606 207 12662
rect 263 12606 275 12662
rect 195 12596 275 12606
rect 379 12662 459 12672
rect 379 12606 391 12662
rect 447 12606 459 12662
rect 379 12596 459 12606
rect 563 12662 643 12672
rect 563 12606 575 12662
rect 631 12606 643 12662
rect 563 12596 643 12606
rect 207 12514 263 12596
rect 195 12512 275 12514
rect 195 12456 207 12512
rect 263 12456 275 12512
rect 195 12454 275 12456
rect 207 12140 263 12454
rect 391 12398 447 12596
rect 379 12396 459 12398
rect 379 12340 391 12396
rect 447 12340 459 12396
rect 379 12338 459 12340
rect 391 12140 447 12338
rect 575 12282 631 12596
rect 708 12398 776 12728
rect 1153 12406 1209 13640
rect 1601 13481 2347 13493
rect 1601 13425 1969 13481
rect 2025 13425 2347 13481
rect 1601 13413 2347 13425
rect 1601 13160 1657 13413
rect 1969 13160 2025 13413
rect 2291 13160 2347 13413
rect 1589 13158 1669 13160
rect 1589 13038 1601 13158
rect 1657 13038 1669 13158
rect 1589 13036 1669 13038
rect 1957 13158 2037 13160
rect 1957 13038 1969 13158
rect 2025 13038 2037 13158
rect 1957 13036 2037 13038
rect 2279 13158 2359 13160
rect 2279 13037 2291 13158
rect 2347 13037 2359 13158
rect 1601 13028 1657 13036
rect 1969 13028 2025 13036
rect 2279 13035 2359 13037
rect 2291 13027 2347 13035
rect 1785 12860 1841 12868
rect 2153 12860 2209 12868
rect 1773 12858 2262 12860
rect 1773 12738 1785 12858
rect 1841 12738 2153 12858
rect 2209 12738 2262 12858
rect 1773 12736 2262 12738
rect 1785 12728 1841 12736
rect 2153 12728 2262 12736
rect 1681 12662 1761 12672
rect 1681 12606 1693 12662
rect 1749 12606 1761 12662
rect 1681 12596 1761 12606
rect 1865 12662 1945 12672
rect 1865 12606 1877 12662
rect 1933 12606 1945 12662
rect 1865 12596 1945 12606
rect 2049 12662 2129 12672
rect 2049 12606 2061 12662
rect 2117 12606 2129 12662
rect 2049 12596 2129 12606
rect 1693 12514 1749 12596
rect 1681 12512 1761 12514
rect 1681 12456 1693 12512
rect 1749 12456 1761 12512
rect 1681 12454 1761 12456
rect 708 12396 788 12398
rect 708 12340 720 12396
rect 776 12340 788 12396
rect 708 12338 788 12340
rect 1151 12396 1211 12406
rect 1151 12340 1153 12396
rect 1209 12340 1211 12396
rect 563 12280 643 12282
rect 563 12224 575 12280
rect 631 12224 643 12280
rect 563 12222 643 12224
rect 575 12140 631 12222
rect 195 12130 275 12140
rect 195 12074 207 12130
rect 263 12074 275 12130
rect 195 12064 275 12074
rect 379 12130 459 12140
rect 379 12074 391 12130
rect 447 12074 459 12130
rect 379 12064 459 12074
rect 563 12130 643 12140
rect 563 12074 575 12130
rect 631 12074 643 12130
rect 563 12064 643 12074
rect 708 12008 776 12338
rect 1151 12328 1211 12340
rect 667 12000 776 12008
rect 655 11998 776 12000
rect 655 11878 667 11998
rect 723 11878 776 11998
rect 655 11876 776 11878
rect 667 11868 723 11876
rect -30 11611 866 11623
rect -30 11555 -18 11611
rect 38 11555 800 11611
rect 856 11555 866 11611
rect -30 11543 866 11555
rect 1153 11385 1209 12328
rect 1693 12140 1749 12454
rect 1877 12398 1933 12596
rect 1865 12396 1945 12398
rect 1865 12340 1877 12396
rect 1933 12340 1945 12396
rect 1865 12338 1945 12340
rect 1877 12140 1933 12338
rect 2061 12282 2117 12596
rect 2194 12398 2262 12728
rect 2194 12396 2274 12398
rect 2194 12340 2206 12396
rect 2262 12340 2274 12396
rect 2194 12338 2274 12340
rect 2461 12396 2531 12408
rect 2461 12340 2463 12396
rect 2519 12340 2787 12396
rect 2049 12280 2129 12282
rect 2049 12224 2061 12280
rect 2117 12224 2129 12280
rect 2049 12222 2129 12224
rect 2061 12140 2117 12222
rect 1681 12130 1761 12140
rect 1681 12074 1693 12130
rect 1749 12074 1761 12130
rect 1681 12064 1761 12074
rect 1865 12130 1945 12140
rect 1865 12074 1877 12130
rect 1933 12074 1945 12130
rect 1865 12064 1945 12074
rect 2049 12130 2129 12140
rect 2049 12074 2061 12130
rect 2117 12074 2129 12130
rect 2049 12064 2129 12074
rect 2194 12008 2262 12338
rect 2461 12330 2531 12340
rect 2153 12000 2262 12008
rect 2141 11998 2262 12000
rect 2141 11878 2153 11998
rect 2209 11878 2262 11998
rect 2141 11876 2262 11878
rect 2153 11868 2209 11876
rect 1456 11611 2352 11623
rect 1456 11555 1468 11611
rect 1524 11555 2286 11611
rect 2342 11555 2352 11611
rect 1456 11543 2352 11555
rect 2463 11386 2519 12330
rect 2627 11494 2707 11504
rect 2627 11438 2639 11494
rect 2695 11438 2707 11494
rect 2627 11436 2707 11438
rect 1151 11383 1221 11385
rect 1151 11327 1153 11383
rect 1209 11327 1221 11383
rect 1151 11315 1221 11327
rect 2451 11384 2531 11386
rect 2451 11328 2463 11384
rect 2519 11328 2531 11384
rect 2451 11316 2531 11328
rect 115 11276 861 11288
rect 115 11220 483 11276
rect 539 11220 861 11276
rect 115 11208 861 11220
rect 115 10955 171 11208
rect 483 10955 539 11208
rect 805 10955 861 11208
rect 1601 11277 2347 11289
rect 1601 11221 1969 11277
rect 2025 11221 2347 11277
rect 1601 11209 2347 11221
rect 1601 10956 1657 11209
rect 1969 10956 2025 11209
rect 2291 10956 2347 11209
rect 103 10953 183 10955
rect 103 10833 115 10953
rect 171 10833 183 10953
rect 103 10831 183 10833
rect 471 10953 551 10955
rect 471 10833 483 10953
rect 539 10833 551 10953
rect 471 10831 551 10833
rect 793 10953 873 10955
rect 793 10832 805 10953
rect 861 10832 873 10953
rect 1589 10954 1669 10956
rect 1589 10834 1601 10954
rect 1657 10834 1669 10954
rect 1589 10832 1669 10834
rect 1957 10954 2037 10956
rect 1957 10834 1969 10954
rect 2025 10834 2037 10954
rect 1957 10832 2037 10834
rect 2279 10954 2359 10956
rect 2279 10833 2291 10954
rect 2347 10833 2359 10954
rect 115 10823 171 10831
rect 483 10823 539 10831
rect 793 10830 873 10832
rect 805 10822 861 10830
rect 1601 10824 1657 10832
rect 1969 10824 2025 10832
rect 2279 10831 2359 10833
rect 2291 10823 2347 10831
rect 299 10655 355 10663
rect 667 10655 723 10663
rect 1785 10656 1841 10664
rect 2153 10656 2209 10664
rect 287 10653 776 10655
rect 287 10533 299 10653
rect 355 10533 667 10653
rect 723 10533 776 10653
rect 287 10531 776 10533
rect 1773 10654 2262 10656
rect 1773 10534 1785 10654
rect 1841 10534 2153 10654
rect 2209 10534 2262 10654
rect 1773 10532 2262 10534
rect 299 10523 355 10531
rect 667 10523 776 10531
rect 1785 10524 1841 10532
rect 2153 10524 2262 10532
rect 195 10457 275 10467
rect 195 10401 207 10457
rect 263 10401 275 10457
rect 195 10391 275 10401
rect 379 10457 459 10467
rect 379 10401 391 10457
rect 447 10401 459 10457
rect 379 10391 459 10401
rect 563 10457 643 10467
rect 563 10401 575 10457
rect 631 10401 643 10457
rect 563 10391 643 10401
rect 207 10309 263 10391
rect 195 10307 275 10309
rect 195 10251 207 10307
rect 263 10251 275 10307
rect 195 10249 275 10251
rect -477 10075 -407 10087
rect -477 10019 -465 10075
rect -409 10019 -407 10075
rect -477 10007 -407 10019
rect 207 9935 263 10249
rect 391 10193 447 10391
rect 379 10191 459 10193
rect 379 10135 391 10191
rect 447 10135 459 10191
rect 379 10133 459 10135
rect 391 9935 447 10133
rect 575 10077 631 10391
rect 708 10193 776 10523
rect 1681 10458 1761 10468
rect 1681 10402 1693 10458
rect 1749 10402 1761 10458
rect 1681 10392 1761 10402
rect 1865 10458 1945 10468
rect 1865 10402 1877 10458
rect 1933 10402 1945 10458
rect 1865 10392 1945 10402
rect 2049 10458 2129 10468
rect 2049 10402 2061 10458
rect 2117 10402 2129 10458
rect 2049 10392 2129 10402
rect 1693 10310 1749 10392
rect 1681 10308 1761 10310
rect 1681 10252 1693 10308
rect 1749 10252 1761 10308
rect 1681 10250 1761 10252
rect 708 10191 788 10193
rect 708 10135 720 10191
rect 776 10135 788 10191
rect 708 10133 788 10135
rect 975 10191 1045 10203
rect 975 10135 977 10191
rect 1033 10135 1045 10191
rect 563 10075 643 10077
rect 563 10019 575 10075
rect 631 10019 643 10075
rect 563 10017 643 10019
rect 575 9935 631 10017
rect 195 9925 275 9935
rect 195 9869 207 9925
rect 263 9869 275 9925
rect 195 9859 275 9869
rect 379 9925 459 9935
rect 379 9869 391 9925
rect 447 9869 459 9925
rect 379 9859 459 9869
rect 563 9925 643 9935
rect 563 9869 575 9925
rect 631 9869 643 9925
rect 563 9859 643 9869
rect 708 9803 776 10133
rect 975 10125 1045 10135
rect 667 9795 776 9803
rect 655 9793 776 9795
rect 655 9673 667 9793
rect 723 9673 776 9793
rect 655 9671 776 9673
rect 667 9663 723 9671
rect -30 9406 866 9418
rect -30 9350 -18 9406
rect 38 9350 800 9406
rect 856 9350 866 9406
rect -30 9338 866 9350
rect 977 9181 1033 10125
rect 1693 9936 1749 10250
rect 1877 10194 1933 10392
rect 1865 10192 1945 10194
rect 1865 10136 1877 10192
rect 1933 10136 1945 10192
rect 1865 10134 1945 10136
rect 1877 9936 1933 10134
rect 2061 10078 2117 10392
rect 2194 10194 2262 10524
rect 2639 10202 2695 11436
rect 2194 10192 2274 10194
rect 2194 10136 2206 10192
rect 2262 10136 2274 10192
rect 2194 10134 2274 10136
rect 2637 10192 2707 10202
rect 2867 10192 2923 24235
rect 3069 21984 3125 25488
rect 3067 21972 3137 21984
rect 3067 21916 3069 21972
rect 3125 21916 3137 21972
rect 3067 21904 3137 21916
rect 3305 21072 3361 25840
rect 4157 25262 4903 25274
rect 4157 25206 4525 25262
rect 4581 25206 4903 25262
rect 4157 25194 4903 25206
rect 4157 24941 4213 25194
rect 4525 24941 4581 25194
rect 4847 24941 4903 25194
rect 4145 24939 4225 24941
rect 4145 24819 4157 24939
rect 4213 24819 4225 24939
rect 4145 24817 4225 24819
rect 4513 24939 4593 24941
rect 4513 24819 4525 24939
rect 4581 24819 4593 24939
rect 4513 24817 4593 24819
rect 4835 24939 4915 24941
rect 4835 24818 4847 24939
rect 4903 24818 4915 24939
rect 4157 24809 4213 24817
rect 4525 24809 4581 24817
rect 4835 24816 4915 24818
rect 4847 24808 4903 24816
rect 4341 24641 4397 24649
rect 4709 24641 4765 24649
rect 4329 24639 4818 24641
rect 4329 24519 4341 24639
rect 4397 24519 4709 24639
rect 4765 24519 4818 24639
rect 4329 24517 4818 24519
rect 4341 24509 4397 24517
rect 4709 24509 4818 24517
rect 4237 24443 4317 24453
rect 4237 24387 4249 24443
rect 4305 24387 4317 24443
rect 4237 24377 4317 24387
rect 4421 24443 4501 24453
rect 4421 24387 4433 24443
rect 4489 24387 4501 24443
rect 4421 24377 4501 24387
rect 4605 24443 4685 24453
rect 4605 24387 4617 24443
rect 4673 24387 4685 24443
rect 4605 24377 4685 24387
rect 4249 24295 4305 24377
rect 4237 24293 4317 24295
rect 4237 24237 4249 24293
rect 4305 24237 4317 24293
rect 4237 24235 4317 24237
rect 3565 24177 3635 24189
rect 3565 24121 3577 24177
rect 3633 24121 3635 24177
rect 3565 24109 3635 24121
rect 3429 21972 3499 21986
rect 3429 21916 3441 21972
rect 3497 21916 3499 21972
rect 3429 21904 3499 21916
rect 3293 21070 3363 21072
rect 3293 21014 3305 21070
rect 3361 21014 3363 21070
rect 3293 21002 3363 21014
rect 3441 17576 3497 21904
rect 3577 19663 3633 24109
rect 4249 23921 4305 24235
rect 4433 24179 4489 24377
rect 4421 24177 4501 24179
rect 4421 24121 4433 24177
rect 4489 24121 4501 24177
rect 4421 24119 4501 24121
rect 4433 23921 4489 24119
rect 4617 24063 4673 24377
rect 4750 24179 4818 24509
rect 6897 24293 6967 24305
rect 6897 24237 6909 24293
rect 6965 24237 6967 24293
rect 6897 24235 6967 24237
rect 4750 24177 4830 24179
rect 4750 24121 4762 24177
rect 4818 24121 4830 24177
rect 4750 24119 4830 24121
rect 5017 24177 5087 24189
rect 5017 24121 5019 24177
rect 5075 24121 5087 24177
rect 4605 24061 4685 24063
rect 4605 24005 4617 24061
rect 4673 24005 4685 24061
rect 4605 24003 4685 24005
rect 4617 23921 4673 24003
rect 4237 23911 4317 23921
rect 4237 23855 4249 23911
rect 4305 23855 4317 23911
rect 4237 23845 4317 23855
rect 4421 23911 4501 23921
rect 4421 23855 4433 23911
rect 4489 23855 4501 23911
rect 4421 23845 4501 23855
rect 4605 23911 4685 23921
rect 4605 23855 4617 23911
rect 4673 23855 4685 23911
rect 4605 23845 4685 23855
rect 4750 23789 4818 24119
rect 5017 24111 5087 24121
rect 4709 23781 4818 23789
rect 4697 23779 4818 23781
rect 4697 23659 4709 23779
rect 4765 23659 4818 23779
rect 4697 23657 4818 23659
rect 4709 23649 4765 23657
rect 4012 23392 4910 23404
rect 4012 23336 4024 23392
rect 4080 23336 4842 23392
rect 4898 23336 4910 23392
rect 4012 23324 4910 23336
rect 5019 23167 5075 24111
rect 5183 23274 5263 23284
rect 5183 23218 5195 23274
rect 5251 23218 5263 23274
rect 5183 23216 5263 23218
rect 5017 23164 5087 23167
rect 5017 23110 5019 23164
rect 5075 23110 5087 23164
rect 5017 23098 5087 23110
rect 4157 23057 4903 23069
rect 4157 23001 4525 23057
rect 4581 23001 4903 23057
rect 4157 22989 4903 23001
rect 4157 22736 4213 22989
rect 4525 22736 4581 22989
rect 4847 22736 4903 22989
rect 4145 22734 4225 22736
rect 4145 22614 4157 22734
rect 4213 22614 4225 22734
rect 4145 22612 4225 22614
rect 4513 22734 4593 22736
rect 4513 22614 4525 22734
rect 4581 22614 4593 22734
rect 4513 22612 4593 22614
rect 4835 22734 4915 22736
rect 4835 22613 4847 22734
rect 4903 22613 4915 22734
rect 4157 22604 4213 22612
rect 4525 22604 4581 22612
rect 4835 22611 4915 22613
rect 4847 22603 4903 22611
rect 4341 22436 4397 22444
rect 4709 22436 4765 22444
rect 4329 22434 4818 22436
rect 4329 22314 4341 22434
rect 4397 22314 4709 22434
rect 4765 22314 4818 22434
rect 4329 22312 4818 22314
rect 4341 22304 4397 22312
rect 4709 22304 4818 22312
rect 4237 22238 4317 22248
rect 4237 22182 4249 22238
rect 4305 22182 4317 22238
rect 4237 22172 4317 22182
rect 4421 22238 4501 22248
rect 4421 22182 4433 22238
rect 4489 22182 4501 22238
rect 4421 22172 4501 22182
rect 4605 22238 4685 22248
rect 4605 22182 4617 22238
rect 4673 22182 4685 22238
rect 4605 22172 4685 22182
rect 4249 22090 4305 22172
rect 4237 22088 4317 22090
rect 4237 22032 4249 22088
rect 4305 22032 4317 22088
rect 4237 22030 4317 22032
rect 4249 21716 4305 22030
rect 4433 21974 4489 22172
rect 4421 21972 4501 21974
rect 4421 21916 4433 21972
rect 4489 21916 4501 21972
rect 4421 21914 4501 21916
rect 4433 21716 4489 21914
rect 4617 21858 4673 22172
rect 4750 21974 4818 22304
rect 5195 21982 5251 23216
rect 5643 23057 6389 23069
rect 5643 23001 6011 23057
rect 6067 23001 6389 23057
rect 5643 22989 6389 23001
rect 5643 22736 5699 22989
rect 6011 22736 6067 22989
rect 6333 22736 6389 22989
rect 5631 22734 5711 22736
rect 5631 22614 5643 22734
rect 5699 22614 5711 22734
rect 5631 22612 5711 22614
rect 5999 22734 6079 22736
rect 5999 22614 6011 22734
rect 6067 22614 6079 22734
rect 5999 22612 6079 22614
rect 6321 22734 6401 22736
rect 6321 22613 6333 22734
rect 6389 22613 6401 22734
rect 5643 22604 5699 22612
rect 6011 22604 6067 22612
rect 6321 22611 6401 22613
rect 6333 22603 6389 22611
rect 5827 22436 5883 22444
rect 6195 22436 6251 22444
rect 5815 22434 6304 22436
rect 5815 22314 5827 22434
rect 5883 22314 6195 22434
rect 6251 22314 6304 22434
rect 5815 22312 6304 22314
rect 5827 22304 5883 22312
rect 6195 22304 6304 22312
rect 5723 22238 5803 22248
rect 5723 22182 5735 22238
rect 5791 22182 5803 22238
rect 5723 22172 5803 22182
rect 5907 22238 5987 22248
rect 5907 22182 5919 22238
rect 5975 22182 5987 22238
rect 5907 22172 5987 22182
rect 6091 22238 6171 22248
rect 6091 22182 6103 22238
rect 6159 22182 6171 22238
rect 6091 22172 6171 22182
rect 5735 22090 5791 22172
rect 5723 22088 5803 22090
rect 5723 22032 5735 22088
rect 5791 22032 5803 22088
rect 5723 22030 5803 22032
rect 4750 21972 4830 21974
rect 4750 21916 4762 21972
rect 4818 21916 4830 21972
rect 4750 21914 4830 21916
rect 5193 21972 5253 21982
rect 5193 21916 5195 21972
rect 5251 21916 5253 21972
rect 4605 21856 4685 21858
rect 4605 21800 4617 21856
rect 4673 21800 4685 21856
rect 4605 21798 4685 21800
rect 4617 21716 4673 21798
rect 4237 21706 4317 21716
rect 4237 21650 4249 21706
rect 4305 21650 4317 21706
rect 4237 21640 4317 21650
rect 4421 21706 4501 21716
rect 4421 21650 4433 21706
rect 4489 21650 4501 21706
rect 4421 21640 4501 21650
rect 4605 21706 4685 21716
rect 4605 21650 4617 21706
rect 4673 21650 4685 21706
rect 4605 21640 4685 21650
rect 4750 21584 4818 21914
rect 5193 21904 5253 21916
rect 4709 21576 4818 21584
rect 4697 21574 4818 21576
rect 4697 21454 4709 21574
rect 4765 21454 4818 21574
rect 4697 21452 4818 21454
rect 4709 21444 4765 21452
rect 4012 21187 4908 21199
rect 4012 21131 4024 21187
rect 4080 21131 4842 21187
rect 4898 21131 4908 21187
rect 4012 21119 4908 21131
rect 5195 20961 5251 21904
rect 5735 21716 5791 22030
rect 5919 21974 5975 22172
rect 5907 21972 5987 21974
rect 5907 21916 5919 21972
rect 5975 21916 5987 21972
rect 5907 21914 5987 21916
rect 5919 21716 5975 21914
rect 6103 21858 6159 22172
rect 6236 21974 6304 22304
rect 6236 21972 6316 21974
rect 6236 21916 6248 21972
rect 6304 21916 6316 21972
rect 6236 21914 6316 21916
rect 6503 21972 6573 21984
rect 6503 21916 6505 21972
rect 6561 21916 6829 21972
rect 6091 21856 6171 21858
rect 6091 21800 6103 21856
rect 6159 21800 6171 21856
rect 6091 21798 6171 21800
rect 6103 21716 6159 21798
rect 5723 21706 5803 21716
rect 5723 21650 5735 21706
rect 5791 21650 5803 21706
rect 5723 21640 5803 21650
rect 5907 21706 5987 21716
rect 5907 21650 5919 21706
rect 5975 21650 5987 21706
rect 5907 21640 5987 21650
rect 6091 21706 6171 21716
rect 6091 21650 6103 21706
rect 6159 21650 6171 21706
rect 6091 21640 6171 21650
rect 6236 21584 6304 21914
rect 6503 21906 6573 21916
rect 6195 21576 6304 21584
rect 6183 21574 6304 21576
rect 6183 21454 6195 21574
rect 6251 21454 6304 21574
rect 6183 21452 6304 21454
rect 6195 21444 6251 21452
rect 5498 21187 6394 21199
rect 5498 21131 5510 21187
rect 5566 21131 6328 21187
rect 6384 21131 6394 21187
rect 5498 21119 6394 21131
rect 6505 20962 6561 21906
rect 6669 21070 6749 21080
rect 6669 21014 6681 21070
rect 6737 21014 6749 21070
rect 6669 21012 6749 21014
rect 5193 20959 5263 20961
rect 5193 20903 5195 20959
rect 5251 20903 5263 20959
rect 5193 20891 5263 20903
rect 6493 20960 6573 20962
rect 6493 20904 6505 20960
rect 6561 20904 6573 20960
rect 6493 20892 6573 20904
rect 4157 20852 4903 20864
rect 4157 20796 4525 20852
rect 4581 20796 4903 20852
rect 4157 20784 4903 20796
rect 4157 20531 4213 20784
rect 4525 20531 4581 20784
rect 4847 20531 4903 20784
rect 5643 20853 6389 20865
rect 5643 20797 6011 20853
rect 6067 20797 6389 20853
rect 5643 20785 6389 20797
rect 5643 20532 5699 20785
rect 6011 20532 6067 20785
rect 6333 20532 6389 20785
rect 4145 20529 4225 20531
rect 4145 20409 4157 20529
rect 4213 20409 4225 20529
rect 4145 20407 4225 20409
rect 4513 20529 4593 20531
rect 4513 20409 4525 20529
rect 4581 20409 4593 20529
rect 4513 20407 4593 20409
rect 4835 20529 4915 20531
rect 4835 20408 4847 20529
rect 4903 20408 4915 20529
rect 5631 20530 5711 20532
rect 5631 20410 5643 20530
rect 5699 20410 5711 20530
rect 5631 20408 5711 20410
rect 5999 20530 6079 20532
rect 5999 20410 6011 20530
rect 6067 20410 6079 20530
rect 5999 20408 6079 20410
rect 6321 20530 6401 20532
rect 6321 20409 6333 20530
rect 6389 20409 6401 20530
rect 4157 20399 4213 20407
rect 4525 20399 4581 20407
rect 4835 20406 4915 20408
rect 4847 20398 4903 20406
rect 5643 20400 5699 20408
rect 6011 20400 6067 20408
rect 6321 20407 6401 20409
rect 6333 20399 6389 20407
rect 4341 20231 4397 20239
rect 4709 20231 4765 20239
rect 5827 20232 5883 20240
rect 6195 20232 6251 20240
rect 4329 20229 4818 20231
rect 4329 20109 4341 20229
rect 4397 20109 4709 20229
rect 4765 20109 4818 20229
rect 4329 20107 4818 20109
rect 5815 20230 6304 20232
rect 5815 20110 5827 20230
rect 5883 20110 6195 20230
rect 6251 20110 6304 20230
rect 5815 20108 6304 20110
rect 4341 20099 4397 20107
rect 4709 20099 4818 20107
rect 5827 20100 5883 20108
rect 6195 20100 6304 20108
rect 4237 20033 4317 20043
rect 4237 19977 4249 20033
rect 4305 19977 4317 20033
rect 4237 19967 4317 19977
rect 4421 20033 4501 20043
rect 4421 19977 4433 20033
rect 4489 19977 4501 20033
rect 4421 19967 4501 19977
rect 4605 20033 4685 20043
rect 4605 19977 4617 20033
rect 4673 19977 4685 20033
rect 4605 19967 4685 19977
rect 4249 19885 4305 19967
rect 4237 19883 4317 19885
rect 4237 19827 4249 19883
rect 4305 19827 4317 19883
rect 4237 19825 4317 19827
rect 3565 19651 3635 19663
rect 3565 19595 3577 19651
rect 3633 19595 3635 19651
rect 3565 19583 3635 19595
rect 4249 19511 4305 19825
rect 4433 19769 4489 19967
rect 4421 19767 4501 19769
rect 4421 19711 4433 19767
rect 4489 19711 4501 19767
rect 4421 19709 4501 19711
rect 4433 19511 4489 19709
rect 4617 19653 4673 19967
rect 4750 19769 4818 20099
rect 5723 20034 5803 20044
rect 5723 19978 5735 20034
rect 5791 19978 5803 20034
rect 5723 19968 5803 19978
rect 5907 20034 5987 20044
rect 5907 19978 5919 20034
rect 5975 19978 5987 20034
rect 5907 19968 5987 19978
rect 6091 20034 6171 20044
rect 6091 19978 6103 20034
rect 6159 19978 6171 20034
rect 6091 19968 6171 19978
rect 5735 19886 5791 19968
rect 5723 19884 5803 19886
rect 5723 19828 5735 19884
rect 5791 19828 5803 19884
rect 5723 19826 5803 19828
rect 4750 19767 4830 19769
rect 4750 19711 4762 19767
rect 4818 19711 4830 19767
rect 4750 19709 4830 19711
rect 5017 19767 5087 19779
rect 5017 19711 5019 19767
rect 5075 19711 5087 19767
rect 4605 19651 4685 19653
rect 4605 19595 4617 19651
rect 4673 19595 4685 19651
rect 4605 19593 4685 19595
rect 4617 19511 4673 19593
rect 4237 19501 4317 19511
rect 4237 19445 4249 19501
rect 4305 19445 4317 19501
rect 4237 19435 4317 19445
rect 4421 19501 4501 19511
rect 4421 19445 4433 19501
rect 4489 19445 4501 19501
rect 4421 19435 4501 19445
rect 4605 19501 4685 19511
rect 4605 19445 4617 19501
rect 4673 19445 4685 19501
rect 4605 19435 4685 19445
rect 4750 19379 4818 19709
rect 5017 19701 5087 19711
rect 4709 19371 4818 19379
rect 4697 19369 4818 19371
rect 4697 19249 4709 19369
rect 4765 19249 4818 19369
rect 4697 19247 4818 19249
rect 4709 19239 4765 19247
rect 4012 18982 4908 18994
rect 4012 18926 4024 18982
rect 4080 18926 4842 18982
rect 4898 18926 4908 18982
rect 4012 18914 4908 18926
rect 5019 18757 5075 19701
rect 5735 19512 5791 19826
rect 5919 19770 5975 19968
rect 5907 19768 5987 19770
rect 5907 19712 5919 19768
rect 5975 19712 5987 19768
rect 5907 19710 5987 19712
rect 5919 19512 5975 19710
rect 6103 19654 6159 19968
rect 6236 19770 6304 20100
rect 6681 19778 6737 21012
rect 6236 19768 6316 19770
rect 6236 19712 6248 19768
rect 6304 19712 6316 19768
rect 6236 19710 6316 19712
rect 6679 19768 6749 19778
rect 6679 19712 6681 19768
rect 6737 19712 6829 19768
rect 6091 19652 6171 19654
rect 6091 19596 6103 19652
rect 6159 19596 6171 19652
rect 6091 19594 6171 19596
rect 6103 19512 6159 19594
rect 5723 19502 5803 19512
rect 5723 19446 5735 19502
rect 5791 19446 5803 19502
rect 5723 19436 5803 19446
rect 5907 19502 5987 19512
rect 5907 19446 5919 19502
rect 5975 19446 5987 19502
rect 5907 19436 5987 19446
rect 6091 19502 6171 19512
rect 6091 19446 6103 19502
rect 6159 19446 6171 19502
rect 6091 19436 6171 19446
rect 6236 19380 6304 19710
rect 6679 19700 6749 19712
rect 6195 19372 6304 19380
rect 6183 19370 6304 19372
rect 6183 19250 6195 19370
rect 6251 19250 6304 19370
rect 6183 19248 6304 19250
rect 6195 19240 6251 19248
rect 5498 18983 6394 18995
rect 5498 18927 5510 18983
rect 5566 18927 6328 18983
rect 6384 18927 6394 18983
rect 5498 18915 6394 18927
rect 5183 18864 5263 18874
rect 5183 18808 5195 18864
rect 5251 18808 5263 18864
rect 5183 18806 5263 18808
rect 5017 18754 5087 18757
rect 5017 18700 5019 18754
rect 5075 18700 5087 18754
rect 5017 18688 5087 18700
rect 4157 18647 4903 18659
rect 4157 18591 4525 18647
rect 4581 18591 4903 18647
rect 4157 18579 4903 18591
rect 4157 18326 4213 18579
rect 4525 18326 4581 18579
rect 4847 18326 4903 18579
rect 4145 18324 4225 18326
rect 4145 18204 4157 18324
rect 4213 18204 4225 18324
rect 4145 18202 4225 18204
rect 4513 18324 4593 18326
rect 4513 18204 4525 18324
rect 4581 18204 4593 18324
rect 4513 18202 4593 18204
rect 4835 18324 4915 18326
rect 4835 18203 4847 18324
rect 4903 18203 4915 18324
rect 4157 18194 4213 18202
rect 4525 18194 4581 18202
rect 4835 18201 4915 18203
rect 4847 18193 4903 18201
rect 4341 18026 4397 18034
rect 4709 18026 4765 18034
rect 4329 18024 4818 18026
rect 4329 17904 4341 18024
rect 4397 17904 4709 18024
rect 4765 17904 4818 18024
rect 4329 17902 4818 17904
rect 4341 17894 4397 17902
rect 4709 17894 4818 17902
rect 4237 17828 4317 17838
rect 4237 17772 4249 17828
rect 4305 17772 4317 17828
rect 4237 17762 4317 17772
rect 4421 17828 4501 17838
rect 4421 17772 4433 17828
rect 4489 17772 4501 17828
rect 4421 17762 4501 17772
rect 4605 17828 4685 17838
rect 4605 17772 4617 17828
rect 4673 17772 4685 17828
rect 4605 17762 4685 17772
rect 4249 17680 4305 17762
rect 4237 17678 4317 17680
rect 4237 17622 4249 17678
rect 4305 17622 4317 17678
rect 4237 17620 4317 17622
rect 3429 17562 3499 17576
rect 3429 17506 3441 17562
rect 3497 17506 3499 17562
rect 3429 17494 3499 17506
rect 3127 16659 3197 16671
rect 3441 16663 3497 17494
rect 4249 17306 4305 17620
rect 4433 17564 4489 17762
rect 4421 17562 4501 17564
rect 4421 17506 4433 17562
rect 4489 17506 4501 17562
rect 4421 17504 4501 17506
rect 4433 17306 4489 17504
rect 4617 17448 4673 17762
rect 4750 17564 4818 17894
rect 5195 17574 5251 18806
rect 4750 17562 4830 17564
rect 4750 17506 4762 17562
rect 4818 17506 4830 17562
rect 4750 17504 4830 17506
rect 5193 17562 5253 17574
rect 5193 17506 5195 17562
rect 5251 17506 5253 17562
rect 4605 17446 4685 17448
rect 4605 17390 4617 17446
rect 4673 17390 4685 17446
rect 4605 17388 4685 17390
rect 4617 17306 4673 17388
rect 4237 17296 4317 17306
rect 4237 17240 4249 17296
rect 4305 17240 4317 17296
rect 4237 17230 4317 17240
rect 4421 17296 4501 17306
rect 4421 17240 4433 17296
rect 4489 17240 4501 17296
rect 4421 17230 4501 17240
rect 4605 17296 4685 17306
rect 4605 17240 4617 17296
rect 4673 17240 4685 17296
rect 4605 17230 4685 17240
rect 4750 17174 4818 17504
rect 5193 17494 5253 17506
rect 6625 17446 6695 17458
rect 6625 17390 6637 17446
rect 6693 17390 6695 17446
rect 6625 17378 6695 17390
rect 4709 17166 4818 17174
rect 4697 17164 4818 17166
rect 4697 17044 4709 17164
rect 4765 17044 4818 17164
rect 4697 17042 4818 17044
rect 4709 17034 4765 17042
rect 4012 16777 4910 16789
rect 4012 16721 4024 16777
rect 4080 16721 4842 16777
rect 4898 16721 4910 16777
rect 4012 16709 4910 16721
rect 3127 16603 3139 16659
rect 3195 16603 3197 16659
rect 3127 16601 3197 16603
rect 3439 16659 3499 16663
rect 3439 16603 3441 16659
rect 3497 16603 3499 16659
rect 3139 15989 3195 16601
rect 3439 16591 3499 16603
rect 6637 16499 6693 17378
rect 6637 16389 6693 16399
rect 2991 11494 3061 11506
rect 2991 11438 3003 11494
rect 3059 11438 3061 11494
rect 2991 11426 3061 11438
rect 2637 10136 2639 10192
rect 2695 10136 2923 10192
rect 2049 10076 2129 10078
rect 2049 10020 2061 10076
rect 2117 10020 2129 10076
rect 2049 10018 2129 10020
rect 2061 9936 2117 10018
rect 1681 9926 1761 9936
rect 1681 9870 1693 9926
rect 1749 9870 1761 9926
rect 1681 9860 1761 9870
rect 1865 9926 1945 9936
rect 1865 9870 1877 9926
rect 1933 9870 1945 9926
rect 1865 9860 1945 9870
rect 2049 9926 2129 9936
rect 2049 9870 2061 9926
rect 2117 9870 2129 9926
rect 2049 9860 2129 9870
rect 2194 9804 2262 10134
rect 2637 10124 2707 10136
rect 2153 9796 2262 9804
rect 2141 9794 2262 9796
rect 2141 9674 2153 9794
rect 2209 9674 2262 9794
rect 2141 9672 2262 9674
rect 2153 9664 2209 9672
rect 1456 9407 2352 9419
rect 1456 9351 1468 9407
rect 1524 9351 2286 9407
rect 2342 9351 2352 9407
rect 1456 9339 2352 9351
rect 1141 9288 1221 9298
rect 1141 9232 1153 9288
rect 1209 9232 1221 9288
rect 1141 9230 1221 9232
rect 975 9178 1045 9181
rect 975 9124 977 9178
rect 1033 9124 1045 9178
rect 975 9112 1045 9124
rect 115 9071 861 9083
rect 115 9015 483 9071
rect 539 9015 861 9071
rect 115 9003 861 9015
rect 115 8750 171 9003
rect 483 8750 539 9003
rect 805 8750 861 9003
rect 103 8748 183 8750
rect 103 8628 115 8748
rect 171 8628 183 8748
rect 103 8626 183 8628
rect 471 8748 551 8750
rect 471 8628 483 8748
rect 539 8628 551 8748
rect 471 8626 551 8628
rect 793 8748 873 8750
rect 793 8627 805 8748
rect 861 8627 873 8748
rect 115 8618 171 8626
rect 483 8618 539 8626
rect 793 8625 873 8627
rect 805 8617 861 8625
rect 299 8450 355 8458
rect 667 8450 723 8458
rect 287 8448 776 8450
rect 287 8328 299 8448
rect 355 8328 667 8448
rect 723 8328 776 8448
rect 287 8326 776 8328
rect 299 8318 355 8326
rect 667 8318 776 8326
rect 195 8252 275 8262
rect 195 8196 207 8252
rect 263 8196 275 8252
rect 195 8186 275 8196
rect 379 8252 459 8262
rect 379 8196 391 8252
rect 447 8196 459 8252
rect 379 8186 459 8196
rect 563 8252 643 8262
rect 563 8196 575 8252
rect 631 8196 643 8252
rect 563 8186 643 8196
rect 207 8104 263 8186
rect 195 8102 275 8104
rect 195 8046 207 8102
rect 263 8046 275 8102
rect 195 8044 275 8046
rect -613 7986 -543 8000
rect -613 7930 -601 7986
rect -545 7930 -543 7986
rect -613 7918 -543 7930
rect -779 7870 -699 7882
rect -779 7814 -767 7870
rect -711 7814 -699 7870
rect -779 7802 -699 7814
rect -915 7083 -845 7095
rect -601 7087 -545 7918
rect 207 7730 263 8044
rect 391 7988 447 8186
rect 379 7986 459 7988
rect 379 7930 391 7986
rect 447 7930 459 7986
rect 379 7928 459 7930
rect 391 7730 447 7928
rect 575 7872 631 8186
rect 708 7988 776 8318
rect 1153 7998 1209 9230
rect 708 7986 788 7988
rect 708 7930 720 7986
rect 776 7930 788 7986
rect 708 7928 788 7930
rect 1151 7986 1211 7998
rect 1151 7930 1153 7986
rect 1209 7930 1211 7986
rect 563 7870 643 7872
rect 563 7814 575 7870
rect 631 7814 643 7870
rect 563 7812 643 7814
rect 575 7730 631 7812
rect 195 7720 275 7730
rect 195 7664 207 7720
rect 263 7664 275 7720
rect 195 7654 275 7664
rect 379 7720 459 7730
rect 379 7664 391 7720
rect 447 7664 459 7720
rect 379 7654 459 7664
rect 563 7720 643 7730
rect 563 7664 575 7720
rect 631 7664 643 7720
rect 563 7654 643 7664
rect 708 7598 776 7928
rect 1151 7918 1211 7930
rect 667 7590 776 7598
rect 655 7588 776 7590
rect 655 7468 667 7588
rect 723 7468 776 7588
rect 655 7466 776 7468
rect 667 7458 723 7466
rect -30 7201 868 7213
rect -30 7145 -18 7201
rect 38 7145 800 7201
rect 856 7145 868 7201
rect -30 7133 868 7145
rect -915 7027 -903 7083
rect -847 7027 -845 7083
rect -915 7015 -845 7027
rect -603 7083 -543 7087
rect -603 7027 -601 7083
rect -545 7027 -543 7083
rect -603 7015 -543 7027
rect -1039 6810 -983 6820
rect 3003 6920 3059 11426
rect 3139 7095 3195 15889
rect 4157 15686 4903 15698
rect 4157 15630 4525 15686
rect 4581 15630 4903 15686
rect 4157 15618 4903 15630
rect 4157 15365 4213 15618
rect 4525 15365 4581 15618
rect 4847 15365 4903 15618
rect 4145 15363 4225 15365
rect 4145 15243 4157 15363
rect 4213 15243 4225 15363
rect 4145 15241 4225 15243
rect 4513 15363 4593 15365
rect 4513 15243 4525 15363
rect 4581 15243 4593 15363
rect 4513 15241 4593 15243
rect 4835 15363 4915 15365
rect 4835 15242 4847 15363
rect 4903 15242 4915 15363
rect 4157 15233 4213 15241
rect 4525 15233 4581 15241
rect 4835 15240 4915 15242
rect 4847 15232 4903 15240
rect 4341 15065 4397 15073
rect 4709 15065 4765 15073
rect 4329 15063 4818 15065
rect 4329 14943 4341 15063
rect 4397 14943 4709 15063
rect 4765 14943 4818 15063
rect 4329 14941 4818 14943
rect 4341 14933 4397 14941
rect 4709 14933 4818 14941
rect 4237 14867 4317 14877
rect 4237 14811 4249 14867
rect 4305 14811 4317 14867
rect 4237 14801 4317 14811
rect 4421 14867 4501 14877
rect 4421 14811 4433 14867
rect 4489 14811 4501 14867
rect 4421 14801 4501 14811
rect 4605 14867 4685 14877
rect 4605 14811 4617 14867
rect 4673 14811 4685 14867
rect 4605 14801 4685 14811
rect 3349 14717 3435 14729
rect 4249 14719 4305 14801
rect 3349 14661 3361 14717
rect 3417 14661 3435 14717
rect 3349 14649 3435 14661
rect 4237 14717 4317 14719
rect 4237 14661 4249 14717
rect 4305 14661 4317 14717
rect 4237 14659 4317 14661
rect 3565 14601 3635 14613
rect 3565 14545 3577 14601
rect 3633 14545 3635 14601
rect 3565 14533 3635 14545
rect 3429 12396 3499 12410
rect 3429 12340 3441 12396
rect 3497 12340 3499 12396
rect 3429 12328 3499 12340
rect 3263 12208 3343 12218
rect 3263 12152 3275 12208
rect 3331 12152 3343 12208
rect 3263 12150 3343 12152
rect 3275 7882 3331 12150
rect 3441 8000 3497 12328
rect 3577 10087 3633 14533
rect 4249 14345 4305 14659
rect 4433 14603 4489 14801
rect 4421 14601 4501 14603
rect 4421 14545 4433 14601
rect 4489 14545 4501 14601
rect 4421 14543 4501 14545
rect 4433 14345 4489 14543
rect 4617 14487 4673 14801
rect 4750 14603 4818 14933
rect 4750 14601 4830 14603
rect 4750 14545 4762 14601
rect 4818 14545 4830 14601
rect 4750 14543 4830 14545
rect 5017 14601 5087 14613
rect 5017 14545 5019 14601
rect 5075 14545 5087 14601
rect 4605 14485 4685 14487
rect 4605 14429 4617 14485
rect 4673 14429 4685 14485
rect 4605 14427 4685 14429
rect 4617 14345 4673 14427
rect 4237 14335 4317 14345
rect 4237 14279 4249 14335
rect 4305 14279 4317 14335
rect 4237 14269 4317 14279
rect 4421 14335 4501 14345
rect 4421 14279 4433 14335
rect 4489 14279 4501 14335
rect 4421 14269 4501 14279
rect 4605 14335 4685 14345
rect 4605 14279 4617 14335
rect 4673 14279 4685 14335
rect 4605 14269 4685 14279
rect 4750 14213 4818 14543
rect 5017 14535 5087 14545
rect 4709 14205 4818 14213
rect 4697 14203 4818 14205
rect 4697 14083 4709 14203
rect 4765 14083 4818 14203
rect 4697 14081 4818 14083
rect 4709 14073 4765 14081
rect 4012 13816 4910 13828
rect 4012 13760 4024 13816
rect 4080 13760 4842 13816
rect 4898 13760 4910 13816
rect 4012 13748 4910 13760
rect 5019 13591 5075 14535
rect 5183 13698 5263 13708
rect 5183 13642 5195 13698
rect 5251 13642 5263 13698
rect 5183 13640 5263 13642
rect 5017 13588 5087 13591
rect 5017 13534 5019 13588
rect 5075 13534 5087 13588
rect 5017 13522 5087 13534
rect 4157 13481 4903 13493
rect 4157 13425 4525 13481
rect 4581 13425 4903 13481
rect 4157 13413 4903 13425
rect 4157 13160 4213 13413
rect 4525 13160 4581 13413
rect 4847 13160 4903 13413
rect 4145 13158 4225 13160
rect 4145 13038 4157 13158
rect 4213 13038 4225 13158
rect 4145 13036 4225 13038
rect 4513 13158 4593 13160
rect 4513 13038 4525 13158
rect 4581 13038 4593 13158
rect 4513 13036 4593 13038
rect 4835 13158 4915 13160
rect 4835 13037 4847 13158
rect 4903 13037 4915 13158
rect 4157 13028 4213 13036
rect 4525 13028 4581 13036
rect 4835 13035 4915 13037
rect 4847 13027 4903 13035
rect 4341 12860 4397 12868
rect 4709 12860 4765 12868
rect 4329 12858 4818 12860
rect 4329 12738 4341 12858
rect 4397 12738 4709 12858
rect 4765 12738 4818 12858
rect 4329 12736 4818 12738
rect 4341 12728 4397 12736
rect 4709 12728 4818 12736
rect 4237 12662 4317 12672
rect 4237 12606 4249 12662
rect 4305 12606 4317 12662
rect 4237 12596 4317 12606
rect 4421 12662 4501 12672
rect 4421 12606 4433 12662
rect 4489 12606 4501 12662
rect 4421 12596 4501 12606
rect 4605 12662 4685 12672
rect 4605 12606 4617 12662
rect 4673 12606 4685 12662
rect 4605 12596 4685 12606
rect 4249 12514 4305 12596
rect 4237 12512 4317 12514
rect 4237 12456 4249 12512
rect 4305 12456 4317 12512
rect 4237 12454 4317 12456
rect 4249 12140 4305 12454
rect 4433 12398 4489 12596
rect 4421 12396 4501 12398
rect 4421 12340 4433 12396
rect 4489 12340 4501 12396
rect 4421 12338 4501 12340
rect 4433 12140 4489 12338
rect 4617 12282 4673 12596
rect 4750 12398 4818 12728
rect 5195 12406 5251 13640
rect 5643 13481 6389 13493
rect 5643 13425 6011 13481
rect 6067 13425 6389 13481
rect 5643 13413 6389 13425
rect 5643 13160 5699 13413
rect 6011 13160 6067 13413
rect 6333 13160 6389 13413
rect 5631 13158 5711 13160
rect 5631 13038 5643 13158
rect 5699 13038 5711 13158
rect 5631 13036 5711 13038
rect 5999 13158 6079 13160
rect 5999 13038 6011 13158
rect 6067 13038 6079 13158
rect 5999 13036 6079 13038
rect 6321 13158 6401 13160
rect 6321 13037 6333 13158
rect 6389 13037 6401 13158
rect 5643 13028 5699 13036
rect 6011 13028 6067 13036
rect 6321 13035 6401 13037
rect 6333 13027 6389 13035
rect 5827 12860 5883 12868
rect 6195 12860 6251 12868
rect 5815 12858 6304 12860
rect 5815 12738 5827 12858
rect 5883 12738 6195 12858
rect 6251 12738 6304 12858
rect 5815 12736 6304 12738
rect 5827 12728 5883 12736
rect 6195 12728 6304 12736
rect 5723 12662 5803 12672
rect 5723 12606 5735 12662
rect 5791 12606 5803 12662
rect 5723 12596 5803 12606
rect 5907 12662 5987 12672
rect 5907 12606 5919 12662
rect 5975 12606 5987 12662
rect 5907 12596 5987 12606
rect 6091 12662 6171 12672
rect 6091 12606 6103 12662
rect 6159 12606 6171 12662
rect 6091 12596 6171 12606
rect 5735 12514 5791 12596
rect 5723 12512 5803 12514
rect 5723 12456 5735 12512
rect 5791 12456 5803 12512
rect 5723 12454 5803 12456
rect 4750 12396 4830 12398
rect 4750 12340 4762 12396
rect 4818 12340 4830 12396
rect 4750 12338 4830 12340
rect 5193 12396 5253 12406
rect 5193 12340 5195 12396
rect 5251 12340 5253 12396
rect 4605 12280 4685 12282
rect 4605 12224 4617 12280
rect 4673 12224 4685 12280
rect 4605 12222 4685 12224
rect 4617 12140 4673 12222
rect 4237 12130 4317 12140
rect 4237 12074 4249 12130
rect 4305 12074 4317 12130
rect 4237 12064 4317 12074
rect 4421 12130 4501 12140
rect 4421 12074 4433 12130
rect 4489 12074 4501 12130
rect 4421 12064 4501 12074
rect 4605 12130 4685 12140
rect 4605 12074 4617 12130
rect 4673 12074 4685 12130
rect 4605 12064 4685 12074
rect 4750 12008 4818 12338
rect 5193 12328 5253 12340
rect 4709 12000 4818 12008
rect 4697 11998 4818 12000
rect 4697 11878 4709 11998
rect 4765 11878 4818 11998
rect 4697 11876 4818 11878
rect 4709 11868 4765 11876
rect 4012 11611 4908 11623
rect 4012 11555 4024 11611
rect 4080 11555 4842 11611
rect 4898 11555 4908 11611
rect 4012 11543 4908 11555
rect 5195 11385 5251 12328
rect 5735 12140 5791 12454
rect 5919 12398 5975 12596
rect 5907 12396 5987 12398
rect 5907 12340 5919 12396
rect 5975 12340 5987 12396
rect 5907 12338 5987 12340
rect 5919 12140 5975 12338
rect 6103 12282 6159 12596
rect 6236 12398 6304 12728
rect 6236 12396 6316 12398
rect 6236 12340 6248 12396
rect 6304 12340 6316 12396
rect 6236 12338 6316 12340
rect 6503 12396 6573 12408
rect 6503 12340 6505 12396
rect 6561 12340 6829 12396
rect 6091 12280 6171 12282
rect 6091 12224 6103 12280
rect 6159 12224 6171 12280
rect 6091 12222 6171 12224
rect 6103 12140 6159 12222
rect 5723 12130 5803 12140
rect 5723 12074 5735 12130
rect 5791 12074 5803 12130
rect 5723 12064 5803 12074
rect 5907 12130 5987 12140
rect 5907 12074 5919 12130
rect 5975 12074 5987 12130
rect 5907 12064 5987 12074
rect 6091 12130 6171 12140
rect 6091 12074 6103 12130
rect 6159 12074 6171 12130
rect 6091 12064 6171 12074
rect 6236 12008 6304 12338
rect 6503 12330 6573 12340
rect 6195 12000 6304 12008
rect 6183 11998 6304 12000
rect 6183 11878 6195 11998
rect 6251 11878 6304 11998
rect 6183 11876 6304 11878
rect 6195 11868 6251 11876
rect 5498 11611 6394 11623
rect 5498 11555 5510 11611
rect 5566 11555 6328 11611
rect 6384 11555 6394 11611
rect 5498 11543 6394 11555
rect 6505 11386 6561 12330
rect 6669 11494 6749 11504
rect 6669 11438 6681 11494
rect 6737 11438 6749 11494
rect 6669 11436 6749 11438
rect 5193 11383 5263 11385
rect 5193 11327 5195 11383
rect 5251 11327 5263 11383
rect 5193 11315 5263 11327
rect 6493 11384 6573 11386
rect 6493 11328 6505 11384
rect 6561 11328 6573 11384
rect 6493 11316 6573 11328
rect 4157 11276 4903 11288
rect 4157 11220 4525 11276
rect 4581 11220 4903 11276
rect 4157 11208 4903 11220
rect 4157 10955 4213 11208
rect 4525 10955 4581 11208
rect 4847 10955 4903 11208
rect 5643 11277 6389 11289
rect 5643 11221 6011 11277
rect 6067 11221 6389 11277
rect 5643 11209 6389 11221
rect 5643 10956 5699 11209
rect 6011 10956 6067 11209
rect 6333 10956 6389 11209
rect 4145 10953 4225 10955
rect 4145 10833 4157 10953
rect 4213 10833 4225 10953
rect 4145 10831 4225 10833
rect 4513 10953 4593 10955
rect 4513 10833 4525 10953
rect 4581 10833 4593 10953
rect 4513 10831 4593 10833
rect 4835 10953 4915 10955
rect 4835 10832 4847 10953
rect 4903 10832 4915 10953
rect 5631 10954 5711 10956
rect 5631 10834 5643 10954
rect 5699 10834 5711 10954
rect 5631 10832 5711 10834
rect 5999 10954 6079 10956
rect 5999 10834 6011 10954
rect 6067 10834 6079 10954
rect 5999 10832 6079 10834
rect 6321 10954 6401 10956
rect 6321 10833 6333 10954
rect 6389 10833 6401 10954
rect 4157 10823 4213 10831
rect 4525 10823 4581 10831
rect 4835 10830 4915 10832
rect 4847 10822 4903 10830
rect 5643 10824 5699 10832
rect 6011 10824 6067 10832
rect 6321 10831 6401 10833
rect 6333 10823 6389 10831
rect 4341 10655 4397 10663
rect 4709 10655 4765 10663
rect 5827 10656 5883 10664
rect 6195 10656 6251 10664
rect 4329 10653 4818 10655
rect 4329 10533 4341 10653
rect 4397 10533 4709 10653
rect 4765 10533 4818 10653
rect 4329 10531 4818 10533
rect 5815 10654 6304 10656
rect 5815 10534 5827 10654
rect 5883 10534 6195 10654
rect 6251 10534 6304 10654
rect 5815 10532 6304 10534
rect 4341 10523 4397 10531
rect 4709 10523 4818 10531
rect 5827 10524 5883 10532
rect 6195 10524 6304 10532
rect 4237 10457 4317 10467
rect 4237 10401 4249 10457
rect 4305 10401 4317 10457
rect 4237 10391 4317 10401
rect 4421 10457 4501 10467
rect 4421 10401 4433 10457
rect 4489 10401 4501 10457
rect 4421 10391 4501 10401
rect 4605 10457 4685 10467
rect 4605 10401 4617 10457
rect 4673 10401 4685 10457
rect 4605 10391 4685 10401
rect 4249 10309 4305 10391
rect 4237 10307 4317 10309
rect 4237 10251 4249 10307
rect 4305 10251 4317 10307
rect 4237 10249 4317 10251
rect 3565 10075 3635 10087
rect 3565 10019 3577 10075
rect 3633 10019 3635 10075
rect 3565 10007 3635 10019
rect 4249 9935 4305 10249
rect 4433 10193 4489 10391
rect 4421 10191 4501 10193
rect 4421 10135 4433 10191
rect 4489 10135 4501 10191
rect 4421 10133 4501 10135
rect 4433 9935 4489 10133
rect 4617 10077 4673 10391
rect 4750 10193 4818 10523
rect 5723 10458 5803 10468
rect 5723 10402 5735 10458
rect 5791 10402 5803 10458
rect 5723 10392 5803 10402
rect 5907 10458 5987 10468
rect 5907 10402 5919 10458
rect 5975 10402 5987 10458
rect 5907 10392 5987 10402
rect 6091 10458 6171 10468
rect 6091 10402 6103 10458
rect 6159 10402 6171 10458
rect 6091 10392 6171 10402
rect 5735 10310 5791 10392
rect 5723 10308 5803 10310
rect 5723 10252 5735 10308
rect 5791 10252 5803 10308
rect 5723 10250 5803 10252
rect 4750 10191 4830 10193
rect 4750 10135 4762 10191
rect 4818 10135 4830 10191
rect 4750 10133 4830 10135
rect 5017 10191 5087 10203
rect 5017 10135 5019 10191
rect 5075 10135 5087 10191
rect 4605 10075 4685 10077
rect 4605 10019 4617 10075
rect 4673 10019 4685 10075
rect 4605 10017 4685 10019
rect 4617 9935 4673 10017
rect 4237 9925 4317 9935
rect 4237 9869 4249 9925
rect 4305 9869 4317 9925
rect 4237 9859 4317 9869
rect 4421 9925 4501 9935
rect 4421 9869 4433 9925
rect 4489 9869 4501 9925
rect 4421 9859 4501 9869
rect 4605 9925 4685 9935
rect 4605 9869 4617 9925
rect 4673 9869 4685 9925
rect 4605 9859 4685 9869
rect 4750 9803 4818 10133
rect 5017 10125 5087 10135
rect 4709 9795 4818 9803
rect 4697 9793 4818 9795
rect 4697 9673 4709 9793
rect 4765 9673 4818 9793
rect 4697 9671 4818 9673
rect 4709 9663 4765 9671
rect 4012 9406 4908 9418
rect 4012 9350 4024 9406
rect 4080 9350 4842 9406
rect 4898 9350 4908 9406
rect 4012 9338 4908 9350
rect 5019 9181 5075 10125
rect 5735 9936 5791 10250
rect 5919 10194 5975 10392
rect 5907 10192 5987 10194
rect 5907 10136 5919 10192
rect 5975 10136 5987 10192
rect 5907 10134 5987 10136
rect 5919 9936 5975 10134
rect 6103 10078 6159 10392
rect 6236 10194 6304 10524
rect 6681 10202 6737 11436
rect 6236 10192 6316 10194
rect 6236 10136 6248 10192
rect 6304 10136 6316 10192
rect 6236 10134 6316 10136
rect 6679 10192 6749 10202
rect 6909 10192 6965 24235
rect 7111 21984 7167 26016
rect 11153 25900 11209 26758
rect 15195 26445 15251 26486
rect 36219 26445 36275 28454
rect 38409 28442 38479 28454
rect 37699 28228 37779 28238
rect 37699 28172 37711 28228
rect 37767 28172 37779 28228
rect 37699 27986 37779 28172
rect 38179 28228 38259 28238
rect 38179 28172 38191 28228
rect 38247 28172 38259 28228
rect 38179 28162 38259 28172
rect 38383 28228 38463 28238
rect 38383 28172 38395 28228
rect 38451 28172 38463 28228
rect 38383 27986 38463 28172
rect 38587 28228 38667 28532
rect 38889 28520 38959 28532
rect 39067 28588 39147 28883
rect 39368 28588 39424 29618
rect 40501 29608 40597 29618
rect 40815 29402 40895 29696
rect 41117 29684 41187 29696
rect 41295 29752 41375 30047
rect 41933 29882 41989 34210
rect 42069 31969 42125 36415
rect 42741 36227 42797 36541
rect 42925 36485 42981 36683
rect 42913 36483 42993 36485
rect 42913 36427 42925 36483
rect 42981 36427 42993 36483
rect 42913 36425 42993 36427
rect 42925 36227 42981 36425
rect 43109 36369 43165 36683
rect 43242 36485 43310 36815
rect 43242 36483 43322 36485
rect 43242 36427 43254 36483
rect 43310 36427 43322 36483
rect 43242 36425 43322 36427
rect 43509 36483 43579 36495
rect 43509 36427 43511 36483
rect 43567 36427 43579 36483
rect 43097 36367 43177 36369
rect 43097 36311 43109 36367
rect 43165 36311 43177 36367
rect 43097 36309 43177 36311
rect 43109 36227 43165 36309
rect 42729 36217 42809 36227
rect 42729 36161 42741 36217
rect 42797 36161 42809 36217
rect 42729 36151 42809 36161
rect 42913 36217 42993 36227
rect 42913 36161 42925 36217
rect 42981 36161 42993 36217
rect 42913 36151 42993 36161
rect 43097 36217 43177 36227
rect 43097 36161 43109 36217
rect 43165 36161 43177 36217
rect 43097 36151 43177 36161
rect 43242 36095 43310 36425
rect 43509 36417 43579 36427
rect 43201 36087 43310 36095
rect 43189 36085 43310 36087
rect 43189 35965 43201 36085
rect 43257 35965 43310 36085
rect 43189 35963 43310 35965
rect 43201 35955 43257 35963
rect 42504 35698 43402 35710
rect 42504 35642 42516 35698
rect 42572 35642 43334 35698
rect 43390 35642 43402 35698
rect 42504 35630 43402 35642
rect 43511 35473 43567 36417
rect 43675 35580 43755 35590
rect 43675 35524 43687 35580
rect 43743 35524 43755 35580
rect 43675 35522 43755 35524
rect 43509 35470 43579 35473
rect 43509 35416 43511 35470
rect 43567 35416 43579 35470
rect 43509 35404 43579 35416
rect 42649 35363 43395 35375
rect 42649 35307 43017 35363
rect 43073 35307 43395 35363
rect 42649 35295 43395 35307
rect 42649 35042 42705 35295
rect 43017 35042 43073 35295
rect 43339 35042 43395 35295
rect 42637 35040 42717 35042
rect 42637 34920 42649 35040
rect 42705 34920 42717 35040
rect 42637 34918 42717 34920
rect 43005 35040 43085 35042
rect 43005 34920 43017 35040
rect 43073 34920 43085 35040
rect 43005 34918 43085 34920
rect 43327 35040 43407 35042
rect 43327 34919 43339 35040
rect 43395 34919 43407 35040
rect 42649 34910 42705 34918
rect 43017 34910 43073 34918
rect 43327 34917 43407 34919
rect 43339 34909 43395 34917
rect 42833 34742 42889 34750
rect 43201 34742 43257 34750
rect 42821 34740 43310 34742
rect 42821 34620 42833 34740
rect 42889 34620 43201 34740
rect 43257 34620 43310 34740
rect 42821 34618 43310 34620
rect 42833 34610 42889 34618
rect 43201 34610 43310 34618
rect 42729 34544 42809 34554
rect 42729 34488 42741 34544
rect 42797 34488 42809 34544
rect 42729 34478 42809 34488
rect 42913 34544 42993 34554
rect 42913 34488 42925 34544
rect 42981 34488 42993 34544
rect 42913 34478 42993 34488
rect 43097 34544 43177 34554
rect 43097 34488 43109 34544
rect 43165 34488 43177 34544
rect 43097 34478 43177 34488
rect 42741 34396 42797 34478
rect 42729 34394 42809 34396
rect 42729 34338 42741 34394
rect 42797 34338 42809 34394
rect 42729 34336 42809 34338
rect 42741 34022 42797 34336
rect 42925 34280 42981 34478
rect 42913 34278 42993 34280
rect 42913 34222 42925 34278
rect 42981 34222 42993 34278
rect 42913 34220 42993 34222
rect 42925 34022 42981 34220
rect 43109 34164 43165 34478
rect 43242 34280 43310 34610
rect 43687 34288 43743 35522
rect 44135 35363 44881 35375
rect 44135 35307 44503 35363
rect 44559 35307 44881 35363
rect 44135 35295 44881 35307
rect 44135 35042 44191 35295
rect 44503 35042 44559 35295
rect 44825 35042 44881 35295
rect 44123 35040 44203 35042
rect 44123 34920 44135 35040
rect 44191 34920 44203 35040
rect 44123 34918 44203 34920
rect 44491 35040 44571 35042
rect 44491 34920 44503 35040
rect 44559 34920 44571 35040
rect 44491 34918 44571 34920
rect 44813 35040 44893 35042
rect 44813 34919 44825 35040
rect 44881 34919 44893 35040
rect 44135 34910 44191 34918
rect 44503 34910 44559 34918
rect 44813 34917 44893 34919
rect 44825 34909 44881 34917
rect 44319 34742 44375 34750
rect 44687 34742 44743 34750
rect 44307 34740 44796 34742
rect 44307 34620 44319 34740
rect 44375 34620 44687 34740
rect 44743 34620 44796 34740
rect 44307 34618 44796 34620
rect 44319 34610 44375 34618
rect 44687 34610 44796 34618
rect 44215 34544 44295 34554
rect 44215 34488 44227 34544
rect 44283 34488 44295 34544
rect 44215 34478 44295 34488
rect 44399 34544 44479 34554
rect 44399 34488 44411 34544
rect 44467 34488 44479 34544
rect 44399 34478 44479 34488
rect 44583 34544 44663 34554
rect 44583 34488 44595 34544
rect 44651 34488 44663 34544
rect 44583 34478 44663 34488
rect 44227 34396 44283 34478
rect 44215 34394 44295 34396
rect 44215 34338 44227 34394
rect 44283 34338 44295 34394
rect 44215 34336 44295 34338
rect 43242 34278 43322 34280
rect 43242 34222 43254 34278
rect 43310 34222 43322 34278
rect 43242 34220 43322 34222
rect 43685 34278 43745 34288
rect 43685 34222 43687 34278
rect 43743 34222 43745 34278
rect 43097 34162 43177 34164
rect 43097 34106 43109 34162
rect 43165 34106 43177 34162
rect 43097 34104 43177 34106
rect 43109 34022 43165 34104
rect 42729 34012 42809 34022
rect 42729 33956 42741 34012
rect 42797 33956 42809 34012
rect 42729 33946 42809 33956
rect 42913 34012 42993 34022
rect 42913 33956 42925 34012
rect 42981 33956 42993 34012
rect 42913 33946 42993 33956
rect 43097 34012 43177 34022
rect 43097 33956 43109 34012
rect 43165 33956 43177 34012
rect 43097 33946 43177 33956
rect 43242 33890 43310 34220
rect 43685 34210 43745 34222
rect 43201 33882 43310 33890
rect 43189 33880 43310 33882
rect 43189 33760 43201 33880
rect 43257 33760 43310 33880
rect 43189 33758 43310 33760
rect 43201 33750 43257 33758
rect 42504 33493 43400 33505
rect 42504 33437 42516 33493
rect 42572 33437 43334 33493
rect 43390 33437 43400 33493
rect 42504 33425 43400 33437
rect 43687 33267 43743 34210
rect 44227 34022 44283 34336
rect 44411 34280 44467 34478
rect 44399 34278 44479 34280
rect 44399 34222 44411 34278
rect 44467 34222 44479 34278
rect 44399 34220 44479 34222
rect 44411 34022 44467 34220
rect 44595 34164 44651 34478
rect 44728 34280 44796 34610
rect 44728 34278 44808 34280
rect 44728 34222 44740 34278
rect 44796 34222 44808 34278
rect 44728 34220 44808 34222
rect 44995 34278 45065 34290
rect 45695 34278 45751 38285
rect 44995 34222 44997 34278
rect 45053 34222 45751 34278
rect 44583 34162 44663 34164
rect 44583 34106 44595 34162
rect 44651 34106 44663 34162
rect 44583 34104 44663 34106
rect 44595 34022 44651 34104
rect 44215 34012 44295 34022
rect 44215 33956 44227 34012
rect 44283 33956 44295 34012
rect 44215 33946 44295 33956
rect 44399 34012 44479 34022
rect 44399 33956 44411 34012
rect 44467 33956 44479 34012
rect 44399 33946 44479 33956
rect 44583 34012 44663 34022
rect 44583 33956 44595 34012
rect 44651 33956 44663 34012
rect 44583 33946 44663 33956
rect 44728 33890 44796 34220
rect 44995 34212 45065 34222
rect 44687 33882 44796 33890
rect 44675 33880 44796 33882
rect 44675 33760 44687 33880
rect 44743 33760 44796 33880
rect 44675 33758 44796 33760
rect 44687 33750 44743 33758
rect 43990 33493 44886 33505
rect 43990 33437 44002 33493
rect 44058 33437 44820 33493
rect 44876 33437 44886 33493
rect 43990 33425 44886 33437
rect 44997 33268 45053 34212
rect 45161 33376 45241 33386
rect 45161 33320 45173 33376
rect 45229 33320 45241 33376
rect 45161 33318 45241 33320
rect 43685 33265 43755 33267
rect 43685 33209 43687 33265
rect 43743 33209 43755 33265
rect 43685 33197 43755 33209
rect 44985 33266 45065 33268
rect 44985 33210 44997 33266
rect 45053 33210 45065 33266
rect 44985 33198 45065 33210
rect 42649 33158 43395 33170
rect 42649 33102 43017 33158
rect 43073 33102 43395 33158
rect 42649 33090 43395 33102
rect 42649 32837 42705 33090
rect 43017 32837 43073 33090
rect 43339 32837 43395 33090
rect 44135 33159 44881 33171
rect 44135 33103 44503 33159
rect 44559 33103 44881 33159
rect 44135 33091 44881 33103
rect 44135 32838 44191 33091
rect 44503 32838 44559 33091
rect 44825 32838 44881 33091
rect 42637 32835 42717 32837
rect 42637 32715 42649 32835
rect 42705 32715 42717 32835
rect 42637 32713 42717 32715
rect 43005 32835 43085 32837
rect 43005 32715 43017 32835
rect 43073 32715 43085 32835
rect 43005 32713 43085 32715
rect 43327 32835 43407 32837
rect 43327 32714 43339 32835
rect 43395 32714 43407 32835
rect 44123 32836 44203 32838
rect 44123 32716 44135 32836
rect 44191 32716 44203 32836
rect 44123 32714 44203 32716
rect 44491 32836 44571 32838
rect 44491 32716 44503 32836
rect 44559 32716 44571 32836
rect 44491 32714 44571 32716
rect 44813 32836 44893 32838
rect 44813 32715 44825 32836
rect 44881 32715 44893 32836
rect 42649 32705 42705 32713
rect 43017 32705 43073 32713
rect 43327 32712 43407 32714
rect 43339 32704 43395 32712
rect 44135 32706 44191 32714
rect 44503 32706 44559 32714
rect 44813 32713 44893 32715
rect 44825 32705 44881 32713
rect 42833 32537 42889 32545
rect 43201 32537 43257 32545
rect 44319 32538 44375 32546
rect 44687 32538 44743 32546
rect 42821 32535 43310 32537
rect 42821 32415 42833 32535
rect 42889 32415 43201 32535
rect 43257 32415 43310 32535
rect 42821 32413 43310 32415
rect 44307 32536 44796 32538
rect 44307 32416 44319 32536
rect 44375 32416 44687 32536
rect 44743 32416 44796 32536
rect 44307 32414 44796 32416
rect 42833 32405 42889 32413
rect 43201 32405 43310 32413
rect 44319 32406 44375 32414
rect 44687 32406 44796 32414
rect 42729 32339 42809 32349
rect 42729 32283 42741 32339
rect 42797 32283 42809 32339
rect 42729 32273 42809 32283
rect 42913 32339 42993 32349
rect 42913 32283 42925 32339
rect 42981 32283 42993 32339
rect 42913 32273 42993 32283
rect 43097 32339 43177 32349
rect 43097 32283 43109 32339
rect 43165 32283 43177 32339
rect 43097 32273 43177 32283
rect 42741 32191 42797 32273
rect 42729 32189 42809 32191
rect 42729 32133 42741 32189
rect 42797 32133 42809 32189
rect 42729 32131 42809 32133
rect 42057 31957 42127 31969
rect 42057 31901 42069 31957
rect 42125 31901 42127 31957
rect 42057 31889 42127 31901
rect 42741 31817 42797 32131
rect 42925 32075 42981 32273
rect 42913 32073 42993 32075
rect 42913 32017 42925 32073
rect 42981 32017 42993 32073
rect 42913 32015 42993 32017
rect 42925 31817 42981 32015
rect 43109 31959 43165 32273
rect 43242 32075 43310 32405
rect 44215 32340 44295 32350
rect 44215 32284 44227 32340
rect 44283 32284 44295 32340
rect 44215 32274 44295 32284
rect 44399 32340 44479 32350
rect 44399 32284 44411 32340
rect 44467 32284 44479 32340
rect 44399 32274 44479 32284
rect 44583 32340 44663 32350
rect 44583 32284 44595 32340
rect 44651 32284 44663 32340
rect 44583 32274 44663 32284
rect 44227 32192 44283 32274
rect 44215 32190 44295 32192
rect 44215 32134 44227 32190
rect 44283 32134 44295 32190
rect 44215 32132 44295 32134
rect 43242 32073 43322 32075
rect 43242 32017 43254 32073
rect 43310 32017 43322 32073
rect 43242 32015 43322 32017
rect 43509 32073 43579 32085
rect 43509 32017 43511 32073
rect 43567 32017 43579 32073
rect 43097 31957 43177 31959
rect 43097 31901 43109 31957
rect 43165 31901 43177 31957
rect 43097 31899 43177 31901
rect 43109 31817 43165 31899
rect 42729 31807 42809 31817
rect 42729 31751 42741 31807
rect 42797 31751 42809 31807
rect 42729 31741 42809 31751
rect 42913 31807 42993 31817
rect 42913 31751 42925 31807
rect 42981 31751 42993 31807
rect 42913 31741 42993 31751
rect 43097 31807 43177 31817
rect 43097 31751 43109 31807
rect 43165 31751 43177 31807
rect 43097 31741 43177 31751
rect 43242 31685 43310 32015
rect 43509 32007 43579 32017
rect 43201 31677 43310 31685
rect 43189 31675 43310 31677
rect 43189 31555 43201 31675
rect 43257 31555 43310 31675
rect 43189 31553 43310 31555
rect 43201 31545 43257 31553
rect 42504 31288 43400 31300
rect 42504 31232 42516 31288
rect 42572 31232 43334 31288
rect 43390 31232 43400 31288
rect 42504 31220 43400 31232
rect 43511 31063 43567 32007
rect 44227 31818 44283 32132
rect 44411 32076 44467 32274
rect 44399 32074 44479 32076
rect 44399 32018 44411 32074
rect 44467 32018 44479 32074
rect 44399 32016 44479 32018
rect 44411 31818 44467 32016
rect 44595 31960 44651 32274
rect 44728 32076 44796 32406
rect 45173 32084 45229 33318
rect 44728 32074 44808 32076
rect 44728 32018 44740 32074
rect 44796 32018 44808 32074
rect 44728 32016 44808 32018
rect 45171 32074 45241 32084
rect 45171 32018 45173 32074
rect 45229 32018 45321 32074
rect 44583 31958 44663 31960
rect 44583 31902 44595 31958
rect 44651 31902 44663 31958
rect 44583 31900 44663 31902
rect 44595 31818 44651 31900
rect 44215 31808 44295 31818
rect 44215 31752 44227 31808
rect 44283 31752 44295 31808
rect 44215 31742 44295 31752
rect 44399 31808 44479 31818
rect 44399 31752 44411 31808
rect 44467 31752 44479 31808
rect 44399 31742 44479 31752
rect 44583 31808 44663 31818
rect 44583 31752 44595 31808
rect 44651 31752 44663 31808
rect 44583 31742 44663 31752
rect 44728 31686 44796 32016
rect 45171 32006 45241 32018
rect 44687 31678 44796 31686
rect 44675 31676 44796 31678
rect 44675 31556 44687 31676
rect 44743 31556 44796 31676
rect 44675 31554 44796 31556
rect 44687 31546 44743 31554
rect 43990 31289 44886 31301
rect 43990 31233 44002 31289
rect 44058 31233 44820 31289
rect 44876 31233 44886 31289
rect 43990 31221 44886 31233
rect 43675 31170 43755 31180
rect 43675 31114 43687 31170
rect 43743 31114 43755 31170
rect 43675 31112 43755 31114
rect 43509 31060 43579 31063
rect 43509 31006 43511 31060
rect 43567 31006 43579 31060
rect 43509 30994 43579 31006
rect 42649 30953 43395 30965
rect 42649 30897 43017 30953
rect 43073 30897 43395 30953
rect 42649 30885 43395 30897
rect 42649 30632 42705 30885
rect 43017 30632 43073 30885
rect 43339 30632 43395 30885
rect 42637 30630 42717 30632
rect 42637 30510 42649 30630
rect 42705 30510 42717 30630
rect 42637 30508 42717 30510
rect 43005 30630 43085 30632
rect 43005 30510 43017 30630
rect 43073 30510 43085 30630
rect 43005 30508 43085 30510
rect 43327 30630 43407 30632
rect 43327 30509 43339 30630
rect 43395 30509 43407 30630
rect 42649 30500 42705 30508
rect 43017 30500 43073 30508
rect 43327 30507 43407 30509
rect 43339 30499 43395 30507
rect 42833 30332 42889 30340
rect 43201 30332 43257 30340
rect 42821 30330 43310 30332
rect 42821 30210 42833 30330
rect 42889 30210 43201 30330
rect 43257 30210 43310 30330
rect 42821 30208 43310 30210
rect 42833 30200 42889 30208
rect 43201 30200 43310 30208
rect 42729 30134 42809 30144
rect 42729 30078 42741 30134
rect 42797 30078 42809 30134
rect 42729 30068 42809 30078
rect 42913 30134 42993 30144
rect 42913 30078 42925 30134
rect 42981 30078 42993 30134
rect 42913 30068 42993 30078
rect 43097 30134 43177 30144
rect 43097 30078 43109 30134
rect 43165 30078 43177 30134
rect 43097 30068 43177 30078
rect 42741 29986 42797 30068
rect 42729 29984 42809 29986
rect 42729 29928 42741 29984
rect 42797 29928 42809 29984
rect 42729 29926 42809 29928
rect 41921 29868 41991 29882
rect 41921 29812 41933 29868
rect 41989 29812 41991 29868
rect 41921 29800 41991 29812
rect 41687 29752 41765 29763
rect 41295 29751 41765 29752
rect 41295 29697 41699 29751
rect 41753 29697 41765 29751
rect 41295 29696 41765 29697
rect 39723 29392 40895 29402
rect 39723 29336 39735 29392
rect 39791 29336 40623 29392
rect 40679 29336 40895 29392
rect 39723 29326 40895 29336
rect 41295 29392 41375 29696
rect 41687 29685 41765 29696
rect 41295 29336 41307 29392
rect 41363 29336 41375 29392
rect 41295 29326 41375 29336
rect 39653 29014 41445 29026
rect 39653 28874 39665 29014
rect 41433 28874 41445 29014
rect 41738 28965 41824 28977
rect 41933 28969 41989 29800
rect 42741 29612 42797 29926
rect 42925 29870 42981 30068
rect 42913 29868 42993 29870
rect 42913 29812 42925 29868
rect 42981 29812 42993 29868
rect 42913 29810 42993 29812
rect 42925 29612 42981 29810
rect 43109 29754 43165 30068
rect 43242 29870 43310 30200
rect 43687 29880 43743 31112
rect 43242 29868 43322 29870
rect 43242 29812 43254 29868
rect 43310 29812 43322 29868
rect 43242 29810 43322 29812
rect 43685 29868 43745 29880
rect 43685 29812 43687 29868
rect 43743 29812 43745 29868
rect 43097 29752 43177 29754
rect 43097 29696 43109 29752
rect 43165 29696 43177 29752
rect 43097 29694 43177 29696
rect 43109 29612 43165 29694
rect 42729 29602 42809 29612
rect 42729 29546 42741 29602
rect 42797 29546 42809 29602
rect 42729 29536 42809 29546
rect 42913 29602 42993 29612
rect 42913 29546 42925 29602
rect 42981 29546 42993 29602
rect 42913 29536 42993 29546
rect 43097 29602 43177 29612
rect 43097 29546 43109 29602
rect 43165 29546 43177 29602
rect 43097 29536 43177 29546
rect 43242 29480 43310 29810
rect 43685 29800 43745 29812
rect 43201 29472 43310 29480
rect 43189 29470 43310 29472
rect 43189 29350 43201 29470
rect 43257 29350 43310 29470
rect 43189 29348 43310 29350
rect 43201 29340 43257 29348
rect 42504 29083 43402 29095
rect 42504 29027 42516 29083
rect 42572 29027 43334 29083
rect 43390 29027 43402 29083
rect 42504 29015 43402 29027
rect 41738 28909 41750 28965
rect 41806 28909 41824 28965
rect 41738 28897 41824 28909
rect 41931 28965 41991 28969
rect 41931 28909 41933 28965
rect 41989 28909 41991 28965
rect 41931 28897 41991 28909
rect 39653 28862 41445 28874
rect 39067 28532 39424 28588
rect 41023 28690 41343 28700
rect 38587 28172 38599 28228
rect 38655 28172 38667 28228
rect 38587 28162 38667 28172
rect 39067 28228 39147 28532
rect 39067 28172 39079 28228
rect 39135 28172 39147 28228
rect 39067 28162 39147 28172
rect 37699 27914 38463 27986
rect 41023 27890 41033 28690
rect 41333 27890 41343 28690
rect 41023 27880 41343 27890
rect 15195 26389 36275 26445
rect 11151 25898 11221 25900
rect 11151 25842 11153 25898
rect 11209 25842 11221 25898
rect 11151 25840 11221 25842
rect 7335 25722 7405 25734
rect 7335 25666 7347 25722
rect 7403 25666 7405 25722
rect 7335 25664 7405 25666
rect 7109 21972 7179 21984
rect 7109 21916 7111 21972
rect 7167 21916 7179 21972
rect 7109 21904 7179 21916
rect 7347 21072 7403 25664
rect 8199 25262 8945 25274
rect 8199 25206 8567 25262
rect 8623 25206 8945 25262
rect 8199 25194 8945 25206
rect 8199 24941 8255 25194
rect 8567 24941 8623 25194
rect 8889 24941 8945 25194
rect 8187 24939 8267 24941
rect 8187 24819 8199 24939
rect 8255 24819 8267 24939
rect 8187 24817 8267 24819
rect 8555 24939 8635 24941
rect 8555 24819 8567 24939
rect 8623 24819 8635 24939
rect 8555 24817 8635 24819
rect 8877 24939 8957 24941
rect 8877 24818 8889 24939
rect 8945 24818 8957 24939
rect 8199 24809 8255 24817
rect 8567 24809 8623 24817
rect 8877 24816 8957 24818
rect 8889 24808 8945 24816
rect 8383 24641 8439 24649
rect 8751 24641 8807 24649
rect 8371 24639 8860 24641
rect 8371 24519 8383 24639
rect 8439 24519 8751 24639
rect 8807 24519 8860 24639
rect 8371 24517 8860 24519
rect 8383 24509 8439 24517
rect 8751 24509 8860 24517
rect 8279 24443 8359 24453
rect 8279 24387 8291 24443
rect 8347 24387 8359 24443
rect 8279 24377 8359 24387
rect 8463 24443 8543 24453
rect 8463 24387 8475 24443
rect 8531 24387 8543 24443
rect 8463 24377 8543 24387
rect 8647 24443 8727 24453
rect 8647 24387 8659 24443
rect 8715 24387 8727 24443
rect 8647 24377 8727 24387
rect 8291 24295 8347 24377
rect 8279 24293 8359 24295
rect 8279 24237 8291 24293
rect 8347 24237 8359 24293
rect 8279 24235 8359 24237
rect 7607 24177 7677 24189
rect 7607 24121 7619 24177
rect 7675 24121 7677 24177
rect 7607 24109 7677 24121
rect 7471 21972 7541 21986
rect 7471 21916 7483 21972
rect 7539 21916 7541 21972
rect 7471 21904 7541 21916
rect 7335 21070 7405 21072
rect 7335 21014 7347 21070
rect 7403 21014 7405 21070
rect 7335 21002 7405 21014
rect 7483 17576 7539 21904
rect 7619 19663 7675 24109
rect 8291 23921 8347 24235
rect 8475 24179 8531 24377
rect 8463 24177 8543 24179
rect 8463 24121 8475 24177
rect 8531 24121 8543 24177
rect 8463 24119 8543 24121
rect 8475 23921 8531 24119
rect 8659 24063 8715 24377
rect 8792 24179 8860 24509
rect 10939 24293 11009 24305
rect 10939 24237 10951 24293
rect 11007 24237 11009 24293
rect 10939 24235 11009 24237
rect 8792 24177 8872 24179
rect 8792 24121 8804 24177
rect 8860 24121 8872 24177
rect 8792 24119 8872 24121
rect 9059 24177 9129 24189
rect 9059 24121 9061 24177
rect 9117 24121 9129 24177
rect 8647 24061 8727 24063
rect 8647 24005 8659 24061
rect 8715 24005 8727 24061
rect 8647 24003 8727 24005
rect 8659 23921 8715 24003
rect 8279 23911 8359 23921
rect 8279 23855 8291 23911
rect 8347 23855 8359 23911
rect 8279 23845 8359 23855
rect 8463 23911 8543 23921
rect 8463 23855 8475 23911
rect 8531 23855 8543 23911
rect 8463 23845 8543 23855
rect 8647 23911 8727 23921
rect 8647 23855 8659 23911
rect 8715 23855 8727 23911
rect 8647 23845 8727 23855
rect 8792 23789 8860 24119
rect 9059 24111 9129 24121
rect 8751 23781 8860 23789
rect 8739 23779 8860 23781
rect 8739 23659 8751 23779
rect 8807 23659 8860 23779
rect 8739 23657 8860 23659
rect 8751 23649 8807 23657
rect 8054 23392 8952 23404
rect 8054 23336 8066 23392
rect 8122 23336 8884 23392
rect 8940 23336 8952 23392
rect 8054 23324 8952 23336
rect 9061 23167 9117 24111
rect 9225 23274 9305 23284
rect 9225 23218 9237 23274
rect 9293 23218 9305 23274
rect 9225 23216 9305 23218
rect 9059 23164 9129 23167
rect 9059 23110 9061 23164
rect 9117 23110 9129 23164
rect 9059 23098 9129 23110
rect 8199 23057 8945 23069
rect 8199 23001 8567 23057
rect 8623 23001 8945 23057
rect 8199 22989 8945 23001
rect 8199 22736 8255 22989
rect 8567 22736 8623 22989
rect 8889 22736 8945 22989
rect 8187 22734 8267 22736
rect 8187 22614 8199 22734
rect 8255 22614 8267 22734
rect 8187 22612 8267 22614
rect 8555 22734 8635 22736
rect 8555 22614 8567 22734
rect 8623 22614 8635 22734
rect 8555 22612 8635 22614
rect 8877 22734 8957 22736
rect 8877 22613 8889 22734
rect 8945 22613 8957 22734
rect 8199 22604 8255 22612
rect 8567 22604 8623 22612
rect 8877 22611 8957 22613
rect 8889 22603 8945 22611
rect 8383 22436 8439 22444
rect 8751 22436 8807 22444
rect 8371 22434 8860 22436
rect 8371 22314 8383 22434
rect 8439 22314 8751 22434
rect 8807 22314 8860 22434
rect 8371 22312 8860 22314
rect 8383 22304 8439 22312
rect 8751 22304 8860 22312
rect 8279 22238 8359 22248
rect 8279 22182 8291 22238
rect 8347 22182 8359 22238
rect 8279 22172 8359 22182
rect 8463 22238 8543 22248
rect 8463 22182 8475 22238
rect 8531 22182 8543 22238
rect 8463 22172 8543 22182
rect 8647 22238 8727 22248
rect 8647 22182 8659 22238
rect 8715 22182 8727 22238
rect 8647 22172 8727 22182
rect 8291 22090 8347 22172
rect 8279 22088 8359 22090
rect 8279 22032 8291 22088
rect 8347 22032 8359 22088
rect 8279 22030 8359 22032
rect 8291 21716 8347 22030
rect 8475 21974 8531 22172
rect 8463 21972 8543 21974
rect 8463 21916 8475 21972
rect 8531 21916 8543 21972
rect 8463 21914 8543 21916
rect 8475 21716 8531 21914
rect 8659 21858 8715 22172
rect 8792 21974 8860 22304
rect 9237 21982 9293 23216
rect 9685 23057 10431 23069
rect 9685 23001 10053 23057
rect 10109 23001 10431 23057
rect 9685 22989 10431 23001
rect 9685 22736 9741 22989
rect 10053 22736 10109 22989
rect 10375 22736 10431 22989
rect 9673 22734 9753 22736
rect 9673 22614 9685 22734
rect 9741 22614 9753 22734
rect 9673 22612 9753 22614
rect 10041 22734 10121 22736
rect 10041 22614 10053 22734
rect 10109 22614 10121 22734
rect 10041 22612 10121 22614
rect 10363 22734 10443 22736
rect 10363 22613 10375 22734
rect 10431 22613 10443 22734
rect 9685 22604 9741 22612
rect 10053 22604 10109 22612
rect 10363 22611 10443 22613
rect 10375 22603 10431 22611
rect 9869 22436 9925 22444
rect 10237 22436 10293 22444
rect 9857 22434 10346 22436
rect 9857 22314 9869 22434
rect 9925 22314 10237 22434
rect 10293 22314 10346 22434
rect 9857 22312 10346 22314
rect 9869 22304 9925 22312
rect 10237 22304 10346 22312
rect 9765 22238 9845 22248
rect 9765 22182 9777 22238
rect 9833 22182 9845 22238
rect 9765 22172 9845 22182
rect 9949 22238 10029 22248
rect 9949 22182 9961 22238
rect 10017 22182 10029 22238
rect 9949 22172 10029 22182
rect 10133 22238 10213 22248
rect 10133 22182 10145 22238
rect 10201 22182 10213 22238
rect 10133 22172 10213 22182
rect 9777 22090 9833 22172
rect 9765 22088 9845 22090
rect 9765 22032 9777 22088
rect 9833 22032 9845 22088
rect 9765 22030 9845 22032
rect 8792 21972 8872 21974
rect 8792 21916 8804 21972
rect 8860 21916 8872 21972
rect 8792 21914 8872 21916
rect 9235 21972 9295 21982
rect 9235 21916 9237 21972
rect 9293 21916 9295 21972
rect 8647 21856 8727 21858
rect 8647 21800 8659 21856
rect 8715 21800 8727 21856
rect 8647 21798 8727 21800
rect 8659 21716 8715 21798
rect 8279 21706 8359 21716
rect 8279 21650 8291 21706
rect 8347 21650 8359 21706
rect 8279 21640 8359 21650
rect 8463 21706 8543 21716
rect 8463 21650 8475 21706
rect 8531 21650 8543 21706
rect 8463 21640 8543 21650
rect 8647 21706 8727 21716
rect 8647 21650 8659 21706
rect 8715 21650 8727 21706
rect 8647 21640 8727 21650
rect 8792 21584 8860 21914
rect 9235 21904 9295 21916
rect 8751 21576 8860 21584
rect 8739 21574 8860 21576
rect 8739 21454 8751 21574
rect 8807 21454 8860 21574
rect 8739 21452 8860 21454
rect 8751 21444 8807 21452
rect 8054 21187 8950 21199
rect 8054 21131 8066 21187
rect 8122 21131 8884 21187
rect 8940 21131 8950 21187
rect 8054 21119 8950 21131
rect 9237 20961 9293 21904
rect 9777 21716 9833 22030
rect 9961 21974 10017 22172
rect 9949 21972 10029 21974
rect 9949 21916 9961 21972
rect 10017 21916 10029 21972
rect 9949 21914 10029 21916
rect 9961 21716 10017 21914
rect 10145 21858 10201 22172
rect 10278 21974 10346 22304
rect 10278 21972 10358 21974
rect 10278 21916 10290 21972
rect 10346 21916 10358 21972
rect 10278 21914 10358 21916
rect 10545 21972 10615 21984
rect 10545 21916 10547 21972
rect 10603 21916 10871 21972
rect 10133 21856 10213 21858
rect 10133 21800 10145 21856
rect 10201 21800 10213 21856
rect 10133 21798 10213 21800
rect 10145 21716 10201 21798
rect 9765 21706 9845 21716
rect 9765 21650 9777 21706
rect 9833 21650 9845 21706
rect 9765 21640 9845 21650
rect 9949 21706 10029 21716
rect 9949 21650 9961 21706
rect 10017 21650 10029 21706
rect 9949 21640 10029 21650
rect 10133 21706 10213 21716
rect 10133 21650 10145 21706
rect 10201 21650 10213 21706
rect 10133 21640 10213 21650
rect 10278 21584 10346 21914
rect 10545 21906 10615 21916
rect 10237 21576 10346 21584
rect 10225 21574 10346 21576
rect 10225 21454 10237 21574
rect 10293 21454 10346 21574
rect 10225 21452 10346 21454
rect 10237 21444 10293 21452
rect 9540 21187 10436 21199
rect 9540 21131 9552 21187
rect 9608 21131 10370 21187
rect 10426 21131 10436 21187
rect 9540 21119 10436 21131
rect 10547 20962 10603 21906
rect 10711 21070 10791 21080
rect 10711 21014 10723 21070
rect 10779 21014 10791 21070
rect 10711 21012 10791 21014
rect 9235 20959 9305 20961
rect 9235 20903 9237 20959
rect 9293 20903 9305 20959
rect 9235 20891 9305 20903
rect 10535 20960 10615 20962
rect 10535 20904 10547 20960
rect 10603 20904 10615 20960
rect 10535 20892 10615 20904
rect 8199 20852 8945 20864
rect 8199 20796 8567 20852
rect 8623 20796 8945 20852
rect 8199 20784 8945 20796
rect 8199 20531 8255 20784
rect 8567 20531 8623 20784
rect 8889 20531 8945 20784
rect 9685 20853 10431 20865
rect 9685 20797 10053 20853
rect 10109 20797 10431 20853
rect 9685 20785 10431 20797
rect 9685 20532 9741 20785
rect 10053 20532 10109 20785
rect 10375 20532 10431 20785
rect 8187 20529 8267 20531
rect 8187 20409 8199 20529
rect 8255 20409 8267 20529
rect 8187 20407 8267 20409
rect 8555 20529 8635 20531
rect 8555 20409 8567 20529
rect 8623 20409 8635 20529
rect 8555 20407 8635 20409
rect 8877 20529 8957 20531
rect 8877 20408 8889 20529
rect 8945 20408 8957 20529
rect 9673 20530 9753 20532
rect 9673 20410 9685 20530
rect 9741 20410 9753 20530
rect 9673 20408 9753 20410
rect 10041 20530 10121 20532
rect 10041 20410 10053 20530
rect 10109 20410 10121 20530
rect 10041 20408 10121 20410
rect 10363 20530 10443 20532
rect 10363 20409 10375 20530
rect 10431 20409 10443 20530
rect 8199 20399 8255 20407
rect 8567 20399 8623 20407
rect 8877 20406 8957 20408
rect 8889 20398 8945 20406
rect 9685 20400 9741 20408
rect 10053 20400 10109 20408
rect 10363 20407 10443 20409
rect 10375 20399 10431 20407
rect 8383 20231 8439 20239
rect 8751 20231 8807 20239
rect 9869 20232 9925 20240
rect 10237 20232 10293 20240
rect 8371 20229 8860 20231
rect 8371 20109 8383 20229
rect 8439 20109 8751 20229
rect 8807 20109 8860 20229
rect 8371 20107 8860 20109
rect 9857 20230 10346 20232
rect 9857 20110 9869 20230
rect 9925 20110 10237 20230
rect 10293 20110 10346 20230
rect 9857 20108 10346 20110
rect 8383 20099 8439 20107
rect 8751 20099 8860 20107
rect 9869 20100 9925 20108
rect 10237 20100 10346 20108
rect 8279 20033 8359 20043
rect 8279 19977 8291 20033
rect 8347 19977 8359 20033
rect 8279 19967 8359 19977
rect 8463 20033 8543 20043
rect 8463 19977 8475 20033
rect 8531 19977 8543 20033
rect 8463 19967 8543 19977
rect 8647 20033 8727 20043
rect 8647 19977 8659 20033
rect 8715 19977 8727 20033
rect 8647 19967 8727 19977
rect 8291 19885 8347 19967
rect 8279 19883 8359 19885
rect 8279 19827 8291 19883
rect 8347 19827 8359 19883
rect 8279 19825 8359 19827
rect 7607 19651 7677 19663
rect 7607 19595 7619 19651
rect 7675 19595 7677 19651
rect 7607 19583 7677 19595
rect 8291 19511 8347 19825
rect 8475 19769 8531 19967
rect 8463 19767 8543 19769
rect 8463 19711 8475 19767
rect 8531 19711 8543 19767
rect 8463 19709 8543 19711
rect 8475 19511 8531 19709
rect 8659 19653 8715 19967
rect 8792 19769 8860 20099
rect 9765 20034 9845 20044
rect 9765 19978 9777 20034
rect 9833 19978 9845 20034
rect 9765 19968 9845 19978
rect 9949 20034 10029 20044
rect 9949 19978 9961 20034
rect 10017 19978 10029 20034
rect 9949 19968 10029 19978
rect 10133 20034 10213 20044
rect 10133 19978 10145 20034
rect 10201 19978 10213 20034
rect 10133 19968 10213 19978
rect 9777 19886 9833 19968
rect 9765 19884 9845 19886
rect 9765 19828 9777 19884
rect 9833 19828 9845 19884
rect 9765 19826 9845 19828
rect 8792 19767 8872 19769
rect 8792 19711 8804 19767
rect 8860 19711 8872 19767
rect 8792 19709 8872 19711
rect 9059 19767 9129 19779
rect 9059 19711 9061 19767
rect 9117 19711 9129 19767
rect 8647 19651 8727 19653
rect 8647 19595 8659 19651
rect 8715 19595 8727 19651
rect 8647 19593 8727 19595
rect 8659 19511 8715 19593
rect 8279 19501 8359 19511
rect 8279 19445 8291 19501
rect 8347 19445 8359 19501
rect 8279 19435 8359 19445
rect 8463 19501 8543 19511
rect 8463 19445 8475 19501
rect 8531 19445 8543 19501
rect 8463 19435 8543 19445
rect 8647 19501 8727 19511
rect 8647 19445 8659 19501
rect 8715 19445 8727 19501
rect 8647 19435 8727 19445
rect 8792 19379 8860 19709
rect 9059 19701 9129 19711
rect 8751 19371 8860 19379
rect 8739 19369 8860 19371
rect 8739 19249 8751 19369
rect 8807 19249 8860 19369
rect 8739 19247 8860 19249
rect 8751 19239 8807 19247
rect 8054 18982 8950 18994
rect 8054 18926 8066 18982
rect 8122 18926 8884 18982
rect 8940 18926 8950 18982
rect 8054 18914 8950 18926
rect 9061 18757 9117 19701
rect 9777 19512 9833 19826
rect 9961 19770 10017 19968
rect 9949 19768 10029 19770
rect 9949 19712 9961 19768
rect 10017 19712 10029 19768
rect 9949 19710 10029 19712
rect 9961 19512 10017 19710
rect 10145 19654 10201 19968
rect 10278 19770 10346 20100
rect 10723 19778 10779 21012
rect 10278 19768 10358 19770
rect 10278 19712 10290 19768
rect 10346 19712 10358 19768
rect 10278 19710 10358 19712
rect 10721 19768 10791 19778
rect 10721 19712 10723 19768
rect 10779 19712 10871 19768
rect 10133 19652 10213 19654
rect 10133 19596 10145 19652
rect 10201 19596 10213 19652
rect 10133 19594 10213 19596
rect 10145 19512 10201 19594
rect 9765 19502 9845 19512
rect 9765 19446 9777 19502
rect 9833 19446 9845 19502
rect 9765 19436 9845 19446
rect 9949 19502 10029 19512
rect 9949 19446 9961 19502
rect 10017 19446 10029 19502
rect 9949 19436 10029 19446
rect 10133 19502 10213 19512
rect 10133 19446 10145 19502
rect 10201 19446 10213 19502
rect 10133 19436 10213 19446
rect 10278 19380 10346 19710
rect 10721 19700 10791 19712
rect 10237 19372 10346 19380
rect 10225 19370 10346 19372
rect 10225 19250 10237 19370
rect 10293 19250 10346 19370
rect 10225 19248 10346 19250
rect 10237 19240 10293 19248
rect 9540 18983 10436 18995
rect 9540 18927 9552 18983
rect 9608 18927 10370 18983
rect 10426 18927 10436 18983
rect 9540 18915 10436 18927
rect 9225 18864 9305 18874
rect 9225 18808 9237 18864
rect 9293 18808 9305 18864
rect 9225 18806 9305 18808
rect 9059 18754 9129 18757
rect 9059 18700 9061 18754
rect 9117 18700 9129 18754
rect 9059 18688 9129 18700
rect 8199 18647 8945 18659
rect 8199 18591 8567 18647
rect 8623 18591 8945 18647
rect 8199 18579 8945 18591
rect 8199 18326 8255 18579
rect 8567 18326 8623 18579
rect 8889 18326 8945 18579
rect 8187 18324 8267 18326
rect 8187 18204 8199 18324
rect 8255 18204 8267 18324
rect 8187 18202 8267 18204
rect 8555 18324 8635 18326
rect 8555 18204 8567 18324
rect 8623 18204 8635 18324
rect 8555 18202 8635 18204
rect 8877 18324 8957 18326
rect 8877 18203 8889 18324
rect 8945 18203 8957 18324
rect 8199 18194 8255 18202
rect 8567 18194 8623 18202
rect 8877 18201 8957 18203
rect 8889 18193 8945 18201
rect 8383 18026 8439 18034
rect 8751 18026 8807 18034
rect 8371 18024 8860 18026
rect 8371 17904 8383 18024
rect 8439 17904 8751 18024
rect 8807 17904 8860 18024
rect 8371 17902 8860 17904
rect 8383 17894 8439 17902
rect 8751 17894 8860 17902
rect 8279 17828 8359 17838
rect 8279 17772 8291 17828
rect 8347 17772 8359 17828
rect 8279 17762 8359 17772
rect 8463 17828 8543 17838
rect 8463 17772 8475 17828
rect 8531 17772 8543 17828
rect 8463 17762 8543 17772
rect 8647 17828 8727 17838
rect 8647 17772 8659 17828
rect 8715 17772 8727 17828
rect 8647 17762 8727 17772
rect 8291 17680 8347 17762
rect 8279 17678 8359 17680
rect 8279 17622 8291 17678
rect 8347 17622 8359 17678
rect 8279 17620 8359 17622
rect 7471 17562 7541 17576
rect 7471 17506 7483 17562
rect 7539 17506 7541 17562
rect 7471 17494 7541 17506
rect 7169 16659 7239 16671
rect 7483 16663 7539 17494
rect 8291 17306 8347 17620
rect 8475 17564 8531 17762
rect 8463 17562 8543 17564
rect 8463 17506 8475 17562
rect 8531 17506 8543 17562
rect 8463 17504 8543 17506
rect 8475 17306 8531 17504
rect 8659 17448 8715 17762
rect 8792 17564 8860 17894
rect 9237 17574 9293 18806
rect 8792 17562 8872 17564
rect 8792 17506 8804 17562
rect 8860 17506 8872 17562
rect 8792 17504 8872 17506
rect 9235 17562 9295 17574
rect 9235 17506 9237 17562
rect 9293 17506 9295 17562
rect 8647 17446 8727 17448
rect 8647 17390 8659 17446
rect 8715 17390 8727 17446
rect 8647 17388 8727 17390
rect 8659 17306 8715 17388
rect 8279 17296 8359 17306
rect 8279 17240 8291 17296
rect 8347 17240 8359 17296
rect 8279 17230 8359 17240
rect 8463 17296 8543 17306
rect 8463 17240 8475 17296
rect 8531 17240 8543 17296
rect 8463 17230 8543 17240
rect 8647 17296 8727 17306
rect 8647 17240 8659 17296
rect 8715 17240 8727 17296
rect 8647 17230 8727 17240
rect 8792 17174 8860 17504
rect 9235 17494 9295 17506
rect 10667 17446 10737 17458
rect 10667 17390 10679 17446
rect 10735 17390 10737 17446
rect 10667 17378 10737 17390
rect 8751 17166 8860 17174
rect 8739 17164 8860 17166
rect 8739 17044 8751 17164
rect 8807 17044 8860 17164
rect 8739 17042 8860 17044
rect 8751 17034 8807 17042
rect 8054 16777 8952 16789
rect 8054 16721 8066 16777
rect 8122 16721 8884 16777
rect 8940 16721 8952 16777
rect 8054 16709 8952 16721
rect 7169 16603 7181 16659
rect 7237 16603 7239 16659
rect 7169 16601 7239 16603
rect 7481 16659 7541 16663
rect 7481 16603 7483 16659
rect 7539 16603 7541 16659
rect 7181 15989 7237 16601
rect 7481 16591 7541 16603
rect 10679 16499 10735 17378
rect 10679 16389 10735 16399
rect 7033 11494 7103 11506
rect 7033 11438 7045 11494
rect 7101 11438 7103 11494
rect 7033 11426 7103 11438
rect 6679 10136 6681 10192
rect 6737 10136 6965 10192
rect 6091 10076 6171 10078
rect 6091 10020 6103 10076
rect 6159 10020 6171 10076
rect 6091 10018 6171 10020
rect 6103 9936 6159 10018
rect 5723 9926 5803 9936
rect 5723 9870 5735 9926
rect 5791 9870 5803 9926
rect 5723 9860 5803 9870
rect 5907 9926 5987 9936
rect 5907 9870 5919 9926
rect 5975 9870 5987 9926
rect 5907 9860 5987 9870
rect 6091 9926 6171 9936
rect 6091 9870 6103 9926
rect 6159 9870 6171 9926
rect 6091 9860 6171 9870
rect 6236 9804 6304 10134
rect 6679 10124 6749 10136
rect 6195 9796 6304 9804
rect 6183 9794 6304 9796
rect 6183 9674 6195 9794
rect 6251 9674 6304 9794
rect 6183 9672 6304 9674
rect 6195 9664 6251 9672
rect 5498 9407 6394 9419
rect 5498 9351 5510 9407
rect 5566 9351 6328 9407
rect 6384 9351 6394 9407
rect 5498 9339 6394 9351
rect 5183 9288 5263 9298
rect 5183 9232 5195 9288
rect 5251 9232 5263 9288
rect 5183 9230 5263 9232
rect 5017 9178 5087 9181
rect 5017 9124 5019 9178
rect 5075 9124 5087 9178
rect 5017 9112 5087 9124
rect 4157 9071 4903 9083
rect 4157 9015 4525 9071
rect 4581 9015 4903 9071
rect 4157 9003 4903 9015
rect 4157 8750 4213 9003
rect 4525 8750 4581 9003
rect 4847 8750 4903 9003
rect 4145 8748 4225 8750
rect 4145 8628 4157 8748
rect 4213 8628 4225 8748
rect 4145 8626 4225 8628
rect 4513 8748 4593 8750
rect 4513 8628 4525 8748
rect 4581 8628 4593 8748
rect 4513 8626 4593 8628
rect 4835 8748 4915 8750
rect 4835 8627 4847 8748
rect 4903 8627 4915 8748
rect 4157 8618 4213 8626
rect 4525 8618 4581 8626
rect 4835 8625 4915 8627
rect 4847 8617 4903 8625
rect 4341 8450 4397 8458
rect 4709 8450 4765 8458
rect 4329 8448 4818 8450
rect 4329 8328 4341 8448
rect 4397 8328 4709 8448
rect 4765 8328 4818 8448
rect 4329 8326 4818 8328
rect 4341 8318 4397 8326
rect 4709 8318 4818 8326
rect 4237 8252 4317 8262
rect 4237 8196 4249 8252
rect 4305 8196 4317 8252
rect 4237 8186 4317 8196
rect 4421 8252 4501 8262
rect 4421 8196 4433 8252
rect 4489 8196 4501 8252
rect 4421 8186 4501 8196
rect 4605 8252 4685 8262
rect 4605 8196 4617 8252
rect 4673 8196 4685 8252
rect 4605 8186 4685 8196
rect 4249 8104 4305 8186
rect 4237 8102 4317 8104
rect 4237 8046 4249 8102
rect 4305 8046 4317 8102
rect 4237 8044 4317 8046
rect 3429 7986 3499 8000
rect 3429 7930 3441 7986
rect 3497 7930 3499 7986
rect 3429 7918 3499 7930
rect 3263 7870 3343 7882
rect 3263 7814 3275 7870
rect 3331 7814 3343 7870
rect 3263 7802 3343 7814
rect 3127 7083 3197 7095
rect 3441 7087 3497 7918
rect 4249 7730 4305 8044
rect 4433 7988 4489 8186
rect 4421 7986 4501 7988
rect 4421 7930 4433 7986
rect 4489 7930 4501 7986
rect 4421 7928 4501 7930
rect 4433 7730 4489 7928
rect 4617 7872 4673 8186
rect 4750 7988 4818 8318
rect 5195 7998 5251 9230
rect 4750 7986 4830 7988
rect 4750 7930 4762 7986
rect 4818 7930 4830 7986
rect 4750 7928 4830 7930
rect 5193 7986 5253 7998
rect 5193 7930 5195 7986
rect 5251 7930 5253 7986
rect 4605 7870 4685 7872
rect 4605 7814 4617 7870
rect 4673 7814 4685 7870
rect 4605 7812 4685 7814
rect 4617 7730 4673 7812
rect 4237 7720 4317 7730
rect 4237 7664 4249 7720
rect 4305 7664 4317 7720
rect 4237 7654 4317 7664
rect 4421 7720 4501 7730
rect 4421 7664 4433 7720
rect 4489 7664 4501 7720
rect 4421 7654 4501 7664
rect 4605 7720 4685 7730
rect 4605 7664 4617 7720
rect 4673 7664 4685 7720
rect 4605 7654 4685 7664
rect 4750 7598 4818 7928
rect 5193 7918 5253 7930
rect 4709 7590 4818 7598
rect 4697 7588 4818 7590
rect 4697 7468 4709 7588
rect 4765 7468 4818 7588
rect 4697 7466 4818 7468
rect 4709 7458 4765 7466
rect 4012 7201 4910 7213
rect 4012 7145 4024 7201
rect 4080 7145 4842 7201
rect 4898 7145 4910 7201
rect 4012 7133 4910 7145
rect 3127 7027 3139 7083
rect 3195 7027 3197 7083
rect 3127 7015 3197 7027
rect 3439 7083 3499 7087
rect 3439 7027 3441 7083
rect 3497 7027 3499 7083
rect 3439 7015 3499 7027
rect 3003 6810 3059 6820
rect 7045 6920 7101 11426
rect 7181 7095 7237 15889
rect 8199 15686 8945 15698
rect 8199 15630 8567 15686
rect 8623 15630 8945 15686
rect 8199 15618 8945 15630
rect 8199 15365 8255 15618
rect 8567 15365 8623 15618
rect 8889 15365 8945 15618
rect 8187 15363 8267 15365
rect 8187 15243 8199 15363
rect 8255 15243 8267 15363
rect 8187 15241 8267 15243
rect 8555 15363 8635 15365
rect 8555 15243 8567 15363
rect 8623 15243 8635 15363
rect 8555 15241 8635 15243
rect 8877 15363 8957 15365
rect 8877 15242 8889 15363
rect 8945 15242 8957 15363
rect 8199 15233 8255 15241
rect 8567 15233 8623 15241
rect 8877 15240 8957 15242
rect 8889 15232 8945 15240
rect 8383 15065 8439 15073
rect 8751 15065 8807 15073
rect 8371 15063 8860 15065
rect 8371 14943 8383 15063
rect 8439 14943 8751 15063
rect 8807 14943 8860 15063
rect 8371 14941 8860 14943
rect 8383 14933 8439 14941
rect 8751 14933 8860 14941
rect 8279 14867 8359 14877
rect 8279 14811 8291 14867
rect 8347 14811 8359 14867
rect 8279 14801 8359 14811
rect 8463 14867 8543 14877
rect 8463 14811 8475 14867
rect 8531 14811 8543 14867
rect 8463 14801 8543 14811
rect 8647 14867 8727 14877
rect 8647 14811 8659 14867
rect 8715 14811 8727 14867
rect 8647 14801 8727 14811
rect 7391 14717 7477 14729
rect 8291 14719 8347 14801
rect 7391 14661 7403 14717
rect 7459 14661 7477 14717
rect 7391 14649 7477 14661
rect 8279 14717 8359 14719
rect 8279 14661 8291 14717
rect 8347 14661 8359 14717
rect 8279 14659 8359 14661
rect 7607 14601 7677 14613
rect 7607 14545 7619 14601
rect 7675 14545 7677 14601
rect 7607 14533 7677 14545
rect 7471 12396 7541 12410
rect 7471 12340 7483 12396
rect 7539 12340 7541 12396
rect 7471 12328 7541 12340
rect 7305 12208 7385 12218
rect 7305 12152 7317 12208
rect 7373 12152 7385 12208
rect 7305 12150 7385 12152
rect 7317 7882 7373 12150
rect 7483 8000 7539 12328
rect 7619 10087 7675 14533
rect 8291 14345 8347 14659
rect 8475 14603 8531 14801
rect 8463 14601 8543 14603
rect 8463 14545 8475 14601
rect 8531 14545 8543 14601
rect 8463 14543 8543 14545
rect 8475 14345 8531 14543
rect 8659 14487 8715 14801
rect 8792 14603 8860 14933
rect 8792 14601 8872 14603
rect 8792 14545 8804 14601
rect 8860 14545 8872 14601
rect 8792 14543 8872 14545
rect 9059 14601 9129 14613
rect 9059 14545 9061 14601
rect 9117 14545 9129 14601
rect 8647 14485 8727 14487
rect 8647 14429 8659 14485
rect 8715 14429 8727 14485
rect 8647 14427 8727 14429
rect 8659 14345 8715 14427
rect 8279 14335 8359 14345
rect 8279 14279 8291 14335
rect 8347 14279 8359 14335
rect 8279 14269 8359 14279
rect 8463 14335 8543 14345
rect 8463 14279 8475 14335
rect 8531 14279 8543 14335
rect 8463 14269 8543 14279
rect 8647 14335 8727 14345
rect 8647 14279 8659 14335
rect 8715 14279 8727 14335
rect 8647 14269 8727 14279
rect 8792 14213 8860 14543
rect 9059 14535 9129 14545
rect 8751 14205 8860 14213
rect 8739 14203 8860 14205
rect 8739 14083 8751 14203
rect 8807 14083 8860 14203
rect 8739 14081 8860 14083
rect 8751 14073 8807 14081
rect 8054 13816 8952 13828
rect 8054 13760 8066 13816
rect 8122 13760 8884 13816
rect 8940 13760 8952 13816
rect 8054 13748 8952 13760
rect 9061 13591 9117 14535
rect 9225 13698 9305 13708
rect 9225 13642 9237 13698
rect 9293 13642 9305 13698
rect 9225 13640 9305 13642
rect 9059 13588 9129 13591
rect 9059 13534 9061 13588
rect 9117 13534 9129 13588
rect 9059 13522 9129 13534
rect 8199 13481 8945 13493
rect 8199 13425 8567 13481
rect 8623 13425 8945 13481
rect 8199 13413 8945 13425
rect 8199 13160 8255 13413
rect 8567 13160 8623 13413
rect 8889 13160 8945 13413
rect 8187 13158 8267 13160
rect 8187 13038 8199 13158
rect 8255 13038 8267 13158
rect 8187 13036 8267 13038
rect 8555 13158 8635 13160
rect 8555 13038 8567 13158
rect 8623 13038 8635 13158
rect 8555 13036 8635 13038
rect 8877 13158 8957 13160
rect 8877 13037 8889 13158
rect 8945 13037 8957 13158
rect 8199 13028 8255 13036
rect 8567 13028 8623 13036
rect 8877 13035 8957 13037
rect 8889 13027 8945 13035
rect 8383 12860 8439 12868
rect 8751 12860 8807 12868
rect 8371 12858 8860 12860
rect 8371 12738 8383 12858
rect 8439 12738 8751 12858
rect 8807 12738 8860 12858
rect 8371 12736 8860 12738
rect 8383 12728 8439 12736
rect 8751 12728 8860 12736
rect 8279 12662 8359 12672
rect 8279 12606 8291 12662
rect 8347 12606 8359 12662
rect 8279 12596 8359 12606
rect 8463 12662 8543 12672
rect 8463 12606 8475 12662
rect 8531 12606 8543 12662
rect 8463 12596 8543 12606
rect 8647 12662 8727 12672
rect 8647 12606 8659 12662
rect 8715 12606 8727 12662
rect 8647 12596 8727 12606
rect 8291 12514 8347 12596
rect 8279 12512 8359 12514
rect 8279 12456 8291 12512
rect 8347 12456 8359 12512
rect 8279 12454 8359 12456
rect 8291 12140 8347 12454
rect 8475 12398 8531 12596
rect 8463 12396 8543 12398
rect 8463 12340 8475 12396
rect 8531 12340 8543 12396
rect 8463 12338 8543 12340
rect 8475 12140 8531 12338
rect 8659 12282 8715 12596
rect 8792 12398 8860 12728
rect 9237 12406 9293 13640
rect 9685 13481 10431 13493
rect 9685 13425 10053 13481
rect 10109 13425 10431 13481
rect 9685 13413 10431 13425
rect 9685 13160 9741 13413
rect 10053 13160 10109 13413
rect 10375 13160 10431 13413
rect 9673 13158 9753 13160
rect 9673 13038 9685 13158
rect 9741 13038 9753 13158
rect 9673 13036 9753 13038
rect 10041 13158 10121 13160
rect 10041 13038 10053 13158
rect 10109 13038 10121 13158
rect 10041 13036 10121 13038
rect 10363 13158 10443 13160
rect 10363 13037 10375 13158
rect 10431 13037 10443 13158
rect 9685 13028 9741 13036
rect 10053 13028 10109 13036
rect 10363 13035 10443 13037
rect 10375 13027 10431 13035
rect 9869 12860 9925 12868
rect 10237 12860 10293 12868
rect 9857 12858 10346 12860
rect 9857 12738 9869 12858
rect 9925 12738 10237 12858
rect 10293 12738 10346 12858
rect 9857 12736 10346 12738
rect 9869 12728 9925 12736
rect 10237 12728 10346 12736
rect 9765 12662 9845 12672
rect 9765 12606 9777 12662
rect 9833 12606 9845 12662
rect 9765 12596 9845 12606
rect 9949 12662 10029 12672
rect 9949 12606 9961 12662
rect 10017 12606 10029 12662
rect 9949 12596 10029 12606
rect 10133 12662 10213 12672
rect 10133 12606 10145 12662
rect 10201 12606 10213 12662
rect 10133 12596 10213 12606
rect 9777 12514 9833 12596
rect 9765 12512 9845 12514
rect 9765 12456 9777 12512
rect 9833 12456 9845 12512
rect 9765 12454 9845 12456
rect 8792 12396 8872 12398
rect 8792 12340 8804 12396
rect 8860 12340 8872 12396
rect 8792 12338 8872 12340
rect 9235 12396 9295 12406
rect 9235 12340 9237 12396
rect 9293 12340 9295 12396
rect 8647 12280 8727 12282
rect 8647 12224 8659 12280
rect 8715 12224 8727 12280
rect 8647 12222 8727 12224
rect 8659 12140 8715 12222
rect 8279 12130 8359 12140
rect 8279 12074 8291 12130
rect 8347 12074 8359 12130
rect 8279 12064 8359 12074
rect 8463 12130 8543 12140
rect 8463 12074 8475 12130
rect 8531 12074 8543 12130
rect 8463 12064 8543 12074
rect 8647 12130 8727 12140
rect 8647 12074 8659 12130
rect 8715 12074 8727 12130
rect 8647 12064 8727 12074
rect 8792 12008 8860 12338
rect 9235 12328 9295 12340
rect 8751 12000 8860 12008
rect 8739 11998 8860 12000
rect 8739 11878 8751 11998
rect 8807 11878 8860 11998
rect 8739 11876 8860 11878
rect 8751 11868 8807 11876
rect 8054 11611 8950 11623
rect 8054 11555 8066 11611
rect 8122 11555 8884 11611
rect 8940 11555 8950 11611
rect 8054 11543 8950 11555
rect 9237 11385 9293 12328
rect 9777 12140 9833 12454
rect 9961 12398 10017 12596
rect 9949 12396 10029 12398
rect 9949 12340 9961 12396
rect 10017 12340 10029 12396
rect 9949 12338 10029 12340
rect 9961 12140 10017 12338
rect 10145 12282 10201 12596
rect 10278 12398 10346 12728
rect 10278 12396 10358 12398
rect 10278 12340 10290 12396
rect 10346 12340 10358 12396
rect 10278 12338 10358 12340
rect 10545 12396 10615 12408
rect 10545 12340 10547 12396
rect 10603 12340 10871 12396
rect 10133 12280 10213 12282
rect 10133 12224 10145 12280
rect 10201 12224 10213 12280
rect 10133 12222 10213 12224
rect 10145 12140 10201 12222
rect 9765 12130 9845 12140
rect 9765 12074 9777 12130
rect 9833 12074 9845 12130
rect 9765 12064 9845 12074
rect 9949 12130 10029 12140
rect 9949 12074 9961 12130
rect 10017 12074 10029 12130
rect 9949 12064 10029 12074
rect 10133 12130 10213 12140
rect 10133 12074 10145 12130
rect 10201 12074 10213 12130
rect 10133 12064 10213 12074
rect 10278 12008 10346 12338
rect 10545 12330 10615 12340
rect 10237 12000 10346 12008
rect 10225 11998 10346 12000
rect 10225 11878 10237 11998
rect 10293 11878 10346 11998
rect 10225 11876 10346 11878
rect 10237 11868 10293 11876
rect 9540 11611 10436 11623
rect 9540 11555 9552 11611
rect 9608 11555 10370 11611
rect 10426 11555 10436 11611
rect 9540 11543 10436 11555
rect 10547 11386 10603 12330
rect 10711 11494 10791 11504
rect 10711 11438 10723 11494
rect 10779 11438 10791 11494
rect 10711 11436 10791 11438
rect 9235 11383 9305 11385
rect 9235 11327 9237 11383
rect 9293 11327 9305 11383
rect 9235 11315 9305 11327
rect 10535 11384 10615 11386
rect 10535 11328 10547 11384
rect 10603 11328 10615 11384
rect 10535 11316 10615 11328
rect 8199 11276 8945 11288
rect 8199 11220 8567 11276
rect 8623 11220 8945 11276
rect 8199 11208 8945 11220
rect 8199 10955 8255 11208
rect 8567 10955 8623 11208
rect 8889 10955 8945 11208
rect 9685 11277 10431 11289
rect 9685 11221 10053 11277
rect 10109 11221 10431 11277
rect 9685 11209 10431 11221
rect 9685 10956 9741 11209
rect 10053 10956 10109 11209
rect 10375 10956 10431 11209
rect 8187 10953 8267 10955
rect 8187 10833 8199 10953
rect 8255 10833 8267 10953
rect 8187 10831 8267 10833
rect 8555 10953 8635 10955
rect 8555 10833 8567 10953
rect 8623 10833 8635 10953
rect 8555 10831 8635 10833
rect 8877 10953 8957 10955
rect 8877 10832 8889 10953
rect 8945 10832 8957 10953
rect 9673 10954 9753 10956
rect 9673 10834 9685 10954
rect 9741 10834 9753 10954
rect 9673 10832 9753 10834
rect 10041 10954 10121 10956
rect 10041 10834 10053 10954
rect 10109 10834 10121 10954
rect 10041 10832 10121 10834
rect 10363 10954 10443 10956
rect 10363 10833 10375 10954
rect 10431 10833 10443 10954
rect 8199 10823 8255 10831
rect 8567 10823 8623 10831
rect 8877 10830 8957 10832
rect 8889 10822 8945 10830
rect 9685 10824 9741 10832
rect 10053 10824 10109 10832
rect 10363 10831 10443 10833
rect 10375 10823 10431 10831
rect 8383 10655 8439 10663
rect 8751 10655 8807 10663
rect 9869 10656 9925 10664
rect 10237 10656 10293 10664
rect 8371 10653 8860 10655
rect 8371 10533 8383 10653
rect 8439 10533 8751 10653
rect 8807 10533 8860 10653
rect 8371 10531 8860 10533
rect 9857 10654 10346 10656
rect 9857 10534 9869 10654
rect 9925 10534 10237 10654
rect 10293 10534 10346 10654
rect 9857 10532 10346 10534
rect 8383 10523 8439 10531
rect 8751 10523 8860 10531
rect 9869 10524 9925 10532
rect 10237 10524 10346 10532
rect 8279 10457 8359 10467
rect 8279 10401 8291 10457
rect 8347 10401 8359 10457
rect 8279 10391 8359 10401
rect 8463 10457 8543 10467
rect 8463 10401 8475 10457
rect 8531 10401 8543 10457
rect 8463 10391 8543 10401
rect 8647 10457 8727 10467
rect 8647 10401 8659 10457
rect 8715 10401 8727 10457
rect 8647 10391 8727 10401
rect 8291 10309 8347 10391
rect 8279 10307 8359 10309
rect 8279 10251 8291 10307
rect 8347 10251 8359 10307
rect 8279 10249 8359 10251
rect 7607 10075 7677 10087
rect 7607 10019 7619 10075
rect 7675 10019 7677 10075
rect 7607 10007 7677 10019
rect 8291 9935 8347 10249
rect 8475 10193 8531 10391
rect 8463 10191 8543 10193
rect 8463 10135 8475 10191
rect 8531 10135 8543 10191
rect 8463 10133 8543 10135
rect 8475 9935 8531 10133
rect 8659 10077 8715 10391
rect 8792 10193 8860 10523
rect 9765 10458 9845 10468
rect 9765 10402 9777 10458
rect 9833 10402 9845 10458
rect 9765 10392 9845 10402
rect 9949 10458 10029 10468
rect 9949 10402 9961 10458
rect 10017 10402 10029 10458
rect 9949 10392 10029 10402
rect 10133 10458 10213 10468
rect 10133 10402 10145 10458
rect 10201 10402 10213 10458
rect 10133 10392 10213 10402
rect 9777 10310 9833 10392
rect 9765 10308 9845 10310
rect 9765 10252 9777 10308
rect 9833 10252 9845 10308
rect 9765 10250 9845 10252
rect 8792 10191 8872 10193
rect 8792 10135 8804 10191
rect 8860 10135 8872 10191
rect 8792 10133 8872 10135
rect 9059 10191 9129 10203
rect 9059 10135 9061 10191
rect 9117 10135 9129 10191
rect 8647 10075 8727 10077
rect 8647 10019 8659 10075
rect 8715 10019 8727 10075
rect 8647 10017 8727 10019
rect 8659 9935 8715 10017
rect 8279 9925 8359 9935
rect 8279 9869 8291 9925
rect 8347 9869 8359 9925
rect 8279 9859 8359 9869
rect 8463 9925 8543 9935
rect 8463 9869 8475 9925
rect 8531 9869 8543 9925
rect 8463 9859 8543 9869
rect 8647 9925 8727 9935
rect 8647 9869 8659 9925
rect 8715 9869 8727 9925
rect 8647 9859 8727 9869
rect 8792 9803 8860 10133
rect 9059 10125 9129 10135
rect 8751 9795 8860 9803
rect 8739 9793 8860 9795
rect 8739 9673 8751 9793
rect 8807 9673 8860 9793
rect 8739 9671 8860 9673
rect 8751 9663 8807 9671
rect 8054 9406 8950 9418
rect 8054 9350 8066 9406
rect 8122 9350 8884 9406
rect 8940 9350 8950 9406
rect 8054 9338 8950 9350
rect 9061 9181 9117 10125
rect 9777 9936 9833 10250
rect 9961 10194 10017 10392
rect 9949 10192 10029 10194
rect 9949 10136 9961 10192
rect 10017 10136 10029 10192
rect 9949 10134 10029 10136
rect 9961 9936 10017 10134
rect 10145 10078 10201 10392
rect 10278 10194 10346 10524
rect 10723 10202 10779 11436
rect 10278 10192 10358 10194
rect 10278 10136 10290 10192
rect 10346 10136 10358 10192
rect 10278 10134 10358 10136
rect 10721 10192 10791 10202
rect 10951 10192 11007 24235
rect 11153 21984 11209 25840
rect 15195 25724 15251 26389
rect 15193 25722 15263 25724
rect 15193 25666 15195 25722
rect 15251 25666 15263 25722
rect 15193 25664 15263 25666
rect 11377 25546 11447 25558
rect 11377 25490 11389 25546
rect 11445 25490 11447 25546
rect 11377 25488 11447 25490
rect 11151 21972 11221 21984
rect 11151 21916 11153 21972
rect 11209 21916 11221 21972
rect 11151 21904 11221 21916
rect 11389 21072 11445 25488
rect 12241 25262 12987 25274
rect 12241 25206 12609 25262
rect 12665 25206 12987 25262
rect 12241 25194 12987 25206
rect 12241 24941 12297 25194
rect 12609 24941 12665 25194
rect 12931 24941 12987 25194
rect 12229 24939 12309 24941
rect 12229 24819 12241 24939
rect 12297 24819 12309 24939
rect 12229 24817 12309 24819
rect 12597 24939 12677 24941
rect 12597 24819 12609 24939
rect 12665 24819 12677 24939
rect 12597 24817 12677 24819
rect 12919 24939 12999 24941
rect 12919 24818 12931 24939
rect 12987 24818 12999 24939
rect 12241 24809 12297 24817
rect 12609 24809 12665 24817
rect 12919 24816 12999 24818
rect 12931 24808 12987 24816
rect 12425 24641 12481 24649
rect 12793 24641 12849 24649
rect 12413 24639 12902 24641
rect 12413 24519 12425 24639
rect 12481 24519 12793 24639
rect 12849 24519 12902 24639
rect 12413 24517 12902 24519
rect 12425 24509 12481 24517
rect 12793 24509 12902 24517
rect 12321 24443 12401 24453
rect 12321 24387 12333 24443
rect 12389 24387 12401 24443
rect 12321 24377 12401 24387
rect 12505 24443 12585 24453
rect 12505 24387 12517 24443
rect 12573 24387 12585 24443
rect 12505 24377 12585 24387
rect 12689 24443 12769 24453
rect 12689 24387 12701 24443
rect 12757 24387 12769 24443
rect 12689 24377 12769 24387
rect 12333 24295 12389 24377
rect 12321 24293 12401 24295
rect 12321 24237 12333 24293
rect 12389 24237 12401 24293
rect 12321 24235 12401 24237
rect 11649 24177 11719 24189
rect 11649 24121 11661 24177
rect 11717 24121 11719 24177
rect 11649 24109 11719 24121
rect 11513 21972 11583 21986
rect 11513 21916 11525 21972
rect 11581 21916 11583 21972
rect 11513 21904 11583 21916
rect 11377 21070 11447 21072
rect 11377 21014 11389 21070
rect 11445 21014 11447 21070
rect 11377 21002 11447 21014
rect 11525 17576 11581 21904
rect 11661 19663 11717 24109
rect 12333 23921 12389 24235
rect 12517 24179 12573 24377
rect 12505 24177 12585 24179
rect 12505 24121 12517 24177
rect 12573 24121 12585 24177
rect 12505 24119 12585 24121
rect 12517 23921 12573 24119
rect 12701 24063 12757 24377
rect 12834 24179 12902 24509
rect 14981 24293 15061 24305
rect 14981 24237 14993 24293
rect 15049 24237 15061 24293
rect 14981 24235 15061 24237
rect 12834 24177 12914 24179
rect 12834 24121 12846 24177
rect 12902 24121 12914 24177
rect 12834 24119 12914 24121
rect 13101 24177 13171 24189
rect 13101 24121 13103 24177
rect 13159 24121 13171 24177
rect 12689 24061 12769 24063
rect 12689 24005 12701 24061
rect 12757 24005 12769 24061
rect 12689 24003 12769 24005
rect 12701 23921 12757 24003
rect 12321 23911 12401 23921
rect 12321 23855 12333 23911
rect 12389 23855 12401 23911
rect 12321 23845 12401 23855
rect 12505 23911 12585 23921
rect 12505 23855 12517 23911
rect 12573 23855 12585 23911
rect 12505 23845 12585 23855
rect 12689 23911 12769 23921
rect 12689 23855 12701 23911
rect 12757 23855 12769 23911
rect 12689 23845 12769 23855
rect 12834 23789 12902 24119
rect 13101 24111 13171 24121
rect 12793 23781 12902 23789
rect 12781 23779 12902 23781
rect 12781 23659 12793 23779
rect 12849 23659 12902 23779
rect 12781 23657 12902 23659
rect 12793 23649 12849 23657
rect 12096 23392 12994 23404
rect 12096 23336 12108 23392
rect 12164 23336 12926 23392
rect 12982 23336 12994 23392
rect 12096 23324 12994 23336
rect 13103 23167 13159 24111
rect 13267 23274 13347 23284
rect 13267 23218 13279 23274
rect 13335 23218 13347 23274
rect 13267 23216 13347 23218
rect 13101 23164 13171 23167
rect 13101 23110 13103 23164
rect 13159 23110 13171 23164
rect 13101 23098 13171 23110
rect 12241 23057 12987 23069
rect 12241 23001 12609 23057
rect 12665 23001 12987 23057
rect 12241 22989 12987 23001
rect 12241 22736 12297 22989
rect 12609 22736 12665 22989
rect 12931 22736 12987 22989
rect 12229 22734 12309 22736
rect 12229 22614 12241 22734
rect 12297 22614 12309 22734
rect 12229 22612 12309 22614
rect 12597 22734 12677 22736
rect 12597 22614 12609 22734
rect 12665 22614 12677 22734
rect 12597 22612 12677 22614
rect 12919 22734 12999 22736
rect 12919 22613 12931 22734
rect 12987 22613 12999 22734
rect 12241 22604 12297 22612
rect 12609 22604 12665 22612
rect 12919 22611 12999 22613
rect 12931 22603 12987 22611
rect 12425 22436 12481 22444
rect 12793 22436 12849 22444
rect 12413 22434 12902 22436
rect 12413 22314 12425 22434
rect 12481 22314 12793 22434
rect 12849 22314 12902 22434
rect 12413 22312 12902 22314
rect 12425 22304 12481 22312
rect 12793 22304 12902 22312
rect 12321 22238 12401 22248
rect 12321 22182 12333 22238
rect 12389 22182 12401 22238
rect 12321 22172 12401 22182
rect 12505 22238 12585 22248
rect 12505 22182 12517 22238
rect 12573 22182 12585 22238
rect 12505 22172 12585 22182
rect 12689 22238 12769 22248
rect 12689 22182 12701 22238
rect 12757 22182 12769 22238
rect 12689 22172 12769 22182
rect 12333 22090 12389 22172
rect 12321 22088 12401 22090
rect 12321 22032 12333 22088
rect 12389 22032 12401 22088
rect 12321 22030 12401 22032
rect 12333 21716 12389 22030
rect 12517 21974 12573 22172
rect 12505 21972 12585 21974
rect 12505 21916 12517 21972
rect 12573 21916 12585 21972
rect 12505 21914 12585 21916
rect 12517 21716 12573 21914
rect 12701 21858 12757 22172
rect 12834 21974 12902 22304
rect 13279 21982 13335 23216
rect 13727 23057 14473 23069
rect 13727 23001 14095 23057
rect 14151 23001 14473 23057
rect 13727 22989 14473 23001
rect 13727 22736 13783 22989
rect 14095 22736 14151 22989
rect 14417 22736 14473 22989
rect 13715 22734 13795 22736
rect 13715 22614 13727 22734
rect 13783 22614 13795 22734
rect 13715 22612 13795 22614
rect 14083 22734 14163 22736
rect 14083 22614 14095 22734
rect 14151 22614 14163 22734
rect 14083 22612 14163 22614
rect 14405 22734 14485 22736
rect 14405 22613 14417 22734
rect 14473 22613 14485 22734
rect 13727 22604 13783 22612
rect 14095 22604 14151 22612
rect 14405 22611 14485 22613
rect 14417 22603 14473 22611
rect 13911 22436 13967 22444
rect 14279 22436 14335 22444
rect 13899 22434 14388 22436
rect 13899 22314 13911 22434
rect 13967 22314 14279 22434
rect 14335 22314 14388 22434
rect 13899 22312 14388 22314
rect 13911 22304 13967 22312
rect 14279 22304 14388 22312
rect 13807 22238 13887 22248
rect 13807 22182 13819 22238
rect 13875 22182 13887 22238
rect 13807 22172 13887 22182
rect 13991 22238 14071 22248
rect 13991 22182 14003 22238
rect 14059 22182 14071 22238
rect 13991 22172 14071 22182
rect 14175 22238 14255 22248
rect 14175 22182 14187 22238
rect 14243 22182 14255 22238
rect 14175 22172 14255 22182
rect 13819 22090 13875 22172
rect 13807 22088 13887 22090
rect 13807 22032 13819 22088
rect 13875 22032 13887 22088
rect 13807 22030 13887 22032
rect 12834 21972 12914 21974
rect 12834 21916 12846 21972
rect 12902 21916 12914 21972
rect 12834 21914 12914 21916
rect 13277 21972 13337 21982
rect 13277 21916 13279 21972
rect 13335 21916 13337 21972
rect 12689 21856 12769 21858
rect 12689 21800 12701 21856
rect 12757 21800 12769 21856
rect 12689 21798 12769 21800
rect 12701 21716 12757 21798
rect 12321 21706 12401 21716
rect 12321 21650 12333 21706
rect 12389 21650 12401 21706
rect 12321 21640 12401 21650
rect 12505 21706 12585 21716
rect 12505 21650 12517 21706
rect 12573 21650 12585 21706
rect 12505 21640 12585 21650
rect 12689 21706 12769 21716
rect 12689 21650 12701 21706
rect 12757 21650 12769 21706
rect 12689 21640 12769 21650
rect 12834 21584 12902 21914
rect 13277 21904 13337 21916
rect 12793 21576 12902 21584
rect 12781 21574 12902 21576
rect 12781 21454 12793 21574
rect 12849 21454 12902 21574
rect 12781 21452 12902 21454
rect 12793 21444 12849 21452
rect 12096 21187 12992 21199
rect 12096 21131 12108 21187
rect 12164 21131 12926 21187
rect 12982 21131 12992 21187
rect 12096 21119 12992 21131
rect 13279 20961 13335 21904
rect 13819 21716 13875 22030
rect 14003 21974 14059 22172
rect 13991 21972 14071 21974
rect 13991 21916 14003 21972
rect 14059 21916 14071 21972
rect 13991 21914 14071 21916
rect 14003 21716 14059 21914
rect 14187 21858 14243 22172
rect 14320 21974 14388 22304
rect 14320 21972 14400 21974
rect 14320 21916 14332 21972
rect 14388 21916 14400 21972
rect 14320 21914 14400 21916
rect 14587 21972 14657 21984
rect 14587 21916 14589 21972
rect 14645 21916 14913 21972
rect 14175 21856 14255 21858
rect 14175 21800 14187 21856
rect 14243 21800 14255 21856
rect 14175 21798 14255 21800
rect 14187 21716 14243 21798
rect 13807 21706 13887 21716
rect 13807 21650 13819 21706
rect 13875 21650 13887 21706
rect 13807 21640 13887 21650
rect 13991 21706 14071 21716
rect 13991 21650 14003 21706
rect 14059 21650 14071 21706
rect 13991 21640 14071 21650
rect 14175 21706 14255 21716
rect 14175 21650 14187 21706
rect 14243 21650 14255 21706
rect 14175 21640 14255 21650
rect 14320 21584 14388 21914
rect 14587 21906 14657 21916
rect 14279 21576 14388 21584
rect 14267 21574 14388 21576
rect 14267 21454 14279 21574
rect 14335 21454 14388 21574
rect 14267 21452 14388 21454
rect 14279 21444 14335 21452
rect 13582 21187 14478 21199
rect 13582 21131 13594 21187
rect 13650 21131 14412 21187
rect 14468 21131 14478 21187
rect 13582 21119 14478 21131
rect 14589 20962 14645 21906
rect 14753 21070 14833 21080
rect 14753 21014 14765 21070
rect 14821 21014 14833 21070
rect 14753 21012 14833 21014
rect 13277 20959 13347 20961
rect 13277 20903 13279 20959
rect 13335 20903 13347 20959
rect 13277 20891 13347 20903
rect 14577 20960 14657 20962
rect 14577 20904 14589 20960
rect 14645 20904 14657 20960
rect 14577 20892 14657 20904
rect 12241 20852 12987 20864
rect 12241 20796 12609 20852
rect 12665 20796 12987 20852
rect 12241 20784 12987 20796
rect 12241 20531 12297 20784
rect 12609 20531 12665 20784
rect 12931 20531 12987 20784
rect 13727 20853 14473 20865
rect 13727 20797 14095 20853
rect 14151 20797 14473 20853
rect 13727 20785 14473 20797
rect 13727 20532 13783 20785
rect 14095 20532 14151 20785
rect 14417 20532 14473 20785
rect 12229 20529 12309 20531
rect 12229 20409 12241 20529
rect 12297 20409 12309 20529
rect 12229 20407 12309 20409
rect 12597 20529 12677 20531
rect 12597 20409 12609 20529
rect 12665 20409 12677 20529
rect 12597 20407 12677 20409
rect 12919 20529 12999 20531
rect 12919 20408 12931 20529
rect 12987 20408 12999 20529
rect 13715 20530 13795 20532
rect 13715 20410 13727 20530
rect 13783 20410 13795 20530
rect 13715 20408 13795 20410
rect 14083 20530 14163 20532
rect 14083 20410 14095 20530
rect 14151 20410 14163 20530
rect 14083 20408 14163 20410
rect 14405 20530 14485 20532
rect 14405 20409 14417 20530
rect 14473 20409 14485 20530
rect 12241 20399 12297 20407
rect 12609 20399 12665 20407
rect 12919 20406 12999 20408
rect 12931 20398 12987 20406
rect 13727 20400 13783 20408
rect 14095 20400 14151 20408
rect 14405 20407 14485 20409
rect 14417 20399 14473 20407
rect 12425 20231 12481 20239
rect 12793 20231 12849 20239
rect 13911 20232 13967 20240
rect 14279 20232 14335 20240
rect 12413 20229 12902 20231
rect 12413 20109 12425 20229
rect 12481 20109 12793 20229
rect 12849 20109 12902 20229
rect 12413 20107 12902 20109
rect 13899 20230 14388 20232
rect 13899 20110 13911 20230
rect 13967 20110 14279 20230
rect 14335 20110 14388 20230
rect 13899 20108 14388 20110
rect 12425 20099 12481 20107
rect 12793 20099 12902 20107
rect 13911 20100 13967 20108
rect 14279 20100 14388 20108
rect 12321 20033 12401 20043
rect 12321 19977 12333 20033
rect 12389 19977 12401 20033
rect 12321 19967 12401 19977
rect 12505 20033 12585 20043
rect 12505 19977 12517 20033
rect 12573 19977 12585 20033
rect 12505 19967 12585 19977
rect 12689 20033 12769 20043
rect 12689 19977 12701 20033
rect 12757 19977 12769 20033
rect 12689 19967 12769 19977
rect 12333 19885 12389 19967
rect 12321 19883 12401 19885
rect 12321 19827 12333 19883
rect 12389 19827 12401 19883
rect 12321 19825 12401 19827
rect 11649 19651 11719 19663
rect 11649 19595 11661 19651
rect 11717 19595 11719 19651
rect 11649 19583 11719 19595
rect 12333 19511 12389 19825
rect 12517 19769 12573 19967
rect 12505 19767 12585 19769
rect 12505 19711 12517 19767
rect 12573 19711 12585 19767
rect 12505 19709 12585 19711
rect 12517 19511 12573 19709
rect 12701 19653 12757 19967
rect 12834 19769 12902 20099
rect 13807 20034 13887 20044
rect 13807 19978 13819 20034
rect 13875 19978 13887 20034
rect 13807 19968 13887 19978
rect 13991 20034 14071 20044
rect 13991 19978 14003 20034
rect 14059 19978 14071 20034
rect 13991 19968 14071 19978
rect 14175 20034 14255 20044
rect 14175 19978 14187 20034
rect 14243 19978 14255 20034
rect 14175 19968 14255 19978
rect 13819 19886 13875 19968
rect 13807 19884 13887 19886
rect 13807 19828 13819 19884
rect 13875 19828 13887 19884
rect 13807 19826 13887 19828
rect 12834 19767 12914 19769
rect 12834 19711 12846 19767
rect 12902 19711 12914 19767
rect 12834 19709 12914 19711
rect 13101 19767 13171 19779
rect 13101 19711 13103 19767
rect 13159 19711 13171 19767
rect 12689 19651 12769 19653
rect 12689 19595 12701 19651
rect 12757 19595 12769 19651
rect 12689 19593 12769 19595
rect 12701 19511 12757 19593
rect 12321 19501 12401 19511
rect 12321 19445 12333 19501
rect 12389 19445 12401 19501
rect 12321 19435 12401 19445
rect 12505 19501 12585 19511
rect 12505 19445 12517 19501
rect 12573 19445 12585 19501
rect 12505 19435 12585 19445
rect 12689 19501 12769 19511
rect 12689 19445 12701 19501
rect 12757 19445 12769 19501
rect 12689 19435 12769 19445
rect 12834 19379 12902 19709
rect 13101 19701 13171 19711
rect 12793 19371 12902 19379
rect 12781 19369 12902 19371
rect 12781 19249 12793 19369
rect 12849 19249 12902 19369
rect 12781 19247 12902 19249
rect 12793 19239 12849 19247
rect 12096 18982 12992 18994
rect 12096 18926 12108 18982
rect 12164 18926 12926 18982
rect 12982 18926 12992 18982
rect 12096 18914 12992 18926
rect 13103 18757 13159 19701
rect 13819 19512 13875 19826
rect 14003 19770 14059 19968
rect 13991 19768 14071 19770
rect 13991 19712 14003 19768
rect 14059 19712 14071 19768
rect 13991 19710 14071 19712
rect 14003 19512 14059 19710
rect 14187 19654 14243 19968
rect 14320 19770 14388 20100
rect 14765 19778 14821 21012
rect 14320 19768 14400 19770
rect 14320 19712 14332 19768
rect 14388 19712 14400 19768
rect 14320 19710 14400 19712
rect 14763 19768 14833 19778
rect 14763 19712 14765 19768
rect 14821 19712 14913 19768
rect 14175 19652 14255 19654
rect 14175 19596 14187 19652
rect 14243 19596 14255 19652
rect 14175 19594 14255 19596
rect 14187 19512 14243 19594
rect 13807 19502 13887 19512
rect 13807 19446 13819 19502
rect 13875 19446 13887 19502
rect 13807 19436 13887 19446
rect 13991 19502 14071 19512
rect 13991 19446 14003 19502
rect 14059 19446 14071 19502
rect 13991 19436 14071 19446
rect 14175 19502 14255 19512
rect 14175 19446 14187 19502
rect 14243 19446 14255 19502
rect 14175 19436 14255 19446
rect 14320 19380 14388 19710
rect 14763 19700 14833 19712
rect 14279 19372 14388 19380
rect 14267 19370 14388 19372
rect 14267 19250 14279 19370
rect 14335 19250 14388 19370
rect 14267 19248 14388 19250
rect 14279 19240 14335 19248
rect 13582 18983 14478 18995
rect 13582 18927 13594 18983
rect 13650 18927 14412 18983
rect 14468 18927 14478 18983
rect 13582 18915 14478 18927
rect 13267 18864 13347 18874
rect 13267 18808 13279 18864
rect 13335 18808 13347 18864
rect 13267 18806 13347 18808
rect 13101 18754 13171 18757
rect 13101 18700 13103 18754
rect 13159 18700 13171 18754
rect 13101 18688 13171 18700
rect 12241 18647 12987 18659
rect 12241 18591 12609 18647
rect 12665 18591 12987 18647
rect 12241 18579 12987 18591
rect 12241 18326 12297 18579
rect 12609 18326 12665 18579
rect 12931 18326 12987 18579
rect 12229 18324 12309 18326
rect 12229 18204 12241 18324
rect 12297 18204 12309 18324
rect 12229 18202 12309 18204
rect 12597 18324 12677 18326
rect 12597 18204 12609 18324
rect 12665 18204 12677 18324
rect 12597 18202 12677 18204
rect 12919 18324 12999 18326
rect 12919 18203 12931 18324
rect 12987 18203 12999 18324
rect 12241 18194 12297 18202
rect 12609 18194 12665 18202
rect 12919 18201 12999 18203
rect 12931 18193 12987 18201
rect 12425 18026 12481 18034
rect 12793 18026 12849 18034
rect 12413 18024 12902 18026
rect 12413 17904 12425 18024
rect 12481 17904 12793 18024
rect 12849 17904 12902 18024
rect 12413 17902 12902 17904
rect 12425 17894 12481 17902
rect 12793 17894 12902 17902
rect 12321 17828 12401 17838
rect 12321 17772 12333 17828
rect 12389 17772 12401 17828
rect 12321 17762 12401 17772
rect 12505 17828 12585 17838
rect 12505 17772 12517 17828
rect 12573 17772 12585 17828
rect 12505 17762 12585 17772
rect 12689 17828 12769 17838
rect 12689 17772 12701 17828
rect 12757 17772 12769 17828
rect 12689 17762 12769 17772
rect 12333 17680 12389 17762
rect 12321 17678 12401 17680
rect 12321 17622 12333 17678
rect 12389 17622 12401 17678
rect 12321 17620 12401 17622
rect 11513 17562 11583 17576
rect 11513 17506 11525 17562
rect 11581 17506 11583 17562
rect 11513 17494 11583 17506
rect 11211 16659 11281 16671
rect 11525 16663 11581 17494
rect 12333 17306 12389 17620
rect 12517 17564 12573 17762
rect 12505 17562 12585 17564
rect 12505 17506 12517 17562
rect 12573 17506 12585 17562
rect 12505 17504 12585 17506
rect 12517 17306 12573 17504
rect 12701 17448 12757 17762
rect 12834 17564 12902 17894
rect 13279 17574 13335 18806
rect 12834 17562 12914 17564
rect 12834 17506 12846 17562
rect 12902 17506 12914 17562
rect 12834 17504 12914 17506
rect 13277 17562 13337 17574
rect 13277 17506 13279 17562
rect 13335 17506 13337 17562
rect 12689 17446 12769 17448
rect 12689 17390 12701 17446
rect 12757 17390 12769 17446
rect 12689 17388 12769 17390
rect 12701 17306 12757 17388
rect 12321 17296 12401 17306
rect 12321 17240 12333 17296
rect 12389 17240 12401 17296
rect 12321 17230 12401 17240
rect 12505 17296 12585 17306
rect 12505 17240 12517 17296
rect 12573 17240 12585 17296
rect 12505 17230 12585 17240
rect 12689 17296 12769 17306
rect 12689 17240 12701 17296
rect 12757 17240 12769 17296
rect 12689 17230 12769 17240
rect 12834 17174 12902 17504
rect 13277 17494 13337 17506
rect 12793 17166 12902 17174
rect 12781 17164 12902 17166
rect 12781 17044 12793 17164
rect 12849 17044 12902 17164
rect 12781 17042 12902 17044
rect 12793 17034 12849 17042
rect 12096 16777 12994 16789
rect 12096 16721 12108 16777
rect 12164 16721 12926 16777
rect 12982 16721 12994 16777
rect 12096 16709 12994 16721
rect 11211 16603 11223 16659
rect 11279 16603 11281 16659
rect 11211 16601 11281 16603
rect 11523 16659 11583 16663
rect 11523 16603 11525 16659
rect 11581 16603 11583 16659
rect 11223 15989 11279 16601
rect 11523 16591 11583 16603
rect 11075 11494 11145 11506
rect 11075 11438 11087 11494
rect 11143 11438 11145 11494
rect 11075 11426 11145 11438
rect 10721 10136 10723 10192
rect 10779 10136 11007 10192
rect 10133 10076 10213 10078
rect 10133 10020 10145 10076
rect 10201 10020 10213 10076
rect 10133 10018 10213 10020
rect 10145 9936 10201 10018
rect 9765 9926 9845 9936
rect 9765 9870 9777 9926
rect 9833 9870 9845 9926
rect 9765 9860 9845 9870
rect 9949 9926 10029 9936
rect 9949 9870 9961 9926
rect 10017 9870 10029 9926
rect 9949 9860 10029 9870
rect 10133 9926 10213 9936
rect 10133 9870 10145 9926
rect 10201 9870 10213 9926
rect 10133 9860 10213 9870
rect 10278 9804 10346 10134
rect 10721 10124 10791 10136
rect 10237 9796 10346 9804
rect 10225 9794 10346 9796
rect 10225 9674 10237 9794
rect 10293 9674 10346 9794
rect 10225 9672 10346 9674
rect 10237 9664 10293 9672
rect 9540 9407 10436 9419
rect 9540 9351 9552 9407
rect 9608 9351 10370 9407
rect 10426 9351 10436 9407
rect 9540 9339 10436 9351
rect 9225 9288 9305 9298
rect 9225 9232 9237 9288
rect 9293 9232 9305 9288
rect 9225 9230 9305 9232
rect 9059 9178 9129 9181
rect 9059 9124 9061 9178
rect 9117 9124 9129 9178
rect 9059 9112 9129 9124
rect 8199 9071 8945 9083
rect 8199 9015 8567 9071
rect 8623 9015 8945 9071
rect 8199 9003 8945 9015
rect 8199 8750 8255 9003
rect 8567 8750 8623 9003
rect 8889 8750 8945 9003
rect 8187 8748 8267 8750
rect 8187 8628 8199 8748
rect 8255 8628 8267 8748
rect 8187 8626 8267 8628
rect 8555 8748 8635 8750
rect 8555 8628 8567 8748
rect 8623 8628 8635 8748
rect 8555 8626 8635 8628
rect 8877 8748 8957 8750
rect 8877 8627 8889 8748
rect 8945 8627 8957 8748
rect 8199 8618 8255 8626
rect 8567 8618 8623 8626
rect 8877 8625 8957 8627
rect 8889 8617 8945 8625
rect 8383 8450 8439 8458
rect 8751 8450 8807 8458
rect 8371 8448 8860 8450
rect 8371 8328 8383 8448
rect 8439 8328 8751 8448
rect 8807 8328 8860 8448
rect 8371 8326 8860 8328
rect 8383 8318 8439 8326
rect 8751 8318 8860 8326
rect 8279 8252 8359 8262
rect 8279 8196 8291 8252
rect 8347 8196 8359 8252
rect 8279 8186 8359 8196
rect 8463 8252 8543 8262
rect 8463 8196 8475 8252
rect 8531 8196 8543 8252
rect 8463 8186 8543 8196
rect 8647 8252 8727 8262
rect 8647 8196 8659 8252
rect 8715 8196 8727 8252
rect 8647 8186 8727 8196
rect 8291 8104 8347 8186
rect 8279 8102 8359 8104
rect 8279 8046 8291 8102
rect 8347 8046 8359 8102
rect 8279 8044 8359 8046
rect 7471 7986 7541 8000
rect 7471 7930 7483 7986
rect 7539 7930 7541 7986
rect 7471 7918 7541 7930
rect 7305 7870 7385 7882
rect 7305 7814 7317 7870
rect 7373 7814 7385 7870
rect 7305 7802 7385 7814
rect 7169 7083 7239 7095
rect 7483 7087 7539 7918
rect 8291 7730 8347 8044
rect 8475 7988 8531 8186
rect 8463 7986 8543 7988
rect 8463 7930 8475 7986
rect 8531 7930 8543 7986
rect 8463 7928 8543 7930
rect 8475 7730 8531 7928
rect 8659 7872 8715 8186
rect 8792 7988 8860 8318
rect 9237 7998 9293 9230
rect 8792 7986 8872 7988
rect 8792 7930 8804 7986
rect 8860 7930 8872 7986
rect 8792 7928 8872 7930
rect 9235 7986 9295 7998
rect 9235 7930 9237 7986
rect 9293 7930 9295 7986
rect 8647 7870 8727 7872
rect 8647 7814 8659 7870
rect 8715 7814 8727 7870
rect 8647 7812 8727 7814
rect 8659 7730 8715 7812
rect 8279 7720 8359 7730
rect 8279 7664 8291 7720
rect 8347 7664 8359 7720
rect 8279 7654 8359 7664
rect 8463 7720 8543 7730
rect 8463 7664 8475 7720
rect 8531 7664 8543 7720
rect 8463 7654 8543 7664
rect 8647 7720 8727 7730
rect 8647 7664 8659 7720
rect 8715 7664 8727 7720
rect 8647 7654 8727 7664
rect 8792 7598 8860 7928
rect 9235 7918 9295 7930
rect 8751 7590 8860 7598
rect 8739 7588 8860 7590
rect 8739 7468 8751 7588
rect 8807 7468 8860 7588
rect 8739 7466 8860 7468
rect 8751 7458 8807 7466
rect 8054 7201 8952 7213
rect 8054 7145 8066 7201
rect 8122 7145 8884 7201
rect 8940 7145 8952 7201
rect 8054 7133 8952 7145
rect 7169 7027 7181 7083
rect 7237 7027 7239 7083
rect 7169 7015 7239 7027
rect 7481 7083 7541 7087
rect 7481 7027 7483 7083
rect 7539 7027 7541 7083
rect 7481 7015 7541 7027
rect 7045 6810 7101 6820
rect 11087 6920 11143 11426
rect 11223 7095 11279 15889
rect 12241 15686 12987 15698
rect 12241 15630 12609 15686
rect 12665 15630 12987 15686
rect 12241 15618 12987 15630
rect 12241 15365 12297 15618
rect 12609 15365 12665 15618
rect 12931 15365 12987 15618
rect 12229 15363 12309 15365
rect 12229 15243 12241 15363
rect 12297 15243 12309 15363
rect 12229 15241 12309 15243
rect 12597 15363 12677 15365
rect 12597 15243 12609 15363
rect 12665 15243 12677 15363
rect 12597 15241 12677 15243
rect 12919 15363 12999 15365
rect 12919 15242 12931 15363
rect 12987 15242 12999 15363
rect 12241 15233 12297 15241
rect 12609 15233 12665 15241
rect 12919 15240 12999 15242
rect 12931 15232 12987 15240
rect 12425 15065 12481 15073
rect 12793 15065 12849 15073
rect 12413 15063 12902 15065
rect 12413 14943 12425 15063
rect 12481 14943 12793 15063
rect 12849 14943 12902 15063
rect 12413 14941 12902 14943
rect 12425 14933 12481 14941
rect 12793 14933 12902 14941
rect 12321 14867 12401 14877
rect 12321 14811 12333 14867
rect 12389 14811 12401 14867
rect 12321 14801 12401 14811
rect 12505 14867 12585 14877
rect 12505 14811 12517 14867
rect 12573 14811 12585 14867
rect 12505 14801 12585 14811
rect 12689 14867 12769 14877
rect 12689 14811 12701 14867
rect 12757 14811 12769 14867
rect 12689 14801 12769 14811
rect 11433 14717 11519 14729
rect 12333 14719 12389 14801
rect 11433 14661 11445 14717
rect 11501 14661 11519 14717
rect 11433 14649 11519 14661
rect 12321 14717 12401 14719
rect 12321 14661 12333 14717
rect 12389 14661 12401 14717
rect 12321 14659 12401 14661
rect 11649 14601 11719 14613
rect 11649 14545 11661 14601
rect 11717 14545 11719 14601
rect 11649 14533 11719 14545
rect 11513 12396 11583 12410
rect 11513 12340 11525 12396
rect 11581 12340 11583 12396
rect 11513 12328 11583 12340
rect 11347 12208 11427 12218
rect 11347 12152 11359 12208
rect 11415 12152 11427 12208
rect 11347 12150 11427 12152
rect 11359 7882 11415 12150
rect 11525 8000 11581 12328
rect 11661 10087 11717 14533
rect 12333 14345 12389 14659
rect 12517 14603 12573 14801
rect 12505 14601 12585 14603
rect 12505 14545 12517 14601
rect 12573 14545 12585 14601
rect 12505 14543 12585 14545
rect 12517 14345 12573 14543
rect 12701 14487 12757 14801
rect 12834 14603 12902 14933
rect 12834 14601 12914 14603
rect 12834 14545 12846 14601
rect 12902 14545 12914 14601
rect 12834 14543 12914 14545
rect 13101 14601 13171 14613
rect 13101 14545 13103 14601
rect 13159 14545 13171 14601
rect 12689 14485 12769 14487
rect 12689 14429 12701 14485
rect 12757 14429 12769 14485
rect 12689 14427 12769 14429
rect 12701 14345 12757 14427
rect 12321 14335 12401 14345
rect 12321 14279 12333 14335
rect 12389 14279 12401 14335
rect 12321 14269 12401 14279
rect 12505 14335 12585 14345
rect 12505 14279 12517 14335
rect 12573 14279 12585 14335
rect 12505 14269 12585 14279
rect 12689 14335 12769 14345
rect 12689 14279 12701 14335
rect 12757 14279 12769 14335
rect 12689 14269 12769 14279
rect 12834 14213 12902 14543
rect 13101 14535 13171 14545
rect 12793 14205 12902 14213
rect 12781 14203 12902 14205
rect 12781 14083 12793 14203
rect 12849 14083 12902 14203
rect 12781 14081 12902 14083
rect 12793 14073 12849 14081
rect 12096 13816 12994 13828
rect 12096 13760 12108 13816
rect 12164 13760 12926 13816
rect 12982 13760 12994 13816
rect 12096 13748 12994 13760
rect 13103 13591 13159 14535
rect 13267 13698 13347 13708
rect 13267 13642 13279 13698
rect 13335 13642 13347 13698
rect 13267 13640 13347 13642
rect 13101 13588 13171 13591
rect 13101 13534 13103 13588
rect 13159 13534 13171 13588
rect 13101 13522 13171 13534
rect 12241 13481 12987 13493
rect 12241 13425 12609 13481
rect 12665 13425 12987 13481
rect 12241 13413 12987 13425
rect 12241 13160 12297 13413
rect 12609 13160 12665 13413
rect 12931 13160 12987 13413
rect 12229 13158 12309 13160
rect 12229 13038 12241 13158
rect 12297 13038 12309 13158
rect 12229 13036 12309 13038
rect 12597 13158 12677 13160
rect 12597 13038 12609 13158
rect 12665 13038 12677 13158
rect 12597 13036 12677 13038
rect 12919 13158 12999 13160
rect 12919 13037 12931 13158
rect 12987 13037 12999 13158
rect 12241 13028 12297 13036
rect 12609 13028 12665 13036
rect 12919 13035 12999 13037
rect 12931 13027 12987 13035
rect 12425 12860 12481 12868
rect 12793 12860 12849 12868
rect 12413 12858 12902 12860
rect 12413 12738 12425 12858
rect 12481 12738 12793 12858
rect 12849 12738 12902 12858
rect 12413 12736 12902 12738
rect 12425 12728 12481 12736
rect 12793 12728 12902 12736
rect 12321 12662 12401 12672
rect 12321 12606 12333 12662
rect 12389 12606 12401 12662
rect 12321 12596 12401 12606
rect 12505 12662 12585 12672
rect 12505 12606 12517 12662
rect 12573 12606 12585 12662
rect 12505 12596 12585 12606
rect 12689 12662 12769 12672
rect 12689 12606 12701 12662
rect 12757 12606 12769 12662
rect 12689 12596 12769 12606
rect 12333 12514 12389 12596
rect 12321 12512 12401 12514
rect 12321 12456 12333 12512
rect 12389 12456 12401 12512
rect 12321 12454 12401 12456
rect 12333 12140 12389 12454
rect 12517 12398 12573 12596
rect 12505 12396 12585 12398
rect 12505 12340 12517 12396
rect 12573 12340 12585 12396
rect 12505 12338 12585 12340
rect 12517 12140 12573 12338
rect 12701 12282 12757 12596
rect 12834 12398 12902 12728
rect 13279 12406 13335 13640
rect 13727 13481 14473 13493
rect 13727 13425 14095 13481
rect 14151 13425 14473 13481
rect 13727 13413 14473 13425
rect 13727 13160 13783 13413
rect 14095 13160 14151 13413
rect 14417 13160 14473 13413
rect 13715 13158 13795 13160
rect 13715 13038 13727 13158
rect 13783 13038 13795 13158
rect 13715 13036 13795 13038
rect 14083 13158 14163 13160
rect 14083 13038 14095 13158
rect 14151 13038 14163 13158
rect 14083 13036 14163 13038
rect 14405 13158 14485 13160
rect 14405 13037 14417 13158
rect 14473 13037 14485 13158
rect 13727 13028 13783 13036
rect 14095 13028 14151 13036
rect 14405 13035 14485 13037
rect 14417 13027 14473 13035
rect 13911 12860 13967 12868
rect 14279 12860 14335 12868
rect 13899 12858 14388 12860
rect 13899 12738 13911 12858
rect 13967 12738 14279 12858
rect 14335 12738 14388 12858
rect 13899 12736 14388 12738
rect 13911 12728 13967 12736
rect 14279 12728 14388 12736
rect 13807 12662 13887 12672
rect 13807 12606 13819 12662
rect 13875 12606 13887 12662
rect 13807 12596 13887 12606
rect 13991 12662 14071 12672
rect 13991 12606 14003 12662
rect 14059 12606 14071 12662
rect 13991 12596 14071 12606
rect 14175 12662 14255 12672
rect 14175 12606 14187 12662
rect 14243 12606 14255 12662
rect 14175 12596 14255 12606
rect 13819 12514 13875 12596
rect 13807 12512 13887 12514
rect 13807 12456 13819 12512
rect 13875 12456 13887 12512
rect 13807 12454 13887 12456
rect 12834 12396 12914 12398
rect 12834 12340 12846 12396
rect 12902 12340 12914 12396
rect 12834 12338 12914 12340
rect 13277 12396 13337 12406
rect 13277 12340 13279 12396
rect 13335 12340 13337 12396
rect 12689 12280 12769 12282
rect 12689 12224 12701 12280
rect 12757 12224 12769 12280
rect 12689 12222 12769 12224
rect 12701 12140 12757 12222
rect 12321 12130 12401 12140
rect 12321 12074 12333 12130
rect 12389 12074 12401 12130
rect 12321 12064 12401 12074
rect 12505 12130 12585 12140
rect 12505 12074 12517 12130
rect 12573 12074 12585 12130
rect 12505 12064 12585 12074
rect 12689 12130 12769 12140
rect 12689 12074 12701 12130
rect 12757 12074 12769 12130
rect 12689 12064 12769 12074
rect 12834 12008 12902 12338
rect 13277 12328 13337 12340
rect 12793 12000 12902 12008
rect 12781 11998 12902 12000
rect 12781 11878 12793 11998
rect 12849 11878 12902 11998
rect 12781 11876 12902 11878
rect 12793 11868 12849 11876
rect 12096 11611 12992 11623
rect 12096 11555 12108 11611
rect 12164 11555 12926 11611
rect 12982 11555 12992 11611
rect 12096 11543 12992 11555
rect 13279 11385 13335 12328
rect 13819 12140 13875 12454
rect 14003 12398 14059 12596
rect 13991 12396 14071 12398
rect 13991 12340 14003 12396
rect 14059 12340 14071 12396
rect 13991 12338 14071 12340
rect 14003 12140 14059 12338
rect 14187 12282 14243 12596
rect 14320 12398 14388 12728
rect 14320 12396 14400 12398
rect 14320 12340 14332 12396
rect 14388 12340 14400 12396
rect 14320 12338 14400 12340
rect 14587 12396 14657 12408
rect 14587 12340 14589 12396
rect 14645 12340 14913 12396
rect 14175 12280 14255 12282
rect 14175 12224 14187 12280
rect 14243 12224 14255 12280
rect 14175 12222 14255 12224
rect 14187 12140 14243 12222
rect 13807 12130 13887 12140
rect 13807 12074 13819 12130
rect 13875 12074 13887 12130
rect 13807 12064 13887 12074
rect 13991 12130 14071 12140
rect 13991 12074 14003 12130
rect 14059 12074 14071 12130
rect 13991 12064 14071 12074
rect 14175 12130 14255 12140
rect 14175 12074 14187 12130
rect 14243 12074 14255 12130
rect 14175 12064 14255 12074
rect 14320 12008 14388 12338
rect 14587 12330 14657 12340
rect 14279 12000 14388 12008
rect 14267 11998 14388 12000
rect 14267 11878 14279 11998
rect 14335 11878 14388 11998
rect 14267 11876 14388 11878
rect 14279 11868 14335 11876
rect 13582 11611 14478 11623
rect 13582 11555 13594 11611
rect 13650 11555 14412 11611
rect 14468 11555 14478 11611
rect 13582 11543 14478 11555
rect 14589 11386 14645 12330
rect 14753 11494 14833 11504
rect 14753 11438 14765 11494
rect 14821 11438 14833 11494
rect 14753 11436 14833 11438
rect 13277 11383 13347 11385
rect 13277 11327 13279 11383
rect 13335 11327 13347 11383
rect 13277 11315 13347 11327
rect 14577 11384 14657 11386
rect 14577 11328 14589 11384
rect 14645 11328 14657 11384
rect 14577 11316 14657 11328
rect 12241 11276 12987 11288
rect 12241 11220 12609 11276
rect 12665 11220 12987 11276
rect 12241 11208 12987 11220
rect 12241 10955 12297 11208
rect 12609 10955 12665 11208
rect 12931 10955 12987 11208
rect 13727 11277 14473 11289
rect 13727 11221 14095 11277
rect 14151 11221 14473 11277
rect 13727 11209 14473 11221
rect 13727 10956 13783 11209
rect 14095 10956 14151 11209
rect 14417 10956 14473 11209
rect 12229 10953 12309 10955
rect 12229 10833 12241 10953
rect 12297 10833 12309 10953
rect 12229 10831 12309 10833
rect 12597 10953 12677 10955
rect 12597 10833 12609 10953
rect 12665 10833 12677 10953
rect 12597 10831 12677 10833
rect 12919 10953 12999 10955
rect 12919 10832 12931 10953
rect 12987 10832 12999 10953
rect 13715 10954 13795 10956
rect 13715 10834 13727 10954
rect 13783 10834 13795 10954
rect 13715 10832 13795 10834
rect 14083 10954 14163 10956
rect 14083 10834 14095 10954
rect 14151 10834 14163 10954
rect 14083 10832 14163 10834
rect 14405 10954 14485 10956
rect 14405 10833 14417 10954
rect 14473 10833 14485 10954
rect 12241 10823 12297 10831
rect 12609 10823 12665 10831
rect 12919 10830 12999 10832
rect 12931 10822 12987 10830
rect 13727 10824 13783 10832
rect 14095 10824 14151 10832
rect 14405 10831 14485 10833
rect 14417 10823 14473 10831
rect 12425 10655 12481 10663
rect 12793 10655 12849 10663
rect 13911 10656 13967 10664
rect 14279 10656 14335 10664
rect 12413 10653 12902 10655
rect 12413 10533 12425 10653
rect 12481 10533 12793 10653
rect 12849 10533 12902 10653
rect 12413 10531 12902 10533
rect 13899 10654 14388 10656
rect 13899 10534 13911 10654
rect 13967 10534 14279 10654
rect 14335 10534 14388 10654
rect 13899 10532 14388 10534
rect 12425 10523 12481 10531
rect 12793 10523 12902 10531
rect 13911 10524 13967 10532
rect 14279 10524 14388 10532
rect 12321 10457 12401 10467
rect 12321 10401 12333 10457
rect 12389 10401 12401 10457
rect 12321 10391 12401 10401
rect 12505 10457 12585 10467
rect 12505 10401 12517 10457
rect 12573 10401 12585 10457
rect 12505 10391 12585 10401
rect 12689 10457 12769 10467
rect 12689 10401 12701 10457
rect 12757 10401 12769 10457
rect 12689 10391 12769 10401
rect 12333 10309 12389 10391
rect 12321 10307 12401 10309
rect 12321 10251 12333 10307
rect 12389 10251 12401 10307
rect 12321 10249 12401 10251
rect 11649 10075 11719 10087
rect 11649 10019 11661 10075
rect 11717 10019 11719 10075
rect 11649 10007 11719 10019
rect 12333 9935 12389 10249
rect 12517 10193 12573 10391
rect 12505 10191 12585 10193
rect 12505 10135 12517 10191
rect 12573 10135 12585 10191
rect 12505 10133 12585 10135
rect 12517 9935 12573 10133
rect 12701 10077 12757 10391
rect 12834 10193 12902 10523
rect 13807 10458 13887 10468
rect 13807 10402 13819 10458
rect 13875 10402 13887 10458
rect 13807 10392 13887 10402
rect 13991 10458 14071 10468
rect 13991 10402 14003 10458
rect 14059 10402 14071 10458
rect 13991 10392 14071 10402
rect 14175 10458 14255 10468
rect 14175 10402 14187 10458
rect 14243 10402 14255 10458
rect 14175 10392 14255 10402
rect 13819 10310 13875 10392
rect 13807 10308 13887 10310
rect 13807 10252 13819 10308
rect 13875 10252 13887 10308
rect 13807 10250 13887 10252
rect 12834 10191 12914 10193
rect 12834 10135 12846 10191
rect 12902 10135 12914 10191
rect 12834 10133 12914 10135
rect 13101 10191 13171 10203
rect 13101 10135 13103 10191
rect 13159 10135 13171 10191
rect 12689 10075 12769 10077
rect 12689 10019 12701 10075
rect 12757 10019 12769 10075
rect 12689 10017 12769 10019
rect 12701 9935 12757 10017
rect 12321 9925 12401 9935
rect 12321 9869 12333 9925
rect 12389 9869 12401 9925
rect 12321 9859 12401 9869
rect 12505 9925 12585 9935
rect 12505 9869 12517 9925
rect 12573 9869 12585 9925
rect 12505 9859 12585 9869
rect 12689 9925 12769 9935
rect 12689 9869 12701 9925
rect 12757 9869 12769 9925
rect 12689 9859 12769 9869
rect 12834 9803 12902 10133
rect 13101 10125 13171 10135
rect 12793 9795 12902 9803
rect 12781 9793 12902 9795
rect 12781 9673 12793 9793
rect 12849 9673 12902 9793
rect 12781 9671 12902 9673
rect 12793 9663 12849 9671
rect 12096 9406 12992 9418
rect 12096 9350 12108 9406
rect 12164 9350 12926 9406
rect 12982 9350 12992 9406
rect 12096 9338 12992 9350
rect 13103 9181 13159 10125
rect 13819 9936 13875 10250
rect 14003 10194 14059 10392
rect 13991 10192 14071 10194
rect 13991 10136 14003 10192
rect 14059 10136 14071 10192
rect 13991 10134 14071 10136
rect 14003 9936 14059 10134
rect 14187 10078 14243 10392
rect 14320 10194 14388 10524
rect 14765 10202 14821 11436
rect 14320 10192 14400 10194
rect 14320 10136 14332 10192
rect 14388 10136 14400 10192
rect 14320 10134 14400 10136
rect 14763 10192 14833 10202
rect 14993 10192 15049 24235
rect 15195 21984 15251 25664
rect 19235 25546 19305 25558
rect 19235 25490 19237 25546
rect 19293 25490 19305 25546
rect 19235 25488 19305 25490
rect 16283 25262 17029 25274
rect 16283 25206 16651 25262
rect 16707 25206 17029 25262
rect 16283 25194 17029 25206
rect 16283 24941 16339 25194
rect 16651 24941 16707 25194
rect 16973 24941 17029 25194
rect 16271 24939 16351 24941
rect 16271 24819 16283 24939
rect 16339 24819 16351 24939
rect 16271 24817 16351 24819
rect 16639 24939 16719 24941
rect 16639 24819 16651 24939
rect 16707 24819 16719 24939
rect 16639 24817 16719 24819
rect 16961 24939 17041 24941
rect 16961 24818 16973 24939
rect 17029 24818 17041 24939
rect 16283 24809 16339 24817
rect 16651 24809 16707 24817
rect 16961 24816 17041 24818
rect 16973 24808 17029 24816
rect 16467 24641 16523 24649
rect 16835 24641 16891 24649
rect 16455 24639 16944 24641
rect 16455 24519 16467 24639
rect 16523 24519 16835 24639
rect 16891 24519 16944 24639
rect 16455 24517 16944 24519
rect 16467 24509 16523 24517
rect 16835 24509 16944 24517
rect 16363 24443 16443 24453
rect 16363 24387 16375 24443
rect 16431 24387 16443 24443
rect 16363 24377 16443 24387
rect 16547 24443 16627 24453
rect 16547 24387 16559 24443
rect 16615 24387 16627 24443
rect 16547 24377 16627 24387
rect 16731 24443 16811 24453
rect 16731 24387 16743 24443
rect 16799 24387 16811 24443
rect 16731 24377 16811 24387
rect 16375 24295 16431 24377
rect 16363 24293 16443 24295
rect 16363 24237 16375 24293
rect 16431 24237 16443 24293
rect 16363 24235 16443 24237
rect 15691 24177 15761 24189
rect 15691 24121 15703 24177
rect 15759 24121 15761 24177
rect 15691 24109 15761 24121
rect 15193 21972 15263 21984
rect 15193 21916 15195 21972
rect 15251 21916 15263 21972
rect 15193 21904 15263 21916
rect 15555 21972 15625 21986
rect 15555 21916 15567 21972
rect 15623 21916 15625 21972
rect 15555 21904 15625 21916
rect 15375 21070 15453 21082
rect 15375 21014 15386 21070
rect 15442 21014 15453 21070
rect 15375 21002 15453 21014
rect 15567 17576 15623 21904
rect 15703 19663 15759 24109
rect 16375 23921 16431 24235
rect 16559 24179 16615 24377
rect 16547 24177 16627 24179
rect 16547 24121 16559 24177
rect 16615 24121 16627 24177
rect 16547 24119 16627 24121
rect 16559 23921 16615 24119
rect 16743 24063 16799 24377
rect 16876 24179 16944 24509
rect 16876 24177 16956 24179
rect 16876 24121 16888 24177
rect 16944 24121 16956 24177
rect 16876 24119 16956 24121
rect 17143 24177 17213 24189
rect 17143 24121 17145 24177
rect 17201 24121 17213 24177
rect 16731 24061 16811 24063
rect 16731 24005 16743 24061
rect 16799 24005 16811 24061
rect 16731 24003 16811 24005
rect 16743 23921 16799 24003
rect 16363 23911 16443 23921
rect 16363 23855 16375 23911
rect 16431 23855 16443 23911
rect 16363 23845 16443 23855
rect 16547 23911 16627 23921
rect 16547 23855 16559 23911
rect 16615 23855 16627 23911
rect 16547 23845 16627 23855
rect 16731 23911 16811 23921
rect 16731 23855 16743 23911
rect 16799 23855 16811 23911
rect 16731 23845 16811 23855
rect 16876 23789 16944 24119
rect 17143 24111 17213 24121
rect 16835 23781 16944 23789
rect 16823 23779 16944 23781
rect 16823 23659 16835 23779
rect 16891 23659 16944 23779
rect 16823 23657 16944 23659
rect 16835 23649 16891 23657
rect 16138 23392 17036 23404
rect 16138 23336 16150 23392
rect 16206 23336 16968 23392
rect 17024 23336 17036 23392
rect 16138 23324 17036 23336
rect 17145 23167 17201 24111
rect 17309 23274 17389 23284
rect 17309 23218 17321 23274
rect 17377 23218 17389 23274
rect 17309 23216 17389 23218
rect 17143 23164 17213 23167
rect 17143 23110 17145 23164
rect 17201 23110 17213 23164
rect 17143 23098 17213 23110
rect 16283 23057 17029 23069
rect 16283 23001 16651 23057
rect 16707 23001 17029 23057
rect 16283 22989 17029 23001
rect 16283 22736 16339 22989
rect 16651 22736 16707 22989
rect 16973 22736 17029 22989
rect 16271 22734 16351 22736
rect 16271 22614 16283 22734
rect 16339 22614 16351 22734
rect 16271 22612 16351 22614
rect 16639 22734 16719 22736
rect 16639 22614 16651 22734
rect 16707 22614 16719 22734
rect 16639 22612 16719 22614
rect 16961 22734 17041 22736
rect 16961 22613 16973 22734
rect 17029 22613 17041 22734
rect 16283 22604 16339 22612
rect 16651 22604 16707 22612
rect 16961 22611 17041 22613
rect 16973 22603 17029 22611
rect 16467 22436 16523 22444
rect 16835 22436 16891 22444
rect 16455 22434 16944 22436
rect 16455 22314 16467 22434
rect 16523 22314 16835 22434
rect 16891 22314 16944 22434
rect 16455 22312 16944 22314
rect 16467 22304 16523 22312
rect 16835 22304 16944 22312
rect 16363 22238 16443 22248
rect 16363 22182 16375 22238
rect 16431 22182 16443 22238
rect 16363 22172 16443 22182
rect 16547 22238 16627 22248
rect 16547 22182 16559 22238
rect 16615 22182 16627 22238
rect 16547 22172 16627 22182
rect 16731 22238 16811 22248
rect 16731 22182 16743 22238
rect 16799 22182 16811 22238
rect 16731 22172 16811 22182
rect 16375 22090 16431 22172
rect 16363 22088 16443 22090
rect 16363 22032 16375 22088
rect 16431 22032 16443 22088
rect 16363 22030 16443 22032
rect 16375 21716 16431 22030
rect 16559 21974 16615 22172
rect 16547 21972 16627 21974
rect 16547 21916 16559 21972
rect 16615 21916 16627 21972
rect 16547 21914 16627 21916
rect 16559 21716 16615 21914
rect 16743 21858 16799 22172
rect 16876 21974 16944 22304
rect 17321 21982 17377 23216
rect 17769 23057 18515 23069
rect 17769 23001 18137 23057
rect 18193 23001 18515 23057
rect 17769 22989 18515 23001
rect 17769 22736 17825 22989
rect 18137 22736 18193 22989
rect 18459 22736 18515 22989
rect 17757 22734 17837 22736
rect 17757 22614 17769 22734
rect 17825 22614 17837 22734
rect 17757 22612 17837 22614
rect 18125 22734 18205 22736
rect 18125 22614 18137 22734
rect 18193 22614 18205 22734
rect 18125 22612 18205 22614
rect 18447 22734 18527 22736
rect 18447 22613 18459 22734
rect 18515 22613 18527 22734
rect 17769 22604 17825 22612
rect 18137 22604 18193 22612
rect 18447 22611 18527 22613
rect 18459 22603 18515 22611
rect 17953 22436 18009 22444
rect 18321 22436 18377 22444
rect 17941 22434 18430 22436
rect 17941 22314 17953 22434
rect 18009 22314 18321 22434
rect 18377 22314 18430 22434
rect 17941 22312 18430 22314
rect 17953 22304 18009 22312
rect 18321 22304 18430 22312
rect 17849 22238 17929 22248
rect 17849 22182 17861 22238
rect 17917 22182 17929 22238
rect 17849 22172 17929 22182
rect 18033 22238 18113 22248
rect 18033 22182 18045 22238
rect 18101 22182 18113 22238
rect 18033 22172 18113 22182
rect 18217 22238 18297 22248
rect 18217 22182 18229 22238
rect 18285 22182 18297 22238
rect 18217 22172 18297 22182
rect 17861 22090 17917 22172
rect 17849 22088 17929 22090
rect 17849 22032 17861 22088
rect 17917 22032 17929 22088
rect 17849 22030 17929 22032
rect 16876 21972 16956 21974
rect 16876 21916 16888 21972
rect 16944 21916 16956 21972
rect 16876 21914 16956 21916
rect 17319 21972 17379 21982
rect 17319 21916 17321 21972
rect 17377 21916 17379 21972
rect 16731 21856 16811 21858
rect 16731 21800 16743 21856
rect 16799 21800 16811 21856
rect 16731 21798 16811 21800
rect 16743 21716 16799 21798
rect 16363 21706 16443 21716
rect 16363 21650 16375 21706
rect 16431 21650 16443 21706
rect 16363 21640 16443 21650
rect 16547 21706 16627 21716
rect 16547 21650 16559 21706
rect 16615 21650 16627 21706
rect 16547 21640 16627 21650
rect 16731 21706 16811 21716
rect 16731 21650 16743 21706
rect 16799 21650 16811 21706
rect 16731 21640 16811 21650
rect 16876 21584 16944 21914
rect 17319 21904 17379 21916
rect 16835 21576 16944 21584
rect 16823 21574 16944 21576
rect 16823 21454 16835 21574
rect 16891 21454 16944 21574
rect 16823 21452 16944 21454
rect 16835 21444 16891 21452
rect 16138 21187 17034 21199
rect 16138 21131 16150 21187
rect 16206 21131 16968 21187
rect 17024 21131 17034 21187
rect 16138 21119 17034 21131
rect 17321 20961 17377 21904
rect 17861 21716 17917 22030
rect 18045 21974 18101 22172
rect 18033 21972 18113 21974
rect 18033 21916 18045 21972
rect 18101 21916 18113 21972
rect 18033 21914 18113 21916
rect 18045 21716 18101 21914
rect 18229 21858 18285 22172
rect 18362 21974 18430 22304
rect 19237 21984 19293 25488
rect 18362 21972 18442 21974
rect 18362 21916 18374 21972
rect 18430 21916 18442 21972
rect 18362 21914 18442 21916
rect 18629 21972 18699 21984
rect 19235 21972 19305 21984
rect 18629 21916 18631 21972
rect 18687 21916 18955 21972
rect 19235 21916 19237 21972
rect 19293 21916 19305 21972
rect 18217 21856 18297 21858
rect 18217 21800 18229 21856
rect 18285 21800 18297 21856
rect 18217 21798 18297 21800
rect 18229 21716 18285 21798
rect 17849 21706 17929 21716
rect 17849 21650 17861 21706
rect 17917 21650 17929 21706
rect 17849 21640 17929 21650
rect 18033 21706 18113 21716
rect 18033 21650 18045 21706
rect 18101 21650 18113 21706
rect 18033 21640 18113 21650
rect 18217 21706 18297 21716
rect 18217 21650 18229 21706
rect 18285 21650 18297 21706
rect 18217 21640 18297 21650
rect 18362 21584 18430 21914
rect 18629 21906 18699 21916
rect 18321 21576 18430 21584
rect 18309 21574 18430 21576
rect 18309 21454 18321 21574
rect 18377 21454 18430 21574
rect 18309 21452 18430 21454
rect 18321 21444 18377 21452
rect 17624 21187 18520 21199
rect 17624 21131 17636 21187
rect 17692 21131 18454 21187
rect 18510 21131 18520 21187
rect 17624 21119 18520 21131
rect 18631 20962 18687 21906
rect 19235 21904 19305 21916
rect 18795 21070 18875 21080
rect 18795 21014 18807 21070
rect 18863 21014 18875 21070
rect 18795 21012 18875 21014
rect 17319 20959 17389 20961
rect 17319 20903 17321 20959
rect 17377 20903 17389 20959
rect 17319 20891 17389 20903
rect 18619 20960 18699 20962
rect 18619 20904 18631 20960
rect 18687 20904 18699 20960
rect 18619 20892 18699 20904
rect 16283 20852 17029 20864
rect 16283 20796 16651 20852
rect 16707 20796 17029 20852
rect 16283 20784 17029 20796
rect 16283 20531 16339 20784
rect 16651 20531 16707 20784
rect 16973 20531 17029 20784
rect 17769 20853 18515 20865
rect 17769 20797 18137 20853
rect 18193 20797 18515 20853
rect 17769 20785 18515 20797
rect 17769 20532 17825 20785
rect 18137 20532 18193 20785
rect 18459 20532 18515 20785
rect 16271 20529 16351 20531
rect 16271 20409 16283 20529
rect 16339 20409 16351 20529
rect 16271 20407 16351 20409
rect 16639 20529 16719 20531
rect 16639 20409 16651 20529
rect 16707 20409 16719 20529
rect 16639 20407 16719 20409
rect 16961 20529 17041 20531
rect 16961 20408 16973 20529
rect 17029 20408 17041 20529
rect 17757 20530 17837 20532
rect 17757 20410 17769 20530
rect 17825 20410 17837 20530
rect 17757 20408 17837 20410
rect 18125 20530 18205 20532
rect 18125 20410 18137 20530
rect 18193 20410 18205 20530
rect 18125 20408 18205 20410
rect 18447 20530 18527 20532
rect 18447 20409 18459 20530
rect 18515 20409 18527 20530
rect 16283 20399 16339 20407
rect 16651 20399 16707 20407
rect 16961 20406 17041 20408
rect 16973 20398 17029 20406
rect 17769 20400 17825 20408
rect 18137 20400 18193 20408
rect 18447 20407 18527 20409
rect 18459 20399 18515 20407
rect 16467 20231 16523 20239
rect 16835 20231 16891 20239
rect 17953 20232 18009 20240
rect 18321 20232 18377 20240
rect 16455 20229 16944 20231
rect 16455 20109 16467 20229
rect 16523 20109 16835 20229
rect 16891 20109 16944 20229
rect 16455 20107 16944 20109
rect 17941 20230 18430 20232
rect 17941 20110 17953 20230
rect 18009 20110 18321 20230
rect 18377 20110 18430 20230
rect 17941 20108 18430 20110
rect 16467 20099 16523 20107
rect 16835 20099 16944 20107
rect 17953 20100 18009 20108
rect 18321 20100 18430 20108
rect 16363 20033 16443 20043
rect 16363 19977 16375 20033
rect 16431 19977 16443 20033
rect 16363 19967 16443 19977
rect 16547 20033 16627 20043
rect 16547 19977 16559 20033
rect 16615 19977 16627 20033
rect 16547 19967 16627 19977
rect 16731 20033 16811 20043
rect 16731 19977 16743 20033
rect 16799 19977 16811 20033
rect 16731 19967 16811 19977
rect 16375 19885 16431 19967
rect 16363 19883 16443 19885
rect 16363 19827 16375 19883
rect 16431 19827 16443 19883
rect 16363 19825 16443 19827
rect 15691 19651 15761 19663
rect 15691 19595 15703 19651
rect 15759 19595 15761 19651
rect 15691 19583 15761 19595
rect 16375 19511 16431 19825
rect 16559 19769 16615 19967
rect 16547 19767 16627 19769
rect 16547 19711 16559 19767
rect 16615 19711 16627 19767
rect 16547 19709 16627 19711
rect 16559 19511 16615 19709
rect 16743 19653 16799 19967
rect 16876 19769 16944 20099
rect 17849 20034 17929 20044
rect 17849 19978 17861 20034
rect 17917 19978 17929 20034
rect 17849 19968 17929 19978
rect 18033 20034 18113 20044
rect 18033 19978 18045 20034
rect 18101 19978 18113 20034
rect 18033 19968 18113 19978
rect 18217 20034 18297 20044
rect 18217 19978 18229 20034
rect 18285 19978 18297 20034
rect 18217 19968 18297 19978
rect 17861 19886 17917 19968
rect 17849 19884 17929 19886
rect 17849 19828 17861 19884
rect 17917 19828 17929 19884
rect 17849 19826 17929 19828
rect 16876 19767 16956 19769
rect 16876 19711 16888 19767
rect 16944 19711 16956 19767
rect 16876 19709 16956 19711
rect 17143 19767 17213 19779
rect 17143 19711 17145 19767
rect 17201 19711 17213 19767
rect 16731 19651 16811 19653
rect 16731 19595 16743 19651
rect 16799 19595 16811 19651
rect 16731 19593 16811 19595
rect 16743 19511 16799 19593
rect 16363 19501 16443 19511
rect 16363 19445 16375 19501
rect 16431 19445 16443 19501
rect 16363 19435 16443 19445
rect 16547 19501 16627 19511
rect 16547 19445 16559 19501
rect 16615 19445 16627 19501
rect 16547 19435 16627 19445
rect 16731 19501 16811 19511
rect 16731 19445 16743 19501
rect 16799 19445 16811 19501
rect 16731 19435 16811 19445
rect 16876 19379 16944 19709
rect 17143 19701 17213 19711
rect 16835 19371 16944 19379
rect 16823 19369 16944 19371
rect 16823 19249 16835 19369
rect 16891 19249 16944 19369
rect 16823 19247 16944 19249
rect 16835 19239 16891 19247
rect 16138 18982 17034 18994
rect 16138 18926 16150 18982
rect 16206 18926 16968 18982
rect 17024 18926 17034 18982
rect 16138 18914 17034 18926
rect 17145 18757 17201 19701
rect 17861 19512 17917 19826
rect 18045 19770 18101 19968
rect 18033 19768 18113 19770
rect 18033 19712 18045 19768
rect 18101 19712 18113 19768
rect 18033 19710 18113 19712
rect 18045 19512 18101 19710
rect 18229 19654 18285 19968
rect 18362 19770 18430 20100
rect 18807 19778 18863 21012
rect 18362 19768 18442 19770
rect 18362 19712 18374 19768
rect 18430 19712 18442 19768
rect 18362 19710 18442 19712
rect 18805 19768 18875 19778
rect 18805 19712 18807 19768
rect 18863 19712 18955 19768
rect 18217 19652 18297 19654
rect 18217 19596 18229 19652
rect 18285 19596 18297 19652
rect 18217 19594 18297 19596
rect 18229 19512 18285 19594
rect 17849 19502 17929 19512
rect 17849 19446 17861 19502
rect 17917 19446 17929 19502
rect 17849 19436 17929 19446
rect 18033 19502 18113 19512
rect 18033 19446 18045 19502
rect 18101 19446 18113 19502
rect 18033 19436 18113 19446
rect 18217 19502 18297 19512
rect 18217 19446 18229 19502
rect 18285 19446 18297 19502
rect 18217 19436 18297 19446
rect 18362 19380 18430 19710
rect 18805 19700 18875 19712
rect 18321 19372 18430 19380
rect 18309 19370 18430 19372
rect 18309 19250 18321 19370
rect 18377 19250 18430 19370
rect 18309 19248 18430 19250
rect 18321 19240 18377 19248
rect 17624 18983 18520 18995
rect 17624 18927 17636 18983
rect 17692 18927 18454 18983
rect 18510 18927 18520 18983
rect 17624 18915 18520 18927
rect 17309 18864 17389 18874
rect 17309 18808 17321 18864
rect 17377 18808 17389 18864
rect 17309 18806 17389 18808
rect 17143 18754 17213 18757
rect 17143 18700 17145 18754
rect 17201 18700 17213 18754
rect 17143 18688 17213 18700
rect 16283 18647 17029 18659
rect 16283 18591 16651 18647
rect 16707 18591 17029 18647
rect 16283 18579 17029 18591
rect 16283 18326 16339 18579
rect 16651 18326 16707 18579
rect 16973 18326 17029 18579
rect 16271 18324 16351 18326
rect 16271 18204 16283 18324
rect 16339 18204 16351 18324
rect 16271 18202 16351 18204
rect 16639 18324 16719 18326
rect 16639 18204 16651 18324
rect 16707 18204 16719 18324
rect 16639 18202 16719 18204
rect 16961 18324 17041 18326
rect 16961 18203 16973 18324
rect 17029 18203 17041 18324
rect 16283 18194 16339 18202
rect 16651 18194 16707 18202
rect 16961 18201 17041 18203
rect 16973 18193 17029 18201
rect 16467 18026 16523 18034
rect 16835 18026 16891 18034
rect 16455 18024 16944 18026
rect 16455 17904 16467 18024
rect 16523 17904 16835 18024
rect 16891 17904 16944 18024
rect 16455 17902 16944 17904
rect 16467 17894 16523 17902
rect 16835 17894 16944 17902
rect 16363 17828 16443 17838
rect 16363 17772 16375 17828
rect 16431 17772 16443 17828
rect 16363 17762 16443 17772
rect 16547 17828 16627 17838
rect 16547 17772 16559 17828
rect 16615 17772 16627 17828
rect 16547 17762 16627 17772
rect 16731 17828 16811 17838
rect 16731 17772 16743 17828
rect 16799 17772 16811 17828
rect 16731 17762 16811 17772
rect 16375 17680 16431 17762
rect 16363 17678 16443 17680
rect 16363 17622 16375 17678
rect 16431 17622 16443 17678
rect 16363 17620 16443 17622
rect 15555 17562 15625 17576
rect 15555 17506 15567 17562
rect 15623 17506 15625 17562
rect 15555 17494 15625 17506
rect 15375 17446 15453 17458
rect 15375 17390 15386 17446
rect 15442 17390 15453 17446
rect 15375 17378 15453 17390
rect 15253 16659 15323 16671
rect 15567 16663 15623 17494
rect 16375 17306 16431 17620
rect 16559 17564 16615 17762
rect 16547 17562 16627 17564
rect 16547 17506 16559 17562
rect 16615 17506 16627 17562
rect 16547 17504 16627 17506
rect 16559 17306 16615 17504
rect 16743 17448 16799 17762
rect 16876 17564 16944 17894
rect 17321 17574 17377 18806
rect 16876 17562 16956 17564
rect 16876 17506 16888 17562
rect 16944 17506 16956 17562
rect 16876 17504 16956 17506
rect 17319 17562 17379 17574
rect 17319 17506 17321 17562
rect 17377 17506 17379 17562
rect 16731 17446 16811 17448
rect 16731 17390 16743 17446
rect 16799 17390 16811 17446
rect 16731 17388 16811 17390
rect 16743 17306 16799 17388
rect 16363 17296 16443 17306
rect 16363 17240 16375 17296
rect 16431 17240 16443 17296
rect 16363 17230 16443 17240
rect 16547 17296 16627 17306
rect 16547 17240 16559 17296
rect 16615 17240 16627 17296
rect 16547 17230 16627 17240
rect 16731 17296 16811 17306
rect 16731 17240 16743 17296
rect 16799 17240 16811 17296
rect 16731 17230 16811 17240
rect 16876 17174 16944 17504
rect 17319 17494 17379 17506
rect 16835 17166 16944 17174
rect 16823 17164 16944 17166
rect 16823 17044 16835 17164
rect 16891 17044 16944 17164
rect 16823 17042 16944 17044
rect 16835 17034 16891 17042
rect 16138 16777 17036 16789
rect 16138 16721 16150 16777
rect 16206 16721 16968 16777
rect 17024 16721 17036 16777
rect 16138 16709 17036 16721
rect 15253 16603 15265 16659
rect 15321 16603 15323 16659
rect 15253 16591 15323 16603
rect 15565 16659 15625 16663
rect 15565 16603 15567 16659
rect 15623 16603 15625 16659
rect 15565 16591 15625 16603
rect 15265 15989 15321 16591
rect 15265 15879 15321 15889
rect 14763 10136 14765 10192
rect 14821 10136 15049 10192
rect 14175 10076 14255 10078
rect 14175 10020 14187 10076
rect 14243 10020 14255 10076
rect 14175 10018 14255 10020
rect 14187 9936 14243 10018
rect 13807 9926 13887 9936
rect 13807 9870 13819 9926
rect 13875 9870 13887 9926
rect 13807 9860 13887 9870
rect 13991 9926 14071 9936
rect 13991 9870 14003 9926
rect 14059 9870 14071 9926
rect 13991 9860 14071 9870
rect 14175 9926 14255 9936
rect 14175 9870 14187 9926
rect 14243 9870 14255 9926
rect 14175 9860 14255 9870
rect 14320 9804 14388 10134
rect 14763 10124 14833 10136
rect 14279 9796 14388 9804
rect 14267 9794 14388 9796
rect 14267 9674 14279 9794
rect 14335 9674 14388 9794
rect 14267 9672 14388 9674
rect 14279 9664 14335 9672
rect 13582 9407 14478 9419
rect 13582 9351 13594 9407
rect 13650 9351 14412 9407
rect 14468 9351 14478 9407
rect 13582 9339 14478 9351
rect 13267 9288 13347 9298
rect 13267 9232 13279 9288
rect 13335 9232 13347 9288
rect 13267 9230 13347 9232
rect 13101 9178 13171 9181
rect 13101 9124 13103 9178
rect 13159 9124 13171 9178
rect 13101 9112 13171 9124
rect 12241 9071 12987 9083
rect 12241 9015 12609 9071
rect 12665 9015 12987 9071
rect 12241 9003 12987 9015
rect 12241 8750 12297 9003
rect 12609 8750 12665 9003
rect 12931 8750 12987 9003
rect 12229 8748 12309 8750
rect 12229 8628 12241 8748
rect 12297 8628 12309 8748
rect 12229 8626 12309 8628
rect 12597 8748 12677 8750
rect 12597 8628 12609 8748
rect 12665 8628 12677 8748
rect 12597 8626 12677 8628
rect 12919 8748 12999 8750
rect 12919 8627 12931 8748
rect 12987 8627 12999 8748
rect 12241 8618 12297 8626
rect 12609 8618 12665 8626
rect 12919 8625 12999 8627
rect 12931 8617 12987 8625
rect 12425 8450 12481 8458
rect 12793 8450 12849 8458
rect 12413 8448 12902 8450
rect 12413 8328 12425 8448
rect 12481 8328 12793 8448
rect 12849 8328 12902 8448
rect 12413 8326 12902 8328
rect 12425 8318 12481 8326
rect 12793 8318 12902 8326
rect 12321 8252 12401 8262
rect 12321 8196 12333 8252
rect 12389 8196 12401 8252
rect 12321 8186 12401 8196
rect 12505 8252 12585 8262
rect 12505 8196 12517 8252
rect 12573 8196 12585 8252
rect 12505 8186 12585 8196
rect 12689 8252 12769 8262
rect 12689 8196 12701 8252
rect 12757 8196 12769 8252
rect 12689 8186 12769 8196
rect 12333 8104 12389 8186
rect 12321 8102 12401 8104
rect 12321 8046 12333 8102
rect 12389 8046 12401 8102
rect 12321 8044 12401 8046
rect 11513 7986 11583 8000
rect 11513 7930 11525 7986
rect 11581 7930 11583 7986
rect 11513 7918 11583 7930
rect 11347 7870 11427 7882
rect 11347 7814 11359 7870
rect 11415 7814 11427 7870
rect 11347 7802 11427 7814
rect 11211 7083 11281 7095
rect 11525 7087 11581 7918
rect 12333 7730 12389 8044
rect 12517 7988 12573 8186
rect 12505 7986 12585 7988
rect 12505 7930 12517 7986
rect 12573 7930 12585 7986
rect 12505 7928 12585 7930
rect 12517 7730 12573 7928
rect 12701 7872 12757 8186
rect 12834 7988 12902 8318
rect 13279 7998 13335 9230
rect 12834 7986 12914 7988
rect 12834 7930 12846 7986
rect 12902 7930 12914 7986
rect 12834 7928 12914 7930
rect 13277 7986 13337 7998
rect 13277 7930 13279 7986
rect 13335 7930 13337 7986
rect 12689 7870 12769 7872
rect 12689 7814 12701 7870
rect 12757 7814 12769 7870
rect 12689 7812 12769 7814
rect 12701 7730 12757 7812
rect 12321 7720 12401 7730
rect 12321 7664 12333 7720
rect 12389 7664 12401 7720
rect 12321 7654 12401 7664
rect 12505 7720 12585 7730
rect 12505 7664 12517 7720
rect 12573 7664 12585 7720
rect 12505 7654 12585 7664
rect 12689 7720 12769 7730
rect 12689 7664 12701 7720
rect 12757 7664 12769 7720
rect 12689 7654 12769 7664
rect 12834 7598 12902 7928
rect 13277 7918 13337 7930
rect 12793 7590 12902 7598
rect 12781 7588 12902 7590
rect 12781 7468 12793 7588
rect 12849 7468 12902 7588
rect 12781 7466 12902 7468
rect 12793 7458 12849 7466
rect 12096 7201 12994 7213
rect 12096 7145 12108 7201
rect 12164 7145 12926 7201
rect 12982 7145 12994 7201
rect 12096 7133 12994 7145
rect 11211 7027 11223 7083
rect 11279 7027 11281 7083
rect 11211 7015 11281 7027
rect 11523 7083 11583 7087
rect 11523 7027 11525 7083
rect 11581 7027 11583 7083
rect 11523 7015 11583 7027
rect 11087 6810 11143 6820
rect -13680 4940 -13603 4954
rect -13894 4939 -13603 4940
rect -13894 4881 -13665 4939
rect -13607 4881 -13603 4939
rect -13894 4880 -13603 4881
rect -13680 4867 -13603 4880
rect -13722 -1177 -13632 -1166
rect -13880 -1179 -13632 -1177
rect -13880 -1252 -13707 -1179
rect -13634 -1252 -13632 -1179
rect -13722 -1266 -13632 -1252
rect -13717 -1502 -13627 -1491
rect -13878 -1504 -13627 -1502
rect -13878 -1577 -13704 -1504
rect -13631 -1577 -13627 -1504
rect -13717 -1591 -13627 -1577
rect -13369 -3000 -13289 6810
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -12380 4940 -12294 4954
rect -10771 4940 -10671 4950
rect -12616 4880 -12366 4940
rect -12306 4936 -10671 4940
rect -12306 4884 -10747 4936
rect -10695 4884 -10671 4936
rect -12306 4880 -10671 4884
rect -12380 4866 -12294 4880
rect -10771 4870 -10671 4880
rect -8339 4795 -8259 4805
rect -8339 4739 -8327 4795
rect -8271 4739 -8259 4795
rect -8339 4729 -8259 4739
rect -8063 4795 -7983 4805
rect -8063 4739 -8051 4795
rect -7995 4739 -7983 4795
rect -8063 4729 -7983 4739
rect -10201 4680 -10121 4690
rect -10211 4676 -10111 4680
rect -10211 4624 -10187 4676
rect -10135 4624 -8820 4676
rect -10211 4620 -8820 4624
rect -10201 4610 -10121 4620
rect -8876 4289 -8820 4620
rect -8327 4537 -8271 4729
rect -8202 4537 -8122 4549
rect -8327 4481 -8189 4537
rect -8133 4481 -8122 4537
rect -8327 4289 -8271 4481
rect -8202 4469 -8122 4481
rect -8201 4399 -8121 4409
rect -8051 4399 -7995 4729
rect -8201 4343 -8189 4399
rect -8133 4343 -7995 4399
rect -8201 4333 -8121 4343
rect -8876 4233 -8271 4289
rect -8327 3985 -8271 4233
rect -8051 4289 -7995 4343
rect -8051 4233 -7451 4289
rect -8051 3985 -7995 4233
rect -8339 3975 -8259 3985
rect -8339 3919 -8327 3975
rect -8271 3919 -8259 3975
rect -8339 3909 -8259 3919
rect -8063 3975 -7983 3985
rect -8063 3919 -8051 3975
rect -7995 3919 -7983 3975
rect -8063 3909 -7983 3919
rect -8431 3799 -8351 3809
rect -8431 3743 -8419 3799
rect -8363 3743 -8351 3799
rect -8431 3733 -8351 3743
rect -7971 3799 -7891 3809
rect -7971 3743 -7959 3799
rect -7903 3743 -7891 3799
rect -7971 3733 -7891 3743
rect -10531 3376 -10437 3388
rect -8419 3378 -8363 3733
rect -7959 3378 -7903 3733
rect -10531 3300 -10519 3376
rect -10439 3300 -10437 3376
rect -10531 3298 -10437 3300
rect -8421 3376 -8349 3378
rect -8421 3300 -8419 3376
rect -8363 3300 -8349 3376
rect -12103 2961 -11990 2978
rect -12103 2883 -12086 2961
rect -12006 2883 -11990 2961
rect -12103 2872 -11990 2883
rect -12086 2417 -12006 2872
rect -11650 2551 -11541 2564
rect -11650 2462 -11642 2551
rect -11551 2462 -11541 2551
rect -11650 2455 -11541 2462
rect -12096 2397 -11996 2417
rect -12096 2317 -12086 2397
rect -12006 2317 -11996 2397
rect -12096 2307 -11996 2317
rect -11642 1079 -11551 2455
rect -11391 2432 -11287 2446
rect -11391 2356 -11379 2432
rect -11299 2356 -11287 2432
rect -11391 2346 -11287 2356
rect -13382 -3004 -13286 -3000
rect -13784 -3082 -13368 -3004
rect -13290 -3082 -13286 -3004
rect -13382 -3096 -13286 -3082
rect -11640 -3421 -11553 1079
rect -11379 -2993 -11299 2346
rect -11051 2123 -10951 2133
rect -11051 2043 -11041 2123
rect -10961 2043 -10951 2123
rect -11051 2033 -10951 2043
rect -10729 2123 -10629 2133
rect -10729 2043 -10719 2123
rect -10639 2043 -10629 2123
rect -10729 2033 -10629 2043
rect -11041 1664 -10961 2033
rect -10845 1666 -10789 1674
rect -11041 1530 -11029 1664
rect -10973 1530 -10961 1664
rect -11041 1528 -10961 1530
rect -10857 1664 -10777 1666
rect -10857 1530 -10845 1664
rect -10789 1530 -10777 1664
rect -11029 1520 -10973 1528
rect -10857 5 -10777 1530
rect -10719 1664 -10639 2033
rect -10719 1530 -10707 1664
rect -10651 1530 -10639 1664
rect -10719 1528 -10639 1530
rect -10707 1520 -10651 1528
rect -10519 1173 -10439 3298
rect -8421 3288 -8349 3300
rect -7973 3376 -7901 3378
rect -7973 3300 -7959 3376
rect -7903 3300 -7901 3376
rect -7973 3288 -7901 3300
rect -5895 3376 -5791 3388
rect -5895 3300 -5883 3376
rect -5803 3300 -5791 3376
rect -5895 3298 -5791 3300
rect -10191 2123 -10091 2133
rect -10191 2043 -10181 2123
rect -10101 2043 -10091 2123
rect -10191 2033 -10091 2043
rect -9869 2123 -9769 2133
rect -9869 2043 -9859 2123
rect -9779 2043 -9769 2123
rect -9869 2033 -9769 2043
rect -9427 2123 -9327 2133
rect -9427 2043 -9417 2123
rect -9337 2043 -9327 2123
rect -9427 2033 -9327 2043
rect -8819 2123 -8719 2133
rect -8819 2043 -8809 2123
rect -8729 2043 -8719 2123
rect -8819 2033 -8719 2043
rect -8211 2123 -8111 2133
rect -8211 2043 -8201 2123
rect -8121 2043 -8111 2123
rect -8211 2033 -8111 2043
rect -7603 2123 -7503 2133
rect -7603 2043 -7593 2123
rect -7513 2043 -7503 2123
rect -7603 2033 -7503 2043
rect -6995 2123 -6895 2133
rect -6995 2043 -6985 2123
rect -6905 2043 -6895 2123
rect -6995 2033 -6895 2043
rect -6553 2123 -6453 2133
rect -6553 2043 -6543 2123
rect -6463 2043 -6453 2123
rect -6553 2033 -6453 2043
rect -6231 2123 -6131 2133
rect -6231 2043 -6221 2123
rect -6141 2043 -6131 2123
rect -6231 2033 -6131 2043
rect -10181 1664 -10101 2033
rect -9985 1666 -9929 1674
rect -10181 1530 -10169 1664
rect -10113 1530 -10101 1664
rect -10181 1528 -10101 1530
rect -9997 1664 -9917 1666
rect -9997 1530 -9985 1664
rect -9929 1530 -9917 1664
rect -10169 1520 -10113 1528
rect -10531 1161 -10427 1173
rect -9997 1171 -9917 1530
rect -9859 1664 -9779 2033
rect -9859 1530 -9847 1664
rect -9791 1530 -9779 1664
rect -9417 1677 -9337 2033
rect -9417 1533 -9405 1677
rect -9349 1533 -9337 1677
rect -8809 1677 -8729 2033
rect -9417 1531 -9337 1533
rect -9113 1576 -9033 1586
rect -9859 1528 -9779 1530
rect -9847 1520 -9791 1528
rect -9405 1523 -9349 1531
rect -9113 1520 -9101 1576
rect -9045 1520 -9033 1576
rect -8809 1533 -8797 1677
rect -8741 1533 -8729 1677
rect -8201 1677 -8121 2033
rect -8809 1531 -8729 1533
rect -8505 1576 -8425 1586
rect -8797 1523 -8741 1531
rect -9113 1510 -9033 1520
rect -8505 1520 -8493 1576
rect -8437 1520 -8425 1576
rect -8201 1533 -8189 1677
rect -8133 1533 -8121 1677
rect -7593 1677 -7513 2033
rect -8201 1531 -8121 1533
rect -7897 1576 -7817 1586
rect -8189 1523 -8133 1531
rect -10531 1077 -10519 1161
rect -10439 1077 -10427 1161
rect -10531 1067 -10427 1077
rect -10009 1161 -9905 1171
rect -8505 1169 -8425 1520
rect -7897 1520 -7885 1576
rect -7829 1520 -7817 1576
rect -7593 1533 -7581 1677
rect -7525 1533 -7513 1677
rect -6985 1677 -6905 2033
rect -7593 1531 -7513 1533
rect -7289 1576 -7209 1586
rect -7581 1523 -7525 1531
rect -8310 1469 -8230 1479
rect -8310 1413 -8298 1469
rect -8242 1413 -8230 1469
rect -8310 1339 -8230 1413
rect -8092 1469 -8012 1479
rect -8092 1413 -8080 1469
rect -8024 1413 -8012 1469
rect -8320 1329 -8220 1339
rect -8320 1249 -8310 1329
rect -8230 1249 -8220 1329
rect -8320 1239 -8220 1249
rect -8092 1169 -8012 1413
rect -7897 1339 -7817 1520
rect -7289 1520 -7277 1576
rect -7221 1520 -7209 1576
rect -6985 1533 -6973 1677
rect -6917 1533 -6905 1677
rect -6985 1531 -6905 1533
rect -6543 1664 -6463 2033
rect -6393 1666 -6337 1674
rect -6973 1523 -6917 1531
rect -6543 1530 -6531 1664
rect -6475 1530 -6463 1664
rect -6543 1528 -6463 1530
rect -6405 1664 -6325 1666
rect -6405 1530 -6393 1664
rect -6337 1530 -6325 1664
rect -6531 1520 -6475 1528
rect -7289 1510 -7209 1520
rect -7907 1329 -7807 1339
rect -7907 1249 -7897 1329
rect -7817 1249 -7807 1329
rect -7907 1239 -7807 1249
rect -7897 1169 -7817 1239
rect -6405 1171 -6325 1530
rect -6221 1664 -6141 2033
rect -6221 1530 -6209 1664
rect -6153 1530 -6141 1664
rect -6221 1528 -6141 1530
rect -6209 1520 -6153 1528
rect -5883 1171 -5803 3298
rect -5696 2887 -5576 2907
rect -5696 2787 -5676 2887
rect -5596 2787 -5576 2887
rect -5696 2767 -5576 2787
rect -4791 2649 -4633 2664
rect -4791 2542 -4764 2649
rect -4655 2542 -4633 2649
rect -4791 2531 -4633 2542
rect -5035 2432 -4931 2444
rect -5035 2356 -5023 2432
rect -4943 2356 -4931 2432
rect -5035 2344 -4931 2356
rect -5693 2123 -5593 2133
rect -5693 2043 -5683 2123
rect -5603 2043 -5593 2123
rect -5693 2033 -5593 2043
rect -5371 2123 -5271 2133
rect -5371 2043 -5361 2123
rect -5281 2043 -5271 2123
rect -5371 2033 -5271 2043
rect -5683 1664 -5603 2033
rect -5533 1666 -5477 1674
rect -5683 1530 -5671 1664
rect -5615 1530 -5603 1664
rect -5683 1528 -5603 1530
rect -5545 1664 -5465 1666
rect -5545 1530 -5533 1664
rect -5477 1530 -5465 1664
rect -5671 1520 -5615 1528
rect -10009 1077 -9997 1161
rect -9917 1077 -9905 1161
rect -10009 1067 -9905 1077
rect -9263 1159 -9159 1169
rect -9263 1079 -9251 1159
rect -9171 1079 -9159 1159
rect -9263 1065 -9159 1079
rect -8655 1159 -8415 1169
rect -8102 1159 -8002 1169
rect -8655 1079 -8643 1159
rect -8563 1079 -8505 1159
rect -8425 1079 -8092 1159
rect -8012 1079 -8002 1159
rect -8655 1065 -8415 1079
rect -8102 1069 -8002 1079
rect -7909 1159 -7667 1169
rect -7909 1079 -7897 1159
rect -7817 1079 -7759 1159
rect -7679 1079 -7667 1159
rect -7909 1065 -7667 1079
rect -7163 1159 -7059 1170
rect -7163 1079 -7151 1159
rect -7071 1079 -7059 1159
rect -7163 1066 -7059 1079
rect -6417 1161 -6313 1171
rect -6417 1077 -6405 1161
rect -6325 1077 -6313 1161
rect -6417 1067 -6313 1077
rect -5895 1161 -5791 1171
rect -5895 1077 -5883 1161
rect -5803 1077 -5791 1161
rect -5895 1067 -5791 1077
rect -9251 721 -9171 1065
rect -8852 865 -8752 875
rect -8852 785 -8842 865
rect -8762 785 -8752 865
rect -8852 775 -8752 785
rect -9251 577 -9239 721
rect -9183 577 -9171 721
rect -9251 575 -9171 577
rect -8643 721 -8563 1065
rect -8643 577 -8631 721
rect -8575 577 -8563 721
rect -8643 575 -8563 577
rect -7759 721 -7679 1065
rect -7570 865 -7470 875
rect -7570 785 -7560 865
rect -7480 785 -7470 865
rect -7570 775 -7470 785
rect -7759 577 -7747 721
rect -7691 577 -7679 721
rect -7759 575 -7679 577
rect -7151 721 -7071 1066
rect -7151 577 -7139 721
rect -7083 577 -7071 721
rect -7151 575 -7071 577
rect -9239 567 -9183 575
rect -8631 567 -8575 575
rect -7747 567 -7691 575
rect -7139 567 -7083 575
rect -9543 507 -9487 515
rect -8935 507 -8879 515
rect -7443 507 -7387 515
rect -6835 507 -6779 515
rect -9555 505 -9475 507
rect -9997 415 -9917 425
rect -10306 271 -9985 415
rect -9929 271 -9917 415
rect -10869 -5 -10765 5
rect -10869 -85 -10857 -5
rect -10777 -85 -10765 -5
rect -10869 -95 -10765 -85
rect -10306 -265 -10202 271
rect -9997 260 -9917 271
rect -9555 361 -9543 505
rect -9487 361 -9475 505
rect -9555 7 -9475 361
rect -8947 505 -8867 507
rect -8947 361 -8935 505
rect -8879 361 -8867 505
rect -8947 7 -8867 361
rect -7455 505 -7375 507
rect -7455 361 -7443 505
rect -7387 361 -7375 505
rect -7455 7 -7375 361
rect -6847 505 -6767 507
rect -6847 361 -6835 505
rect -6779 361 -6767 505
rect -6847 7 -6767 361
rect -6405 415 -6325 425
rect -6405 271 -6393 415
rect -6337 271 -6016 415
rect -6405 260 -6325 271
rect -9733 -5 -9629 7
rect -9733 -85 -9721 -5
rect -9641 -85 -9629 -5
rect -9733 -97 -9629 -85
rect -9567 -5 -9463 7
rect -9567 -85 -9555 -5
rect -9475 -85 -9463 -5
rect -9567 -97 -9463 -85
rect -8959 -5 -8855 7
rect -8959 -85 -8947 -5
rect -8867 -85 -8855 -5
rect -8959 -97 -8855 -85
rect -7467 -5 -7363 7
rect -7467 -85 -7455 -5
rect -7375 -85 -7363 -5
rect -7467 -97 -7363 -85
rect -6859 -5 -6755 7
rect -6859 -85 -6847 -5
rect -6767 -85 -6755 -5
rect -6859 -97 -6755 -85
rect -6693 -5 -6589 7
rect -6693 -85 -6681 -5
rect -6601 -85 -6589 -5
rect -6693 -97 -6589 -85
rect -10647 -369 -10202 -265
rect -11391 -3003 -11287 -2993
rect -11391 -3083 -11379 -3003
rect -11299 -3083 -11287 -3003
rect -11391 -3093 -11287 -3083
rect -10639 -3123 -10550 -369
rect -10306 -403 -10202 -369
rect -10306 -564 -10304 -403
rect -10204 -564 -10202 -403
rect -10306 -576 -10202 -564
rect -9721 -813 -9641 -97
rect -6681 -575 -6601 -97
rect -9721 -974 -9709 -813
rect -9653 -974 -9641 -813
rect -9113 -631 -6601 -575
rect -6120 -256 -6016 271
rect -5545 5 -5465 1530
rect -5361 1664 -5281 2033
rect -5361 1530 -5349 1664
rect -5293 1530 -5281 1664
rect -5361 1528 -5281 1530
rect -5349 1520 -5293 1528
rect -5557 -5 -5453 5
rect -5557 -85 -5545 -5
rect -5465 -85 -5453 -5
rect -5557 -95 -5453 -85
rect -6120 -360 -5550 -256
rect -6120 -403 -6016 -360
rect -6120 -564 -6118 -403
rect -6018 -564 -6016 -403
rect -6120 -576 -6016 -564
rect -9113 -777 -9033 -631
rect -9721 -984 -9641 -974
rect -9417 -861 -9337 -851
rect -9417 -1022 -9405 -861
rect -9349 -1022 -9337 -861
rect -9113 -994 -9101 -777
rect -9045 -994 -9033 -777
rect -8505 -777 -8425 -767
rect -8505 -833 -8493 -777
rect -8437 -833 -8425 -777
rect -8505 -843 -8425 -833
rect -7897 -777 -7817 -631
rect -7897 -833 -7885 -777
rect -7829 -833 -7817 -777
rect -7897 -843 -7817 -833
rect -7289 -777 -7209 -767
rect -9113 -1002 -9033 -994
rect -8809 -861 -8729 -851
rect -9417 -1352 -9337 -1022
rect -8809 -1022 -8797 -861
rect -8741 -1022 -8729 -861
rect -9276 -1068 -8871 -1058
rect -9276 -1128 -9261 -1068
rect -9191 -1128 -8956 -1068
rect -8886 -1128 -8871 -1068
rect -9276 -1138 -8871 -1128
rect -9266 -1226 -9186 -1216
rect -9266 -1282 -9254 -1226
rect -9198 -1282 -9186 -1226
rect -9266 -1292 -9186 -1282
rect -8809 -1352 -8729 -1022
rect -8201 -861 -8121 -851
rect -8201 -1022 -8189 -861
rect -8133 -1022 -8121 -861
rect -8201 -1352 -8121 -1022
rect -7593 -861 -7513 -851
rect -7593 -1022 -7581 -861
rect -7525 -1022 -7513 -861
rect -8061 -1068 -7656 -1058
rect -8061 -1128 -8046 -1068
rect -7976 -1128 -7741 -1068
rect -7671 -1128 -7656 -1068
rect -8061 -1138 -7656 -1128
rect -8051 -1226 -7971 -1216
rect -8051 -1282 -8039 -1226
rect -7983 -1282 -7971 -1226
rect -8051 -1292 -7971 -1282
rect -7593 -1352 -7513 -1022
rect -7289 -1022 -7277 -777
rect -7221 -1022 -7209 -777
rect -6681 -813 -6601 -631
rect -7289 -1032 -7209 -1022
rect -6985 -861 -6905 -851
rect -6985 -1022 -6973 -861
rect -6917 -1022 -6905 -861
rect -6681 -974 -6669 -813
rect -6613 -974 -6601 -813
rect -6681 -984 -6601 -974
rect -6985 -1352 -6905 -1022
rect -6841 -1068 -6741 -1058
rect -6547 -1068 -6321 -1067
rect -6841 -1128 -6826 -1068
rect -6756 -1127 -6321 -1068
rect -6756 -1128 -6582 -1127
rect -6841 -1138 -6741 -1128
rect -6526 -1193 -6441 -1183
rect -6526 -1253 -6511 -1193
rect -6451 -1253 -6441 -1193
rect -6526 -1268 -6441 -1253
rect -9417 -1408 -6905 -1352
rect -9417 -1732 -9337 -1408
rect -8961 -1474 -8881 -1464
rect -8961 -1530 -8949 -1474
rect -8893 -1530 -8881 -1474
rect -8961 -1540 -8881 -1530
rect -9276 -1628 -8871 -1618
rect -9276 -1688 -9261 -1628
rect -9191 -1688 -8956 -1628
rect -8886 -1688 -8871 -1628
rect -9276 -1698 -8871 -1688
rect -9417 -1893 -9405 -1732
rect -9349 -1893 -9337 -1732
rect -8809 -1732 -8729 -1408
rect -9721 -1921 -9641 -1911
rect -9721 -1977 -9709 -1921
rect -9653 -1977 -9641 -1921
rect -9721 -1987 -9641 -1977
rect -10306 -2187 -10202 -2175
rect -10306 -2348 -10304 -2187
rect -10204 -2348 -10202 -2187
rect -9417 -2239 -9337 -1893
rect -9113 -1766 -9033 -1756
rect -9113 -1977 -9101 -1766
rect -9045 -1977 -9033 -1766
rect -8809 -1893 -8797 -1732
rect -8741 -1893 -8729 -1732
rect -8809 -1903 -8729 -1893
rect -8505 -1732 -8425 -1722
rect -9113 -2123 -9033 -1977
rect -8505 -1977 -8493 -1732
rect -8437 -1977 -8425 -1732
rect -8201 -1732 -8121 -1408
rect -7746 -1474 -7666 -1464
rect -7746 -1530 -7734 -1474
rect -7678 -1530 -7666 -1474
rect -7746 -1540 -7666 -1530
rect -8061 -1628 -7656 -1618
rect -8061 -1688 -8046 -1628
rect -7976 -1688 -7741 -1628
rect -7671 -1688 -7656 -1628
rect -8061 -1698 -7656 -1688
rect -8201 -1893 -8189 -1732
rect -8133 -1893 -8121 -1732
rect -7593 -1732 -7513 -1408
rect -8201 -1903 -8121 -1893
rect -7897 -1766 -7817 -1756
rect -8505 -1987 -8425 -1977
rect -7897 -1977 -7885 -1766
rect -7829 -1977 -7817 -1766
rect -7593 -1893 -7581 -1732
rect -7525 -1893 -7513 -1732
rect -7593 -1903 -7513 -1893
rect -7289 -1732 -7209 -1722
rect -7897 -2123 -7817 -1977
rect -7289 -1977 -7277 -1732
rect -7221 -1977 -7209 -1732
rect -7289 -1987 -7209 -1977
rect -6985 -1732 -6905 -1408
rect -6511 -1408 -6451 -1268
rect -6381 -1288 -6321 -1127
rect -6381 -1348 -6191 -1288
rect -6511 -1468 -6321 -1408
rect -6841 -1628 -6741 -1618
rect -6381 -1628 -6321 -1468
rect -6251 -1493 -6191 -1348
rect -6261 -1503 -6181 -1493
rect -6261 -1563 -6251 -1503
rect -6191 -1563 -6181 -1503
rect -6261 -1573 -6181 -1563
rect -6841 -1688 -6826 -1628
rect -6756 -1688 -6321 -1628
rect -6841 -1698 -6741 -1688
rect -6985 -1977 -6973 -1732
rect -6917 -1977 -6905 -1732
rect -6985 -1987 -6905 -1977
rect -6681 -1920 -6601 -1910
rect -6681 -1977 -6669 -1920
rect -6613 -1977 -6601 -1920
rect -6681 -2123 -6601 -1977
rect -9113 -2179 -6601 -2123
rect -6143 -2160 -6002 -2144
rect -9417 -2250 -6895 -2239
rect -9417 -2306 -6985 -2250
rect -6905 -2306 -6895 -2250
rect -6143 -2297 -6129 -2160
rect -9417 -2316 -6895 -2306
rect -10306 -2650 -10202 -2348
rect -10306 -2652 -8213 -2650
rect -10306 -2774 -8603 -2652
rect -8547 -2774 -8281 -2652
rect -8225 -2774 -8213 -2652
rect -10306 -2776 -8213 -2774
rect -8109 -2652 -8029 -2316
rect -6144 -2370 -6129 -2297
rect -6024 -2308 -6002 -2160
rect -6024 -2370 -6007 -2308
rect -6144 -2388 -6007 -2370
rect -8109 -2774 -8097 -2652
rect -8041 -2774 -8029 -2652
rect -8109 -2776 -8029 -2774
rect -10665 -3376 -10513 -3123
rect -10078 -3372 -9728 -2776
rect -6126 -3311 -6027 -2388
rect -6126 -3356 -6009 -3311
rect -6136 -3367 -6009 -3356
rect -11664 -3443 -11529 -3421
rect -11664 -3530 -11640 -3443
rect -11555 -3530 -11529 -3443
rect -10665 -3463 -10639 -3376
rect -10550 -3463 -10513 -3376
rect -10665 -3496 -10513 -3463
rect -10097 -3381 -9707 -3372
rect -11664 -3545 -11529 -3530
rect -10097 -3592 -10083 -3381
rect -9728 -3592 -9707 -3381
rect -10097 -3613 -9707 -3592
rect -6136 -3375 -6010 -3367
rect -6136 -3578 -6132 -3375
rect -6018 -3578 -6010 -3375
rect -5654 -3419 -5550 -360
rect -5023 -2993 -4943 2344
rect -5035 -3003 -4931 -2993
rect -5035 -3083 -5023 -3003
rect -4943 -3083 -4931 -3003
rect -5035 -3093 -4931 -3083
rect -5665 -3429 -5537 -3419
rect -5665 -3531 -5654 -3429
rect -5550 -3531 -5537 -3429
rect -4764 -3439 -4655 2531
rect -4464 -3363 -2407 -3321
rect -5665 -3565 -5537 -3531
rect -4774 -3451 -4646 -3439
rect -4774 -3558 -4764 -3451
rect -4655 -3558 -4646 -3451
rect -6136 -3597 -6010 -3578
rect -4774 -3580 -4646 -3558
rect -4464 -3663 -4454 -3363
rect -2454 -3663 -2407 -3363
rect -4464 -3701 -2407 -3663
<< via2 >>
rect 40739 39093 40957 39167
rect 40737 37749 40955 37823
rect -4343 37511 -4287 37567
rect 5129 37511 5185 37567
rect 14601 37512 14657 37568
rect 24073 37512 24129 37568
rect 33545 37512 33601 37568
rect 43017 37512 43073 37568
rect -5507 36542 -5451 36598
rect -8093 33316 -8037 33372
rect -5707 33319 -5651 33375
rect -10199 30949 -10143 31005
rect -9169 30511 -9113 30567
rect -6327 31169 -6027 31969
rect -8761 30511 -8705 30567
rect -9985 30090 -9905 30166
rect -8755 30059 -8155 30199
rect -7695 30833 -5927 30973
rect -8755 29659 -8155 29799
rect -11830 27521 -11774 27577
rect -11592 27488 -11536 27608
rect -9169 28171 -9113 28227
rect 3965 36542 4021 36598
rect -4844 35641 -4788 35697
rect -4026 35641 -3970 35697
rect -4343 35306 -4287 35362
rect -2857 35306 -2801 35362
rect -4844 33436 -4788 33492
rect -4026 33436 -3970 33492
rect -3358 33436 -3302 33492
rect -2540 33436 -2484 33492
rect -4343 33101 -4287 33157
rect -2857 33102 -2801 33158
rect -4844 31231 -4788 31287
rect -4026 31231 -3970 31287
rect -3358 31232 -3302 31288
rect -2540 31232 -2484 31288
rect -4343 30896 -4287 30952
rect -7695 28873 -5927 29013
rect 3765 33319 3821 33375
rect -1245 31169 -1045 31969
rect 303 30511 359 30567
rect 3145 31169 3445 31969
rect 711 30511 767 30567
rect 717 30059 1317 30199
rect 1777 30833 3545 30973
rect -4844 29026 -4788 29082
rect -4026 29026 -3970 29082
rect -5610 28908 -5554 28964
rect -8761 28171 -8705 28227
rect -6327 27889 -6027 28689
rect 717 29659 1317 29799
rect -2064 27489 -2008 27609
rect 303 28171 359 28227
rect 13437 36543 13493 36599
rect 4628 35641 4684 35697
rect 5446 35641 5502 35697
rect 5129 35306 5185 35362
rect 6615 35306 6671 35362
rect 4628 33436 4684 33492
rect 5446 33436 5502 33492
rect 6114 33436 6170 33492
rect 6932 33436 6988 33492
rect 5129 33101 5185 33157
rect 6615 33102 6671 33158
rect 4628 31231 4684 31287
rect 5446 31231 5502 31287
rect 6114 31232 6170 31288
rect 6932 31232 6988 31288
rect 5129 30896 5185 30952
rect 1777 28873 3545 29013
rect 13237 33320 13293 33376
rect 8227 31170 8427 31970
rect 9775 30512 9831 30568
rect 12617 31170 12917 31970
rect 10183 30512 10239 30568
rect 10189 30060 10789 30200
rect 11249 30834 13017 30974
rect 4628 29026 4684 29082
rect 5446 29026 5502 29082
rect 3862 28908 3918 28964
rect 711 28171 767 28227
rect 3145 27889 3445 28689
rect 10189 29660 10789 29800
rect 7408 27489 7464 27609
rect 9775 28172 9831 28228
rect 22909 36543 22965 36599
rect 14100 35642 14156 35698
rect 14918 35642 14974 35698
rect 14601 35307 14657 35363
rect 16087 35307 16143 35363
rect 14100 33437 14156 33493
rect 14918 33437 14974 33493
rect 15586 33437 15642 33493
rect 16404 33437 16460 33493
rect 14601 33102 14657 33158
rect 16087 33103 16143 33159
rect 14100 31232 14156 31288
rect 14918 31232 14974 31288
rect 15586 31233 15642 31289
rect 16404 31233 16460 31289
rect 14601 30897 14657 30953
rect 11249 28874 13017 29014
rect 22709 33320 22765 33376
rect 17699 31170 17899 31970
rect 19247 30512 19303 30568
rect 22089 31170 22389 31970
rect 19655 30512 19711 30568
rect 19661 30060 20261 30200
rect 20721 30834 22489 30974
rect 14100 29027 14156 29083
rect 14918 29027 14974 29083
rect 13334 28909 13390 28965
rect 10183 28172 10239 28228
rect 12617 27890 12917 28690
rect 19661 29660 20261 29800
rect 16880 27490 16936 27610
rect -12833 16399 -12777 16499
rect -9501 16399 -9445 16499
rect -12833 15889 -12777 15989
rect -11613 15630 -11557 15686
rect -12114 13760 -12058 13816
rect -11296 13760 -11240 13816
rect -11613 13425 -11557 13481
rect -10127 13425 -10071 13481
rect -12114 11555 -12058 11611
rect -11296 11555 -11240 11611
rect -10628 11555 -10572 11611
rect -9810 11555 -9754 11611
rect -11613 11220 -11557 11276
rect -10127 11221 -10071 11277
rect -12114 9350 -12058 9406
rect -11296 9350 -11240 9406
rect -7601 25209 -7545 25265
rect -8102 23339 -8046 23395
rect -7284 23339 -7228 23395
rect -7601 23004 -7545 23060
rect -6115 23004 -6059 23060
rect -8102 21134 -8046 21190
rect -7284 21134 -7228 21190
rect -6616 21134 -6560 21190
rect -5798 21134 -5742 21190
rect -7601 20799 -7545 20855
rect -6115 20800 -6059 20856
rect -8102 18929 -8046 18985
rect -7284 18929 -7228 18985
rect -6616 18930 -6560 18986
rect -5798 18930 -5742 18986
rect -7601 18594 -7545 18650
rect -8102 16724 -8046 16780
rect -7284 16724 -7228 16780
rect -5489 16399 -5433 16499
rect -8957 15892 -8901 15992
rect -10628 9351 -10572 9407
rect -9810 9351 -9754 9407
rect -11613 9015 -11557 9071
rect -12896 7814 -12840 7870
rect -12114 7145 -12058 7201
rect -11296 7145 -11240 7201
rect -12896 7027 -12840 7083
rect -13105 6820 -13049 6920
rect -7601 15630 -7545 15686
rect -8765 14661 -8709 14717
rect -8102 13760 -8046 13816
rect -7284 13760 -7228 13816
rect -7601 13425 -7545 13481
rect -6115 13425 -6059 13481
rect -8102 11555 -8046 11611
rect -7284 11555 -7228 11611
rect -6616 11555 -6560 11611
rect -5798 11555 -5742 11611
rect -7601 11220 -7545 11276
rect -6115 11221 -6059 11277
rect -8102 9350 -8046 9406
rect -7284 9350 -7228 9406
rect -3559 25206 -3503 25262
rect -4060 23336 -4004 23392
rect -3242 23336 -3186 23392
rect -3559 23001 -3503 23057
rect -2073 23001 -2017 23057
rect -4060 21131 -4004 21187
rect -3242 21131 -3186 21187
rect -2574 21131 -2518 21187
rect -1756 21131 -1700 21187
rect -3559 20796 -3503 20852
rect -2073 20797 -2017 20853
rect -4060 18926 -4004 18982
rect -3242 18926 -3186 18982
rect -2574 18927 -2518 18983
rect -1756 18927 -1700 18983
rect -3559 18591 -3503 18647
rect -4060 16721 -4004 16777
rect -3242 16721 -3186 16777
rect -1447 16399 -1391 16499
rect -4945 15889 -4889 15989
rect -6616 9351 -6560 9407
rect -5798 9351 -5742 9407
rect -7601 9015 -7545 9071
rect -8102 7145 -8046 7201
rect -7284 7145 -7228 7201
rect -9093 6820 -9037 6920
rect -3559 15630 -3503 15686
rect -4723 14661 -4667 14717
rect -4060 13760 -4004 13816
rect -3242 13760 -3186 13816
rect -3559 13425 -3503 13481
rect -2073 13425 -2017 13481
rect -4060 11555 -4004 11611
rect -3242 11555 -3186 11611
rect -2574 11555 -2518 11611
rect -1756 11555 -1700 11611
rect -3559 11220 -3503 11276
rect -2073 11221 -2017 11277
rect -4060 9350 -4004 9406
rect -3242 9350 -3186 9406
rect 19247 28172 19303 28228
rect 32381 36543 32437 36599
rect 23572 35642 23628 35698
rect 24390 35642 24446 35698
rect 24073 35307 24129 35363
rect 25559 35307 25615 35363
rect 23572 33437 23628 33493
rect 24390 33437 24446 33493
rect 25058 33437 25114 33493
rect 25876 33437 25932 33493
rect 24073 33102 24129 33158
rect 25559 33103 25615 33159
rect 23572 31232 23628 31288
rect 24390 31232 24446 31288
rect 25058 31233 25114 31289
rect 25876 31233 25932 31289
rect 24073 30897 24129 30953
rect 20721 28874 22489 29014
rect 32181 33320 32237 33376
rect 27171 31170 27371 31970
rect 28719 30512 28775 30568
rect 31561 31170 31861 31970
rect 29127 30512 29183 30568
rect 29133 30060 29733 30200
rect 30193 30834 31961 30974
rect 23572 29027 23628 29083
rect 24390 29027 24446 29083
rect 22806 28909 22862 28965
rect 19655 28172 19711 28228
rect 22089 27890 22389 28690
rect 29133 29660 29733 29800
rect 26352 27490 26408 27610
rect 28719 28172 28775 28228
rect 41853 36543 41909 36599
rect 33044 35642 33100 35698
rect 33862 35642 33918 35698
rect 33545 35307 33601 35363
rect 35031 35307 35087 35363
rect 33044 33437 33100 33493
rect 33862 33437 33918 33493
rect 34530 33437 34586 33493
rect 35348 33437 35404 33493
rect 33545 33102 33601 33158
rect 35031 33103 35087 33159
rect 33044 31232 33100 31288
rect 33862 31232 33918 31288
rect 34530 31233 34586 31289
rect 35348 31233 35404 31289
rect 33545 30897 33601 30953
rect 30193 28874 31961 29014
rect 41653 33320 41709 33376
rect 36643 31170 36843 31970
rect 38191 30512 38247 30568
rect 41033 31170 41333 31970
rect 38599 30512 38655 30568
rect 38605 30060 39205 30200
rect 39665 30834 41433 30974
rect 33044 29027 33100 29083
rect 33862 29027 33918 29083
rect 32278 28909 32334 28965
rect 29127 28172 29183 28228
rect 31561 27890 31861 28690
rect 38605 29660 39205 29800
rect 35824 27490 35880 27610
rect 483 25206 539 25262
rect -18 23336 38 23392
rect 800 23336 856 23392
rect 483 23001 539 23057
rect 1969 23001 2025 23057
rect -18 21131 38 21187
rect 800 21131 856 21187
rect 1468 21131 1524 21187
rect 2286 21131 2342 21187
rect 483 20796 539 20852
rect 1969 20797 2025 20853
rect -18 18926 38 18982
rect 800 18926 856 18982
rect 1468 18927 1524 18983
rect 2286 18927 2342 18983
rect 483 18591 539 18647
rect -18 16721 38 16777
rect 800 16721 856 16777
rect 2595 16399 2651 16499
rect -903 15889 -847 15989
rect -2574 9351 -2518 9407
rect -1756 9351 -1700 9407
rect -3559 9015 -3503 9071
rect -4060 7145 -4004 7201
rect -3242 7145 -3186 7201
rect -5081 6820 -5025 6920
rect 483 15630 539 15686
rect -681 14661 -625 14717
rect -18 13760 38 13816
rect 800 13760 856 13816
rect 483 13425 539 13481
rect 1969 13425 2025 13481
rect -18 11555 38 11611
rect 800 11555 856 11611
rect 1468 11555 1524 11611
rect 2286 11555 2342 11611
rect 483 11220 539 11276
rect 1969 11221 2025 11277
rect -18 9350 38 9406
rect 800 9350 856 9406
rect 4525 25206 4581 25262
rect 4024 23336 4080 23392
rect 4842 23336 4898 23392
rect 4525 23001 4581 23057
rect 6011 23001 6067 23057
rect 4024 21131 4080 21187
rect 4842 21131 4898 21187
rect 5510 21131 5566 21187
rect 6328 21131 6384 21187
rect 4525 20796 4581 20852
rect 6011 20797 6067 20853
rect 4024 18926 4080 18982
rect 4842 18926 4898 18982
rect 5510 18927 5566 18983
rect 6328 18927 6384 18983
rect 4525 18591 4581 18647
rect 4024 16721 4080 16777
rect 4842 16721 4898 16777
rect 6637 16399 6693 16499
rect 3139 15889 3195 15989
rect 1468 9351 1524 9407
rect 2286 9351 2342 9407
rect 483 9015 539 9071
rect -18 7145 38 7201
rect 800 7145 856 7201
rect -1039 6820 -983 6920
rect 4525 15630 4581 15686
rect 3361 14661 3417 14717
rect 4024 13760 4080 13816
rect 4842 13760 4898 13816
rect 4525 13425 4581 13481
rect 6011 13425 6067 13481
rect 4024 11555 4080 11611
rect 4842 11555 4898 11611
rect 5510 11555 5566 11611
rect 6328 11555 6384 11611
rect 4525 11220 4581 11276
rect 6011 11221 6067 11277
rect 4024 9350 4080 9406
rect 4842 9350 4898 9406
rect 38191 28172 38247 28228
rect 42516 35642 42572 35698
rect 43334 35642 43390 35698
rect 43017 35307 43073 35363
rect 44503 35307 44559 35363
rect 42516 33437 42572 33493
rect 43334 33437 43390 33493
rect 44002 33437 44058 33493
rect 44820 33437 44876 33493
rect 43017 33102 43073 33158
rect 44503 33103 44559 33159
rect 42516 31232 42572 31288
rect 43334 31232 43390 31288
rect 44002 31233 44058 31289
rect 44820 31233 44876 31289
rect 43017 30897 43073 30953
rect 39665 28874 41433 29014
rect 42516 29027 42572 29083
rect 43334 29027 43390 29083
rect 41750 28909 41806 28965
rect 38599 28172 38655 28228
rect 41033 27890 41333 28690
rect 8567 25206 8623 25262
rect 8066 23336 8122 23392
rect 8884 23336 8940 23392
rect 8567 23001 8623 23057
rect 10053 23001 10109 23057
rect 8066 21131 8122 21187
rect 8884 21131 8940 21187
rect 9552 21131 9608 21187
rect 10370 21131 10426 21187
rect 8567 20796 8623 20852
rect 10053 20797 10109 20853
rect 8066 18926 8122 18982
rect 8884 18926 8940 18982
rect 9552 18927 9608 18983
rect 10370 18927 10426 18983
rect 8567 18591 8623 18647
rect 8066 16721 8122 16777
rect 8884 16721 8940 16777
rect 10679 16399 10735 16499
rect 7181 15889 7237 15989
rect 5510 9351 5566 9407
rect 6328 9351 6384 9407
rect 4525 9015 4581 9071
rect 4024 7145 4080 7201
rect 4842 7145 4898 7201
rect 3003 6820 3059 6920
rect 8567 15630 8623 15686
rect 7403 14661 7459 14717
rect 8066 13760 8122 13816
rect 8884 13760 8940 13816
rect 8567 13425 8623 13481
rect 10053 13425 10109 13481
rect 8066 11555 8122 11611
rect 8884 11555 8940 11611
rect 9552 11555 9608 11611
rect 10370 11555 10426 11611
rect 8567 11220 8623 11276
rect 10053 11221 10109 11277
rect 8066 9350 8122 9406
rect 8884 9350 8940 9406
rect 12609 25206 12665 25262
rect 12108 23336 12164 23392
rect 12926 23336 12982 23392
rect 12609 23001 12665 23057
rect 14095 23001 14151 23057
rect 12108 21131 12164 21187
rect 12926 21131 12982 21187
rect 13594 21131 13650 21187
rect 14412 21131 14468 21187
rect 12609 20796 12665 20852
rect 14095 20797 14151 20853
rect 12108 18926 12164 18982
rect 12926 18926 12982 18982
rect 13594 18927 13650 18983
rect 14412 18927 14468 18983
rect 12609 18591 12665 18647
rect 12108 16721 12164 16777
rect 12926 16721 12982 16777
rect 11223 15889 11279 15989
rect 9552 9351 9608 9407
rect 10370 9351 10426 9407
rect 8567 9015 8623 9071
rect 8066 7145 8122 7201
rect 8884 7145 8940 7201
rect 7045 6820 7101 6920
rect 12609 15630 12665 15686
rect 11445 14661 11501 14717
rect 12108 13760 12164 13816
rect 12926 13760 12982 13816
rect 12609 13425 12665 13481
rect 14095 13425 14151 13481
rect 12108 11555 12164 11611
rect 12926 11555 12982 11611
rect 13594 11555 13650 11611
rect 14412 11555 14468 11611
rect 12609 11220 12665 11276
rect 14095 11221 14151 11277
rect 12108 9350 12164 9406
rect 12926 9350 12982 9406
rect 16651 25206 16707 25262
rect 15386 21014 15442 21070
rect 16150 23336 16206 23392
rect 16968 23336 17024 23392
rect 16651 23001 16707 23057
rect 18137 23001 18193 23057
rect 16150 21131 16206 21187
rect 16968 21131 17024 21187
rect 17636 21131 17692 21187
rect 18454 21131 18510 21187
rect 16651 20796 16707 20852
rect 18137 20797 18193 20853
rect 16150 18926 16206 18982
rect 16968 18926 17024 18982
rect 17636 18927 17692 18983
rect 18454 18927 18510 18983
rect 16651 18591 16707 18647
rect 15386 17390 15442 17446
rect 16150 16721 16206 16777
rect 16968 16721 17024 16777
rect 15265 15889 15321 15989
rect 13594 9351 13650 9407
rect 14412 9351 14468 9407
rect 12609 9015 12665 9071
rect 12108 7145 12164 7201
rect 12926 7145 12982 7201
rect 11087 6820 11143 6920
rect -4454 6134 -2454 6434
rect -12086 2317 -12006 2397
rect -11041 2043 -10961 2123
rect -10719 2043 -10639 2123
rect -10181 2043 -10101 2123
rect -9859 2043 -9779 2123
rect -9417 2043 -9337 2123
rect -8809 2043 -8729 2123
rect -8201 2043 -8121 2123
rect -7593 2043 -7513 2123
rect -6985 2043 -6905 2123
rect -6543 2043 -6463 2123
rect -6221 2043 -6141 2123
rect -9101 1520 -9045 1576
rect -8493 1520 -8437 1576
rect -8310 1249 -8230 1329
rect -7277 1520 -7221 1576
rect -7897 1249 -7817 1329
rect -5676 2847 -5596 2887
rect -5676 2807 -5596 2847
rect -5683 2043 -5603 2123
rect -5361 2043 -5281 2123
rect -8092 1079 -8012 1159
rect -8842 785 -8762 865
rect -7560 785 -7480 865
rect -9709 -974 -9653 -813
rect -9101 -994 -9045 -938
rect -8493 -833 -8437 -777
rect -8949 -1126 -8893 -1070
rect -9254 -1282 -9198 -1226
rect -7734 -1126 -7678 -1070
rect -8039 -1282 -7983 -1226
rect -7277 -1022 -7221 -777
rect -6669 -974 -6613 -813
rect -8949 -1530 -8893 -1474
rect -9254 -1686 -9198 -1630
rect -9709 -1977 -9653 -1921
rect -9101 -1822 -9045 -1766
rect -8493 -1977 -8437 -1732
rect -7734 -1530 -7678 -1474
rect -8039 -1686 -7983 -1630
rect -7885 -1822 -7829 -1766
rect -7277 -1977 -7221 -1732
rect -6973 -1977 -6917 -1732
rect -6985 -2306 -6905 -2250
rect -4454 -3663 -2454 -3363
<< metal3 >>
rect 40726 39167 40972 39180
rect 40726 39093 40739 39167
rect 40957 39093 40972 39167
rect 40726 39080 40972 39093
rect 40723 37823 40967 37836
rect 40723 37749 40737 37823
rect 40955 37749 40967 37823
rect 40723 37737 40967 37749
rect -4355 37567 -4269 37571
rect -4355 37511 -4343 37567
rect -4287 37511 -4269 37567
rect -4355 37499 -4269 37511
rect 5117 37567 5203 37571
rect 5117 37511 5129 37567
rect 5185 37511 5203 37567
rect 5117 37499 5203 37511
rect 14589 37568 14675 37572
rect 14589 37512 14601 37568
rect 14657 37512 14675 37568
rect 14589 37500 14675 37512
rect 24061 37568 24147 37572
rect 24061 37512 24073 37568
rect 24129 37512 24147 37568
rect 24061 37500 24147 37512
rect 33533 37568 33619 37572
rect 33533 37512 33545 37568
rect 33601 37512 33619 37568
rect 33533 37500 33619 37512
rect 43005 37568 43091 37572
rect 43005 37512 43017 37568
rect 43073 37512 43091 37568
rect 43005 37500 43091 37512
rect -5521 36598 -5433 36610
rect -5521 36542 -5507 36598
rect -5451 36542 -5433 36598
rect -5521 36530 -5433 36542
rect 3951 36598 4039 36610
rect 3951 36542 3965 36598
rect 4021 36542 4039 36598
rect 3951 36530 4039 36542
rect 13423 36599 13511 36611
rect 13423 36543 13437 36599
rect 13493 36543 13511 36599
rect 13423 36531 13511 36543
rect 22895 36599 22983 36611
rect 22895 36543 22909 36599
rect 22965 36543 22983 36599
rect 22895 36531 22983 36543
rect 32367 36599 32455 36611
rect 32367 36543 32381 36599
rect 32437 36543 32455 36599
rect 32367 36531 32455 36543
rect 41839 36599 41927 36611
rect 41839 36543 41853 36599
rect 41909 36543 41927 36599
rect 41839 36531 41927 36543
rect -4856 35697 -4776 35709
rect -4856 35641 -4844 35697
rect -4788 35641 -4776 35697
rect -4856 35629 -4776 35641
rect -4038 35697 -3958 35709
rect -4038 35641 -4026 35697
rect -3970 35641 -3958 35697
rect -4038 35629 -3958 35641
rect 4616 35697 4696 35709
rect 4616 35641 4628 35697
rect 4684 35641 4696 35697
rect 4616 35629 4696 35641
rect 5434 35697 5514 35709
rect 5434 35641 5446 35697
rect 5502 35641 5514 35697
rect 5434 35629 5514 35641
rect 14088 35698 14168 35710
rect 14088 35642 14100 35698
rect 14156 35642 14168 35698
rect 14088 35630 14168 35642
rect 14906 35698 14986 35710
rect 14906 35642 14918 35698
rect 14974 35642 14986 35698
rect 14906 35630 14986 35642
rect 23560 35698 23640 35710
rect 23560 35642 23572 35698
rect 23628 35642 23640 35698
rect 23560 35630 23640 35642
rect 24378 35698 24458 35710
rect 24378 35642 24390 35698
rect 24446 35642 24458 35698
rect 24378 35630 24458 35642
rect 33032 35698 33112 35710
rect 33032 35642 33044 35698
rect 33100 35642 33112 35698
rect 33032 35630 33112 35642
rect 33850 35698 33930 35710
rect 33850 35642 33862 35698
rect 33918 35642 33930 35698
rect 33850 35630 33930 35642
rect 42504 35698 42584 35710
rect 42504 35642 42516 35698
rect 42572 35642 42584 35698
rect 42504 35630 42584 35642
rect 43322 35698 43402 35710
rect 43322 35642 43334 35698
rect 43390 35642 43402 35698
rect 43322 35630 43402 35642
rect -4355 35362 -4269 35366
rect -4355 35306 -4343 35362
rect -4287 35306 -4269 35362
rect -4355 35294 -4269 35306
rect -2869 35362 -2783 35366
rect -2869 35306 -2857 35362
rect -2801 35306 -2783 35362
rect -2869 35294 -2783 35306
rect 5117 35362 5203 35366
rect 5117 35306 5129 35362
rect 5185 35306 5203 35362
rect 5117 35294 5203 35306
rect 6603 35362 6689 35366
rect 6603 35306 6615 35362
rect 6671 35306 6689 35362
rect 6603 35294 6689 35306
rect 14589 35363 14675 35367
rect 14589 35307 14601 35363
rect 14657 35307 14675 35363
rect 14589 35295 14675 35307
rect 16075 35363 16161 35367
rect 16075 35307 16087 35363
rect 16143 35307 16161 35363
rect 16075 35295 16161 35307
rect 24061 35363 24147 35367
rect 24061 35307 24073 35363
rect 24129 35307 24147 35363
rect 24061 35295 24147 35307
rect 25547 35363 25633 35367
rect 25547 35307 25559 35363
rect 25615 35307 25633 35363
rect 25547 35295 25633 35307
rect 33533 35363 33619 35367
rect 33533 35307 33545 35363
rect 33601 35307 33619 35363
rect 33533 35295 33619 35307
rect 35019 35363 35105 35367
rect 35019 35307 35031 35363
rect 35087 35307 35105 35363
rect 35019 35295 35105 35307
rect 43005 35363 43091 35367
rect 43005 35307 43017 35363
rect 43073 35307 43091 35363
rect 43005 35295 43091 35307
rect 44491 35363 44577 35367
rect 44491 35307 44503 35363
rect 44559 35307 44577 35363
rect 44491 35295 44577 35307
rect -4856 33492 -4776 33504
rect -4856 33436 -4844 33492
rect -4788 33436 -4776 33492
rect -4856 33424 -4776 33436
rect -4038 33492 -3958 33504
rect -4038 33436 -4026 33492
rect -3970 33436 -3958 33492
rect -4038 33424 -3958 33436
rect -3370 33492 -3290 33504
rect -3370 33436 -3358 33492
rect -3302 33436 -3290 33492
rect -3370 33424 -3290 33436
rect -2552 33492 -2472 33504
rect -2552 33436 -2540 33492
rect -2484 33436 -2472 33492
rect -2552 33424 -2472 33436
rect 4616 33492 4696 33504
rect 4616 33436 4628 33492
rect 4684 33436 4696 33492
rect 4616 33424 4696 33436
rect 5434 33492 5514 33504
rect 5434 33436 5446 33492
rect 5502 33436 5514 33492
rect 5434 33424 5514 33436
rect 6102 33492 6182 33504
rect 6102 33436 6114 33492
rect 6170 33436 6182 33492
rect 6102 33424 6182 33436
rect 6920 33492 7000 33504
rect 6920 33436 6932 33492
rect 6988 33436 7000 33492
rect 6920 33424 7000 33436
rect 14088 33493 14168 33505
rect 14088 33437 14100 33493
rect 14156 33437 14168 33493
rect 14088 33425 14168 33437
rect 14906 33493 14986 33505
rect 14906 33437 14918 33493
rect 14974 33437 14986 33493
rect 14906 33425 14986 33437
rect 15574 33493 15654 33505
rect 15574 33437 15586 33493
rect 15642 33437 15654 33493
rect 15574 33425 15654 33437
rect 16392 33493 16472 33505
rect 16392 33437 16404 33493
rect 16460 33437 16472 33493
rect 16392 33425 16472 33437
rect 23560 33493 23640 33505
rect 23560 33437 23572 33493
rect 23628 33437 23640 33493
rect 23560 33425 23640 33437
rect 24378 33493 24458 33505
rect 24378 33437 24390 33493
rect 24446 33437 24458 33493
rect 24378 33425 24458 33437
rect 25046 33493 25126 33505
rect 25046 33437 25058 33493
rect 25114 33437 25126 33493
rect 25046 33425 25126 33437
rect 25864 33493 25944 33505
rect 25864 33437 25876 33493
rect 25932 33437 25944 33493
rect 25864 33425 25944 33437
rect 33032 33493 33112 33505
rect 33032 33437 33044 33493
rect 33100 33437 33112 33493
rect 33032 33425 33112 33437
rect 33850 33493 33930 33505
rect 33850 33437 33862 33493
rect 33918 33437 33930 33493
rect 33850 33425 33930 33437
rect 34518 33493 34598 33505
rect 34518 33437 34530 33493
rect 34586 33437 34598 33493
rect 34518 33425 34598 33437
rect 35336 33493 35416 33505
rect 35336 33437 35348 33493
rect 35404 33437 35416 33493
rect 35336 33425 35416 33437
rect 42504 33493 42584 33505
rect 42504 33437 42516 33493
rect 42572 33437 42584 33493
rect 42504 33425 42584 33437
rect 43322 33493 43402 33505
rect 43322 33437 43334 33493
rect 43390 33437 43402 33493
rect 43322 33425 43402 33437
rect 43990 33493 44070 33505
rect 43990 33437 44002 33493
rect 44058 33437 44070 33493
rect 43990 33425 44070 33437
rect 44808 33493 44888 33505
rect 44808 33437 44820 33493
rect 44876 33437 44888 33493
rect 44808 33425 44888 33437
rect -8103 33375 -8027 33382
rect -5721 33375 -5639 33387
rect -8103 33372 -5707 33375
rect -8103 33316 -8093 33372
rect -8037 33319 -5707 33372
rect -5651 33368 -5639 33375
rect 3751 33375 3833 33387
rect 3751 33368 3765 33375
rect -5651 33319 3765 33368
rect 3821 33368 3833 33375
rect 13223 33376 13305 33388
rect 13223 33368 13237 33376
rect 3821 33320 13237 33368
rect 13293 33368 13305 33376
rect 22695 33376 22777 33388
rect 22695 33368 22709 33376
rect 13293 33320 22709 33368
rect 22765 33368 22777 33376
rect 32167 33376 32249 33388
rect 32167 33368 32181 33376
rect 22765 33320 32181 33368
rect 32237 33368 32249 33376
rect 41639 33376 41721 33388
rect 41639 33368 41653 33376
rect 32237 33320 41653 33368
rect 41709 33320 41721 33376
rect 3821 33319 41721 33320
rect -8037 33316 41721 33319
rect -8103 33314 41721 33316
rect -8103 33306 -8027 33314
rect -5721 33308 41721 33314
rect -5721 33307 41639 33308
rect -4355 33157 -4269 33161
rect -4355 33101 -4343 33157
rect -4287 33101 -4269 33157
rect -4355 33089 -4269 33101
rect -2869 33158 -2783 33162
rect -2869 33102 -2857 33158
rect -2801 33102 -2783 33158
rect -2869 33090 -2783 33102
rect 5117 33157 5203 33161
rect 5117 33101 5129 33157
rect 5185 33101 5203 33157
rect 5117 33089 5203 33101
rect 6603 33158 6689 33162
rect 6603 33102 6615 33158
rect 6671 33102 6689 33158
rect 6603 33090 6689 33102
rect 14589 33158 14675 33162
rect 14589 33102 14601 33158
rect 14657 33102 14675 33158
rect 14589 33090 14675 33102
rect 16075 33159 16161 33163
rect 16075 33103 16087 33159
rect 16143 33103 16161 33159
rect 16075 33091 16161 33103
rect 24061 33158 24147 33162
rect 24061 33102 24073 33158
rect 24129 33102 24147 33158
rect 24061 33090 24147 33102
rect 25547 33159 25633 33163
rect 25547 33103 25559 33159
rect 25615 33103 25633 33159
rect 25547 33091 25633 33103
rect 33533 33158 33619 33162
rect 33533 33102 33545 33158
rect 33601 33102 33619 33158
rect 33533 33090 33619 33102
rect 35019 33159 35105 33163
rect 35019 33103 35031 33159
rect 35087 33103 35105 33159
rect 35019 33091 35105 33103
rect 43005 33158 43091 33162
rect 43005 33102 43017 33158
rect 43073 33102 43091 33158
rect 43005 33090 43091 33102
rect 44491 33159 44577 33163
rect 44491 33103 44503 33159
rect 44559 33103 44577 33159
rect 44491 33091 44577 33103
rect -6337 31969 -6017 31979
rect -6337 31169 -6327 31969
rect -6027 31169 -6017 31969
rect -1255 31969 -1035 31979
rect -4856 31287 -4776 31299
rect -4856 31231 -4844 31287
rect -4788 31231 -4776 31287
rect -4856 31219 -4776 31231
rect -4038 31287 -3958 31299
rect -4038 31231 -4026 31287
rect -3970 31231 -3958 31287
rect -4038 31219 -3958 31231
rect -3370 31288 -3290 31300
rect -3370 31232 -3358 31288
rect -3302 31232 -3290 31288
rect -3370 31220 -3290 31232
rect -2552 31288 -2472 31300
rect -2552 31232 -2540 31288
rect -2484 31232 -2472 31288
rect -2552 31220 -2472 31232
rect -6337 31159 -6017 31169
rect -1255 31169 -1245 31969
rect -1045 31169 -1035 31969
rect -1255 31159 -1035 31169
rect 3135 31969 3455 31979
rect 3135 31169 3145 31969
rect 3445 31169 3455 31969
rect 8217 31970 8437 31980
rect 4616 31287 4696 31299
rect 4616 31231 4628 31287
rect 4684 31231 4696 31287
rect 4616 31219 4696 31231
rect 5434 31287 5514 31299
rect 5434 31231 5446 31287
rect 5502 31231 5514 31287
rect 5434 31219 5514 31231
rect 6102 31288 6182 31300
rect 6102 31232 6114 31288
rect 6170 31232 6182 31288
rect 6102 31220 6182 31232
rect 6920 31288 7000 31300
rect 6920 31232 6932 31288
rect 6988 31232 7000 31288
rect 6920 31220 7000 31232
rect 3135 31159 3455 31169
rect 8217 31170 8227 31970
rect 8427 31170 8437 31970
rect 8217 31160 8437 31170
rect 12607 31970 12927 31980
rect 12607 31170 12617 31970
rect 12917 31170 12927 31970
rect 17689 31970 17909 31980
rect 14088 31288 14168 31300
rect 14088 31232 14100 31288
rect 14156 31232 14168 31288
rect 14088 31220 14168 31232
rect 14906 31288 14986 31300
rect 14906 31232 14918 31288
rect 14974 31232 14986 31288
rect 14906 31220 14986 31232
rect 15574 31289 15654 31301
rect 15574 31233 15586 31289
rect 15642 31233 15654 31289
rect 15574 31221 15654 31233
rect 16392 31289 16472 31301
rect 16392 31233 16404 31289
rect 16460 31233 16472 31289
rect 16392 31221 16472 31233
rect 12607 31160 12927 31170
rect 17689 31170 17699 31970
rect 17899 31170 17909 31970
rect 17689 31160 17909 31170
rect 22079 31970 22399 31980
rect 22079 31170 22089 31970
rect 22389 31170 22399 31970
rect 27161 31970 27381 31980
rect 23560 31288 23640 31300
rect 23560 31232 23572 31288
rect 23628 31232 23640 31288
rect 23560 31220 23640 31232
rect 24378 31288 24458 31300
rect 24378 31232 24390 31288
rect 24446 31232 24458 31288
rect 24378 31220 24458 31232
rect 25046 31289 25126 31301
rect 25046 31233 25058 31289
rect 25114 31233 25126 31289
rect 25046 31221 25126 31233
rect 25864 31289 25944 31301
rect 25864 31233 25876 31289
rect 25932 31233 25944 31289
rect 25864 31221 25944 31233
rect 22079 31160 22399 31170
rect 27161 31170 27171 31970
rect 27371 31170 27381 31970
rect 27161 31160 27381 31170
rect 31551 31970 31871 31980
rect 31551 31170 31561 31970
rect 31861 31170 31871 31970
rect 36633 31970 36853 31980
rect 33032 31288 33112 31300
rect 33032 31232 33044 31288
rect 33100 31232 33112 31288
rect 33032 31220 33112 31232
rect 33850 31288 33930 31300
rect 33850 31232 33862 31288
rect 33918 31232 33930 31288
rect 33850 31220 33930 31232
rect 34518 31289 34598 31301
rect 34518 31233 34530 31289
rect 34586 31233 34598 31289
rect 34518 31221 34598 31233
rect 35336 31289 35416 31301
rect 35336 31233 35348 31289
rect 35404 31233 35416 31289
rect 35336 31221 35416 31233
rect 31551 31160 31871 31170
rect 36633 31170 36643 31970
rect 36843 31170 36853 31970
rect 36633 31160 36853 31170
rect 41023 31970 41343 31980
rect 41023 31170 41033 31970
rect 41333 31170 41343 31970
rect 42504 31288 42584 31300
rect 42504 31232 42516 31288
rect 42572 31232 42584 31288
rect 42504 31220 42584 31232
rect 43322 31288 43402 31300
rect 43322 31232 43334 31288
rect 43390 31232 43402 31288
rect 43322 31220 43402 31232
rect 43990 31289 44070 31301
rect 43990 31233 44002 31289
rect 44058 31233 44070 31289
rect 43990 31221 44070 31233
rect 44808 31289 44888 31301
rect 44808 31233 44820 31289
rect 44876 31233 44888 31289
rect 44808 31221 44888 31233
rect 41023 31160 41343 31170
rect -10211 31005 -10131 31015
rect -10211 30949 -10199 31005
rect -10143 30949 -10131 31005
rect -10211 30176 -10131 30949
rect -7707 30973 -5915 30985
rect -7707 30833 -7695 30973
rect -5927 30833 -5915 30973
rect 1765 30973 3557 30985
rect -4355 30952 -4269 30956
rect -4355 30896 -4343 30952
rect -4287 30896 -4269 30952
rect -4355 30884 -4269 30896
rect -9181 30567 -8693 30577
rect -9181 30511 -9169 30567
rect -9113 30511 -8761 30567
rect -8705 30511 -8693 30567
rect -9181 30501 -8693 30511
rect -8767 30199 -8143 30211
rect -10211 30166 -9895 30176
rect -10211 30090 -9985 30166
rect -9905 30090 -9895 30166
rect -10211 30080 -9895 30090
rect -8767 30059 -8755 30199
rect -8155 30059 -8143 30199
rect -8767 30047 -8143 30059
rect -7707 29811 -5915 30833
rect 1765 30833 1777 30973
rect 3545 30833 3557 30973
rect 11237 30974 13029 30986
rect 5117 30952 5203 30956
rect 5117 30896 5129 30952
rect 5185 30896 5203 30952
rect 5117 30884 5203 30896
rect 291 30567 779 30577
rect 291 30511 303 30567
rect 359 30511 711 30567
rect 767 30511 779 30567
rect 291 30501 779 30511
rect 705 30199 1329 30211
rect 705 30059 717 30199
rect 1317 30059 1329 30199
rect 705 30047 1329 30059
rect 1765 29811 3557 30833
rect 11237 30834 11249 30974
rect 13017 30834 13029 30974
rect 20709 30974 22501 30986
rect 14589 30953 14675 30957
rect 14589 30897 14601 30953
rect 14657 30897 14675 30953
rect 14589 30885 14675 30897
rect 9763 30568 10251 30578
rect 9763 30512 9775 30568
rect 9831 30512 10183 30568
rect 10239 30512 10251 30568
rect 9763 30502 10251 30512
rect 10177 30200 10801 30212
rect 10177 30060 10189 30200
rect 10789 30060 10801 30200
rect 10177 30048 10801 30060
rect 11237 29812 13029 30834
rect 20709 30834 20721 30974
rect 22489 30834 22501 30974
rect 30181 30974 31973 30986
rect 24061 30953 24147 30957
rect 24061 30897 24073 30953
rect 24129 30897 24147 30953
rect 24061 30885 24147 30897
rect 19235 30568 19723 30578
rect 19235 30512 19247 30568
rect 19303 30512 19655 30568
rect 19711 30512 19723 30568
rect 19235 30502 19723 30512
rect 19649 30200 20273 30212
rect 19649 30060 19661 30200
rect 20261 30060 20273 30200
rect 19649 30048 20273 30060
rect 20709 29812 22501 30834
rect 30181 30834 30193 30974
rect 31961 30834 31973 30974
rect 39653 30974 41445 30986
rect 33533 30953 33619 30957
rect 33533 30897 33545 30953
rect 33601 30897 33619 30953
rect 33533 30885 33619 30897
rect 28707 30568 29195 30578
rect 28707 30512 28719 30568
rect 28775 30512 29127 30568
rect 29183 30512 29195 30568
rect 28707 30502 29195 30512
rect 29121 30200 29745 30212
rect 29121 30060 29133 30200
rect 29733 30060 29745 30200
rect 29121 30048 29745 30060
rect 30181 29812 31973 30834
rect 39653 30834 39665 30974
rect 41433 30834 41445 30974
rect 43005 30953 43091 30957
rect 43005 30897 43017 30953
rect 43073 30897 43091 30953
rect 43005 30885 43091 30897
rect 38179 30568 38667 30578
rect 38179 30512 38191 30568
rect 38247 30512 38599 30568
rect 38655 30512 38667 30568
rect 38179 30502 38667 30512
rect 38593 30200 39217 30212
rect 38593 30060 38605 30200
rect 39205 30060 39217 30200
rect 38593 30048 39217 30060
rect 39653 29812 41445 30834
rect -8767 29799 -5915 29811
rect -8767 29659 -8755 29799
rect -8155 29659 -5915 29799
rect -8767 29647 -5915 29659
rect 705 29799 3557 29811
rect 705 29659 717 29799
rect 1317 29659 3557 29799
rect 705 29647 3557 29659
rect 10177 29800 13029 29812
rect 10177 29660 10189 29800
rect 10789 29660 13029 29800
rect 10177 29648 13029 29660
rect 19649 29800 22501 29812
rect 19649 29660 19661 29800
rect 20261 29660 22501 29800
rect 19649 29648 22501 29660
rect 29121 29800 31973 29812
rect 29121 29660 29133 29800
rect 29733 29660 31973 29800
rect 29121 29648 31973 29660
rect 38593 29800 41445 29812
rect 38593 29660 38605 29800
rect 39205 29660 41445 29800
rect 38593 29648 41445 29660
rect -4856 29082 -4776 29094
rect -4856 29026 -4844 29082
rect -4788 29026 -4776 29082
rect -7707 29013 -5915 29025
rect -4856 29014 -4776 29026
rect -4038 29082 -3958 29094
rect -4038 29026 -4026 29082
rect -3970 29026 -3958 29082
rect -4038 29014 -3958 29026
rect 4616 29082 4696 29094
rect 4616 29026 4628 29082
rect 4684 29026 4696 29082
rect -7707 28873 -7695 29013
rect -5927 28873 -5915 29013
rect 1765 29013 3557 29025
rect 4616 29014 4696 29026
rect 5434 29082 5514 29094
rect 5434 29026 5446 29082
rect 5502 29026 5514 29082
rect 14088 29083 14168 29095
rect 14088 29027 14100 29083
rect 14156 29027 14168 29083
rect 5434 29014 5514 29026
rect 11237 29014 13029 29026
rect 14088 29015 14168 29027
rect 14906 29083 14986 29095
rect 14906 29027 14918 29083
rect 14974 29027 14986 29083
rect 14906 29015 14986 29027
rect 23560 29083 23640 29095
rect 23560 29027 23572 29083
rect 23628 29027 23640 29083
rect -5622 28964 -5536 28976
rect -5622 28908 -5610 28964
rect -5554 28908 -5536 28964
rect -5622 28896 -5536 28908
rect -7707 28861 -5915 28873
rect 1765 28873 1777 29013
rect 3545 28873 3557 29013
rect 3850 28964 3936 28976
rect 3850 28908 3862 28964
rect 3918 28908 3936 28964
rect 3850 28896 3936 28908
rect 1765 28861 3557 28873
rect 11237 28874 11249 29014
rect 13017 28874 13029 29014
rect 20709 29014 22501 29026
rect 23560 29015 23640 29027
rect 24378 29083 24458 29095
rect 24378 29027 24390 29083
rect 24446 29027 24458 29083
rect 24378 29015 24458 29027
rect 33032 29083 33112 29095
rect 33032 29027 33044 29083
rect 33100 29027 33112 29083
rect 13322 28965 13408 28977
rect 13322 28909 13334 28965
rect 13390 28909 13408 28965
rect 13322 28897 13408 28909
rect 11237 28862 13029 28874
rect 20709 28874 20721 29014
rect 22489 28874 22501 29014
rect 30181 29014 31973 29026
rect 33032 29015 33112 29027
rect 33850 29083 33930 29095
rect 33850 29027 33862 29083
rect 33918 29027 33930 29083
rect 33850 29015 33930 29027
rect 42504 29083 42584 29095
rect 42504 29027 42516 29083
rect 42572 29027 42584 29083
rect 22794 28965 22880 28977
rect 22794 28909 22806 28965
rect 22862 28909 22880 28965
rect 22794 28897 22880 28909
rect 20709 28862 22501 28874
rect 30181 28874 30193 29014
rect 31961 28874 31973 29014
rect 39653 29014 41445 29026
rect 42504 29015 42584 29027
rect 43322 29083 43402 29095
rect 43322 29027 43334 29083
rect 43390 29027 43402 29083
rect 43322 29015 43402 29027
rect 32266 28965 32352 28977
rect 32266 28909 32278 28965
rect 32334 28909 32352 28965
rect 32266 28897 32352 28909
rect 30181 28862 31973 28874
rect 39653 28874 39665 29014
rect 41433 28874 41445 29014
rect 41738 28965 41824 28977
rect 41738 28909 41750 28965
rect 41806 28909 41824 28965
rect 41738 28897 41824 28909
rect 39653 28862 41445 28874
rect -6337 28689 -6017 28699
rect -9181 28227 -8693 28237
rect -9181 28171 -9169 28227
rect -9113 28171 -8761 28227
rect -8705 28171 -8693 28227
rect -9181 28161 -8693 28171
rect -6337 27889 -6327 28689
rect -6027 27889 -6017 28689
rect 3135 28689 3455 28699
rect 291 28227 779 28237
rect 291 28171 303 28227
rect 359 28171 711 28227
rect 767 28171 779 28227
rect 291 28161 779 28171
rect -6337 27879 -6017 27889
rect 3135 27889 3145 28689
rect 3445 27889 3455 28689
rect 12607 28690 12927 28700
rect 9763 28228 10251 28238
rect 9763 28172 9775 28228
rect 9831 28172 10183 28228
rect 10239 28172 10251 28228
rect 9763 28162 10251 28172
rect 3135 27879 3455 27889
rect 12607 27890 12617 28690
rect 12917 27890 12927 28690
rect 22079 28690 22399 28700
rect 19235 28228 19723 28238
rect 19235 28172 19247 28228
rect 19303 28172 19655 28228
rect 19711 28172 19723 28228
rect 19235 28162 19723 28172
rect 12607 27880 12927 27890
rect 22079 27890 22089 28690
rect 22389 27890 22399 28690
rect 31551 28690 31871 28700
rect 28707 28228 29195 28238
rect 28707 28172 28719 28228
rect 28775 28172 29127 28228
rect 29183 28172 29195 28228
rect 28707 28162 29195 28172
rect 22079 27880 22399 27890
rect 31551 27890 31561 28690
rect 31861 27890 31871 28690
rect 41023 28690 41343 28700
rect 38179 28228 38667 28238
rect 38179 28172 38191 28228
rect 38247 28172 38599 28228
rect 38655 28172 38667 28228
rect 38179 28162 38667 28172
rect 31551 27880 31871 27890
rect 41023 27890 41033 28690
rect 41333 27890 41343 28690
rect 41023 27880 41343 27890
rect -2074 27608 -2064 27609
rect -11840 27577 -11592 27608
rect -11840 27521 -11830 27577
rect -11774 27521 -11592 27577
rect -11840 27490 -11592 27521
rect -11602 27488 -11592 27490
rect -11536 27490 -2064 27608
rect -11536 27488 -11526 27490
rect -2074 27489 -2064 27490
rect -2008 27608 -1998 27609
rect 7398 27608 7408 27609
rect -2008 27490 7408 27608
rect -2008 27489 -1998 27490
rect 7398 27489 7408 27490
rect 7464 27608 7474 27609
rect 16870 27608 16880 27610
rect 7464 27490 16880 27608
rect 16936 27608 16946 27610
rect 26342 27608 26352 27610
rect 16936 27490 26352 27608
rect 26408 27608 26418 27610
rect 35814 27608 35824 27610
rect 26408 27490 35824 27608
rect 35880 27490 35890 27610
rect 7464 27489 7474 27490
rect -7613 25265 -7527 25269
rect -7613 25209 -7601 25265
rect -7545 25209 -7527 25265
rect -7613 25197 -7527 25209
rect -3571 25262 -3485 25266
rect -3571 25206 -3559 25262
rect -3503 25206 -3485 25262
rect -3571 25194 -3485 25206
rect 471 25262 557 25266
rect 471 25206 483 25262
rect 539 25206 557 25262
rect 471 25194 557 25206
rect 4513 25262 4599 25266
rect 4513 25206 4525 25262
rect 4581 25206 4599 25262
rect 4513 25194 4599 25206
rect 8555 25262 8641 25266
rect 8555 25206 8567 25262
rect 8623 25206 8641 25262
rect 8555 25194 8641 25206
rect 12597 25262 12683 25266
rect 12597 25206 12609 25262
rect 12665 25206 12683 25262
rect 12597 25194 12683 25206
rect 16639 25262 16725 25266
rect 16639 25206 16651 25262
rect 16707 25206 16725 25262
rect 16639 25194 16725 25206
rect -8114 23395 -8034 23407
rect -8114 23339 -8102 23395
rect -8046 23339 -8034 23395
rect -8114 23327 -8034 23339
rect -7296 23395 -7216 23407
rect -7296 23339 -7284 23395
rect -7228 23339 -7216 23395
rect -7296 23327 -7216 23339
rect -4072 23392 -3992 23404
rect -4072 23336 -4060 23392
rect -4004 23336 -3992 23392
rect -4072 23324 -3992 23336
rect -3254 23392 -3174 23404
rect -3254 23336 -3242 23392
rect -3186 23336 -3174 23392
rect -3254 23324 -3174 23336
rect -30 23392 50 23404
rect -30 23336 -18 23392
rect 38 23336 50 23392
rect -30 23324 50 23336
rect 788 23392 868 23404
rect 788 23336 800 23392
rect 856 23336 868 23392
rect 788 23324 868 23336
rect 4012 23392 4092 23404
rect 4012 23336 4024 23392
rect 4080 23336 4092 23392
rect 4012 23324 4092 23336
rect 4830 23392 4910 23404
rect 4830 23336 4842 23392
rect 4898 23336 4910 23392
rect 4830 23324 4910 23336
rect 8054 23392 8134 23404
rect 8054 23336 8066 23392
rect 8122 23336 8134 23392
rect 8054 23324 8134 23336
rect 8872 23392 8952 23404
rect 8872 23336 8884 23392
rect 8940 23336 8952 23392
rect 8872 23324 8952 23336
rect 12096 23392 12176 23404
rect 12096 23336 12108 23392
rect 12164 23336 12176 23392
rect 12096 23324 12176 23336
rect 12914 23392 12994 23404
rect 12914 23336 12926 23392
rect 12982 23336 12994 23392
rect 12914 23324 12994 23336
rect 16138 23392 16218 23404
rect 16138 23336 16150 23392
rect 16206 23336 16218 23392
rect 16138 23324 16218 23336
rect 16956 23392 17036 23404
rect 16956 23336 16968 23392
rect 17024 23336 17036 23392
rect 16956 23324 17036 23336
rect -7613 23060 -7527 23064
rect -7613 23004 -7601 23060
rect -7545 23004 -7527 23060
rect -7613 22992 -7527 23004
rect -6127 23060 -6041 23064
rect -6127 23004 -6115 23060
rect -6059 23004 -6041 23060
rect -6127 22992 -6041 23004
rect -3571 23057 -3485 23061
rect -3571 23001 -3559 23057
rect -3503 23001 -3485 23057
rect -3571 22989 -3485 23001
rect -2085 23057 -1999 23061
rect -2085 23001 -2073 23057
rect -2017 23001 -1999 23057
rect -2085 22989 -1999 23001
rect 471 23057 557 23061
rect 471 23001 483 23057
rect 539 23001 557 23057
rect 471 22989 557 23001
rect 1957 23057 2043 23061
rect 1957 23001 1969 23057
rect 2025 23001 2043 23057
rect 1957 22989 2043 23001
rect 4513 23057 4599 23061
rect 4513 23001 4525 23057
rect 4581 23001 4599 23057
rect 4513 22989 4599 23001
rect 5999 23057 6085 23061
rect 5999 23001 6011 23057
rect 6067 23001 6085 23057
rect 5999 22989 6085 23001
rect 8555 23057 8641 23061
rect 8555 23001 8567 23057
rect 8623 23001 8641 23057
rect 8555 22989 8641 23001
rect 10041 23057 10127 23061
rect 10041 23001 10053 23057
rect 10109 23001 10127 23057
rect 10041 22989 10127 23001
rect 12597 23057 12683 23061
rect 12597 23001 12609 23057
rect 12665 23001 12683 23057
rect 12597 22989 12683 23001
rect 14083 23057 14169 23061
rect 14083 23001 14095 23057
rect 14151 23001 14169 23057
rect 14083 22989 14169 23001
rect 16639 23057 16725 23061
rect 16639 23001 16651 23057
rect 16707 23001 16725 23057
rect 16639 22989 16725 23001
rect 18125 23057 18211 23061
rect 18125 23001 18137 23057
rect 18193 23001 18211 23057
rect 18125 22989 18211 23001
rect -8114 21190 -8034 21202
rect -8114 21134 -8102 21190
rect -8046 21134 -8034 21190
rect -8114 21122 -8034 21134
rect -7296 21190 -7216 21202
rect -7296 21134 -7284 21190
rect -7228 21134 -7216 21190
rect -7296 21122 -7216 21134
rect -6628 21190 -6548 21202
rect -6628 21134 -6616 21190
rect -6560 21134 -6548 21190
rect -6628 21122 -6548 21134
rect -5810 21190 -5730 21202
rect -5810 21134 -5798 21190
rect -5742 21134 -5730 21190
rect -5810 21122 -5730 21134
rect -4072 21187 -3992 21199
rect -4072 21131 -4060 21187
rect -4004 21131 -3992 21187
rect -4072 21119 -3992 21131
rect -3254 21187 -3174 21199
rect -3254 21131 -3242 21187
rect -3186 21131 -3174 21187
rect -3254 21119 -3174 21131
rect -2586 21187 -2506 21199
rect -2586 21131 -2574 21187
rect -2518 21131 -2506 21187
rect -2586 21119 -2506 21131
rect -1768 21187 -1688 21199
rect -1768 21131 -1756 21187
rect -1700 21131 -1688 21187
rect -1768 21119 -1688 21131
rect -30 21187 50 21199
rect -30 21131 -18 21187
rect 38 21131 50 21187
rect -30 21119 50 21131
rect 788 21187 868 21199
rect 788 21131 800 21187
rect 856 21131 868 21187
rect 788 21119 868 21131
rect 1456 21187 1536 21199
rect 1456 21131 1468 21187
rect 1524 21131 1536 21187
rect 1456 21119 1536 21131
rect 2274 21187 2354 21199
rect 2274 21131 2286 21187
rect 2342 21131 2354 21187
rect 2274 21119 2354 21131
rect 4012 21187 4092 21199
rect 4012 21131 4024 21187
rect 4080 21131 4092 21187
rect 4012 21119 4092 21131
rect 4830 21187 4910 21199
rect 4830 21131 4842 21187
rect 4898 21131 4910 21187
rect 4830 21119 4910 21131
rect 5498 21187 5578 21199
rect 5498 21131 5510 21187
rect 5566 21131 5578 21187
rect 5498 21119 5578 21131
rect 6316 21187 6396 21199
rect 6316 21131 6328 21187
rect 6384 21131 6396 21187
rect 6316 21119 6396 21131
rect 8054 21187 8134 21199
rect 8054 21131 8066 21187
rect 8122 21131 8134 21187
rect 8054 21119 8134 21131
rect 8872 21187 8952 21199
rect 8872 21131 8884 21187
rect 8940 21131 8952 21187
rect 8872 21119 8952 21131
rect 9540 21187 9620 21199
rect 9540 21131 9552 21187
rect 9608 21131 9620 21187
rect 9540 21119 9620 21131
rect 10358 21187 10438 21199
rect 10358 21131 10370 21187
rect 10426 21131 10438 21187
rect 10358 21119 10438 21131
rect 12096 21187 12176 21199
rect 12096 21131 12108 21187
rect 12164 21131 12176 21187
rect 12096 21119 12176 21131
rect 12914 21187 12994 21199
rect 12914 21131 12926 21187
rect 12982 21131 12994 21187
rect 12914 21119 12994 21131
rect 13582 21187 13662 21199
rect 13582 21131 13594 21187
rect 13650 21131 13662 21187
rect 13582 21119 13662 21131
rect 14400 21187 14480 21199
rect 14400 21131 14412 21187
rect 14468 21131 14480 21187
rect 14400 21119 14480 21131
rect 16138 21187 16218 21199
rect 16138 21131 16150 21187
rect 16206 21131 16218 21187
rect 16138 21119 16218 21131
rect 16956 21187 17036 21199
rect 16956 21131 16968 21187
rect 17024 21131 17036 21187
rect 16956 21119 17036 21131
rect 17624 21187 17704 21199
rect 17624 21131 17636 21187
rect 17692 21131 17704 21187
rect 17624 21119 17704 21131
rect 18442 21187 18522 21199
rect 18442 21131 18454 21187
rect 18510 21131 18522 21187
rect 18442 21119 18522 21131
rect 15375 21070 15453 21082
rect 15375 21014 15386 21070
rect 15442 21014 15453 21070
rect 15375 21002 15453 21014
rect -7613 20855 -7527 20859
rect -7613 20799 -7601 20855
rect -7545 20799 -7527 20855
rect -7613 20787 -7527 20799
rect -6127 20856 -6041 20860
rect -6127 20800 -6115 20856
rect -6059 20800 -6041 20856
rect -6127 20788 -6041 20800
rect -3571 20852 -3485 20856
rect -3571 20796 -3559 20852
rect -3503 20796 -3485 20852
rect -3571 20784 -3485 20796
rect -2085 20853 -1999 20857
rect -2085 20797 -2073 20853
rect -2017 20797 -1999 20853
rect -2085 20785 -1999 20797
rect 471 20852 557 20856
rect 471 20796 483 20852
rect 539 20796 557 20852
rect 471 20784 557 20796
rect 1957 20853 2043 20857
rect 1957 20797 1969 20853
rect 2025 20797 2043 20853
rect 1957 20785 2043 20797
rect 4513 20852 4599 20856
rect 4513 20796 4525 20852
rect 4581 20796 4599 20852
rect 4513 20784 4599 20796
rect 5999 20853 6085 20857
rect 5999 20797 6011 20853
rect 6067 20797 6085 20853
rect 5999 20785 6085 20797
rect 8555 20852 8641 20856
rect 8555 20796 8567 20852
rect 8623 20796 8641 20852
rect 8555 20784 8641 20796
rect 10041 20853 10127 20857
rect 10041 20797 10053 20853
rect 10109 20797 10127 20853
rect 10041 20785 10127 20797
rect 12597 20852 12683 20856
rect 12597 20796 12609 20852
rect 12665 20796 12683 20852
rect 12597 20784 12683 20796
rect 14083 20853 14169 20857
rect 14083 20797 14095 20853
rect 14151 20797 14169 20853
rect 14083 20785 14169 20797
rect 16639 20852 16725 20856
rect 16639 20796 16651 20852
rect 16707 20796 16725 20852
rect 16639 20784 16725 20796
rect 18125 20853 18211 20857
rect 18125 20797 18137 20853
rect 18193 20797 18211 20853
rect 18125 20785 18211 20797
rect -8114 18985 -8034 18997
rect -8114 18929 -8102 18985
rect -8046 18929 -8034 18985
rect -8114 18917 -8034 18929
rect -7296 18985 -7216 18997
rect -7296 18929 -7284 18985
rect -7228 18929 -7216 18985
rect -7296 18917 -7216 18929
rect -6628 18986 -6548 18998
rect -6628 18930 -6616 18986
rect -6560 18930 -6548 18986
rect -6628 18918 -6548 18930
rect -5810 18986 -5730 18998
rect -5810 18930 -5798 18986
rect -5742 18930 -5730 18986
rect -5810 18918 -5730 18930
rect -4072 18982 -3992 18994
rect -4072 18926 -4060 18982
rect -4004 18926 -3992 18982
rect -4072 18914 -3992 18926
rect -3254 18982 -3174 18994
rect -3254 18926 -3242 18982
rect -3186 18926 -3174 18982
rect -3254 18914 -3174 18926
rect -2586 18983 -2506 18995
rect -2586 18927 -2574 18983
rect -2518 18927 -2506 18983
rect -2586 18915 -2506 18927
rect -1768 18983 -1688 18995
rect -1768 18927 -1756 18983
rect -1700 18927 -1688 18983
rect -1768 18915 -1688 18927
rect -30 18982 50 18994
rect -30 18926 -18 18982
rect 38 18926 50 18982
rect -30 18914 50 18926
rect 788 18982 868 18994
rect 788 18926 800 18982
rect 856 18926 868 18982
rect 788 18914 868 18926
rect 1456 18983 1536 18995
rect 1456 18927 1468 18983
rect 1524 18927 1536 18983
rect 1456 18915 1536 18927
rect 2274 18983 2354 18995
rect 2274 18927 2286 18983
rect 2342 18927 2354 18983
rect 2274 18915 2354 18927
rect 4012 18982 4092 18994
rect 4012 18926 4024 18982
rect 4080 18926 4092 18982
rect 4012 18914 4092 18926
rect 4830 18982 4910 18994
rect 4830 18926 4842 18982
rect 4898 18926 4910 18982
rect 4830 18914 4910 18926
rect 5498 18983 5578 18995
rect 5498 18927 5510 18983
rect 5566 18927 5578 18983
rect 5498 18915 5578 18927
rect 6316 18983 6396 18995
rect 6316 18927 6328 18983
rect 6384 18927 6396 18983
rect 6316 18915 6396 18927
rect 8054 18982 8134 18994
rect 8054 18926 8066 18982
rect 8122 18926 8134 18982
rect 8054 18914 8134 18926
rect 8872 18982 8952 18994
rect 8872 18926 8884 18982
rect 8940 18926 8952 18982
rect 8872 18914 8952 18926
rect 9540 18983 9620 18995
rect 9540 18927 9552 18983
rect 9608 18927 9620 18983
rect 9540 18915 9620 18927
rect 10358 18983 10438 18995
rect 10358 18927 10370 18983
rect 10426 18927 10438 18983
rect 10358 18915 10438 18927
rect 12096 18982 12176 18994
rect 12096 18926 12108 18982
rect 12164 18926 12176 18982
rect 12096 18914 12176 18926
rect 12914 18982 12994 18994
rect 12914 18926 12926 18982
rect 12982 18926 12994 18982
rect 12914 18914 12994 18926
rect 13582 18983 13662 18995
rect 13582 18927 13594 18983
rect 13650 18927 13662 18983
rect 13582 18915 13662 18927
rect 14400 18983 14480 18995
rect 14400 18927 14412 18983
rect 14468 18927 14480 18983
rect 14400 18915 14480 18927
rect 16138 18982 16218 18994
rect 16138 18926 16150 18982
rect 16206 18926 16218 18982
rect 16138 18914 16218 18926
rect 16956 18982 17036 18994
rect 16956 18926 16968 18982
rect 17024 18926 17036 18982
rect 16956 18914 17036 18926
rect 17624 18983 17704 18995
rect 17624 18927 17636 18983
rect 17692 18927 17704 18983
rect 17624 18915 17704 18927
rect 18442 18983 18522 18995
rect 18442 18927 18454 18983
rect 18510 18927 18522 18983
rect 18442 18915 18522 18927
rect -7613 18650 -7527 18654
rect -7613 18594 -7601 18650
rect -7545 18594 -7527 18650
rect -7613 18582 -7527 18594
rect -3571 18647 -3485 18651
rect -3571 18591 -3559 18647
rect -3503 18591 -3485 18647
rect -3571 18579 -3485 18591
rect 471 18647 557 18651
rect 471 18591 483 18647
rect 539 18591 557 18647
rect 471 18579 557 18591
rect 4513 18647 4599 18651
rect 4513 18591 4525 18647
rect 4581 18591 4599 18647
rect 4513 18579 4599 18591
rect 8555 18647 8641 18651
rect 8555 18591 8567 18647
rect 8623 18591 8641 18647
rect 8555 18579 8641 18591
rect 12597 18647 12683 18651
rect 12597 18591 12609 18647
rect 12665 18591 12683 18647
rect 12597 18579 12683 18591
rect 16639 18647 16725 18651
rect 16639 18591 16651 18647
rect 16707 18591 16725 18647
rect 16639 18579 16725 18591
rect 15375 17446 15453 17458
rect 15375 17390 15386 17446
rect 15442 17390 15453 17446
rect 15375 17378 15453 17390
rect -8114 16780 -8034 16792
rect -8114 16724 -8102 16780
rect -8046 16724 -8034 16780
rect -8114 16712 -8034 16724
rect -7296 16780 -7216 16792
rect -7296 16724 -7284 16780
rect -7228 16724 -7216 16780
rect -7296 16712 -7216 16724
rect -4072 16777 -3992 16789
rect -4072 16721 -4060 16777
rect -4004 16721 -3992 16777
rect -4072 16709 -3992 16721
rect -3254 16777 -3174 16789
rect -3254 16721 -3242 16777
rect -3186 16721 -3174 16777
rect -3254 16709 -3174 16721
rect -30 16777 50 16789
rect -30 16721 -18 16777
rect 38 16721 50 16777
rect -30 16709 50 16721
rect 788 16777 868 16789
rect 788 16721 800 16777
rect 856 16721 868 16777
rect 788 16709 868 16721
rect 4012 16777 4092 16789
rect 4012 16721 4024 16777
rect 4080 16721 4092 16777
rect 4012 16709 4092 16721
rect 4830 16777 4910 16789
rect 4830 16721 4842 16777
rect 4898 16721 4910 16777
rect 4830 16709 4910 16721
rect 8054 16777 8134 16789
rect 8054 16721 8066 16777
rect 8122 16721 8134 16777
rect 8054 16709 8134 16721
rect 8872 16777 8952 16789
rect 8872 16721 8884 16777
rect 8940 16721 8952 16777
rect 8872 16709 8952 16721
rect 12096 16777 12176 16789
rect 12096 16721 12108 16777
rect 12164 16721 12176 16777
rect 12096 16709 12176 16721
rect 12914 16777 12994 16789
rect 12914 16721 12926 16777
rect 12982 16721 12994 16777
rect 12914 16709 12994 16721
rect 16138 16777 16218 16789
rect 16138 16721 16150 16777
rect 16206 16721 16218 16777
rect 16138 16709 16218 16721
rect 16956 16777 17036 16789
rect 16956 16721 16968 16777
rect 17024 16721 17036 16777
rect 16956 16709 17036 16721
rect -12843 16399 -12833 16499
rect -12777 16399 -9501 16499
rect -9445 16399 -5489 16499
rect -5433 16399 -1447 16499
rect -1391 16399 2595 16499
rect 2651 16399 6637 16499
rect 6693 16399 10679 16499
rect 10735 16399 10745 16499
rect -8967 15989 -8957 15992
rect -12843 15889 -12833 15989
rect -12777 15892 -8957 15989
rect -8901 15989 -8891 15992
rect -8901 15892 -4945 15989
rect -12777 15889 -4945 15892
rect -4889 15889 -903 15989
rect -847 15889 3139 15989
rect 3195 15889 7181 15989
rect 7237 15889 11223 15989
rect 11279 15889 15265 15989
rect 15321 15889 15331 15989
rect -11625 15686 -11539 15690
rect -11625 15630 -11613 15686
rect -11557 15630 -11539 15686
rect -11625 15618 -11539 15630
rect -7613 15686 -7527 15690
rect -7613 15630 -7601 15686
rect -7545 15630 -7527 15686
rect -7613 15618 -7527 15630
rect -3571 15686 -3485 15690
rect -3571 15630 -3559 15686
rect -3503 15630 -3485 15686
rect -3571 15618 -3485 15630
rect 471 15686 557 15690
rect 471 15630 483 15686
rect 539 15630 557 15686
rect 471 15618 557 15630
rect 4513 15686 4599 15690
rect 4513 15630 4525 15686
rect 4581 15630 4599 15686
rect 4513 15618 4599 15630
rect 8555 15686 8641 15690
rect 8555 15630 8567 15686
rect 8623 15630 8641 15686
rect 8555 15618 8641 15630
rect 12597 15686 12683 15690
rect 12597 15630 12609 15686
rect 12665 15630 12683 15686
rect 12597 15618 12683 15630
rect -8777 14717 -8691 14729
rect -8777 14661 -8765 14717
rect -8709 14661 -8691 14717
rect -8777 14649 -8691 14661
rect -4735 14717 -4649 14729
rect -4735 14661 -4723 14717
rect -4667 14661 -4649 14717
rect -4735 14649 -4649 14661
rect -693 14717 -607 14729
rect -693 14661 -681 14717
rect -625 14661 -607 14717
rect -693 14649 -607 14661
rect 3349 14717 3435 14729
rect 3349 14661 3361 14717
rect 3417 14661 3435 14717
rect 3349 14649 3435 14661
rect 7391 14717 7477 14729
rect 7391 14661 7403 14717
rect 7459 14661 7477 14717
rect 7391 14649 7477 14661
rect 11433 14717 11519 14729
rect 11433 14661 11445 14717
rect 11501 14661 11519 14717
rect 11433 14649 11519 14661
rect -12126 13816 -12046 13828
rect -12126 13760 -12114 13816
rect -12058 13760 -12046 13816
rect -12126 13748 -12046 13760
rect -11308 13816 -11228 13828
rect -11308 13760 -11296 13816
rect -11240 13760 -11228 13816
rect -11308 13748 -11228 13760
rect -8114 13816 -8034 13828
rect -8114 13760 -8102 13816
rect -8046 13760 -8034 13816
rect -8114 13748 -8034 13760
rect -7296 13816 -7216 13828
rect -7296 13760 -7284 13816
rect -7228 13760 -7216 13816
rect -7296 13748 -7216 13760
rect -4072 13816 -3992 13828
rect -4072 13760 -4060 13816
rect -4004 13760 -3992 13816
rect -4072 13748 -3992 13760
rect -3254 13816 -3174 13828
rect -3254 13760 -3242 13816
rect -3186 13760 -3174 13816
rect -3254 13748 -3174 13760
rect -30 13816 50 13828
rect -30 13760 -18 13816
rect 38 13760 50 13816
rect -30 13748 50 13760
rect 788 13816 868 13828
rect 788 13760 800 13816
rect 856 13760 868 13816
rect 788 13748 868 13760
rect 4012 13816 4092 13828
rect 4012 13760 4024 13816
rect 4080 13760 4092 13816
rect 4012 13748 4092 13760
rect 4830 13816 4910 13828
rect 4830 13760 4842 13816
rect 4898 13760 4910 13816
rect 4830 13748 4910 13760
rect 8054 13816 8134 13828
rect 8054 13760 8066 13816
rect 8122 13760 8134 13816
rect 8054 13748 8134 13760
rect 8872 13816 8952 13828
rect 8872 13760 8884 13816
rect 8940 13760 8952 13816
rect 8872 13748 8952 13760
rect 12096 13816 12176 13828
rect 12096 13760 12108 13816
rect 12164 13760 12176 13816
rect 12096 13748 12176 13760
rect 12914 13816 12994 13828
rect 12914 13760 12926 13816
rect 12982 13760 12994 13816
rect 12914 13748 12994 13760
rect -11625 13481 -11539 13485
rect -11625 13425 -11613 13481
rect -11557 13425 -11539 13481
rect -11625 13413 -11539 13425
rect -10139 13481 -10053 13485
rect -10139 13425 -10127 13481
rect -10071 13425 -10053 13481
rect -10139 13413 -10053 13425
rect -7613 13481 -7527 13485
rect -7613 13425 -7601 13481
rect -7545 13425 -7527 13481
rect -7613 13413 -7527 13425
rect -6127 13481 -6041 13485
rect -6127 13425 -6115 13481
rect -6059 13425 -6041 13481
rect -6127 13413 -6041 13425
rect -3571 13481 -3485 13485
rect -3571 13425 -3559 13481
rect -3503 13425 -3485 13481
rect -3571 13413 -3485 13425
rect -2085 13481 -1999 13485
rect -2085 13425 -2073 13481
rect -2017 13425 -1999 13481
rect -2085 13413 -1999 13425
rect 471 13481 557 13485
rect 471 13425 483 13481
rect 539 13425 557 13481
rect 471 13413 557 13425
rect 1957 13481 2043 13485
rect 1957 13425 1969 13481
rect 2025 13425 2043 13481
rect 1957 13413 2043 13425
rect 4513 13481 4599 13485
rect 4513 13425 4525 13481
rect 4581 13425 4599 13481
rect 4513 13413 4599 13425
rect 5999 13481 6085 13485
rect 5999 13425 6011 13481
rect 6067 13425 6085 13481
rect 5999 13413 6085 13425
rect 8555 13481 8641 13485
rect 8555 13425 8567 13481
rect 8623 13425 8641 13481
rect 8555 13413 8641 13425
rect 10041 13481 10127 13485
rect 10041 13425 10053 13481
rect 10109 13425 10127 13481
rect 10041 13413 10127 13425
rect 12597 13481 12683 13485
rect 12597 13425 12609 13481
rect 12665 13425 12683 13481
rect 12597 13413 12683 13425
rect 14083 13481 14169 13485
rect 14083 13425 14095 13481
rect 14151 13425 14169 13481
rect 14083 13413 14169 13425
rect -12126 11611 -12046 11623
rect -12126 11555 -12114 11611
rect -12058 11555 -12046 11611
rect -12126 11543 -12046 11555
rect -11308 11611 -11228 11623
rect -11308 11555 -11296 11611
rect -11240 11555 -11228 11611
rect -11308 11543 -11228 11555
rect -10640 11611 -10560 11623
rect -10640 11555 -10628 11611
rect -10572 11555 -10560 11611
rect -10640 11543 -10560 11555
rect -9822 11611 -9742 11623
rect -9822 11555 -9810 11611
rect -9754 11555 -9742 11611
rect -9822 11543 -9742 11555
rect -8114 11611 -8034 11623
rect -8114 11555 -8102 11611
rect -8046 11555 -8034 11611
rect -8114 11543 -8034 11555
rect -7296 11611 -7216 11623
rect -7296 11555 -7284 11611
rect -7228 11555 -7216 11611
rect -7296 11543 -7216 11555
rect -6628 11611 -6548 11623
rect -6628 11555 -6616 11611
rect -6560 11555 -6548 11611
rect -6628 11543 -6548 11555
rect -5810 11611 -5730 11623
rect -5810 11555 -5798 11611
rect -5742 11555 -5730 11611
rect -5810 11543 -5730 11555
rect -4072 11611 -3992 11623
rect -4072 11555 -4060 11611
rect -4004 11555 -3992 11611
rect -4072 11543 -3992 11555
rect -3254 11611 -3174 11623
rect -3254 11555 -3242 11611
rect -3186 11555 -3174 11611
rect -3254 11543 -3174 11555
rect -2586 11611 -2506 11623
rect -2586 11555 -2574 11611
rect -2518 11555 -2506 11611
rect -2586 11543 -2506 11555
rect -1768 11611 -1688 11623
rect -1768 11555 -1756 11611
rect -1700 11555 -1688 11611
rect -1768 11543 -1688 11555
rect -30 11611 50 11623
rect -30 11555 -18 11611
rect 38 11555 50 11611
rect -30 11543 50 11555
rect 788 11611 868 11623
rect 788 11555 800 11611
rect 856 11555 868 11611
rect 788 11543 868 11555
rect 1456 11611 1536 11623
rect 1456 11555 1468 11611
rect 1524 11555 1536 11611
rect 1456 11543 1536 11555
rect 2274 11611 2354 11623
rect 2274 11555 2286 11611
rect 2342 11555 2354 11611
rect 2274 11543 2354 11555
rect 4012 11611 4092 11623
rect 4012 11555 4024 11611
rect 4080 11555 4092 11611
rect 4012 11543 4092 11555
rect 4830 11611 4910 11623
rect 4830 11555 4842 11611
rect 4898 11555 4910 11611
rect 4830 11543 4910 11555
rect 5498 11611 5578 11623
rect 5498 11555 5510 11611
rect 5566 11555 5578 11611
rect 5498 11543 5578 11555
rect 6316 11611 6396 11623
rect 6316 11555 6328 11611
rect 6384 11555 6396 11611
rect 6316 11543 6396 11555
rect 8054 11611 8134 11623
rect 8054 11555 8066 11611
rect 8122 11555 8134 11611
rect 8054 11543 8134 11555
rect 8872 11611 8952 11623
rect 8872 11555 8884 11611
rect 8940 11555 8952 11611
rect 8872 11543 8952 11555
rect 9540 11611 9620 11623
rect 9540 11555 9552 11611
rect 9608 11555 9620 11611
rect 9540 11543 9620 11555
rect 10358 11611 10438 11623
rect 10358 11555 10370 11611
rect 10426 11555 10438 11611
rect 10358 11543 10438 11555
rect 12096 11611 12176 11623
rect 12096 11555 12108 11611
rect 12164 11555 12176 11611
rect 12096 11543 12176 11555
rect 12914 11611 12994 11623
rect 12914 11555 12926 11611
rect 12982 11555 12994 11611
rect 12914 11543 12994 11555
rect 13582 11611 13662 11623
rect 13582 11555 13594 11611
rect 13650 11555 13662 11611
rect 13582 11543 13662 11555
rect 14400 11611 14480 11623
rect 14400 11555 14412 11611
rect 14468 11555 14480 11611
rect 14400 11543 14480 11555
rect -11625 11276 -11539 11280
rect -11625 11220 -11613 11276
rect -11557 11220 -11539 11276
rect -11625 11208 -11539 11220
rect -10139 11277 -10053 11281
rect -10139 11221 -10127 11277
rect -10071 11221 -10053 11277
rect -10139 11209 -10053 11221
rect -7613 11276 -7527 11280
rect -7613 11220 -7601 11276
rect -7545 11220 -7527 11276
rect -7613 11208 -7527 11220
rect -6127 11277 -6041 11281
rect -6127 11221 -6115 11277
rect -6059 11221 -6041 11277
rect -6127 11209 -6041 11221
rect -3571 11276 -3485 11280
rect -3571 11220 -3559 11276
rect -3503 11220 -3485 11276
rect -3571 11208 -3485 11220
rect -2085 11277 -1999 11281
rect -2085 11221 -2073 11277
rect -2017 11221 -1999 11277
rect -2085 11209 -1999 11221
rect 471 11276 557 11280
rect 471 11220 483 11276
rect 539 11220 557 11276
rect 471 11208 557 11220
rect 1957 11277 2043 11281
rect 1957 11221 1969 11277
rect 2025 11221 2043 11277
rect 1957 11209 2043 11221
rect 4513 11276 4599 11280
rect 4513 11220 4525 11276
rect 4581 11220 4599 11276
rect 4513 11208 4599 11220
rect 5999 11277 6085 11281
rect 5999 11221 6011 11277
rect 6067 11221 6085 11277
rect 5999 11209 6085 11221
rect 8555 11276 8641 11280
rect 8555 11220 8567 11276
rect 8623 11220 8641 11276
rect 8555 11208 8641 11220
rect 10041 11277 10127 11281
rect 10041 11221 10053 11277
rect 10109 11221 10127 11277
rect 10041 11209 10127 11221
rect 12597 11276 12683 11280
rect 12597 11220 12609 11276
rect 12665 11220 12683 11276
rect 12597 11208 12683 11220
rect 14083 11277 14169 11281
rect 14083 11221 14095 11277
rect 14151 11221 14169 11277
rect 14083 11209 14169 11221
rect -12126 9406 -12046 9418
rect -12126 9350 -12114 9406
rect -12058 9350 -12046 9406
rect -12126 9338 -12046 9350
rect -11308 9406 -11228 9418
rect -11308 9350 -11296 9406
rect -11240 9350 -11228 9406
rect -11308 9338 -11228 9350
rect -10640 9407 -10560 9419
rect -10640 9351 -10628 9407
rect -10572 9351 -10560 9407
rect -10640 9339 -10560 9351
rect -9822 9407 -9742 9419
rect -9822 9351 -9810 9407
rect -9754 9351 -9742 9407
rect -9822 9339 -9742 9351
rect -8114 9406 -8034 9418
rect -8114 9350 -8102 9406
rect -8046 9350 -8034 9406
rect -8114 9338 -8034 9350
rect -7296 9406 -7216 9418
rect -7296 9350 -7284 9406
rect -7228 9350 -7216 9406
rect -7296 9338 -7216 9350
rect -6628 9407 -6548 9419
rect -6628 9351 -6616 9407
rect -6560 9351 -6548 9407
rect -6628 9339 -6548 9351
rect -5810 9407 -5730 9419
rect -5810 9351 -5798 9407
rect -5742 9351 -5730 9407
rect -5810 9339 -5730 9351
rect -4072 9406 -3992 9418
rect -4072 9350 -4060 9406
rect -4004 9350 -3992 9406
rect -4072 9338 -3992 9350
rect -3254 9406 -3174 9418
rect -3254 9350 -3242 9406
rect -3186 9350 -3174 9406
rect -3254 9338 -3174 9350
rect -2586 9407 -2506 9419
rect -2586 9351 -2574 9407
rect -2518 9351 -2506 9407
rect -2586 9339 -2506 9351
rect -1768 9407 -1688 9419
rect -1768 9351 -1756 9407
rect -1700 9351 -1688 9407
rect -1768 9339 -1688 9351
rect -30 9406 50 9418
rect -30 9350 -18 9406
rect 38 9350 50 9406
rect -30 9338 50 9350
rect 788 9406 868 9418
rect 788 9350 800 9406
rect 856 9350 868 9406
rect 788 9338 868 9350
rect 1456 9407 1536 9419
rect 1456 9351 1468 9407
rect 1524 9351 1536 9407
rect 1456 9339 1536 9351
rect 2274 9407 2354 9419
rect 2274 9351 2286 9407
rect 2342 9351 2354 9407
rect 2274 9339 2354 9351
rect 4012 9406 4092 9418
rect 4012 9350 4024 9406
rect 4080 9350 4092 9406
rect 4012 9338 4092 9350
rect 4830 9406 4910 9418
rect 4830 9350 4842 9406
rect 4898 9350 4910 9406
rect 4830 9338 4910 9350
rect 5498 9407 5578 9419
rect 5498 9351 5510 9407
rect 5566 9351 5578 9407
rect 5498 9339 5578 9351
rect 6316 9407 6396 9419
rect 6316 9351 6328 9407
rect 6384 9351 6396 9407
rect 6316 9339 6396 9351
rect 8054 9406 8134 9418
rect 8054 9350 8066 9406
rect 8122 9350 8134 9406
rect 8054 9338 8134 9350
rect 8872 9406 8952 9418
rect 8872 9350 8884 9406
rect 8940 9350 8952 9406
rect 8872 9338 8952 9350
rect 9540 9407 9620 9419
rect 9540 9351 9552 9407
rect 9608 9351 9620 9407
rect 9540 9339 9620 9351
rect 10358 9407 10438 9419
rect 10358 9351 10370 9407
rect 10426 9351 10438 9407
rect 10358 9339 10438 9351
rect 12096 9406 12176 9418
rect 12096 9350 12108 9406
rect 12164 9350 12176 9406
rect 12096 9338 12176 9350
rect 12914 9406 12994 9418
rect 12914 9350 12926 9406
rect 12982 9350 12994 9406
rect 12914 9338 12994 9350
rect 13582 9407 13662 9419
rect 13582 9351 13594 9407
rect 13650 9351 13662 9407
rect 13582 9339 13662 9351
rect 14400 9407 14480 9419
rect 14400 9351 14412 9407
rect 14468 9351 14480 9407
rect 14400 9339 14480 9351
rect -11625 9071 -11539 9075
rect -11625 9015 -11613 9071
rect -11557 9015 -11539 9071
rect -11625 9003 -11539 9015
rect -7613 9071 -7527 9075
rect -7613 9015 -7601 9071
rect -7545 9015 -7527 9071
rect -7613 9003 -7527 9015
rect -3571 9071 -3485 9075
rect -3571 9015 -3559 9071
rect -3503 9015 -3485 9071
rect -3571 9003 -3485 9015
rect 471 9071 557 9075
rect 471 9015 483 9071
rect 539 9015 557 9071
rect 471 9003 557 9015
rect 4513 9071 4599 9075
rect 4513 9015 4525 9071
rect 4581 9015 4599 9071
rect 4513 9003 4599 9015
rect 8555 9071 8641 9075
rect 8555 9015 8567 9071
rect 8623 9015 8641 9071
rect 8555 9003 8641 9015
rect 12597 9071 12683 9075
rect 12597 9015 12609 9071
rect 12665 9015 12683 9071
rect 12597 9003 12683 9015
rect -12908 7870 -12828 7882
rect -12908 7814 -12896 7870
rect -12840 7814 -12828 7870
rect -12908 7802 -12828 7814
rect -12126 7201 -12046 7213
rect -12126 7145 -12114 7201
rect -12058 7145 -12046 7201
rect -12126 7133 -12046 7145
rect -11308 7201 -11228 7213
rect -11308 7145 -11296 7201
rect -11240 7145 -11228 7201
rect -11308 7133 -11228 7145
rect -8114 7201 -8034 7213
rect -8114 7145 -8102 7201
rect -8046 7145 -8034 7201
rect -8114 7133 -8034 7145
rect -7296 7201 -7216 7213
rect -7296 7145 -7284 7201
rect -7228 7145 -7216 7201
rect -7296 7133 -7216 7145
rect -4072 7201 -3992 7213
rect -4072 7145 -4060 7201
rect -4004 7145 -3992 7201
rect -4072 7133 -3992 7145
rect -3254 7201 -3174 7213
rect -3254 7145 -3242 7201
rect -3186 7145 -3174 7201
rect -3254 7133 -3174 7145
rect -30 7201 50 7213
rect -30 7145 -18 7201
rect 38 7145 50 7201
rect -30 7133 50 7145
rect 788 7201 868 7213
rect 788 7145 800 7201
rect 856 7145 868 7201
rect 788 7133 868 7145
rect 4012 7201 4092 7213
rect 4012 7145 4024 7201
rect 4080 7145 4092 7201
rect 4012 7133 4092 7145
rect 4830 7201 4910 7213
rect 4830 7145 4842 7201
rect 4898 7145 4910 7201
rect 4830 7133 4910 7145
rect 8054 7201 8134 7213
rect 8054 7145 8066 7201
rect 8122 7145 8134 7201
rect 8054 7133 8134 7145
rect 8872 7201 8952 7213
rect 8872 7145 8884 7201
rect 8940 7145 8952 7201
rect 8872 7133 8952 7145
rect 12096 7201 12176 7213
rect 12096 7145 12108 7201
rect 12164 7145 12176 7201
rect 12096 7133 12176 7145
rect 12914 7201 12994 7213
rect 12914 7145 12926 7201
rect 12982 7145 12994 7201
rect 12914 7133 12994 7145
rect -12908 7083 -12822 7095
rect -12908 7027 -12896 7083
rect -12840 7027 -12822 7083
rect -12908 7015 -12822 7027
rect -13115 6820 -13105 6920
rect -13049 6820 -9093 6920
rect -9037 6820 -5081 6920
rect -5025 6820 -1039 6920
rect -983 6820 3003 6920
rect 3059 6820 7045 6920
rect 7101 6820 11087 6920
rect 11143 6820 11153 6920
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -5696 2887 -5576 2907
rect -5696 2807 -5676 2887
rect -5596 2807 -5576 2887
rect -5696 2787 -5576 2807
rect -12096 2397 -11996 2417
rect -12096 2317 -12086 2397
rect -12006 2317 -11996 2397
rect -12096 2307 -11996 2317
rect -12086 2123 -12006 2307
rect -11051 2123 -10951 2133
rect -10729 2123 -10629 2133
rect -10191 2123 -10091 2133
rect -9869 2123 -9769 2133
rect -9427 2123 -9327 2133
rect -8211 2123 -8111 2243
rect -5676 2133 -5596 2787
rect -7603 2123 -7503 2133
rect -6995 2123 -6895 2133
rect -6553 2123 -6453 2133
rect -6231 2123 -6131 2133
rect -5693 2123 -5593 2133
rect -5371 2123 -5271 2133
rect -12086 2043 -11041 2123
rect -10961 2043 -10719 2123
rect -10639 2043 -10181 2123
rect -10101 2043 -9859 2123
rect -9779 2043 -9417 2123
rect -9337 2043 -8809 2123
rect -8729 2043 -8201 2123
rect -8121 2043 -7593 2123
rect -7513 2043 -6985 2123
rect -6905 2043 -6543 2123
rect -6463 2043 -6221 2123
rect -6141 2043 -5683 2123
rect -5603 2043 -5361 2123
rect -5281 2043 -5271 2123
rect -11051 2033 -10951 2043
rect -10729 2033 -10629 2043
rect -10191 2033 -10091 2043
rect -9869 2033 -9769 2043
rect -9427 2033 -9327 2043
rect -8819 2033 -8719 2043
rect -8211 2033 -8111 2043
rect -7603 2033 -7503 2043
rect -6995 2033 -6895 2043
rect -6553 2033 -6453 2043
rect -6231 2033 -6131 2043
rect -5693 2033 -5593 2043
rect -5371 2033 -5271 2043
rect -9113 1576 -9033 1586
rect -9113 1520 -9101 1576
rect -9045 1520 -9033 1576
rect -9113 1510 -9033 1520
rect -8505 1576 -8425 1586
rect -7289 1576 -7209 1586
rect -8505 1520 -8493 1576
rect -8437 1520 -7277 1576
rect -7221 1520 -7209 1576
rect -8505 1510 -8425 1520
rect -7289 1510 -7209 1520
rect -9101 1329 -9045 1510
rect -8320 1329 -8220 1339
rect -7907 1329 -7807 1339
rect -9101 1249 -8310 1329
rect -8230 1249 -7897 1329
rect -7817 1249 -7807 1329
rect -8852 865 -8752 1249
rect -8320 1239 -8220 1249
rect -7907 1239 -7807 1249
rect -8102 1159 -8002 1169
rect -8102 1079 -8092 1159
rect -8012 1079 -8002 1159
rect -8102 1031 -8002 1079
rect -8102 951 -7480 1031
rect -7560 875 -7480 951
rect -8852 785 -8842 865
rect -8762 785 -8752 865
rect -8852 775 -8752 785
rect -7570 865 -7470 875
rect -7570 785 -7560 865
rect -7480 785 -7470 865
rect -7570 775 -7470 785
rect -9721 -777 -7209 -767
rect -9721 -813 -8493 -777
rect -9721 -974 -9709 -813
rect -9653 -833 -8493 -813
rect -8437 -833 -7277 -777
rect -9653 -843 -7277 -833
rect -9653 -974 -9641 -843
rect -9721 -984 -9641 -974
rect -9113 -938 -9033 -928
rect -9714 -1408 -9649 -984
rect -9113 -994 -9101 -938
rect -9045 -994 -9033 -938
rect -9266 -1226 -9186 -1216
rect -9266 -1282 -9254 -1226
rect -9198 -1282 -9186 -1226
rect -9266 -1292 -9186 -1282
rect -9113 -1292 -9033 -994
rect -7289 -1022 -7277 -843
rect -7221 -1022 -7209 -777
rect -6681 -813 -6601 -803
rect -6681 -974 -6669 -813
rect -6613 -974 -6601 -813
rect -6681 -984 -6601 -974
rect -8971 -1070 -8871 -1058
rect -8971 -1126 -8949 -1070
rect -8893 -1126 -8871 -1070
rect -8971 -1138 -8871 -1126
rect -7756 -1070 -7656 -1058
rect -7756 -1126 -7734 -1070
rect -7678 -1126 -7656 -1070
rect -7756 -1138 -7656 -1126
rect -8051 -1226 -7971 -1216
rect -8051 -1282 -8039 -1226
rect -7983 -1282 -7971 -1226
rect -8051 -1292 -7971 -1282
rect -7289 -1292 -7209 -1022
rect -9113 -1352 -8425 -1292
rect -9714 -1468 -9033 -1408
rect -9276 -1630 -9176 -1618
rect -9276 -1686 -9254 -1630
rect -9198 -1686 -9176 -1630
rect -9276 -1698 -9176 -1686
rect -9113 -1766 -9033 -1468
rect -8961 -1474 -8881 -1464
rect -8961 -1530 -8949 -1474
rect -8893 -1530 -8881 -1474
rect -8961 -1540 -8881 -1530
rect -9113 -1822 -9101 -1766
rect -9045 -1822 -9033 -1766
rect -9113 -1832 -9033 -1822
rect -8505 -1732 -8425 -1352
rect -7897 -1352 -7209 -1292
rect -8061 -1630 -7961 -1618
rect -8061 -1686 -8039 -1630
rect -7983 -1686 -7961 -1630
rect -8061 -1698 -7961 -1686
rect -8505 -1911 -8493 -1732
rect -9721 -1921 -8493 -1911
rect -9721 -1977 -9709 -1921
rect -9653 -1977 -8493 -1921
rect -8437 -1911 -8425 -1732
rect -7897 -1766 -7817 -1352
rect -6674 -1408 -6609 -984
rect -7746 -1474 -7666 -1464
rect -7746 -1530 -7734 -1474
rect -7678 -1530 -7666 -1474
rect -7746 -1540 -7666 -1530
rect -7289 -1468 -6609 -1408
rect -7897 -1822 -7885 -1766
rect -7829 -1822 -7817 -1766
rect -7897 -1832 -7817 -1822
rect -7289 -1732 -7209 -1468
rect -7289 -1911 -7277 -1732
rect -8437 -1977 -7277 -1911
rect -7221 -1977 -7209 -1732
rect -9721 -1987 -7209 -1977
rect -6985 -1732 -6905 -1722
rect -6985 -1977 -6973 -1732
rect -6917 -1977 -6905 -1732
rect -6985 -2239 -6905 -1977
rect -6995 -2250 -6895 -2239
rect -6995 -2306 -6985 -2250
rect -6905 -2306 -6895 -2250
rect -6995 -2316 -6895 -2306
rect -4464 -3363 -2407 -3321
rect -4464 -3663 -4454 -3363
rect -2454 -3663 -2407 -3363
rect -4464 -3701 -2407 -3663
<< via3 >>
rect 40739 39093 40957 39167
rect 40737 37749 40955 37823
rect -4343 37511 -4287 37567
rect 5129 37511 5185 37567
rect 14601 37512 14657 37568
rect 24073 37512 24129 37568
rect 33545 37512 33601 37568
rect 43017 37512 43073 37568
rect -5507 36542 -5451 36598
rect 3965 36542 4021 36598
rect 13437 36543 13493 36599
rect 22909 36543 22965 36599
rect 32381 36543 32437 36599
rect 41853 36543 41909 36599
rect -4844 35641 -4788 35697
rect -4026 35641 -3970 35697
rect 4628 35641 4684 35697
rect 5446 35641 5502 35697
rect 14100 35642 14156 35698
rect 14918 35642 14974 35698
rect 23572 35642 23628 35698
rect 24390 35642 24446 35698
rect 33044 35642 33100 35698
rect 33862 35642 33918 35698
rect 42516 35642 42572 35698
rect 43334 35642 43390 35698
rect -4343 35306 -4287 35362
rect -2857 35306 -2801 35362
rect 5129 35306 5185 35362
rect 6615 35306 6671 35362
rect 14601 35307 14657 35363
rect 16087 35307 16143 35363
rect 24073 35307 24129 35363
rect 25559 35307 25615 35363
rect 33545 35307 33601 35363
rect 35031 35307 35087 35363
rect 43017 35307 43073 35363
rect 44503 35307 44559 35363
rect -4844 33436 -4788 33492
rect -4026 33436 -3970 33492
rect -3358 33436 -3302 33492
rect -2540 33436 -2484 33492
rect 4628 33436 4684 33492
rect 5446 33436 5502 33492
rect 6114 33436 6170 33492
rect 6932 33436 6988 33492
rect 14100 33437 14156 33493
rect 14918 33437 14974 33493
rect 15586 33437 15642 33493
rect 16404 33437 16460 33493
rect 23572 33437 23628 33493
rect 24390 33437 24446 33493
rect 25058 33437 25114 33493
rect 25876 33437 25932 33493
rect 33044 33437 33100 33493
rect 33862 33437 33918 33493
rect 34530 33437 34586 33493
rect 35348 33437 35404 33493
rect 42516 33437 42572 33493
rect 43334 33437 43390 33493
rect 44002 33437 44058 33493
rect 44820 33437 44876 33493
rect -4343 33101 -4287 33157
rect -2857 33102 -2801 33158
rect 5129 33101 5185 33157
rect 6615 33102 6671 33158
rect 14601 33102 14657 33158
rect 16087 33103 16143 33159
rect 24073 33102 24129 33158
rect 25559 33103 25615 33159
rect 33545 33102 33601 33158
rect 35031 33103 35087 33159
rect 43017 33102 43073 33158
rect 44503 33103 44559 33159
rect -6327 31169 -6027 31969
rect -4844 31231 -4788 31287
rect -4026 31231 -3970 31287
rect -3358 31232 -3302 31288
rect -2540 31232 -2484 31288
rect -1245 31169 -1045 31969
rect 3145 31169 3445 31969
rect 4628 31231 4684 31287
rect 5446 31231 5502 31287
rect 6114 31232 6170 31288
rect 6932 31232 6988 31288
rect 8227 31170 8427 31970
rect 12617 31170 12917 31970
rect 14100 31232 14156 31288
rect 14918 31232 14974 31288
rect 15586 31233 15642 31289
rect 16404 31233 16460 31289
rect 17699 31170 17899 31970
rect 22089 31170 22389 31970
rect 23572 31232 23628 31288
rect 24390 31232 24446 31288
rect 25058 31233 25114 31289
rect 25876 31233 25932 31289
rect 27171 31170 27371 31970
rect 31561 31170 31861 31970
rect 33044 31232 33100 31288
rect 33862 31232 33918 31288
rect 34530 31233 34586 31289
rect 35348 31233 35404 31289
rect 36643 31170 36843 31970
rect 41033 31170 41333 31970
rect 42516 31232 42572 31288
rect 43334 31232 43390 31288
rect 44002 31233 44058 31289
rect 44820 31233 44876 31289
rect -4343 30896 -4287 30952
rect -8755 30059 -8155 30199
rect 5129 30896 5185 30952
rect 717 30059 1317 30199
rect 14601 30897 14657 30953
rect 10189 30060 10789 30200
rect 24073 30897 24129 30953
rect 19661 30060 20261 30200
rect 33545 30897 33601 30953
rect 29133 30060 29733 30200
rect 43017 30897 43073 30953
rect 38605 30060 39205 30200
rect -4844 29026 -4788 29082
rect -4026 29026 -3970 29082
rect 4628 29026 4684 29082
rect -7695 28873 -5927 29013
rect 5446 29026 5502 29082
rect 14100 29027 14156 29083
rect 14918 29027 14974 29083
rect 23572 29027 23628 29083
rect -5610 28908 -5554 28964
rect 1777 28873 3545 29013
rect 3862 28908 3918 28964
rect 11249 28874 13017 29014
rect 24390 29027 24446 29083
rect 33044 29027 33100 29083
rect 13334 28909 13390 28965
rect 20721 28874 22489 29014
rect 33862 29027 33918 29083
rect 42516 29027 42572 29083
rect 22806 28909 22862 28965
rect 30193 28874 31961 29014
rect 43334 29027 43390 29083
rect 32278 28909 32334 28965
rect 39665 28874 41433 29014
rect 41750 28909 41806 28965
rect -6327 27889 -6027 28689
rect 3145 27889 3445 28689
rect 12617 27890 12917 28690
rect 22089 27890 22389 28690
rect 31561 27890 31861 28690
rect 41033 27890 41333 28690
rect -7601 25209 -7545 25265
rect -3559 25206 -3503 25262
rect 483 25206 539 25262
rect 4525 25206 4581 25262
rect 8567 25206 8623 25262
rect 12609 25206 12665 25262
rect 16651 25206 16707 25262
rect -8102 23339 -8046 23395
rect -7284 23339 -7228 23395
rect -4060 23336 -4004 23392
rect -3242 23336 -3186 23392
rect -18 23336 38 23392
rect 800 23336 856 23392
rect 4024 23336 4080 23392
rect 4842 23336 4898 23392
rect 8066 23336 8122 23392
rect 8884 23336 8940 23392
rect 12108 23336 12164 23392
rect 12926 23336 12982 23392
rect 16150 23336 16206 23392
rect 16968 23336 17024 23392
rect -7601 23004 -7545 23060
rect -6115 23004 -6059 23060
rect -3559 23001 -3503 23057
rect -2073 23001 -2017 23057
rect 483 23001 539 23057
rect 1969 23001 2025 23057
rect 4525 23001 4581 23057
rect 6011 23001 6067 23057
rect 8567 23001 8623 23057
rect 10053 23001 10109 23057
rect 12609 23001 12665 23057
rect 14095 23001 14151 23057
rect 16651 23001 16707 23057
rect 18137 23001 18193 23057
rect -8102 21134 -8046 21190
rect -7284 21134 -7228 21190
rect -6616 21134 -6560 21190
rect -5798 21134 -5742 21190
rect -4060 21131 -4004 21187
rect -3242 21131 -3186 21187
rect -2574 21131 -2518 21187
rect -1756 21131 -1700 21187
rect -18 21131 38 21187
rect 800 21131 856 21187
rect 1468 21131 1524 21187
rect 2286 21131 2342 21187
rect 4024 21131 4080 21187
rect 4842 21131 4898 21187
rect 5510 21131 5566 21187
rect 6328 21131 6384 21187
rect 8066 21131 8122 21187
rect 8884 21131 8940 21187
rect 9552 21131 9608 21187
rect 10370 21131 10426 21187
rect 12108 21131 12164 21187
rect 12926 21131 12982 21187
rect 13594 21131 13650 21187
rect 14412 21131 14468 21187
rect 16150 21131 16206 21187
rect 16968 21131 17024 21187
rect 17636 21131 17692 21187
rect 18454 21131 18510 21187
rect 15386 21014 15442 21070
rect -7601 20799 -7545 20855
rect -6115 20800 -6059 20856
rect -3559 20796 -3503 20852
rect -2073 20797 -2017 20853
rect 483 20796 539 20852
rect 1969 20797 2025 20853
rect 4525 20796 4581 20852
rect 6011 20797 6067 20853
rect 8567 20796 8623 20852
rect 10053 20797 10109 20853
rect 12609 20796 12665 20852
rect 14095 20797 14151 20853
rect 16651 20796 16707 20852
rect 18137 20797 18193 20853
rect -8102 18929 -8046 18985
rect -7284 18929 -7228 18985
rect -6616 18930 -6560 18986
rect -5798 18930 -5742 18986
rect -4060 18926 -4004 18982
rect -3242 18926 -3186 18982
rect -2574 18927 -2518 18983
rect -1756 18927 -1700 18983
rect -18 18926 38 18982
rect 800 18926 856 18982
rect 1468 18927 1524 18983
rect 2286 18927 2342 18983
rect 4024 18926 4080 18982
rect 4842 18926 4898 18982
rect 5510 18927 5566 18983
rect 6328 18927 6384 18983
rect 8066 18926 8122 18982
rect 8884 18926 8940 18982
rect 9552 18927 9608 18983
rect 10370 18927 10426 18983
rect 12108 18926 12164 18982
rect 12926 18926 12982 18982
rect 13594 18927 13650 18983
rect 14412 18927 14468 18983
rect 16150 18926 16206 18982
rect 16968 18926 17024 18982
rect 17636 18927 17692 18983
rect 18454 18927 18510 18983
rect -7601 18594 -7545 18650
rect -3559 18591 -3503 18647
rect 483 18591 539 18647
rect 4525 18591 4581 18647
rect 8567 18591 8623 18647
rect 12609 18591 12665 18647
rect 16651 18591 16707 18647
rect 15386 17390 15442 17446
rect -8102 16724 -8046 16780
rect -7284 16724 -7228 16780
rect -4060 16721 -4004 16777
rect -3242 16721 -3186 16777
rect -18 16721 38 16777
rect 800 16721 856 16777
rect 4024 16721 4080 16777
rect 4842 16721 4898 16777
rect 8066 16721 8122 16777
rect 8884 16721 8940 16777
rect 12108 16721 12164 16777
rect 12926 16721 12982 16777
rect 16150 16721 16206 16777
rect 16968 16721 17024 16777
rect -11613 15630 -11557 15686
rect -7601 15630 -7545 15686
rect -3559 15630 -3503 15686
rect 483 15630 539 15686
rect 4525 15630 4581 15686
rect 8567 15630 8623 15686
rect 12609 15630 12665 15686
rect -8765 14661 -8709 14717
rect -4723 14661 -4667 14717
rect -681 14661 -625 14717
rect 3361 14661 3417 14717
rect 7403 14661 7459 14717
rect 11445 14661 11501 14717
rect -12114 13760 -12058 13816
rect -11296 13760 -11240 13816
rect -8102 13760 -8046 13816
rect -7284 13760 -7228 13816
rect -4060 13760 -4004 13816
rect -3242 13760 -3186 13816
rect -18 13760 38 13816
rect 800 13760 856 13816
rect 4024 13760 4080 13816
rect 4842 13760 4898 13816
rect 8066 13760 8122 13816
rect 8884 13760 8940 13816
rect 12108 13760 12164 13816
rect 12926 13760 12982 13816
rect -11613 13425 -11557 13481
rect -10127 13425 -10071 13481
rect -7601 13425 -7545 13481
rect -6115 13425 -6059 13481
rect -3559 13425 -3503 13481
rect -2073 13425 -2017 13481
rect 483 13425 539 13481
rect 1969 13425 2025 13481
rect 4525 13425 4581 13481
rect 6011 13425 6067 13481
rect 8567 13425 8623 13481
rect 10053 13425 10109 13481
rect 12609 13425 12665 13481
rect 14095 13425 14151 13481
rect -12114 11555 -12058 11611
rect -11296 11555 -11240 11611
rect -10628 11555 -10572 11611
rect -9810 11555 -9754 11611
rect -8102 11555 -8046 11611
rect -7284 11555 -7228 11611
rect -6616 11555 -6560 11611
rect -5798 11555 -5742 11611
rect -4060 11555 -4004 11611
rect -3242 11555 -3186 11611
rect -2574 11555 -2518 11611
rect -1756 11555 -1700 11611
rect -18 11555 38 11611
rect 800 11555 856 11611
rect 1468 11555 1524 11611
rect 2286 11555 2342 11611
rect 4024 11555 4080 11611
rect 4842 11555 4898 11611
rect 5510 11555 5566 11611
rect 6328 11555 6384 11611
rect 8066 11555 8122 11611
rect 8884 11555 8940 11611
rect 9552 11555 9608 11611
rect 10370 11555 10426 11611
rect 12108 11555 12164 11611
rect 12926 11555 12982 11611
rect 13594 11555 13650 11611
rect 14412 11555 14468 11611
rect -11613 11220 -11557 11276
rect -10127 11221 -10071 11277
rect -7601 11220 -7545 11276
rect -6115 11221 -6059 11277
rect -3559 11220 -3503 11276
rect -2073 11221 -2017 11277
rect 483 11220 539 11276
rect 1969 11221 2025 11277
rect 4525 11220 4581 11276
rect 6011 11221 6067 11277
rect 8567 11220 8623 11276
rect 10053 11221 10109 11277
rect 12609 11220 12665 11276
rect 14095 11221 14151 11277
rect -12114 9350 -12058 9406
rect -11296 9350 -11240 9406
rect -10628 9351 -10572 9407
rect -9810 9351 -9754 9407
rect -8102 9350 -8046 9406
rect -7284 9350 -7228 9406
rect -6616 9351 -6560 9407
rect -5798 9351 -5742 9407
rect -4060 9350 -4004 9406
rect -3242 9350 -3186 9406
rect -2574 9351 -2518 9407
rect -1756 9351 -1700 9407
rect -18 9350 38 9406
rect 800 9350 856 9406
rect 1468 9351 1524 9407
rect 2286 9351 2342 9407
rect 4024 9350 4080 9406
rect 4842 9350 4898 9406
rect 5510 9351 5566 9407
rect 6328 9351 6384 9407
rect 8066 9350 8122 9406
rect 8884 9350 8940 9406
rect 9552 9351 9608 9407
rect 10370 9351 10426 9407
rect 12108 9350 12164 9406
rect 12926 9350 12982 9406
rect 13594 9351 13650 9407
rect 14412 9351 14468 9407
rect -11613 9015 -11557 9071
rect -7601 9015 -7545 9071
rect -3559 9015 -3503 9071
rect 483 9015 539 9071
rect 4525 9015 4581 9071
rect 8567 9015 8623 9071
rect 12609 9015 12665 9071
rect -12896 7814 -12840 7870
rect -12114 7145 -12058 7201
rect -11296 7145 -11240 7201
rect -8102 7145 -8046 7201
rect -7284 7145 -7228 7201
rect -4060 7145 -4004 7201
rect -3242 7145 -3186 7201
rect -18 7145 38 7201
rect 800 7145 856 7201
rect 4024 7145 4080 7201
rect 4842 7145 4898 7201
rect 8066 7145 8122 7201
rect 8884 7145 8940 7201
rect 12108 7145 12164 7201
rect 12926 7145 12982 7201
rect -12896 7027 -12840 7083
rect -4454 6134 -2454 6434
rect -9254 -1282 -9198 -1226
rect -8949 -1126 -8893 -1070
rect -7734 -1126 -7678 -1070
rect -8039 -1282 -7983 -1226
rect -9254 -1686 -9198 -1630
rect -8949 -1530 -8893 -1474
rect -8039 -1686 -7983 -1630
rect -7734 -1530 -7678 -1474
rect -4454 -3663 -2454 -3363
<< metal4 >>
rect 40726 39167 40972 39180
rect 40726 39093 40739 39167
rect 40957 39093 40972 39167
rect 40726 39080 40972 39093
rect 40723 37823 40967 37836
rect 40723 37749 40737 37823
rect 40955 37749 40967 37823
rect -4355 37567 -4269 37571
rect -4355 37511 -4343 37567
rect -4287 37511 -4269 37567
rect -4355 37499 -4269 37511
rect 5117 37567 5203 37571
rect 5117 37511 5129 37567
rect 5185 37511 5203 37567
rect 5117 37499 5203 37511
rect 14589 37568 14675 37572
rect 14589 37512 14601 37568
rect 14657 37512 14675 37568
rect 14589 37500 14675 37512
rect 24061 37568 24147 37572
rect 24061 37512 24073 37568
rect 24129 37512 24147 37568
rect 24061 37500 24147 37512
rect 33533 37568 33619 37572
rect 33533 37512 33545 37568
rect 33601 37512 33619 37568
rect 33533 37500 33619 37512
rect 40723 37364 40967 37749
rect 43005 37568 43091 37572
rect 43005 37512 43017 37568
rect 43073 37512 43091 37568
rect 43005 37500 43091 37512
rect -5521 36598 -5433 36610
rect -5521 36542 -5507 36598
rect -5451 36542 -5433 36598
rect -5521 36530 -5433 36542
rect -5369 35697 -2069 37363
rect 3951 36598 4039 36610
rect 3951 36542 3965 36598
rect 4021 36542 4039 36598
rect 3951 36530 4039 36542
rect -5369 35641 -4844 35697
rect -4788 35641 -4026 35697
rect -3970 35641 -2069 35697
rect -5369 35523 -2069 35641
rect -5369 35158 -4537 35523
rect -4355 35362 -4269 35366
rect -4355 35306 -4343 35362
rect -4287 35306 -4269 35362
rect -4355 35294 -4269 35306
rect -4087 35158 -3051 35523
rect -2869 35362 -2783 35366
rect -2869 35306 -2857 35362
rect -2801 35306 -2783 35362
rect -2869 35294 -2783 35306
rect -2601 35158 -2069 35523
rect -5369 33492 -2069 35158
rect -5369 33436 -4844 33492
rect -4788 33436 -4026 33492
rect -3970 33436 -3358 33492
rect -3302 33436 -2540 33492
rect -2484 33436 -2069 33492
rect -5369 33318 -2069 33436
rect -5369 32953 -4537 33318
rect -4355 33157 -4269 33161
rect -4355 33101 -4343 33157
rect -4287 33101 -4269 33157
rect -4355 33089 -4269 33101
rect -4087 32953 -3051 33318
rect -2869 33158 -2783 33162
rect -2869 33102 -2857 33158
rect -2801 33102 -2783 33158
rect -2869 33090 -2783 33102
rect -2601 32953 -2069 33318
rect -6337 31969 -6017 31979
rect -6337 31169 -6327 31969
rect -6027 31169 -6017 31969
rect -6337 31159 -6017 31169
rect -5369 31288 -2069 32953
rect 4103 35697 7403 37363
rect 13423 36599 13511 36611
rect 13423 36543 13437 36599
rect 13493 36543 13511 36599
rect 13423 36531 13511 36543
rect 4103 35641 4628 35697
rect 4684 35641 5446 35697
rect 5502 35641 7403 35697
rect 4103 35523 7403 35641
rect 4103 35158 4935 35523
rect 5117 35362 5203 35366
rect 5117 35306 5129 35362
rect 5185 35306 5203 35362
rect 5117 35294 5203 35306
rect 5385 35158 6421 35523
rect 6603 35362 6689 35366
rect 6603 35306 6615 35362
rect 6671 35306 6689 35362
rect 6603 35294 6689 35306
rect 6871 35158 7403 35523
rect 4103 33492 7403 35158
rect 4103 33436 4628 33492
rect 4684 33436 5446 33492
rect 5502 33436 6114 33492
rect 6170 33436 6932 33492
rect 6988 33436 7403 33492
rect 4103 33318 7403 33436
rect 4103 32953 4935 33318
rect 5117 33157 5203 33161
rect 5117 33101 5129 33157
rect 5185 33101 5203 33157
rect 5117 33089 5203 33101
rect 5385 32953 6421 33318
rect 6603 33158 6689 33162
rect 6603 33102 6615 33158
rect 6671 33102 6689 33158
rect 6603 33090 6689 33102
rect 6871 32953 7403 33318
rect -5369 31287 -3358 31288
rect -5369 31231 -4844 31287
rect -4788 31231 -4026 31287
rect -3970 31232 -3358 31287
rect -3302 31232 -2540 31288
rect -2484 31232 -2069 31288
rect -3970 31231 -2069 31232
rect -5369 31113 -2069 31231
rect -1255 31969 -1035 31979
rect -1255 31169 -1245 31969
rect -1045 31169 -1035 31969
rect -1255 31159 -1035 31169
rect 3135 31969 3455 31979
rect 3135 31169 3145 31969
rect 3445 31169 3455 31969
rect 3135 31159 3455 31169
rect 4103 31288 7403 32953
rect 13575 35698 16875 37364
rect 22895 36599 22983 36611
rect 22895 36543 22909 36599
rect 22965 36543 22983 36599
rect 22895 36531 22983 36543
rect 13575 35642 14100 35698
rect 14156 35642 14918 35698
rect 14974 35642 16875 35698
rect 13575 35524 16875 35642
rect 13575 35159 14407 35524
rect 14589 35363 14675 35367
rect 14589 35307 14601 35363
rect 14657 35307 14675 35363
rect 14589 35295 14675 35307
rect 14857 35159 15893 35524
rect 16075 35363 16161 35367
rect 16075 35307 16087 35363
rect 16143 35307 16161 35363
rect 16075 35295 16161 35307
rect 16343 35159 16875 35524
rect 13575 33493 16875 35159
rect 13575 33437 14100 33493
rect 14156 33437 14918 33493
rect 14974 33437 15586 33493
rect 15642 33437 16404 33493
rect 16460 33437 16875 33493
rect 13575 33319 16875 33437
rect 13575 32954 14407 33319
rect 14589 33158 14675 33162
rect 14589 33102 14601 33158
rect 14657 33102 14675 33158
rect 14589 33090 14675 33102
rect 14857 32954 15893 33319
rect 16075 33159 16161 33163
rect 16075 33103 16087 33159
rect 16143 33103 16161 33159
rect 16075 33091 16161 33103
rect 16343 32954 16875 33319
rect 4103 31287 6114 31288
rect 4103 31231 4628 31287
rect 4684 31231 5446 31287
rect 5502 31232 6114 31287
rect 6170 31232 6932 31288
rect 6988 31232 7403 31288
rect 5502 31231 7403 31232
rect -5369 30748 -4537 31113
rect -4355 30952 -4269 30956
rect -4355 30896 -4343 30952
rect -4287 30896 -4269 30952
rect -4355 30884 -4269 30896
rect -4087 30748 -2069 31113
rect -8767 30199 -5915 30211
rect -8767 30059 -8755 30199
rect -8155 30059 -5915 30199
rect -8767 30047 -5915 30059
rect -7707 29013 -5915 30047
rect -7707 28873 -7695 29013
rect -5927 28873 -5915 29013
rect -5369 29082 -2069 30748
rect 4103 31113 7403 31231
rect 8217 31970 8437 31980
rect 8217 31170 8227 31970
rect 8427 31170 8437 31970
rect 8217 31160 8437 31170
rect 12607 31970 12927 31980
rect 12607 31170 12617 31970
rect 12917 31170 12927 31970
rect 12607 31160 12927 31170
rect 13575 31289 16875 32954
rect 23047 35698 26347 37364
rect 32367 36599 32455 36611
rect 32367 36543 32381 36599
rect 32437 36543 32455 36599
rect 32367 36531 32455 36543
rect 23047 35642 23572 35698
rect 23628 35642 24390 35698
rect 24446 35642 26347 35698
rect 23047 35524 26347 35642
rect 23047 35159 23879 35524
rect 24061 35363 24147 35367
rect 24061 35307 24073 35363
rect 24129 35307 24147 35363
rect 24061 35295 24147 35307
rect 24329 35159 25365 35524
rect 25547 35363 25633 35367
rect 25547 35307 25559 35363
rect 25615 35307 25633 35363
rect 25547 35295 25633 35307
rect 25815 35159 26347 35524
rect 23047 33493 26347 35159
rect 23047 33437 23572 33493
rect 23628 33437 24390 33493
rect 24446 33437 25058 33493
rect 25114 33437 25876 33493
rect 25932 33437 26347 33493
rect 23047 33319 26347 33437
rect 23047 32954 23879 33319
rect 24061 33158 24147 33162
rect 24061 33102 24073 33158
rect 24129 33102 24147 33158
rect 24061 33090 24147 33102
rect 24329 32954 25365 33319
rect 25547 33159 25633 33163
rect 25547 33103 25559 33159
rect 25615 33103 25633 33159
rect 25547 33091 25633 33103
rect 25815 32954 26347 33319
rect 13575 31288 15586 31289
rect 13575 31232 14100 31288
rect 14156 31232 14918 31288
rect 14974 31233 15586 31288
rect 15642 31233 16404 31289
rect 16460 31233 16875 31289
rect 14974 31232 16875 31233
rect 4103 30748 4935 31113
rect 5117 30952 5203 30956
rect 5117 30896 5129 30952
rect 5185 30896 5203 30952
rect 5117 30884 5203 30896
rect 5385 30748 7403 31113
rect 705 30199 3557 30211
rect 705 30059 717 30199
rect 1317 30059 3557 30199
rect 705 30047 3557 30059
rect -5369 29026 -4844 29082
rect -4788 29026 -4026 29082
rect -3970 29026 -2069 29082
rect -5622 28964 -5536 28976
rect -5622 28908 -5610 28964
rect -5554 28908 -5536 28964
rect -5622 28896 -5536 28908
rect -5369 28896 -2069 29026
rect 1765 29013 3557 30047
rect -7707 28861 -5915 28873
rect -5369 28699 -4073 28896
rect 1765 28873 1777 29013
rect 3545 28873 3557 29013
rect 4103 29082 7403 30748
rect 13575 31114 16875 31232
rect 17689 31970 17909 31980
rect 17689 31170 17699 31970
rect 17899 31170 17909 31970
rect 17689 31160 17909 31170
rect 22079 31970 22399 31980
rect 22079 31170 22089 31970
rect 22389 31170 22399 31970
rect 22079 31160 22399 31170
rect 23047 31289 26347 32954
rect 32519 35698 35819 37364
rect 40723 36844 45291 37364
rect 41839 36599 41927 36611
rect 41839 36543 41853 36599
rect 41909 36543 41927 36599
rect 41839 36531 41927 36543
rect 32519 35642 33044 35698
rect 33100 35642 33862 35698
rect 33918 35642 35819 35698
rect 32519 35524 35819 35642
rect 32519 35159 33351 35524
rect 33533 35363 33619 35367
rect 33533 35307 33545 35363
rect 33601 35307 33619 35363
rect 33533 35295 33619 35307
rect 33801 35159 34837 35524
rect 35019 35363 35105 35367
rect 35019 35307 35031 35363
rect 35087 35307 35105 35363
rect 35019 35295 35105 35307
rect 35287 35159 35819 35524
rect 32519 33493 35819 35159
rect 32519 33437 33044 33493
rect 33100 33437 33862 33493
rect 33918 33437 34530 33493
rect 34586 33437 35348 33493
rect 35404 33437 35819 33493
rect 32519 33319 35819 33437
rect 32519 32954 33351 33319
rect 33533 33158 33619 33162
rect 33533 33102 33545 33158
rect 33601 33102 33619 33158
rect 33533 33090 33619 33102
rect 33801 32954 34837 33319
rect 35019 33159 35105 33163
rect 35019 33103 35031 33159
rect 35087 33103 35105 33159
rect 35019 33091 35105 33103
rect 35287 32954 35819 33319
rect 23047 31288 25058 31289
rect 23047 31232 23572 31288
rect 23628 31232 24390 31288
rect 24446 31233 25058 31288
rect 25114 31233 25876 31289
rect 25932 31233 26347 31289
rect 24446 31232 26347 31233
rect 13575 30749 14407 31114
rect 14589 30953 14675 30957
rect 14589 30897 14601 30953
rect 14657 30897 14675 30953
rect 14589 30885 14675 30897
rect 14857 30749 16875 31114
rect 10177 30200 13029 30212
rect 10177 30060 10189 30200
rect 10789 30060 13029 30200
rect 10177 30048 13029 30060
rect 4103 29026 4628 29082
rect 4684 29026 5446 29082
rect 5502 29026 7403 29082
rect 3850 28964 3936 28976
rect 3850 28908 3862 28964
rect 3918 28908 3936 28964
rect 3850 28896 3936 28908
rect 4103 28896 7403 29026
rect 11237 29014 13029 30048
rect 1765 28861 3557 28873
rect 4103 28699 5399 28896
rect 11237 28874 11249 29014
rect 13017 28874 13029 29014
rect 13575 29083 16875 30749
rect 23047 31114 26347 31232
rect 27161 31970 27381 31980
rect 27161 31170 27171 31970
rect 27371 31170 27381 31970
rect 27161 31160 27381 31170
rect 31551 31970 31871 31980
rect 31551 31170 31561 31970
rect 31861 31170 31871 31970
rect 31551 31160 31871 31170
rect 32519 31289 35819 32954
rect 41991 35698 45291 36844
rect 41991 35642 42516 35698
rect 42572 35642 43334 35698
rect 43390 35642 45291 35698
rect 41991 35524 45291 35642
rect 41991 35159 42823 35524
rect 43005 35363 43091 35367
rect 43005 35307 43017 35363
rect 43073 35307 43091 35363
rect 43005 35295 43091 35307
rect 43273 35159 44309 35524
rect 44491 35363 44577 35367
rect 44491 35307 44503 35363
rect 44559 35307 44577 35363
rect 44491 35295 44577 35307
rect 44759 35159 45291 35524
rect 41991 33493 45291 35159
rect 41991 33437 42516 33493
rect 42572 33437 43334 33493
rect 43390 33437 44002 33493
rect 44058 33437 44820 33493
rect 44876 33437 45291 33493
rect 41991 33319 45291 33437
rect 41991 32954 42823 33319
rect 43005 33158 43091 33162
rect 43005 33102 43017 33158
rect 43073 33102 43091 33158
rect 43005 33090 43091 33102
rect 43273 32954 44309 33319
rect 44491 33159 44577 33163
rect 44491 33103 44503 33159
rect 44559 33103 44577 33159
rect 44491 33091 44577 33103
rect 44759 32954 45291 33319
rect 32519 31288 34530 31289
rect 32519 31232 33044 31288
rect 33100 31232 33862 31288
rect 33918 31233 34530 31288
rect 34586 31233 35348 31289
rect 35404 31233 35819 31289
rect 33918 31232 35819 31233
rect 23047 30749 23879 31114
rect 24061 30953 24147 30957
rect 24061 30897 24073 30953
rect 24129 30897 24147 30953
rect 24061 30885 24147 30897
rect 24329 30749 26347 31114
rect 19649 30200 22501 30212
rect 19649 30060 19661 30200
rect 20261 30060 22501 30200
rect 19649 30048 22501 30060
rect 13575 29027 14100 29083
rect 14156 29027 14918 29083
rect 14974 29027 16875 29083
rect 13322 28965 13408 28977
rect 13322 28909 13334 28965
rect 13390 28909 13408 28965
rect 13322 28897 13408 28909
rect 13575 28897 16875 29027
rect 20709 29014 22501 30048
rect 11237 28862 13029 28874
rect 13575 28700 14871 28897
rect 20709 28874 20721 29014
rect 22489 28874 22501 29014
rect 23047 29083 26347 30749
rect 32519 31114 35819 31232
rect 36633 31970 36853 31980
rect 36633 31170 36643 31970
rect 36843 31170 36853 31970
rect 36633 31160 36853 31170
rect 41023 31970 41343 31980
rect 41023 31170 41033 31970
rect 41333 31170 41343 31970
rect 41023 31160 41343 31170
rect 41991 31289 45291 32954
rect 41991 31288 44002 31289
rect 41991 31232 42516 31288
rect 42572 31232 43334 31288
rect 43390 31233 44002 31288
rect 44058 31233 44820 31289
rect 44876 31233 45291 31289
rect 43390 31232 45291 31233
rect 32519 30749 33351 31114
rect 33533 30953 33619 30957
rect 33533 30897 33545 30953
rect 33601 30897 33619 30953
rect 33533 30885 33619 30897
rect 33801 30749 35819 31114
rect 29121 30200 31973 30212
rect 29121 30060 29133 30200
rect 29733 30060 31973 30200
rect 29121 30048 31973 30060
rect 23047 29027 23572 29083
rect 23628 29027 24390 29083
rect 24446 29027 26347 29083
rect 22794 28965 22880 28977
rect 22794 28909 22806 28965
rect 22862 28909 22880 28965
rect 22794 28897 22880 28909
rect 23047 28897 26347 29027
rect 30181 29014 31973 30048
rect 20709 28862 22501 28874
rect 23047 28700 24343 28897
rect 30181 28874 30193 29014
rect 31961 28874 31973 29014
rect 32519 29083 35819 30749
rect 41991 31114 45291 31232
rect 41991 30749 42823 31114
rect 43005 30953 43091 30957
rect 43005 30897 43017 30953
rect 43073 30897 43091 30953
rect 43005 30885 43091 30897
rect 43273 30749 45291 31114
rect 38593 30200 41445 30212
rect 38593 30060 38605 30200
rect 39205 30060 41445 30200
rect 38593 30048 41445 30060
rect 32519 29027 33044 29083
rect 33100 29027 33862 29083
rect 33918 29027 35819 29083
rect 32266 28965 32352 28977
rect 32266 28909 32278 28965
rect 32334 28909 32352 28965
rect 32266 28897 32352 28909
rect 30181 28862 31973 28874
rect 32519 28700 35819 29027
rect 39653 29014 41445 30048
rect 39653 28874 39665 29014
rect 41433 28874 41445 29014
rect 41991 29083 45291 30749
rect 41991 29027 42516 29083
rect 42572 29027 43334 29083
rect 43390 29027 45291 29083
rect 41738 28965 41824 28977
rect 41738 28909 41750 28965
rect 41806 28909 41824 28965
rect 41738 28897 41824 28909
rect 41991 28897 45291 29027
rect 39653 28862 41445 28874
rect 41991 28700 43287 28897
rect -6337 28689 -4073 28699
rect -6337 27889 -6327 28689
rect -6027 27889 -4073 28689
rect -6337 27880 -4073 27889
rect 3135 28689 5399 28699
rect 3135 27889 3145 28689
rect 3445 27889 5399 28689
rect 3135 27880 5399 27889
rect 12607 28690 14871 28700
rect 12607 27890 12617 28690
rect 12917 27890 14871 28690
rect 12607 27880 14871 27890
rect 22079 28690 24343 28700
rect 22079 27890 22089 28690
rect 22389 27890 24343 28690
rect 22079 27880 24343 27890
rect 31551 28690 35819 28700
rect 31551 27890 31561 28690
rect 31861 27890 35819 28690
rect 31551 27880 35819 27890
rect 41023 28690 43287 28700
rect 41023 27890 41033 28690
rect 41333 27890 43287 28690
rect 41023 27880 43287 27890
rect -8627 25373 24343 27880
rect 32519 26106 35819 27880
rect 41533 26106 43287 27880
rect -5327 25370 18925 25373
rect -7613 25265 -7527 25269
rect -7613 25209 -7601 25265
rect -7545 25209 -7527 25265
rect -7613 25197 -7527 25209
rect -5327 25061 -4585 25370
rect -3571 25262 -3485 25266
rect -3571 25206 -3559 25262
rect -3503 25206 -3485 25262
rect -3571 25194 -3485 25206
rect -8627 25058 -4585 25061
rect -1285 25058 -543 25370
rect 471 25262 557 25266
rect 471 25206 483 25262
rect 539 25206 557 25262
rect 471 25194 557 25206
rect 2757 25058 3499 25370
rect 4513 25262 4599 25266
rect 4513 25206 4525 25262
rect 4581 25206 4599 25262
rect 4513 25194 4599 25206
rect 6799 25058 7541 25370
rect 8555 25262 8641 25266
rect 8555 25206 8567 25262
rect 8623 25206 8641 25262
rect 8555 25194 8641 25206
rect 10841 25058 11583 25370
rect 12597 25262 12683 25266
rect 12597 25206 12609 25262
rect 12665 25206 12683 25262
rect 12597 25194 12683 25206
rect 14883 25058 15625 25370
rect 16639 25262 16725 25266
rect 16639 25206 16651 25262
rect 16707 25206 16725 25262
rect 16639 25194 16725 25206
rect -8627 23395 18925 25058
rect -8627 23339 -8102 23395
rect -8046 23339 -7284 23395
rect -7228 23392 18925 23395
rect -7228 23339 -4060 23392
rect -8627 23336 -4060 23339
rect -4004 23336 -3242 23392
rect -3186 23336 -18 23392
rect 38 23336 800 23392
rect 856 23336 4024 23392
rect 4080 23336 4842 23392
rect 4898 23336 8066 23392
rect 8122 23336 8884 23392
rect 8940 23336 12108 23392
rect 12164 23336 12926 23392
rect 12982 23336 16150 23392
rect 16206 23336 16968 23392
rect 17024 23336 18925 23392
rect -8627 23221 18925 23336
rect -8627 22856 -7795 23221
rect -7613 23060 -7527 23064
rect -7613 23004 -7601 23060
rect -7545 23004 -7527 23060
rect -7613 22992 -7527 23004
rect -7345 22856 -6309 23221
rect -5859 23218 18925 23221
rect -6127 23060 -6041 23064
rect -6127 23004 -6115 23060
rect -6059 23004 -6041 23060
rect -6127 22992 -6041 23004
rect -5859 22856 -3753 23218
rect -3571 23057 -3485 23061
rect -3571 23001 -3559 23057
rect -3503 23001 -3485 23057
rect -3571 22989 -3485 23001
rect -8627 22853 -3753 22856
rect -3303 22853 -2267 23218
rect -2085 23057 -1999 23061
rect -2085 23001 -2073 23057
rect -2017 23001 -1999 23057
rect -2085 22989 -1999 23001
rect -1817 22853 289 23218
rect 471 23057 557 23061
rect 471 23001 483 23057
rect 539 23001 557 23057
rect 471 22989 557 23001
rect 739 22853 1775 23218
rect 1957 23057 2043 23061
rect 1957 23001 1969 23057
rect 2025 23001 2043 23057
rect 1957 22989 2043 23001
rect 2225 22853 4331 23218
rect 4513 23057 4599 23061
rect 4513 23001 4525 23057
rect 4581 23001 4599 23057
rect 4513 22989 4599 23001
rect 4781 22853 5817 23218
rect 5999 23057 6085 23061
rect 5999 23001 6011 23057
rect 6067 23001 6085 23057
rect 5999 22989 6085 23001
rect 6267 22853 8373 23218
rect 8555 23057 8641 23061
rect 8555 23001 8567 23057
rect 8623 23001 8641 23057
rect 8555 22989 8641 23001
rect 8823 22853 9859 23218
rect 10041 23057 10127 23061
rect 10041 23001 10053 23057
rect 10109 23001 10127 23057
rect 10041 22989 10127 23001
rect 10309 22853 12415 23218
rect 12597 23057 12683 23061
rect 12597 23001 12609 23057
rect 12665 23001 12683 23057
rect 12597 22989 12683 23001
rect 12865 22853 13901 23218
rect 14083 23057 14169 23061
rect 14083 23001 14095 23057
rect 14151 23001 14169 23057
rect 14083 22989 14169 23001
rect 14351 22853 16457 23218
rect 16639 23057 16725 23061
rect 16639 23001 16651 23057
rect 16707 23001 16725 23057
rect 16639 22989 16725 23001
rect 16907 22853 17943 23218
rect 18125 23057 18211 23061
rect 18125 23001 18137 23057
rect 18193 23001 18211 23057
rect 18125 22989 18211 23001
rect 18393 22853 18925 23218
rect -8627 21190 18925 22853
rect -8627 21134 -8102 21190
rect -8046 21134 -7284 21190
rect -7228 21134 -6616 21190
rect -6560 21134 -5798 21190
rect -5742 21187 18925 21190
rect -5742 21134 -4060 21187
rect -8627 21131 -4060 21134
rect -4004 21131 -3242 21187
rect -3186 21131 -2574 21187
rect -2518 21131 -1756 21187
rect -1700 21131 -18 21187
rect 38 21131 800 21187
rect 856 21131 1468 21187
rect 1524 21131 2286 21187
rect 2342 21131 4024 21187
rect 4080 21131 4842 21187
rect 4898 21131 5510 21187
rect 5566 21131 6328 21187
rect 6384 21131 8066 21187
rect 8122 21131 8884 21187
rect 8940 21131 9552 21187
rect 9608 21131 10370 21187
rect 10426 21131 12108 21187
rect 12164 21131 12926 21187
rect 12982 21131 13594 21187
rect 13650 21131 14412 21187
rect 14468 21131 16150 21187
rect 16206 21131 16968 21187
rect 17024 21131 17636 21187
rect 17692 21131 18454 21187
rect 18510 21131 18925 21187
rect -8627 21070 18925 21131
rect -8627 21016 15386 21070
rect -8627 20651 -7795 21016
rect -7613 20855 -7527 20859
rect -7613 20799 -7601 20855
rect -7545 20799 -7527 20855
rect -7613 20787 -7527 20799
rect -7345 20651 -6309 21016
rect -5859 21014 15386 21016
rect 15442 21014 18925 21070
rect -5859 21013 18925 21014
rect -6127 20856 -6041 20860
rect -6127 20800 -6115 20856
rect -6059 20800 -6041 20856
rect -6127 20788 -6041 20800
rect -5859 20651 -3753 21013
rect -3571 20852 -3485 20856
rect -3571 20796 -3559 20852
rect -3503 20796 -3485 20852
rect -3571 20784 -3485 20796
rect -8627 20648 -3753 20651
rect -3303 20648 -2267 21013
rect -2085 20853 -1999 20857
rect -2085 20797 -2073 20853
rect -2017 20797 -1999 20853
rect -2085 20785 -1999 20797
rect -1817 20648 289 21013
rect 471 20852 557 20856
rect 471 20796 483 20852
rect 539 20796 557 20852
rect 471 20784 557 20796
rect 739 20648 1775 21013
rect 1957 20853 2043 20857
rect 1957 20797 1969 20853
rect 2025 20797 2043 20853
rect 1957 20785 2043 20797
rect 2225 20648 4331 21013
rect 4513 20852 4599 20856
rect 4513 20796 4525 20852
rect 4581 20796 4599 20852
rect 4513 20784 4599 20796
rect 4781 20648 5817 21013
rect 5999 20853 6085 20857
rect 5999 20797 6011 20853
rect 6067 20797 6085 20853
rect 5999 20785 6085 20797
rect 6267 20648 8373 21013
rect 8555 20852 8641 20856
rect 8555 20796 8567 20852
rect 8623 20796 8641 20852
rect 8555 20784 8641 20796
rect 8823 20648 9859 21013
rect 10041 20853 10127 20857
rect 10041 20797 10053 20853
rect 10109 20797 10127 20853
rect 10041 20785 10127 20797
rect 10309 20648 12415 21013
rect 12597 20852 12683 20856
rect 12597 20796 12609 20852
rect 12665 20796 12683 20852
rect 12597 20784 12683 20796
rect 12865 20648 13901 21013
rect 14083 20853 14169 20857
rect 14083 20797 14095 20853
rect 14151 20797 14169 20853
rect 14083 20785 14169 20797
rect 14351 20648 16457 21013
rect 16639 20852 16725 20856
rect 16639 20796 16651 20852
rect 16707 20796 16725 20852
rect 16639 20784 16725 20796
rect 16907 20648 17943 21013
rect 18125 20853 18211 20857
rect 18125 20797 18137 20853
rect 18193 20797 18211 20853
rect 18125 20785 18211 20797
rect 18393 20648 18925 21013
rect -8627 18986 18925 20648
rect -8627 18985 -6616 18986
rect -8627 18929 -8102 18985
rect -8046 18929 -7284 18985
rect -7228 18930 -6616 18985
rect -6560 18930 -5798 18986
rect -5742 18983 18925 18986
rect -5742 18982 -2574 18983
rect -5742 18930 -4060 18982
rect -7228 18929 -4060 18930
rect -8627 18926 -4060 18929
rect -4004 18926 -3242 18982
rect -3186 18927 -2574 18982
rect -2518 18927 -1756 18983
rect -1700 18982 1468 18983
rect -1700 18927 -18 18982
rect -3186 18926 -18 18927
rect 38 18926 800 18982
rect 856 18927 1468 18982
rect 1524 18927 2286 18983
rect 2342 18982 5510 18983
rect 2342 18927 4024 18982
rect 856 18926 4024 18927
rect 4080 18926 4842 18982
rect 4898 18927 5510 18982
rect 5566 18927 6328 18983
rect 6384 18982 9552 18983
rect 6384 18927 8066 18982
rect 4898 18926 8066 18927
rect 8122 18926 8884 18982
rect 8940 18927 9552 18982
rect 9608 18927 10370 18983
rect 10426 18982 13594 18983
rect 10426 18927 12108 18982
rect 8940 18926 12108 18927
rect 12164 18926 12926 18982
rect 12982 18927 13594 18982
rect 13650 18927 14412 18983
rect 14468 18982 17636 18983
rect 14468 18927 16150 18982
rect 12982 18926 16150 18927
rect 16206 18926 16968 18982
rect 17024 18927 17636 18982
rect 17692 18927 18454 18983
rect 18510 18927 18925 18983
rect 17024 18926 18925 18927
rect -8627 18811 18925 18926
rect -8627 18446 -7795 18811
rect -7345 18808 18925 18811
rect -7613 18650 -7527 18654
rect -7613 18594 -7601 18650
rect -7545 18594 -7527 18650
rect -7613 18582 -7527 18594
rect -7345 18446 -3753 18808
rect -3571 18647 -3485 18651
rect -3571 18591 -3559 18647
rect -3503 18591 -3485 18647
rect -3571 18579 -3485 18591
rect -8627 18443 -3753 18446
rect -3303 18443 289 18808
rect 471 18647 557 18651
rect 471 18591 483 18647
rect 539 18591 557 18647
rect 471 18579 557 18591
rect 739 18443 4331 18808
rect 4513 18647 4599 18651
rect 4513 18591 4525 18647
rect 4581 18591 4599 18647
rect 4513 18579 4599 18591
rect 4781 18443 8373 18808
rect 8555 18647 8641 18651
rect 8555 18591 8567 18647
rect 8623 18591 8641 18647
rect 8555 18579 8641 18591
rect 8823 18443 12415 18808
rect 12597 18647 12683 18651
rect 12597 18591 12609 18647
rect 12665 18591 12683 18647
rect 12597 18579 12683 18591
rect 12865 18443 16457 18808
rect 16639 18647 16725 18651
rect 16639 18591 16651 18647
rect 16707 18591 16725 18647
rect 16639 18579 16725 18591
rect 16907 18443 18925 18808
rect -8627 17446 18925 18443
rect -8627 17390 15386 17446
rect 15442 17390 18925 17446
rect -8627 16780 18925 17390
rect -8627 16724 -8102 16780
rect -8046 16724 -7284 16780
rect -7228 16777 18925 16780
rect -7228 16724 -4060 16777
rect -8627 16721 -4060 16724
rect -4004 16721 -3242 16777
rect -3186 16721 -18 16777
rect 38 16721 800 16777
rect 856 16721 4024 16777
rect 4080 16721 4842 16777
rect 4898 16721 8066 16777
rect 8122 16721 8884 16777
rect 8940 16721 12108 16777
rect 12164 16721 12926 16777
rect 12982 16721 16150 16777
rect 16206 16721 16968 16777
rect 17024 16721 18925 16777
rect -8627 16594 18925 16721
rect -8687 16591 18925 16594
rect 32519 22673 43287 26106
rect -8687 15794 14943 16591
rect -11625 15686 -11539 15690
rect -11625 15630 -11613 15686
rect -11557 15630 -11539 15686
rect -11625 15618 -11539 15630
rect -9339 15482 -8627 15794
rect -7613 15686 -7527 15690
rect -7613 15630 -7601 15686
rect -7545 15630 -7527 15686
rect -7613 15618 -7527 15630
rect -5327 15482 -4585 15794
rect -3571 15686 -3485 15690
rect -3571 15630 -3559 15686
rect -3503 15630 -3485 15686
rect -3571 15618 -3485 15630
rect -1285 15482 -543 15794
rect 471 15686 557 15690
rect 471 15630 483 15686
rect 539 15630 557 15686
rect 471 15618 557 15630
rect 2757 15482 3499 15794
rect 4513 15686 4599 15690
rect 4513 15630 4525 15686
rect 4581 15630 4599 15686
rect 4513 15618 4599 15630
rect 6799 15482 7541 15794
rect 8555 15686 8641 15690
rect 8555 15630 8567 15686
rect 8623 15630 8641 15686
rect 8555 15618 8641 15630
rect 10841 15482 11583 15794
rect 12597 15686 12683 15690
rect 12597 15630 12609 15686
rect 12665 15630 12683 15686
rect 12597 15618 12683 15630
rect -12639 14809 14883 15482
rect -12639 14569 -8857 14809
rect -8777 14717 -8691 14729
rect -8777 14661 -8765 14717
rect -8709 14661 -8691 14717
rect -8777 14649 -8691 14661
rect -8627 14569 -4815 14809
rect -4735 14717 -4649 14729
rect -4735 14661 -4723 14717
rect -4667 14661 -4649 14717
rect -4735 14649 -4649 14661
rect -4585 14569 -773 14809
rect -693 14717 -607 14729
rect -693 14661 -681 14717
rect -625 14661 -607 14717
rect -693 14649 -607 14661
rect -543 14569 3269 14809
rect 3349 14717 3435 14729
rect 3349 14661 3361 14717
rect 3417 14661 3435 14717
rect 3349 14649 3435 14661
rect 3499 14569 7311 14809
rect 7391 14717 7477 14729
rect 7391 14661 7403 14717
rect 7459 14661 7477 14717
rect 7391 14649 7477 14661
rect 7541 14569 11353 14809
rect 11433 14717 11519 14729
rect 11433 14661 11445 14717
rect 11501 14661 11519 14717
rect 11433 14649 11519 14661
rect 11583 14569 14883 14809
rect -12639 13816 14883 14569
rect -12639 13760 -12114 13816
rect -12058 13760 -11296 13816
rect -11240 13760 -8102 13816
rect -8046 13760 -7284 13816
rect -7228 13760 -4060 13816
rect -4004 13760 -3242 13816
rect -3186 13760 -18 13816
rect 38 13760 800 13816
rect 856 13760 4024 13816
rect 4080 13760 4842 13816
rect 4898 13760 8066 13816
rect 8122 13760 8884 13816
rect 8940 13760 12108 13816
rect 12164 13760 12926 13816
rect 12982 13760 14883 13816
rect -12639 13642 14883 13760
rect -12639 13277 -11807 13642
rect -11625 13481 -11539 13485
rect -11625 13425 -11613 13481
rect -11557 13425 -11539 13481
rect -11625 13413 -11539 13425
rect -11357 13277 -10321 13642
rect -10139 13481 -10053 13485
rect -10139 13425 -10127 13481
rect -10071 13425 -10053 13481
rect -10139 13413 -10053 13425
rect -9871 13277 -7795 13642
rect -7613 13481 -7527 13485
rect -7613 13425 -7601 13481
rect -7545 13425 -7527 13481
rect -7613 13413 -7527 13425
rect -7345 13277 -6309 13642
rect -6127 13481 -6041 13485
rect -6127 13425 -6115 13481
rect -6059 13425 -6041 13481
rect -6127 13413 -6041 13425
rect -5859 13277 -3753 13642
rect -3571 13481 -3485 13485
rect -3571 13425 -3559 13481
rect -3503 13425 -3485 13481
rect -3571 13413 -3485 13425
rect -3303 13277 -2267 13642
rect -2085 13481 -1999 13485
rect -2085 13425 -2073 13481
rect -2017 13425 -1999 13481
rect -2085 13413 -1999 13425
rect -1817 13277 289 13642
rect 471 13481 557 13485
rect 471 13425 483 13481
rect 539 13425 557 13481
rect 471 13413 557 13425
rect 739 13277 1775 13642
rect 1957 13481 2043 13485
rect 1957 13425 1969 13481
rect 2025 13425 2043 13481
rect 1957 13413 2043 13425
rect 2225 13277 4331 13642
rect 4513 13481 4599 13485
rect 4513 13425 4525 13481
rect 4581 13425 4599 13481
rect 4513 13413 4599 13425
rect 4781 13277 5817 13642
rect 5999 13481 6085 13485
rect 5999 13425 6011 13481
rect 6067 13425 6085 13481
rect 5999 13413 6085 13425
rect 6267 13277 8373 13642
rect 8555 13481 8641 13485
rect 8555 13425 8567 13481
rect 8623 13425 8641 13481
rect 8555 13413 8641 13425
rect 8823 13277 9859 13642
rect 10041 13481 10127 13485
rect 10041 13425 10053 13481
rect 10109 13425 10127 13481
rect 10041 13413 10127 13425
rect 10309 13277 12415 13642
rect 12597 13481 12683 13485
rect 12597 13425 12609 13481
rect 12665 13425 12683 13481
rect 12597 13413 12683 13425
rect 12865 13277 13901 13642
rect 14083 13481 14169 13485
rect 14083 13425 14095 13481
rect 14151 13425 14169 13481
rect 14083 13413 14169 13425
rect 14351 13277 14883 13642
rect -12639 11611 14883 13277
rect -12639 11555 -12114 11611
rect -12058 11555 -11296 11611
rect -11240 11555 -10628 11611
rect -10572 11555 -9810 11611
rect -9754 11555 -8102 11611
rect -8046 11555 -7284 11611
rect -7228 11555 -6616 11611
rect -6560 11555 -5798 11611
rect -5742 11555 -4060 11611
rect -4004 11555 -3242 11611
rect -3186 11555 -2574 11611
rect -2518 11555 -1756 11611
rect -1700 11555 -18 11611
rect 38 11555 800 11611
rect 856 11555 1468 11611
rect 1524 11555 2286 11611
rect 2342 11555 4024 11611
rect 4080 11555 4842 11611
rect 4898 11555 5510 11611
rect 5566 11555 6328 11611
rect 6384 11555 8066 11611
rect 8122 11555 8884 11611
rect 8940 11555 9552 11611
rect 9608 11555 10370 11611
rect 10426 11555 12108 11611
rect 12164 11555 12926 11611
rect 12982 11555 13594 11611
rect 13650 11555 14412 11611
rect 14468 11555 14883 11611
rect -12639 11437 14883 11555
rect -12639 11072 -11807 11437
rect -11625 11276 -11539 11280
rect -11625 11220 -11613 11276
rect -11557 11220 -11539 11276
rect -11625 11208 -11539 11220
rect -11357 11072 -10321 11437
rect -10139 11277 -10053 11281
rect -10139 11221 -10127 11277
rect -10071 11221 -10053 11277
rect -10139 11209 -10053 11221
rect -9871 11072 -7795 11437
rect -7613 11276 -7527 11280
rect -7613 11220 -7601 11276
rect -7545 11220 -7527 11276
rect -7613 11208 -7527 11220
rect -7345 11072 -6309 11437
rect -6127 11277 -6041 11281
rect -6127 11221 -6115 11277
rect -6059 11221 -6041 11277
rect -6127 11209 -6041 11221
rect -5859 11072 -3753 11437
rect -3571 11276 -3485 11280
rect -3571 11220 -3559 11276
rect -3503 11220 -3485 11276
rect -3571 11208 -3485 11220
rect -3303 11072 -2267 11437
rect -2085 11277 -1999 11281
rect -2085 11221 -2073 11277
rect -2017 11221 -1999 11277
rect -2085 11209 -1999 11221
rect -1817 11072 289 11437
rect 471 11276 557 11280
rect 471 11220 483 11276
rect 539 11220 557 11276
rect 471 11208 557 11220
rect 739 11072 1775 11437
rect 1957 11277 2043 11281
rect 1957 11221 1969 11277
rect 2025 11221 2043 11277
rect 1957 11209 2043 11221
rect 2225 11072 4331 11437
rect 4513 11276 4599 11280
rect 4513 11220 4525 11276
rect 4581 11220 4599 11276
rect 4513 11208 4599 11220
rect 4781 11072 5817 11437
rect 5999 11277 6085 11281
rect 5999 11221 6011 11277
rect 6067 11221 6085 11277
rect 5999 11209 6085 11221
rect 6267 11072 8373 11437
rect 8555 11276 8641 11280
rect 8555 11220 8567 11276
rect 8623 11220 8641 11276
rect 8555 11208 8641 11220
rect 8823 11072 9859 11437
rect 10041 11277 10127 11281
rect 10041 11221 10053 11277
rect 10109 11221 10127 11277
rect 10041 11209 10127 11221
rect 10309 11072 12415 11437
rect 12597 11276 12683 11280
rect 12597 11220 12609 11276
rect 12665 11220 12683 11276
rect 12597 11208 12683 11220
rect 12865 11072 13901 11437
rect 14083 11277 14169 11281
rect 14083 11221 14095 11277
rect 14151 11221 14169 11277
rect 14083 11209 14169 11221
rect 14351 11072 14883 11437
rect -12639 9407 14883 11072
rect -12639 9406 -10628 9407
rect -12639 9350 -12114 9406
rect -12058 9350 -11296 9406
rect -11240 9351 -10628 9406
rect -10572 9351 -9810 9407
rect -9754 9406 -6616 9407
rect -9754 9351 -8102 9406
rect -11240 9350 -8102 9351
rect -8046 9350 -7284 9406
rect -7228 9351 -6616 9406
rect -6560 9351 -5798 9407
rect -5742 9406 -2574 9407
rect -5742 9351 -4060 9406
rect -7228 9350 -4060 9351
rect -4004 9350 -3242 9406
rect -3186 9351 -2574 9406
rect -2518 9351 -1756 9407
rect -1700 9406 1468 9407
rect -1700 9351 -18 9406
rect -3186 9350 -18 9351
rect 38 9350 800 9406
rect 856 9351 1468 9406
rect 1524 9351 2286 9407
rect 2342 9406 5510 9407
rect 2342 9351 4024 9406
rect 856 9350 4024 9351
rect 4080 9350 4842 9406
rect 4898 9351 5510 9406
rect 5566 9351 6328 9407
rect 6384 9406 9552 9407
rect 6384 9351 8066 9406
rect 4898 9350 8066 9351
rect 8122 9350 8884 9406
rect 8940 9351 9552 9406
rect 9608 9351 10370 9407
rect 10426 9406 13594 9407
rect 10426 9351 12108 9406
rect 8940 9350 12108 9351
rect 12164 9350 12926 9406
rect 12982 9351 13594 9406
rect 13650 9351 14412 9407
rect 14468 9351 14883 9407
rect 12982 9350 14883 9351
rect -12639 9232 14883 9350
rect -12639 8867 -11807 9232
rect -11625 9071 -11539 9075
rect -11625 9015 -11613 9071
rect -11557 9015 -11539 9071
rect -11625 9003 -11539 9015
rect -11357 8867 -7795 9232
rect -7613 9071 -7527 9075
rect -7613 9015 -7601 9071
rect -7545 9015 -7527 9071
rect -7613 9003 -7527 9015
rect -7345 8867 -3753 9232
rect -3571 9071 -3485 9075
rect -3571 9015 -3559 9071
rect -3503 9015 -3485 9071
rect -3571 9003 -3485 9015
rect -3303 8867 289 9232
rect 471 9071 557 9075
rect 471 9015 483 9071
rect 539 9015 557 9071
rect 471 9003 557 9015
rect 739 8867 4331 9232
rect 4513 9071 4599 9075
rect 4513 9015 4525 9071
rect 4581 9015 4599 9071
rect 4513 9003 4599 9015
rect 4781 8867 8373 9232
rect 8555 9071 8641 9075
rect 8555 9015 8567 9071
rect 8623 9015 8641 9071
rect 8555 9003 8641 9015
rect 8823 8867 12415 9232
rect 12597 9071 12683 9075
rect 12597 9015 12609 9071
rect 12665 9015 12683 9071
rect 12597 9003 12683 9015
rect 12865 8867 14883 9232
rect -12639 7882 14883 8867
rect -12908 7870 14883 7882
rect -12908 7814 -12896 7870
rect -12840 7814 14883 7870
rect -12908 7722 14883 7814
rect -12639 7201 14883 7722
rect -12639 7145 -12114 7201
rect -12058 7145 -11296 7201
rect -11240 7145 -8102 7201
rect -8046 7145 -7284 7201
rect -7228 7145 -4060 7201
rect -4004 7145 -3242 7201
rect -3186 7145 -18 7201
rect 38 7145 800 7201
rect 856 7145 4024 7201
rect 4080 7145 4842 7201
rect 4898 7145 8066 7201
rect 8122 7145 8884 7201
rect 8940 7145 12108 7201
rect 12164 7145 12926 7201
rect 12982 7145 14883 7201
rect -12908 7083 -12822 7095
rect -12908 7027 -12896 7083
rect -12840 7027 -12822 7083
rect -12908 7015 -12822 7027
rect -12639 7015 14883 7145
rect -4464 6434 -2430 6477
rect -4464 6134 -4454 6434
rect -2454 6134 -2430 6434
rect -4464 6097 -2430 6134
rect -8971 -1070 -8871 -1058
rect -8971 -1126 -8949 -1070
rect -8893 -1126 -8871 -1070
rect -8971 -1138 -8871 -1126
rect -7756 -1070 -7656 -1058
rect -7756 -1126 -7734 -1070
rect -7678 -1126 -7656 -1070
rect -7756 -1138 -7656 -1126
rect -9266 -1226 -9186 -1216
rect -9266 -1282 -9254 -1226
rect -9198 -1282 -9186 -1226
rect -9266 -1292 -9186 -1282
rect -9254 -1618 -9198 -1292
rect -8949 -1464 -8893 -1138
rect -8051 -1226 -7971 -1216
rect -8051 -1282 -8039 -1226
rect -7983 -1282 -7971 -1226
rect -8051 -1292 -7971 -1282
rect -8961 -1474 -8881 -1464
rect -8961 -1530 -8949 -1474
rect -8893 -1530 -8881 -1474
rect -8961 -1540 -8881 -1530
rect -8039 -1618 -7983 -1292
rect -7734 -1464 -7678 -1138
rect -7746 -1474 -7666 -1464
rect -7746 -1530 -7734 -1474
rect -7678 -1530 -7666 -1474
rect -7746 -1540 -7666 -1530
rect -9276 -1630 -9176 -1618
rect -9276 -1686 -9254 -1630
rect -9198 -1686 -9176 -1630
rect -9276 -1698 -9176 -1686
rect -8061 -1630 -7961 -1618
rect -8061 -1686 -8039 -1630
rect -7983 -1686 -7961 -1630
rect -8061 -1698 -7961 -1686
rect -4464 -3322 30646 -3321
rect 32519 -3322 35819 22673
rect -4464 -3363 35819 -3322
rect -4464 -3663 -4454 -3363
rect -2454 -3663 35819 -3363
rect -4464 -3701 35819 -3663
rect 30646 -3702 35819 -3701
<< via4 >>
rect 40739 39093 40957 39167
rect -4343 37511 -4287 37567
rect 5129 37511 5185 37567
rect 14601 37512 14657 37568
rect 24073 37512 24129 37568
rect 33545 37512 33601 37568
rect 43017 37512 43073 37568
rect -5507 36542 -5451 36598
rect 3965 36542 4021 36598
rect -4343 35306 -4287 35362
rect -2857 35306 -2801 35362
rect -4343 33101 -4287 33157
rect -2857 33102 -2801 33158
rect -6327 31169 -6027 31969
rect 13437 36543 13493 36599
rect 5129 35306 5185 35362
rect 6615 35306 6671 35362
rect 5129 33101 5185 33157
rect 6615 33102 6671 33158
rect -1245 31169 -1045 31969
rect 3145 31169 3445 31969
rect 22909 36543 22965 36599
rect 14601 35307 14657 35363
rect 16087 35307 16143 35363
rect 14601 33102 14657 33158
rect 16087 33103 16143 33159
rect -4343 30896 -4287 30952
rect 8227 31170 8427 31970
rect 12617 31170 12917 31970
rect 32381 36543 32437 36599
rect 24073 35307 24129 35363
rect 25559 35307 25615 35363
rect 24073 33102 24129 33158
rect 25559 33103 25615 33159
rect 5129 30896 5185 30952
rect -5610 28908 -5554 28964
rect 17699 31170 17899 31970
rect 22089 31170 22389 31970
rect 41853 36543 41909 36599
rect 33545 35307 33601 35363
rect 35031 35307 35087 35363
rect 33545 33102 33601 33158
rect 35031 33103 35087 33159
rect 14601 30897 14657 30953
rect 3862 28908 3918 28964
rect 27171 31170 27371 31970
rect 31561 31170 31861 31970
rect 43017 35307 43073 35363
rect 44503 35307 44559 35363
rect 43017 33102 43073 33158
rect 44503 33103 44559 33159
rect 24073 30897 24129 30953
rect 13334 28909 13390 28965
rect 36643 31170 36843 31970
rect 41033 31170 41333 31970
rect 33545 30897 33601 30953
rect 22806 28909 22862 28965
rect 43017 30897 43073 30953
rect 32278 28909 32334 28965
rect 41750 28909 41806 28965
rect -7601 25209 -7545 25265
rect -3559 25206 -3503 25262
rect 483 25206 539 25262
rect 4525 25206 4581 25262
rect 8567 25206 8623 25262
rect 12609 25206 12665 25262
rect 16651 25206 16707 25262
rect -7601 23004 -7545 23060
rect -6115 23004 -6059 23060
rect -3559 23001 -3503 23057
rect -2073 23001 -2017 23057
rect 483 23001 539 23057
rect 1969 23001 2025 23057
rect 4525 23001 4581 23057
rect 6011 23001 6067 23057
rect 8567 23001 8623 23057
rect 10053 23001 10109 23057
rect 12609 23001 12665 23057
rect 14095 23001 14151 23057
rect 16651 23001 16707 23057
rect 18137 23001 18193 23057
rect -7601 20799 -7545 20855
rect -6115 20800 -6059 20856
rect -3559 20796 -3503 20852
rect -2073 20797 -2017 20853
rect 483 20796 539 20852
rect 1969 20797 2025 20853
rect 4525 20796 4581 20852
rect 6011 20797 6067 20853
rect 8567 20796 8623 20852
rect 10053 20797 10109 20853
rect 12609 20796 12665 20852
rect 14095 20797 14151 20853
rect 16651 20796 16707 20852
rect 18137 20797 18193 20853
rect -7601 18594 -7545 18650
rect -3559 18591 -3503 18647
rect 483 18591 539 18647
rect 4525 18591 4581 18647
rect 8567 18591 8623 18647
rect 12609 18591 12665 18647
rect 16651 18591 16707 18647
rect -11613 15630 -11557 15686
rect -7601 15630 -7545 15686
rect -3559 15630 -3503 15686
rect 483 15630 539 15686
rect 4525 15630 4581 15686
rect 8567 15630 8623 15686
rect 12609 15630 12665 15686
rect -8765 14661 -8709 14717
rect -4723 14661 -4667 14717
rect -681 14661 -625 14717
rect 3361 14661 3417 14717
rect 7403 14661 7459 14717
rect 11445 14661 11501 14717
rect -11613 13425 -11557 13481
rect -10127 13425 -10071 13481
rect -7601 13425 -7545 13481
rect -6115 13425 -6059 13481
rect -3559 13425 -3503 13481
rect -2073 13425 -2017 13481
rect 483 13425 539 13481
rect 1969 13425 2025 13481
rect 4525 13425 4581 13481
rect 6011 13425 6067 13481
rect 8567 13425 8623 13481
rect 10053 13425 10109 13481
rect 12609 13425 12665 13481
rect 14095 13425 14151 13481
rect -11613 11220 -11557 11276
rect -10127 11221 -10071 11277
rect -7601 11220 -7545 11276
rect -6115 11221 -6059 11277
rect -3559 11220 -3503 11276
rect -2073 11221 -2017 11277
rect 483 11220 539 11276
rect 1969 11221 2025 11277
rect 4525 11220 4581 11276
rect 6011 11221 6067 11277
rect 8567 11220 8623 11276
rect 10053 11221 10109 11277
rect 12609 11220 12665 11276
rect 14095 11221 14151 11277
rect -11613 9015 -11557 9071
rect -7601 9015 -7545 9071
rect -3559 9015 -3503 9071
rect 483 9015 539 9071
rect 4525 9015 4581 9071
rect 8567 9015 8623 9071
rect 12609 9015 12665 9071
rect -12896 7027 -12840 7083
rect -4454 6134 -2454 6434
<< metal5 >>
rect 4441 37675 7099 39882
rect 40726 39167 42468 39280
rect 40726 39093 40739 39167
rect 40957 39093 42468 39167
rect 40726 39080 42468 39093
rect 41991 37676 42468 39080
rect -5369 37567 -2069 37675
rect -5369 37511 -4343 37567
rect -4287 37511 -2069 37567
rect -5369 36801 -2069 37511
rect 4103 37567 7403 37675
rect 4103 37511 5129 37567
rect 5185 37511 7403 37567
rect 4103 36801 7403 37511
rect 13575 37568 16875 37676
rect 13575 37512 14601 37568
rect 14657 37512 16875 37568
rect 13575 36801 16875 37512
rect 23047 37568 26347 37676
rect 23047 37512 24073 37568
rect 24129 37512 26347 37568
rect 23047 36801 26347 37512
rect 32519 37568 35819 37676
rect 32519 37512 33545 37568
rect 33601 37512 35819 37568
rect 32519 36801 35819 37512
rect -5369 36791 35819 36801
rect 41991 37568 45291 37676
rect 41991 37512 43017 37568
rect 43073 37512 45291 37568
rect 41991 36791 45291 37512
rect -5369 36690 45291 36791
rect -5521 36599 45291 36690
rect -5521 36598 13437 36599
rect -5521 36542 -5507 36598
rect -5451 36542 3965 36598
rect 4021 36543 13437 36598
rect 13493 36543 22909 36599
rect 22965 36543 32381 36599
rect 32437 36543 41853 36599
rect 41909 36543 45291 36599
rect 4021 36542 45291 36543
rect -5521 36530 45291 36542
rect -5369 35723 45291 36530
rect -5369 35362 -2069 35723
rect -5369 35306 -4343 35362
rect -4287 35306 -2857 35362
rect -2801 35306 -2069 35362
rect -5369 33158 -2069 35306
rect -5369 33157 -2857 33158
rect -5369 33101 -4343 33157
rect -4287 33102 -2857 33157
rect -2801 33102 -2069 33158
rect -4287 33101 -2069 33102
rect -5369 31979 -2069 33101
rect 4103 35362 7403 35723
rect 4103 35306 5129 35362
rect 5185 35306 6615 35362
rect 6671 35306 7403 35362
rect 4103 33158 7403 35306
rect 4103 33157 6615 33158
rect 4103 33101 5129 33157
rect 5185 33102 6615 33157
rect 6671 33102 7403 33158
rect 5185 33101 7403 33102
rect 4103 31980 7403 33101
rect 13575 35363 16875 35723
rect 13575 35307 14601 35363
rect 14657 35307 16087 35363
rect 16143 35307 16875 35363
rect 13575 33159 16875 35307
rect 13575 33158 16087 33159
rect 13575 33102 14601 33158
rect 14657 33103 16087 33158
rect 16143 33103 16875 33159
rect 14657 33102 16875 33103
rect 13575 31980 16875 33102
rect 23047 35363 26347 35723
rect 23047 35307 24073 35363
rect 24129 35307 25559 35363
rect 25615 35307 26347 35363
rect 23047 33159 26347 35307
rect 23047 33158 25559 33159
rect 23047 33102 24073 33158
rect 24129 33103 25559 33158
rect 25615 33103 26347 33159
rect 24129 33102 26347 33103
rect 23047 31980 26347 33102
rect 32519 35713 45291 35723
rect 32519 35363 35819 35713
rect 32519 35307 33545 35363
rect 33601 35307 35031 35363
rect 35087 35307 35819 35363
rect 32519 33159 35819 35307
rect 32519 33158 35031 33159
rect 32519 33102 33545 33158
rect 33601 33103 35031 33158
rect 35087 33103 35819 33159
rect 33601 33102 35819 33103
rect 32519 31980 35819 33102
rect 41991 35363 45291 35713
rect 41991 35307 43017 35363
rect 43073 35307 44503 35363
rect 44559 35307 45291 35363
rect 41991 33159 45291 35307
rect 41991 33158 44503 33159
rect 41991 33102 43017 33158
rect 43073 33103 44503 33158
rect 44559 33103 45291 33159
rect 43073 33102 45291 33103
rect 41991 31980 45291 33102
rect 4103 31979 8437 31980
rect -6337 31969 -1035 31979
rect -6337 31169 -6327 31969
rect -6027 31169 -1245 31969
rect -1045 31169 -1035 31969
rect -6337 31159 -1035 31169
rect 3135 31970 8437 31979
rect 3135 31969 8227 31970
rect 3135 31169 3145 31969
rect 3445 31170 8227 31969
rect 8427 31170 8437 31970
rect 3445 31169 8437 31170
rect 3135 31160 8437 31169
rect 12607 31970 17909 31980
rect 12607 31170 12617 31970
rect 12917 31170 17699 31970
rect 17899 31170 17909 31970
rect 12607 31160 17909 31170
rect 22079 31970 27381 31980
rect 22079 31170 22089 31970
rect 22389 31170 27171 31970
rect 27371 31170 27381 31970
rect 22079 31160 27381 31170
rect 31551 31970 36853 31980
rect 31551 31170 31561 31970
rect 31861 31170 36643 31970
rect 36843 31170 36853 31970
rect 31551 31160 36853 31170
rect 41023 31970 45291 31980
rect 41023 31170 41033 31970
rect 41333 31170 45291 31970
rect 41023 31160 45291 31170
rect 3135 31159 7403 31160
rect -5369 30952 -2069 31159
rect -5369 30896 -4343 30952
rect -4287 30896 -2069 30952
rect -5369 29056 -2069 30896
rect 4103 30952 7403 31159
rect 4103 30896 5129 30952
rect 5185 30896 7403 30952
rect 4103 29056 7403 30896
rect 13575 30953 16875 31160
rect 13575 30897 14601 30953
rect 14657 30897 16875 30953
rect 13575 29057 16875 30897
rect 23047 30953 26347 31160
rect 23047 30897 24073 30953
rect 24129 30897 26347 30953
rect 23047 29057 26347 30897
rect 32519 30953 35819 31160
rect 32519 30897 33545 30953
rect 33601 30897 35819 30953
rect 32519 29057 35819 30897
rect 41991 30953 45291 31160
rect 41991 30897 43017 30953
rect 43073 30897 45291 30953
rect 41991 29057 45291 30897
rect -5622 28964 -2069 29056
rect -5622 28908 -5610 28964
rect -5554 28908 -2069 28964
rect -5622 28896 -2069 28908
rect 3850 28964 7403 29056
rect 3850 28908 3862 28964
rect 3918 28908 7403 28964
rect 3850 28896 7403 28908
rect 13322 28965 16875 29057
rect 13322 28909 13334 28965
rect 13390 28909 16875 28965
rect 13322 28897 16875 28909
rect 22794 28965 26347 29057
rect 22794 28909 22806 28965
rect 22862 28909 26347 28965
rect 22794 28897 26347 28909
rect 32266 28965 35819 29057
rect 32266 28909 32278 28965
rect 32334 28909 35819 28965
rect 32266 28897 35819 28909
rect 41738 28965 45291 29057
rect 41738 28909 41750 28965
rect 41806 28909 45291 28965
rect 41738 28897 45291 28909
rect -5369 25373 -2069 28896
rect -8627 25370 -2069 25373
rect 4103 25370 7403 28896
rect 13575 25370 16875 28897
rect 23047 25370 26347 28897
rect -8627 25265 26347 25370
rect -8627 25209 -7601 25265
rect -7545 25262 26347 25265
rect -7545 25209 -3559 25262
rect -8627 25206 -3559 25209
rect -3503 25206 483 25262
rect 539 25206 4525 25262
rect 4581 25206 8567 25262
rect 8623 25206 12609 25262
rect 12665 25206 16651 25262
rect 16707 25206 26347 25262
rect -8627 23060 26347 25206
rect -8627 23004 -7601 23060
rect -7545 23004 -6115 23060
rect -6059 23057 26347 23060
rect -6059 23004 -3559 23057
rect -8627 23001 -3559 23004
rect -3503 23001 -2073 23057
rect -2017 23001 483 23057
rect 539 23001 1969 23057
rect 2025 23001 4525 23057
rect 4581 23001 6011 23057
rect 6067 23001 8567 23057
rect 8623 23001 10053 23057
rect 10109 23001 12609 23057
rect 12665 23001 14095 23057
rect 14151 23001 16651 23057
rect 16707 23001 18137 23057
rect 18193 23001 26347 23057
rect -8627 21844 26347 23001
rect -8627 21162 18925 21844
rect -8627 20922 15295 21162
rect 15533 20922 18925 21162
rect -8627 20856 18925 20922
rect -8627 20855 -6115 20856
rect -8627 20799 -7601 20855
rect -7545 20800 -6115 20855
rect -6059 20853 18925 20856
rect -6059 20852 -2073 20853
rect -6059 20800 -3559 20852
rect -7545 20799 -3559 20800
rect -8627 20796 -3559 20799
rect -3503 20797 -2073 20852
rect -2017 20852 1969 20853
rect -2017 20797 483 20852
rect -3503 20796 483 20797
rect 539 20797 1969 20852
rect 2025 20852 6011 20853
rect 2025 20797 4525 20852
rect 539 20796 4525 20797
rect 4581 20797 6011 20852
rect 6067 20852 10053 20853
rect 6067 20797 8567 20852
rect 4581 20796 8567 20797
rect 8623 20797 10053 20852
rect 10109 20852 14095 20853
rect 10109 20797 12609 20852
rect 8623 20796 12609 20797
rect 12665 20797 14095 20852
rect 14151 20852 18137 20853
rect 14151 20797 16651 20852
rect 12665 20796 16651 20797
rect 16707 20797 18137 20852
rect 18193 20797 18925 20853
rect 16707 20796 18925 20797
rect -8627 18650 18925 20796
rect -8627 18594 -7601 18650
rect -7545 18647 18925 18650
rect -7545 18594 -3559 18647
rect -8627 18591 -3559 18594
rect -3503 18591 483 18647
rect 539 18591 4525 18647
rect 4581 18591 8567 18647
rect 8623 18591 12609 18647
rect 12665 18591 16651 18647
rect 16707 18591 18925 18647
rect -8627 17538 18925 18591
rect -8627 17298 15293 17538
rect 15535 17298 18925 17538
rect -8627 16594 18925 17298
rect -8687 16591 18925 16594
rect -8687 15794 14943 16591
rect -12639 15686 14883 15794
rect -12639 15630 -11613 15686
rect -11557 15630 -7601 15686
rect -7545 15630 -3559 15686
rect -3503 15630 483 15686
rect 539 15630 4525 15686
rect 4581 15630 8567 15686
rect 8623 15630 12609 15686
rect 12665 15630 14883 15686
rect -12639 14717 14883 15630
rect -12639 14661 -8765 14717
rect -8709 14661 -4723 14717
rect -4667 14661 -681 14717
rect -625 14661 3361 14717
rect 3417 14661 7403 14717
rect 7459 14661 11445 14717
rect 11501 14661 14883 14717
rect -12639 13481 14883 14661
rect -12639 13425 -11613 13481
rect -11557 13425 -10127 13481
rect -10071 13425 -7601 13481
rect -7545 13425 -6115 13481
rect -6059 13425 -3559 13481
rect -3503 13425 -2073 13481
rect -2017 13425 483 13481
rect 539 13425 1969 13481
rect 2025 13425 4525 13481
rect 4581 13425 6011 13481
rect 6067 13425 8567 13481
rect 8623 13425 10053 13481
rect 10109 13425 12609 13481
rect 12665 13425 14095 13481
rect 14151 13425 14883 13481
rect -12639 11277 14883 13425
rect -12639 11276 -10127 11277
rect -12639 11220 -11613 11276
rect -11557 11221 -10127 11276
rect -10071 11276 -6115 11277
rect -10071 11221 -7601 11276
rect -11557 11220 -7601 11221
rect -7545 11221 -6115 11276
rect -6059 11276 -2073 11277
rect -6059 11221 -3559 11276
rect -7545 11220 -3559 11221
rect -3503 11221 -2073 11276
rect -2017 11276 1969 11277
rect -2017 11221 483 11276
rect -3503 11220 483 11221
rect 539 11221 1969 11276
rect 2025 11276 6011 11277
rect 2025 11221 4525 11276
rect 539 11220 4525 11221
rect 4581 11221 6011 11276
rect 6067 11276 10053 11277
rect 6067 11221 8567 11276
rect 4581 11220 8567 11221
rect 8623 11221 10053 11276
rect 10109 11276 14095 11277
rect 10109 11221 12609 11276
rect 8623 11220 12609 11221
rect 12665 11221 14095 11276
rect 14151 11221 14883 11277
rect 12665 11220 14883 11221
rect -12639 9071 14883 11220
rect -12639 9015 -11613 9071
rect -11557 9015 -7601 9071
rect -7545 9015 -3559 9071
rect -3503 9015 483 9071
rect 539 9015 4525 9071
rect 4581 9015 8567 9071
rect 8623 9015 12609 9071
rect 12665 9015 14883 9071
rect -12639 7175 14883 9015
rect -12908 7083 14883 7175
rect -12908 7027 -12896 7083
rect -12840 7027 14883 7083
rect -12908 7015 14883 7027
rect 22821 6477 26347 21844
rect -4464 6434 26347 6477
rect -4464 6134 -4454 6434
rect -2454 6134 26347 6434
rect -4464 6097 26347 6134
rect 22821 -3206 26347 6097
<< labels >>
rlabel metal2 -13784 -3047 -13784 -3047 7 Clk
port 2 w
rlabel metal2 -13233 15938 -13233 15938 7 Reset
port 6 w
rlabel metal2 -13224 16448 -13224 16448 7 SAR_in
port 7 w
rlabel metal2 -13170 27549 -13170 27549 7 Load
port 8 w
rlabel metal2 -8063 38726 -8063 38726 1 Clk_piso
port 9 n
rlabel metal5 24711 -3206 24711 -3206 5 Vdd
port 0 s
rlabel metal4 34239 -3702 34239 -3702 5 Vss
port 1 s
rlabel metal2 -13880 -1213 -13880 -1213 7 Vin1
port 3 w
rlabel metal2 -13878 -1540 -13878 -1540 7 Vin2
port 4 w
rlabel metal2 -13894 4909 -13894 4909 7 Comp_out
port 5 w
rlabel metal1 -12861 6283 -12861 6283 7 comparator_no_offsetcal_0.VDD
rlabel metal1 -13302 -3521 -13302 -3521 7 comparator_no_offsetcal_0.VSS
rlabel metal1 -12776 -3043 -12776 -3043 7 comparator_no_offsetcal_0.CLK
rlabel metal1 -12871 -1218 -12871 -1218 7 comparator_no_offsetcal_0.Vin1
rlabel metal1 -12871 -1540 -12871 -1540 7 comparator_no_offsetcal_0.Vin2
rlabel metal2 -12616 4912 -12616 4912 7 comparator_no_offsetcal_0.Vout
rlabel metal2 -8799 -2720 -8799 -2720 7 comparator_no_offsetcal_0.no_offsetLatch_0.VSS
rlabel metal2 -10478 2277 -10478 2277 1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout1
rlabel metal2 -5842 2277 -5842 2277 1 comparator_no_offsetcal_0.no_offsetLatch_0.Vout2
rlabel metal1 -8163 2432 -8163 2432 1 comparator_no_offsetcal_0.no_offsetLatch_0.Clk
rlabel metal1 -6031 -1539 -6031 -1539 3 comparator_no_offsetcal_0.no_offsetLatch_0.Vin2
rlabel metal1 -6031 -1218 -6031 -1218 3 comparator_no_offsetcal_0.no_offsetLatch_0.Vin1
rlabel metal1 -9937 -5 -9937 -5 1 comparator_no_offsetcal_0.no_offsetLatch_0.Vp
rlabel metal1 -6338 -5 -6338 -5 1 comparator_no_offsetcal_0.no_offsetLatch_0.Vq
rlabel metal3 -8162 2243 -8162 2243 1 comparator_no_offsetcal_0.no_offsetLatch_0.VDD
rlabel metal1 -6729 4454 -6729 4454 3 comparator_no_offsetcal_0.x5.avdd
rlabel metal1 -6733 2598 -6733 2598 3 comparator_no_offsetcal_0.x5.avss
rlabel metal1 -6933 3326 -6933 3326 3 comparator_no_offsetcal_0.x5.in
rlabel metal1 -7085 3330 -7085 3330 3 comparator_no_offsetcal_0.x5.out
rlabel metal2 -10161 4650 -10161 4650 6 comparator_no_offsetcal_0.x4.A
rlabel metal2 -10721 4910 -10721 4910 6 comparator_no_offsetcal_0.x4.Y
rlabel metal1 -10031 5330 -10031 5330 6 comparator_no_offsetcal_0.x4.VDD
rlabel metal1 -10031 4250 -10031 4250 6 comparator_no_offsetcal_0.x4.VSS
rlabel metal1 -9593 4454 -9593 4454 7 comparator_no_offsetcal_0.x3.avdd
rlabel metal1 -9589 2598 -9589 2598 7 comparator_no_offsetcal_0.x3.avss
rlabel metal1 -9389 3326 -9389 3326 7 comparator_no_offsetcal_0.x3.in
rlabel metal1 -9237 3330 -9237 3330 7 comparator_no_offsetcal_0.x3.out
rlabel metal1 -8163 5157 -8163 5157 1 comparator_no_offsetcal_0.x2.VDD
rlabel metal2 -8871 4259 -8871 4259 7 comparator_no_offsetcal_0.x2.Vout1
rlabel metal2 -7451 4259 -7451 4259 3 comparator_no_offsetcal_0.x2.Vout2
rlabel metal2 -8391 3399 -8391 3399 5 comparator_no_offsetcal_0.x2.Vin1
rlabel metal2 -7930 3399 -7930 3399 5 comparator_no_offsetcal_0.x2.Vin2
rlabel metal1 -8158 3557 -8158 3557 5 comparator_no_offsetcal_0.x2.VSS
rlabel metal2 -13260 6872 -13260 6872 7 SARlogic_0.clk
rlabel metal2 -12988 15939 -12988 15939 7 SARlogic_0.reset
rlabel metal2 -12988 16447 -12988 16447 7 SARlogic_0.comp_in
rlabel metal2 -5053 26489 -5053 26489 1 SARlogic_0.d5
rlabel metal2 -998 26486 -998 26486 1 SARlogic_0.d4
rlabel metal2 3098 26486 3098 26486 1 SARlogic_0.d3
rlabel metal2 7139 26486 7139 26486 1 SARlogic_0.d2
rlabel metal2 11181 26489 11181 26489 1 SARlogic_0.d1
rlabel metal2 15225 26486 15225 26486 1 SARlogic_0.d0
rlabel metal5 6843 25370 6843 25370 1 SARlogic_0.vdd
rlabel metal4 2791 7015 2791 7015 5 SARlogic_0.vss
rlabel metal1 -8765 14689 -8765 14689 7 SARlogic_0.dffrs_0.setb
rlabel metal1 -8765 11466 -8765 11466 7 SARlogic_0.dffrs_0.clk
rlabel metal1 -8765 7841 -8765 7841 7 SARlogic_0.dffrs_0.d
rlabel metal1 -8748 7054 -8748 7054 7 SARlogic_0.dffrs_0.resetb
rlabel metal2 -5297 12368 -5297 12368 3 SARlogic_0.dffrs_0.Q
rlabel metal2 -5297 10163 -5297 10163 3 SARlogic_0.dffrs_0.Qb
rlabel metal5 -6657 15794 -6657 15794 1 SARlogic_0.dffrs_0.vdd
rlabel metal4 -6549 7015 -6549 7015 5 SARlogic_0.dffrs_0.vss
rlabel metal2 -7601 9083 -7601 9083 1 SARlogic_0.dffrs_0.nand3_8.VDD
rlabel metal1 -7191 7957 -7191 7957 3 SARlogic_0.dffrs_0.nand3_8.Z
rlabel metal1 -8277 7839 -8277 7839 7 SARlogic_0.dffrs_0.nand3_8.A
rlabel metal1 -8277 7958 -8277 7958 7 SARlogic_0.dffrs_0.nand3_8.B
rlabel metal1 -8277 8074 -8277 8074 7 SARlogic_0.dffrs_0.nand3_8.C
rlabel metal2 -7673 7133 -7673 7133 5 SARlogic_0.dffrs_0.nand3_8.VSS
rlabel metal2 -6115 11289 -6115 11289 1 SARlogic_0.dffrs_0.nand3_7.VDD
rlabel metal1 -5705 10163 -5705 10163 3 SARlogic_0.dffrs_0.nand3_7.Z
rlabel metal1 -6791 10045 -6791 10045 7 SARlogic_0.dffrs_0.nand3_7.A
rlabel metal1 -6791 10164 -6791 10164 7 SARlogic_0.dffrs_0.nand3_7.B
rlabel metal1 -6791 10280 -6791 10280 7 SARlogic_0.dffrs_0.nand3_7.C
rlabel metal2 -6187 9339 -6187 9339 5 SARlogic_0.dffrs_0.nand3_7.VSS
rlabel metal2 -7601 11288 -7601 11288 1 SARlogic_0.dffrs_0.nand3_6.VDD
rlabel metal1 -7191 10162 -7191 10162 3 SARlogic_0.dffrs_0.nand3_6.Z
rlabel metal1 -8277 10044 -8277 10044 7 SARlogic_0.dffrs_0.nand3_6.A
rlabel metal1 -8277 10163 -8277 10163 7 SARlogic_0.dffrs_0.nand3_6.B
rlabel metal1 -8277 10279 -8277 10279 7 SARlogic_0.dffrs_0.nand3_6.C
rlabel metal2 -7673 9338 -7673 9338 5 SARlogic_0.dffrs_0.nand3_6.VSS
rlabel metal2 -6115 13493 -6115 13493 1 SARlogic_0.dffrs_0.nand3_2.VDD
rlabel metal1 -5705 12367 -5705 12367 3 SARlogic_0.dffrs_0.nand3_2.Z
rlabel metal1 -6791 12249 -6791 12249 7 SARlogic_0.dffrs_0.nand3_2.A
rlabel metal1 -6791 12368 -6791 12368 7 SARlogic_0.dffrs_0.nand3_2.B
rlabel metal1 -6791 12484 -6791 12484 7 SARlogic_0.dffrs_0.nand3_2.C
rlabel metal2 -6187 11543 -6187 11543 5 SARlogic_0.dffrs_0.nand3_2.VSS
rlabel metal2 -7601 13493 -7601 13493 1 SARlogic_0.dffrs_0.nand3_1.VDD
rlabel metal1 -7191 12367 -7191 12367 3 SARlogic_0.dffrs_0.nand3_1.Z
rlabel metal1 -8277 12249 -8277 12249 7 SARlogic_0.dffrs_0.nand3_1.A
rlabel metal1 -8277 12368 -8277 12368 7 SARlogic_0.dffrs_0.nand3_1.B
rlabel metal1 -8277 12484 -8277 12484 7 SARlogic_0.dffrs_0.nand3_1.C
rlabel metal2 -7673 11543 -7673 11543 5 SARlogic_0.dffrs_0.nand3_1.VSS
rlabel metal2 -7601 15698 -7601 15698 1 SARlogic_0.dffrs_0.nand3_0.VDD
rlabel metal1 -7191 14572 -7191 14572 3 SARlogic_0.dffrs_0.nand3_0.Z
rlabel metal1 -8277 14454 -8277 14454 7 SARlogic_0.dffrs_0.nand3_0.A
rlabel metal1 -8277 14573 -8277 14573 7 SARlogic_0.dffrs_0.nand3_0.B
rlabel metal1 -8277 14689 -8277 14689 7 SARlogic_0.dffrs_0.nand3_0.C
rlabel metal2 -7673 13748 -7673 13748 5 SARlogic_0.dffrs_0.nand3_0.VSS
rlabel metal1 -12777 14689 -12777 14689 7 SARlogic_0.dffrs_13.setb
rlabel metal1 -12777 11466 -12777 11466 7 SARlogic_0.dffrs_13.clk
rlabel metal1 -12777 7841 -12777 7841 7 SARlogic_0.dffrs_13.d
rlabel metal1 -12760 7054 -12760 7054 7 SARlogic_0.dffrs_13.resetb
rlabel metal2 -9309 12368 -9309 12368 3 SARlogic_0.dffrs_13.Q
rlabel metal2 -9309 10163 -9309 10163 3 SARlogic_0.dffrs_13.Qb
rlabel metal5 -10669 15794 -10669 15794 1 SARlogic_0.dffrs_13.vdd
rlabel metal4 -10561 7015 -10561 7015 5 SARlogic_0.dffrs_13.vss
rlabel metal2 -11613 9083 -11613 9083 1 SARlogic_0.dffrs_13.nand3_8.VDD
rlabel metal1 -11203 7957 -11203 7957 3 SARlogic_0.dffrs_13.nand3_8.Z
rlabel metal1 -12289 7839 -12289 7839 7 SARlogic_0.dffrs_13.nand3_8.A
rlabel metal1 -12289 7958 -12289 7958 7 SARlogic_0.dffrs_13.nand3_8.B
rlabel metal1 -12289 8074 -12289 8074 7 SARlogic_0.dffrs_13.nand3_8.C
rlabel metal2 -11685 7133 -11685 7133 5 SARlogic_0.dffrs_13.nand3_8.VSS
rlabel metal2 -10127 11289 -10127 11289 1 SARlogic_0.dffrs_13.nand3_7.VDD
rlabel metal1 -9717 10163 -9717 10163 3 SARlogic_0.dffrs_13.nand3_7.Z
rlabel metal1 -10803 10045 -10803 10045 7 SARlogic_0.dffrs_13.nand3_7.A
rlabel metal1 -10803 10164 -10803 10164 7 SARlogic_0.dffrs_13.nand3_7.B
rlabel metal1 -10803 10280 -10803 10280 7 SARlogic_0.dffrs_13.nand3_7.C
rlabel metal2 -10199 9339 -10199 9339 5 SARlogic_0.dffrs_13.nand3_7.VSS
rlabel metal2 -11613 11288 -11613 11288 1 SARlogic_0.dffrs_13.nand3_6.VDD
rlabel metal1 -11203 10162 -11203 10162 3 SARlogic_0.dffrs_13.nand3_6.Z
rlabel metal1 -12289 10044 -12289 10044 7 SARlogic_0.dffrs_13.nand3_6.A
rlabel metal1 -12289 10163 -12289 10163 7 SARlogic_0.dffrs_13.nand3_6.B
rlabel metal1 -12289 10279 -12289 10279 7 SARlogic_0.dffrs_13.nand3_6.C
rlabel metal2 -11685 9338 -11685 9338 5 SARlogic_0.dffrs_13.nand3_6.VSS
rlabel metal2 -10127 13493 -10127 13493 1 SARlogic_0.dffrs_13.nand3_2.VDD
rlabel metal1 -9717 12367 -9717 12367 3 SARlogic_0.dffrs_13.nand3_2.Z
rlabel metal1 -10803 12249 -10803 12249 7 SARlogic_0.dffrs_13.nand3_2.A
rlabel metal1 -10803 12368 -10803 12368 7 SARlogic_0.dffrs_13.nand3_2.B
rlabel metal1 -10803 12484 -10803 12484 7 SARlogic_0.dffrs_13.nand3_2.C
rlabel metal2 -10199 11543 -10199 11543 5 SARlogic_0.dffrs_13.nand3_2.VSS
rlabel metal2 -11613 13493 -11613 13493 1 SARlogic_0.dffrs_13.nand3_1.VDD
rlabel metal1 -11203 12367 -11203 12367 3 SARlogic_0.dffrs_13.nand3_1.Z
rlabel metal1 -12289 12249 -12289 12249 7 SARlogic_0.dffrs_13.nand3_1.A
rlabel metal1 -12289 12368 -12289 12368 7 SARlogic_0.dffrs_13.nand3_1.B
rlabel metal1 -12289 12484 -12289 12484 7 SARlogic_0.dffrs_13.nand3_1.C
rlabel metal2 -11685 11543 -11685 11543 5 SARlogic_0.dffrs_13.nand3_1.VSS
rlabel metal2 -11613 15698 -11613 15698 1 SARlogic_0.dffrs_13.nand3_0.VDD
rlabel metal1 -11203 14572 -11203 14572 3 SARlogic_0.dffrs_13.nand3_0.Z
rlabel metal1 -12289 14454 -12289 14454 7 SARlogic_0.dffrs_13.nand3_0.A
rlabel metal1 -12289 14573 -12289 14573 7 SARlogic_0.dffrs_13.nand3_0.B
rlabel metal1 -12289 14689 -12289 14689 7 SARlogic_0.dffrs_13.nand3_0.C
rlabel metal2 -11685 13748 -11685 13748 5 SARlogic_0.dffrs_13.nand3_0.VSS
rlabel metal1 -681 14689 -681 14689 7 SARlogic_0.dffrs_2.setb
rlabel metal1 -681 11466 -681 11466 7 SARlogic_0.dffrs_2.clk
rlabel metal1 -681 7841 -681 7841 7 SARlogic_0.dffrs_2.d
rlabel metal1 -664 7054 -664 7054 7 SARlogic_0.dffrs_2.resetb
rlabel metal2 2787 12368 2787 12368 3 SARlogic_0.dffrs_2.Q
rlabel metal2 2787 10163 2787 10163 3 SARlogic_0.dffrs_2.Qb
rlabel metal5 1427 15794 1427 15794 1 SARlogic_0.dffrs_2.vdd
rlabel metal4 1535 7015 1535 7015 5 SARlogic_0.dffrs_2.vss
rlabel metal2 483 9083 483 9083 1 SARlogic_0.dffrs_2.nand3_8.VDD
rlabel metal1 893 7957 893 7957 3 SARlogic_0.dffrs_2.nand3_8.Z
rlabel metal1 -193 7839 -193 7839 7 SARlogic_0.dffrs_2.nand3_8.A
rlabel metal1 -193 7958 -193 7958 7 SARlogic_0.dffrs_2.nand3_8.B
rlabel metal1 -193 8074 -193 8074 7 SARlogic_0.dffrs_2.nand3_8.C
rlabel metal2 411 7133 411 7133 5 SARlogic_0.dffrs_2.nand3_8.VSS
rlabel metal2 1969 11289 1969 11289 1 SARlogic_0.dffrs_2.nand3_7.VDD
rlabel metal1 2379 10163 2379 10163 3 SARlogic_0.dffrs_2.nand3_7.Z
rlabel metal1 1293 10045 1293 10045 7 SARlogic_0.dffrs_2.nand3_7.A
rlabel metal1 1293 10164 1293 10164 7 SARlogic_0.dffrs_2.nand3_7.B
rlabel metal1 1293 10280 1293 10280 7 SARlogic_0.dffrs_2.nand3_7.C
rlabel metal2 1897 9339 1897 9339 5 SARlogic_0.dffrs_2.nand3_7.VSS
rlabel metal2 483 11288 483 11288 1 SARlogic_0.dffrs_2.nand3_6.VDD
rlabel metal1 893 10162 893 10162 3 SARlogic_0.dffrs_2.nand3_6.Z
rlabel metal1 -193 10044 -193 10044 7 SARlogic_0.dffrs_2.nand3_6.A
rlabel metal1 -193 10163 -193 10163 7 SARlogic_0.dffrs_2.nand3_6.B
rlabel metal1 -193 10279 -193 10279 7 SARlogic_0.dffrs_2.nand3_6.C
rlabel metal2 411 9338 411 9338 5 SARlogic_0.dffrs_2.nand3_6.VSS
rlabel metal2 1969 13493 1969 13493 1 SARlogic_0.dffrs_2.nand3_2.VDD
rlabel metal1 2379 12367 2379 12367 3 SARlogic_0.dffrs_2.nand3_2.Z
rlabel metal1 1293 12249 1293 12249 7 SARlogic_0.dffrs_2.nand3_2.A
rlabel metal1 1293 12368 1293 12368 7 SARlogic_0.dffrs_2.nand3_2.B
rlabel metal1 1293 12484 1293 12484 7 SARlogic_0.dffrs_2.nand3_2.C
rlabel metal2 1897 11543 1897 11543 5 SARlogic_0.dffrs_2.nand3_2.VSS
rlabel metal2 483 13493 483 13493 1 SARlogic_0.dffrs_2.nand3_1.VDD
rlabel metal1 893 12367 893 12367 3 SARlogic_0.dffrs_2.nand3_1.Z
rlabel metal1 -193 12249 -193 12249 7 SARlogic_0.dffrs_2.nand3_1.A
rlabel metal1 -193 12368 -193 12368 7 SARlogic_0.dffrs_2.nand3_1.B
rlabel metal1 -193 12484 -193 12484 7 SARlogic_0.dffrs_2.nand3_1.C
rlabel metal2 411 11543 411 11543 5 SARlogic_0.dffrs_2.nand3_1.VSS
rlabel metal2 483 15698 483 15698 1 SARlogic_0.dffrs_2.nand3_0.VDD
rlabel metal1 893 14572 893 14572 3 SARlogic_0.dffrs_2.nand3_0.Z
rlabel metal1 -193 14454 -193 14454 7 SARlogic_0.dffrs_2.nand3_0.A
rlabel metal1 -193 14573 -193 14573 7 SARlogic_0.dffrs_2.nand3_0.B
rlabel metal1 -193 14689 -193 14689 7 SARlogic_0.dffrs_2.nand3_0.C
rlabel metal2 411 13748 411 13748 5 SARlogic_0.dffrs_2.nand3_0.VSS
rlabel metal1 -4723 14689 -4723 14689 7 SARlogic_0.dffrs_1.setb
rlabel metal1 -4723 11466 -4723 11466 7 SARlogic_0.dffrs_1.clk
rlabel metal1 -4723 7841 -4723 7841 7 SARlogic_0.dffrs_1.d
rlabel metal1 -4706 7054 -4706 7054 7 SARlogic_0.dffrs_1.resetb
rlabel metal2 -1255 12368 -1255 12368 3 SARlogic_0.dffrs_1.Q
rlabel metal2 -1255 10163 -1255 10163 3 SARlogic_0.dffrs_1.Qb
rlabel metal5 -2615 15794 -2615 15794 1 SARlogic_0.dffrs_1.vdd
rlabel metal4 -2507 7015 -2507 7015 5 SARlogic_0.dffrs_1.vss
rlabel metal2 -3559 9083 -3559 9083 1 SARlogic_0.dffrs_1.nand3_8.VDD
rlabel metal1 -3149 7957 -3149 7957 3 SARlogic_0.dffrs_1.nand3_8.Z
rlabel metal1 -4235 7839 -4235 7839 7 SARlogic_0.dffrs_1.nand3_8.A
rlabel metal1 -4235 7958 -4235 7958 7 SARlogic_0.dffrs_1.nand3_8.B
rlabel metal1 -4235 8074 -4235 8074 7 SARlogic_0.dffrs_1.nand3_8.C
rlabel metal2 -3631 7133 -3631 7133 5 SARlogic_0.dffrs_1.nand3_8.VSS
rlabel metal2 -2073 11289 -2073 11289 1 SARlogic_0.dffrs_1.nand3_7.VDD
rlabel metal1 -1663 10163 -1663 10163 3 SARlogic_0.dffrs_1.nand3_7.Z
rlabel metal1 -2749 10045 -2749 10045 7 SARlogic_0.dffrs_1.nand3_7.A
rlabel metal1 -2749 10164 -2749 10164 7 SARlogic_0.dffrs_1.nand3_7.B
rlabel metal1 -2749 10280 -2749 10280 7 SARlogic_0.dffrs_1.nand3_7.C
rlabel metal2 -2145 9339 -2145 9339 5 SARlogic_0.dffrs_1.nand3_7.VSS
rlabel metal2 -3559 11288 -3559 11288 1 SARlogic_0.dffrs_1.nand3_6.VDD
rlabel metal1 -3149 10162 -3149 10162 3 SARlogic_0.dffrs_1.nand3_6.Z
rlabel metal1 -4235 10044 -4235 10044 7 SARlogic_0.dffrs_1.nand3_6.A
rlabel metal1 -4235 10163 -4235 10163 7 SARlogic_0.dffrs_1.nand3_6.B
rlabel metal1 -4235 10279 -4235 10279 7 SARlogic_0.dffrs_1.nand3_6.C
rlabel metal2 -3631 9338 -3631 9338 5 SARlogic_0.dffrs_1.nand3_6.VSS
rlabel metal2 -2073 13493 -2073 13493 1 SARlogic_0.dffrs_1.nand3_2.VDD
rlabel metal1 -1663 12367 -1663 12367 3 SARlogic_0.dffrs_1.nand3_2.Z
rlabel metal1 -2749 12249 -2749 12249 7 SARlogic_0.dffrs_1.nand3_2.A
rlabel metal1 -2749 12368 -2749 12368 7 SARlogic_0.dffrs_1.nand3_2.B
rlabel metal1 -2749 12484 -2749 12484 7 SARlogic_0.dffrs_1.nand3_2.C
rlabel metal2 -2145 11543 -2145 11543 5 SARlogic_0.dffrs_1.nand3_2.VSS
rlabel metal2 -3559 13493 -3559 13493 1 SARlogic_0.dffrs_1.nand3_1.VDD
rlabel metal1 -3149 12367 -3149 12367 3 SARlogic_0.dffrs_1.nand3_1.Z
rlabel metal1 -4235 12249 -4235 12249 7 SARlogic_0.dffrs_1.nand3_1.A
rlabel metal1 -4235 12368 -4235 12368 7 SARlogic_0.dffrs_1.nand3_1.B
rlabel metal1 -4235 12484 -4235 12484 7 SARlogic_0.dffrs_1.nand3_1.C
rlabel metal2 -3631 11543 -3631 11543 5 SARlogic_0.dffrs_1.nand3_1.VSS
rlabel metal2 -3559 15698 -3559 15698 1 SARlogic_0.dffrs_1.nand3_0.VDD
rlabel metal1 -3149 14572 -3149 14572 3 SARlogic_0.dffrs_1.nand3_0.Z
rlabel metal1 -4235 14454 -4235 14454 7 SARlogic_0.dffrs_1.nand3_0.A
rlabel metal1 -4235 14573 -4235 14573 7 SARlogic_0.dffrs_1.nand3_0.B
rlabel metal1 -4235 14689 -4235 14689 7 SARlogic_0.dffrs_1.nand3_0.C
rlabel metal2 -3631 13748 -3631 13748 5 SARlogic_0.dffrs_1.nand3_0.VSS
rlabel metal1 7403 14689 7403 14689 7 SARlogic_0.dffrs_4.setb
rlabel metal1 7403 11466 7403 11466 7 SARlogic_0.dffrs_4.clk
rlabel metal1 7403 7841 7403 7841 7 SARlogic_0.dffrs_4.d
rlabel metal1 7420 7054 7420 7054 7 SARlogic_0.dffrs_4.resetb
rlabel metal2 10871 12368 10871 12368 3 SARlogic_0.dffrs_4.Q
rlabel metal2 10871 10163 10871 10163 3 SARlogic_0.dffrs_4.Qb
rlabel metal5 9511 15794 9511 15794 1 SARlogic_0.dffrs_4.vdd
rlabel metal4 9619 7015 9619 7015 5 SARlogic_0.dffrs_4.vss
rlabel metal2 8567 9083 8567 9083 1 SARlogic_0.dffrs_4.nand3_8.VDD
rlabel metal1 8977 7957 8977 7957 3 SARlogic_0.dffrs_4.nand3_8.Z
rlabel metal1 7891 7839 7891 7839 7 SARlogic_0.dffrs_4.nand3_8.A
rlabel metal1 7891 7958 7891 7958 7 SARlogic_0.dffrs_4.nand3_8.B
rlabel metal1 7891 8074 7891 8074 7 SARlogic_0.dffrs_4.nand3_8.C
rlabel metal2 8495 7133 8495 7133 5 SARlogic_0.dffrs_4.nand3_8.VSS
rlabel metal2 10053 11289 10053 11289 1 SARlogic_0.dffrs_4.nand3_7.VDD
rlabel metal1 10463 10163 10463 10163 3 SARlogic_0.dffrs_4.nand3_7.Z
rlabel metal1 9377 10045 9377 10045 7 SARlogic_0.dffrs_4.nand3_7.A
rlabel metal1 9377 10164 9377 10164 7 SARlogic_0.dffrs_4.nand3_7.B
rlabel metal1 9377 10280 9377 10280 7 SARlogic_0.dffrs_4.nand3_7.C
rlabel metal2 9981 9339 9981 9339 5 SARlogic_0.dffrs_4.nand3_7.VSS
rlabel metal2 8567 11288 8567 11288 1 SARlogic_0.dffrs_4.nand3_6.VDD
rlabel metal1 8977 10162 8977 10162 3 SARlogic_0.dffrs_4.nand3_6.Z
rlabel metal1 7891 10044 7891 10044 7 SARlogic_0.dffrs_4.nand3_6.A
rlabel metal1 7891 10163 7891 10163 7 SARlogic_0.dffrs_4.nand3_6.B
rlabel metal1 7891 10279 7891 10279 7 SARlogic_0.dffrs_4.nand3_6.C
rlabel metal2 8495 9338 8495 9338 5 SARlogic_0.dffrs_4.nand3_6.VSS
rlabel metal2 10053 13493 10053 13493 1 SARlogic_0.dffrs_4.nand3_2.VDD
rlabel metal1 10463 12367 10463 12367 3 SARlogic_0.dffrs_4.nand3_2.Z
rlabel metal1 9377 12249 9377 12249 7 SARlogic_0.dffrs_4.nand3_2.A
rlabel metal1 9377 12368 9377 12368 7 SARlogic_0.dffrs_4.nand3_2.B
rlabel metal1 9377 12484 9377 12484 7 SARlogic_0.dffrs_4.nand3_2.C
rlabel metal2 9981 11543 9981 11543 5 SARlogic_0.dffrs_4.nand3_2.VSS
rlabel metal2 8567 13493 8567 13493 1 SARlogic_0.dffrs_4.nand3_1.VDD
rlabel metal1 8977 12367 8977 12367 3 SARlogic_0.dffrs_4.nand3_1.Z
rlabel metal1 7891 12249 7891 12249 7 SARlogic_0.dffrs_4.nand3_1.A
rlabel metal1 7891 12368 7891 12368 7 SARlogic_0.dffrs_4.nand3_1.B
rlabel metal1 7891 12484 7891 12484 7 SARlogic_0.dffrs_4.nand3_1.C
rlabel metal2 8495 11543 8495 11543 5 SARlogic_0.dffrs_4.nand3_1.VSS
rlabel metal2 8567 15698 8567 15698 1 SARlogic_0.dffrs_4.nand3_0.VDD
rlabel metal1 8977 14572 8977 14572 3 SARlogic_0.dffrs_4.nand3_0.Z
rlabel metal1 7891 14454 7891 14454 7 SARlogic_0.dffrs_4.nand3_0.A
rlabel metal1 7891 14573 7891 14573 7 SARlogic_0.dffrs_4.nand3_0.B
rlabel metal1 7891 14689 7891 14689 7 SARlogic_0.dffrs_4.nand3_0.C
rlabel metal2 8495 13748 8495 13748 5 SARlogic_0.dffrs_4.nand3_0.VSS
rlabel metal1 3361 14689 3361 14689 7 SARlogic_0.dffrs_3.setb
rlabel metal1 3361 11466 3361 11466 7 SARlogic_0.dffrs_3.clk
rlabel metal1 3361 7841 3361 7841 7 SARlogic_0.dffrs_3.d
rlabel metal1 3378 7054 3378 7054 7 SARlogic_0.dffrs_3.resetb
rlabel metal2 6829 12368 6829 12368 3 SARlogic_0.dffrs_3.Q
rlabel metal2 6829 10163 6829 10163 3 SARlogic_0.dffrs_3.Qb
rlabel metal5 5469 15794 5469 15794 1 SARlogic_0.dffrs_3.vdd
rlabel metal4 5577 7015 5577 7015 5 SARlogic_0.dffrs_3.vss
rlabel metal2 4525 9083 4525 9083 1 SARlogic_0.dffrs_3.nand3_8.VDD
rlabel metal1 4935 7957 4935 7957 3 SARlogic_0.dffrs_3.nand3_8.Z
rlabel metal1 3849 7839 3849 7839 7 SARlogic_0.dffrs_3.nand3_8.A
rlabel metal1 3849 7958 3849 7958 7 SARlogic_0.dffrs_3.nand3_8.B
rlabel metal1 3849 8074 3849 8074 7 SARlogic_0.dffrs_3.nand3_8.C
rlabel metal2 4453 7133 4453 7133 5 SARlogic_0.dffrs_3.nand3_8.VSS
rlabel metal2 6011 11289 6011 11289 1 SARlogic_0.dffrs_3.nand3_7.VDD
rlabel metal1 6421 10163 6421 10163 3 SARlogic_0.dffrs_3.nand3_7.Z
rlabel metal1 5335 10045 5335 10045 7 SARlogic_0.dffrs_3.nand3_7.A
rlabel metal1 5335 10164 5335 10164 7 SARlogic_0.dffrs_3.nand3_7.B
rlabel metal1 5335 10280 5335 10280 7 SARlogic_0.dffrs_3.nand3_7.C
rlabel metal2 5939 9339 5939 9339 5 SARlogic_0.dffrs_3.nand3_7.VSS
rlabel metal2 4525 11288 4525 11288 1 SARlogic_0.dffrs_3.nand3_6.VDD
rlabel metal1 4935 10162 4935 10162 3 SARlogic_0.dffrs_3.nand3_6.Z
rlabel metal1 3849 10044 3849 10044 7 SARlogic_0.dffrs_3.nand3_6.A
rlabel metal1 3849 10163 3849 10163 7 SARlogic_0.dffrs_3.nand3_6.B
rlabel metal1 3849 10279 3849 10279 7 SARlogic_0.dffrs_3.nand3_6.C
rlabel metal2 4453 9338 4453 9338 5 SARlogic_0.dffrs_3.nand3_6.VSS
rlabel metal2 6011 13493 6011 13493 1 SARlogic_0.dffrs_3.nand3_2.VDD
rlabel metal1 6421 12367 6421 12367 3 SARlogic_0.dffrs_3.nand3_2.Z
rlabel metal1 5335 12249 5335 12249 7 SARlogic_0.dffrs_3.nand3_2.A
rlabel metal1 5335 12368 5335 12368 7 SARlogic_0.dffrs_3.nand3_2.B
rlabel metal1 5335 12484 5335 12484 7 SARlogic_0.dffrs_3.nand3_2.C
rlabel metal2 5939 11543 5939 11543 5 SARlogic_0.dffrs_3.nand3_2.VSS
rlabel metal2 4525 13493 4525 13493 1 SARlogic_0.dffrs_3.nand3_1.VDD
rlabel metal1 4935 12367 4935 12367 3 SARlogic_0.dffrs_3.nand3_1.Z
rlabel metal1 3849 12249 3849 12249 7 SARlogic_0.dffrs_3.nand3_1.A
rlabel metal1 3849 12368 3849 12368 7 SARlogic_0.dffrs_3.nand3_1.B
rlabel metal1 3849 12484 3849 12484 7 SARlogic_0.dffrs_3.nand3_1.C
rlabel metal2 4453 11543 4453 11543 5 SARlogic_0.dffrs_3.nand3_1.VSS
rlabel metal2 4525 15698 4525 15698 1 SARlogic_0.dffrs_3.nand3_0.VDD
rlabel metal1 4935 14572 4935 14572 3 SARlogic_0.dffrs_3.nand3_0.Z
rlabel metal1 3849 14454 3849 14454 7 SARlogic_0.dffrs_3.nand3_0.A
rlabel metal1 3849 14573 3849 14573 7 SARlogic_0.dffrs_3.nand3_0.B
rlabel metal1 3849 14689 3849 14689 7 SARlogic_0.dffrs_3.nand3_0.C
rlabel metal2 4453 13748 4453 13748 5 SARlogic_0.dffrs_3.nand3_0.VSS
rlabel metal1 11445 14689 11445 14689 7 SARlogic_0.dffrs_5.setb
rlabel metal1 11445 11466 11445 11466 7 SARlogic_0.dffrs_5.clk
rlabel metal1 11445 7841 11445 7841 7 SARlogic_0.dffrs_5.d
rlabel metal1 11462 7054 11462 7054 7 SARlogic_0.dffrs_5.resetb
rlabel metal2 14913 12368 14913 12368 3 SARlogic_0.dffrs_5.Q
rlabel metal2 14913 10163 14913 10163 3 SARlogic_0.dffrs_5.Qb
rlabel metal5 13553 15794 13553 15794 1 SARlogic_0.dffrs_5.vdd
rlabel metal4 13661 7015 13661 7015 5 SARlogic_0.dffrs_5.vss
rlabel metal2 12609 9083 12609 9083 1 SARlogic_0.dffrs_5.nand3_8.VDD
rlabel metal1 13019 7957 13019 7957 3 SARlogic_0.dffrs_5.nand3_8.Z
rlabel metal1 11933 7839 11933 7839 7 SARlogic_0.dffrs_5.nand3_8.A
rlabel metal1 11933 7958 11933 7958 7 SARlogic_0.dffrs_5.nand3_8.B
rlabel metal1 11933 8074 11933 8074 7 SARlogic_0.dffrs_5.nand3_8.C
rlabel metal2 12537 7133 12537 7133 5 SARlogic_0.dffrs_5.nand3_8.VSS
rlabel metal2 14095 11289 14095 11289 1 SARlogic_0.dffrs_5.nand3_7.VDD
rlabel metal1 14505 10163 14505 10163 3 SARlogic_0.dffrs_5.nand3_7.Z
rlabel metal1 13419 10045 13419 10045 7 SARlogic_0.dffrs_5.nand3_7.A
rlabel metal1 13419 10164 13419 10164 7 SARlogic_0.dffrs_5.nand3_7.B
rlabel metal1 13419 10280 13419 10280 7 SARlogic_0.dffrs_5.nand3_7.C
rlabel metal2 14023 9339 14023 9339 5 SARlogic_0.dffrs_5.nand3_7.VSS
rlabel metal2 12609 11288 12609 11288 1 SARlogic_0.dffrs_5.nand3_6.VDD
rlabel metal1 13019 10162 13019 10162 3 SARlogic_0.dffrs_5.nand3_6.Z
rlabel metal1 11933 10044 11933 10044 7 SARlogic_0.dffrs_5.nand3_6.A
rlabel metal1 11933 10163 11933 10163 7 SARlogic_0.dffrs_5.nand3_6.B
rlabel metal1 11933 10279 11933 10279 7 SARlogic_0.dffrs_5.nand3_6.C
rlabel metal2 12537 9338 12537 9338 5 SARlogic_0.dffrs_5.nand3_6.VSS
rlabel metal2 14095 13493 14095 13493 1 SARlogic_0.dffrs_5.nand3_2.VDD
rlabel metal1 14505 12367 14505 12367 3 SARlogic_0.dffrs_5.nand3_2.Z
rlabel metal1 13419 12249 13419 12249 7 SARlogic_0.dffrs_5.nand3_2.A
rlabel metal1 13419 12368 13419 12368 7 SARlogic_0.dffrs_5.nand3_2.B
rlabel metal1 13419 12484 13419 12484 7 SARlogic_0.dffrs_5.nand3_2.C
rlabel metal2 14023 11543 14023 11543 5 SARlogic_0.dffrs_5.nand3_2.VSS
rlabel metal2 12609 13493 12609 13493 1 SARlogic_0.dffrs_5.nand3_1.VDD
rlabel metal1 13019 12367 13019 12367 3 SARlogic_0.dffrs_5.nand3_1.Z
rlabel metal1 11933 12249 11933 12249 7 SARlogic_0.dffrs_5.nand3_1.A
rlabel metal1 11933 12368 11933 12368 7 SARlogic_0.dffrs_5.nand3_1.B
rlabel metal1 11933 12484 11933 12484 7 SARlogic_0.dffrs_5.nand3_1.C
rlabel metal2 12537 11543 12537 11543 5 SARlogic_0.dffrs_5.nand3_1.VSS
rlabel metal2 12609 15698 12609 15698 1 SARlogic_0.dffrs_5.nand3_0.VDD
rlabel metal1 13019 14572 13019 14572 3 SARlogic_0.dffrs_5.nand3_0.Z
rlabel metal1 11933 14454 11933 14454 7 SARlogic_0.dffrs_5.nand3_0.A
rlabel metal1 11933 14573 11933 14573 7 SARlogic_0.dffrs_5.nand3_0.B
rlabel metal1 11933 14689 11933 14689 7 SARlogic_0.dffrs_5.nand3_0.C
rlabel metal2 12537 13748 12537 13748 5 SARlogic_0.dffrs_5.nand3_0.VSS
rlabel metal1 -8765 24268 -8765 24268 7 SARlogic_0.dffrs_14.setb
rlabel metal1 -8765 21045 -8765 21045 7 SARlogic_0.dffrs_14.clk
rlabel metal1 -8765 17420 -8765 17420 7 SARlogic_0.dffrs_14.d
rlabel metal1 -8748 16633 -8748 16633 7 SARlogic_0.dffrs_14.resetb
rlabel metal2 -5297 21947 -5297 21947 3 SARlogic_0.dffrs_14.Q
rlabel metal2 -5297 19742 -5297 19742 3 SARlogic_0.dffrs_14.Qb
rlabel metal5 -6657 25373 -6657 25373 1 SARlogic_0.dffrs_14.vdd
rlabel metal4 -6549 16594 -6549 16594 5 SARlogic_0.dffrs_14.vss
rlabel metal2 -7601 18662 -7601 18662 1 SARlogic_0.dffrs_14.nand3_8.VDD
rlabel metal1 -7191 17536 -7191 17536 3 SARlogic_0.dffrs_14.nand3_8.Z
rlabel metal1 -8277 17418 -8277 17418 7 SARlogic_0.dffrs_14.nand3_8.A
rlabel metal1 -8277 17537 -8277 17537 7 SARlogic_0.dffrs_14.nand3_8.B
rlabel metal1 -8277 17653 -8277 17653 7 SARlogic_0.dffrs_14.nand3_8.C
rlabel metal2 -7673 16712 -7673 16712 5 SARlogic_0.dffrs_14.nand3_8.VSS
rlabel metal2 -6115 20868 -6115 20868 1 SARlogic_0.dffrs_14.nand3_7.VDD
rlabel metal1 -5705 19742 -5705 19742 3 SARlogic_0.dffrs_14.nand3_7.Z
rlabel metal1 -6791 19624 -6791 19624 7 SARlogic_0.dffrs_14.nand3_7.A
rlabel metal1 -6791 19743 -6791 19743 7 SARlogic_0.dffrs_14.nand3_7.B
rlabel metal1 -6791 19859 -6791 19859 7 SARlogic_0.dffrs_14.nand3_7.C
rlabel metal2 -6187 18918 -6187 18918 5 SARlogic_0.dffrs_14.nand3_7.VSS
rlabel metal2 -7601 20867 -7601 20867 1 SARlogic_0.dffrs_14.nand3_6.VDD
rlabel metal1 -7191 19741 -7191 19741 3 SARlogic_0.dffrs_14.nand3_6.Z
rlabel metal1 -8277 19623 -8277 19623 7 SARlogic_0.dffrs_14.nand3_6.A
rlabel metal1 -8277 19742 -8277 19742 7 SARlogic_0.dffrs_14.nand3_6.B
rlabel metal1 -8277 19858 -8277 19858 7 SARlogic_0.dffrs_14.nand3_6.C
rlabel metal2 -7673 18917 -7673 18917 5 SARlogic_0.dffrs_14.nand3_6.VSS
rlabel metal2 -6115 23072 -6115 23072 1 SARlogic_0.dffrs_14.nand3_2.VDD
rlabel metal1 -5705 21946 -5705 21946 3 SARlogic_0.dffrs_14.nand3_2.Z
rlabel metal1 -6791 21828 -6791 21828 7 SARlogic_0.dffrs_14.nand3_2.A
rlabel metal1 -6791 21947 -6791 21947 7 SARlogic_0.dffrs_14.nand3_2.B
rlabel metal1 -6791 22063 -6791 22063 7 SARlogic_0.dffrs_14.nand3_2.C
rlabel metal2 -6187 21122 -6187 21122 5 SARlogic_0.dffrs_14.nand3_2.VSS
rlabel metal2 -7601 23072 -7601 23072 1 SARlogic_0.dffrs_14.nand3_1.VDD
rlabel metal1 -7191 21946 -7191 21946 3 SARlogic_0.dffrs_14.nand3_1.Z
rlabel metal1 -8277 21828 -8277 21828 7 SARlogic_0.dffrs_14.nand3_1.A
rlabel metal1 -8277 21947 -8277 21947 7 SARlogic_0.dffrs_14.nand3_1.B
rlabel metal1 -8277 22063 -8277 22063 7 SARlogic_0.dffrs_14.nand3_1.C
rlabel metal2 -7673 21122 -7673 21122 5 SARlogic_0.dffrs_14.nand3_1.VSS
rlabel metal2 -7601 25277 -7601 25277 1 SARlogic_0.dffrs_14.nand3_0.VDD
rlabel metal1 -7191 24151 -7191 24151 3 SARlogic_0.dffrs_14.nand3_0.Z
rlabel metal1 -8277 24033 -8277 24033 7 SARlogic_0.dffrs_14.nand3_0.A
rlabel metal1 -8277 24152 -8277 24152 7 SARlogic_0.dffrs_14.nand3_0.B
rlabel metal1 -8277 24268 -8277 24268 7 SARlogic_0.dffrs_14.nand3_0.C
rlabel metal2 -7673 23327 -7673 23327 5 SARlogic_0.dffrs_14.nand3_0.VSS
rlabel metal1 -681 24265 -681 24265 7 SARlogic_0.dffrs_8.setb
rlabel metal1 -681 21042 -681 21042 7 SARlogic_0.dffrs_8.clk
rlabel metal1 -681 17417 -681 17417 7 SARlogic_0.dffrs_8.d
rlabel metal1 -664 16630 -664 16630 7 SARlogic_0.dffrs_8.resetb
rlabel metal2 2787 21944 2787 21944 3 SARlogic_0.dffrs_8.Q
rlabel metal2 2787 19739 2787 19739 3 SARlogic_0.dffrs_8.Qb
rlabel metal5 1427 25370 1427 25370 1 SARlogic_0.dffrs_8.vdd
rlabel metal4 1535 16591 1535 16591 5 SARlogic_0.dffrs_8.vss
rlabel metal2 483 18659 483 18659 1 SARlogic_0.dffrs_8.nand3_8.VDD
rlabel metal1 893 17533 893 17533 3 SARlogic_0.dffrs_8.nand3_8.Z
rlabel metal1 -193 17415 -193 17415 7 SARlogic_0.dffrs_8.nand3_8.A
rlabel metal1 -193 17534 -193 17534 7 SARlogic_0.dffrs_8.nand3_8.B
rlabel metal1 -193 17650 -193 17650 7 SARlogic_0.dffrs_8.nand3_8.C
rlabel metal2 411 16709 411 16709 5 SARlogic_0.dffrs_8.nand3_8.VSS
rlabel metal2 1969 20865 1969 20865 1 SARlogic_0.dffrs_8.nand3_7.VDD
rlabel metal1 2379 19739 2379 19739 3 SARlogic_0.dffrs_8.nand3_7.Z
rlabel metal1 1293 19621 1293 19621 7 SARlogic_0.dffrs_8.nand3_7.A
rlabel metal1 1293 19740 1293 19740 7 SARlogic_0.dffrs_8.nand3_7.B
rlabel metal1 1293 19856 1293 19856 7 SARlogic_0.dffrs_8.nand3_7.C
rlabel metal2 1897 18915 1897 18915 5 SARlogic_0.dffrs_8.nand3_7.VSS
rlabel metal2 483 20864 483 20864 1 SARlogic_0.dffrs_8.nand3_6.VDD
rlabel metal1 893 19738 893 19738 3 SARlogic_0.dffrs_8.nand3_6.Z
rlabel metal1 -193 19620 -193 19620 7 SARlogic_0.dffrs_8.nand3_6.A
rlabel metal1 -193 19739 -193 19739 7 SARlogic_0.dffrs_8.nand3_6.B
rlabel metal1 -193 19855 -193 19855 7 SARlogic_0.dffrs_8.nand3_6.C
rlabel metal2 411 18914 411 18914 5 SARlogic_0.dffrs_8.nand3_6.VSS
rlabel metal2 1969 23069 1969 23069 1 SARlogic_0.dffrs_8.nand3_2.VDD
rlabel metal1 2379 21943 2379 21943 3 SARlogic_0.dffrs_8.nand3_2.Z
rlabel metal1 1293 21825 1293 21825 7 SARlogic_0.dffrs_8.nand3_2.A
rlabel metal1 1293 21944 1293 21944 7 SARlogic_0.dffrs_8.nand3_2.B
rlabel metal1 1293 22060 1293 22060 7 SARlogic_0.dffrs_8.nand3_2.C
rlabel metal2 1897 21119 1897 21119 5 SARlogic_0.dffrs_8.nand3_2.VSS
rlabel metal2 483 23069 483 23069 1 SARlogic_0.dffrs_8.nand3_1.VDD
rlabel metal1 893 21943 893 21943 3 SARlogic_0.dffrs_8.nand3_1.Z
rlabel metal1 -193 21825 -193 21825 7 SARlogic_0.dffrs_8.nand3_1.A
rlabel metal1 -193 21944 -193 21944 7 SARlogic_0.dffrs_8.nand3_1.B
rlabel metal1 -193 22060 -193 22060 7 SARlogic_0.dffrs_8.nand3_1.C
rlabel metal2 411 21119 411 21119 5 SARlogic_0.dffrs_8.nand3_1.VSS
rlabel metal2 483 25274 483 25274 1 SARlogic_0.dffrs_8.nand3_0.VDD
rlabel metal1 893 24148 893 24148 3 SARlogic_0.dffrs_8.nand3_0.Z
rlabel metal1 -193 24030 -193 24030 7 SARlogic_0.dffrs_8.nand3_0.A
rlabel metal1 -193 24149 -193 24149 7 SARlogic_0.dffrs_8.nand3_0.B
rlabel metal1 -193 24265 -193 24265 7 SARlogic_0.dffrs_8.nand3_0.C
rlabel metal2 411 23324 411 23324 5 SARlogic_0.dffrs_8.nand3_0.VSS
rlabel metal1 -4723 24265 -4723 24265 7 SARlogic_0.dffrs_7.setb
rlabel metal1 -4723 21042 -4723 21042 7 SARlogic_0.dffrs_7.clk
rlabel metal1 -4723 17417 -4723 17417 7 SARlogic_0.dffrs_7.d
rlabel metal1 -4706 16630 -4706 16630 7 SARlogic_0.dffrs_7.resetb
rlabel metal2 -1255 21944 -1255 21944 3 SARlogic_0.dffrs_7.Q
rlabel metal2 -1255 19739 -1255 19739 3 SARlogic_0.dffrs_7.Qb
rlabel metal5 -2615 25370 -2615 25370 1 SARlogic_0.dffrs_7.vdd
rlabel metal4 -2507 16591 -2507 16591 5 SARlogic_0.dffrs_7.vss
rlabel metal2 -3559 18659 -3559 18659 1 SARlogic_0.dffrs_7.nand3_8.VDD
rlabel metal1 -3149 17533 -3149 17533 3 SARlogic_0.dffrs_7.nand3_8.Z
rlabel metal1 -4235 17415 -4235 17415 7 SARlogic_0.dffrs_7.nand3_8.A
rlabel metal1 -4235 17534 -4235 17534 7 SARlogic_0.dffrs_7.nand3_8.B
rlabel metal1 -4235 17650 -4235 17650 7 SARlogic_0.dffrs_7.nand3_8.C
rlabel metal2 -3631 16709 -3631 16709 5 SARlogic_0.dffrs_7.nand3_8.VSS
rlabel metal2 -2073 20865 -2073 20865 1 SARlogic_0.dffrs_7.nand3_7.VDD
rlabel metal1 -1663 19739 -1663 19739 3 SARlogic_0.dffrs_7.nand3_7.Z
rlabel metal1 -2749 19621 -2749 19621 7 SARlogic_0.dffrs_7.nand3_7.A
rlabel metal1 -2749 19740 -2749 19740 7 SARlogic_0.dffrs_7.nand3_7.B
rlabel metal1 -2749 19856 -2749 19856 7 SARlogic_0.dffrs_7.nand3_7.C
rlabel metal2 -2145 18915 -2145 18915 5 SARlogic_0.dffrs_7.nand3_7.VSS
rlabel metal2 -3559 20864 -3559 20864 1 SARlogic_0.dffrs_7.nand3_6.VDD
rlabel metal1 -3149 19738 -3149 19738 3 SARlogic_0.dffrs_7.nand3_6.Z
rlabel metal1 -4235 19620 -4235 19620 7 SARlogic_0.dffrs_7.nand3_6.A
rlabel metal1 -4235 19739 -4235 19739 7 SARlogic_0.dffrs_7.nand3_6.B
rlabel metal1 -4235 19855 -4235 19855 7 SARlogic_0.dffrs_7.nand3_6.C
rlabel metal2 -3631 18914 -3631 18914 5 SARlogic_0.dffrs_7.nand3_6.VSS
rlabel metal2 -2073 23069 -2073 23069 1 SARlogic_0.dffrs_7.nand3_2.VDD
rlabel metal1 -1663 21943 -1663 21943 3 SARlogic_0.dffrs_7.nand3_2.Z
rlabel metal1 -2749 21825 -2749 21825 7 SARlogic_0.dffrs_7.nand3_2.A
rlabel metal1 -2749 21944 -2749 21944 7 SARlogic_0.dffrs_7.nand3_2.B
rlabel metal1 -2749 22060 -2749 22060 7 SARlogic_0.dffrs_7.nand3_2.C
rlabel metal2 -2145 21119 -2145 21119 5 SARlogic_0.dffrs_7.nand3_2.VSS
rlabel metal2 -3559 23069 -3559 23069 1 SARlogic_0.dffrs_7.nand3_1.VDD
rlabel metal1 -3149 21943 -3149 21943 3 SARlogic_0.dffrs_7.nand3_1.Z
rlabel metal1 -4235 21825 -4235 21825 7 SARlogic_0.dffrs_7.nand3_1.A
rlabel metal1 -4235 21944 -4235 21944 7 SARlogic_0.dffrs_7.nand3_1.B
rlabel metal1 -4235 22060 -4235 22060 7 SARlogic_0.dffrs_7.nand3_1.C
rlabel metal2 -3631 21119 -3631 21119 5 SARlogic_0.dffrs_7.nand3_1.VSS
rlabel metal2 -3559 25274 -3559 25274 1 SARlogic_0.dffrs_7.nand3_0.VDD
rlabel metal1 -3149 24148 -3149 24148 3 SARlogic_0.dffrs_7.nand3_0.Z
rlabel metal1 -4235 24030 -4235 24030 7 SARlogic_0.dffrs_7.nand3_0.A
rlabel metal1 -4235 24149 -4235 24149 7 SARlogic_0.dffrs_7.nand3_0.B
rlabel metal1 -4235 24265 -4235 24265 7 SARlogic_0.dffrs_7.nand3_0.C
rlabel metal2 -3631 23324 -3631 23324 5 SARlogic_0.dffrs_7.nand3_0.VSS
rlabel metal1 7403 24265 7403 24265 7 SARlogic_0.dffrs_10.setb
rlabel metal1 7403 21042 7403 21042 7 SARlogic_0.dffrs_10.clk
rlabel metal1 7403 17417 7403 17417 7 SARlogic_0.dffrs_10.d
rlabel metal1 7420 16630 7420 16630 7 SARlogic_0.dffrs_10.resetb
rlabel metal2 10871 21944 10871 21944 3 SARlogic_0.dffrs_10.Q
rlabel metal2 10871 19739 10871 19739 3 SARlogic_0.dffrs_10.Qb
rlabel metal5 9511 25370 9511 25370 1 SARlogic_0.dffrs_10.vdd
rlabel metal4 9619 16591 9619 16591 5 SARlogic_0.dffrs_10.vss
rlabel metal2 8567 18659 8567 18659 1 SARlogic_0.dffrs_10.nand3_8.VDD
rlabel metal1 8977 17533 8977 17533 3 SARlogic_0.dffrs_10.nand3_8.Z
rlabel metal1 7891 17415 7891 17415 7 SARlogic_0.dffrs_10.nand3_8.A
rlabel metal1 7891 17534 7891 17534 7 SARlogic_0.dffrs_10.nand3_8.B
rlabel metal1 7891 17650 7891 17650 7 SARlogic_0.dffrs_10.nand3_8.C
rlabel metal2 8495 16709 8495 16709 5 SARlogic_0.dffrs_10.nand3_8.VSS
rlabel metal2 10053 20865 10053 20865 1 SARlogic_0.dffrs_10.nand3_7.VDD
rlabel metal1 10463 19739 10463 19739 3 SARlogic_0.dffrs_10.nand3_7.Z
rlabel metal1 9377 19621 9377 19621 7 SARlogic_0.dffrs_10.nand3_7.A
rlabel metal1 9377 19740 9377 19740 7 SARlogic_0.dffrs_10.nand3_7.B
rlabel metal1 9377 19856 9377 19856 7 SARlogic_0.dffrs_10.nand3_7.C
rlabel metal2 9981 18915 9981 18915 5 SARlogic_0.dffrs_10.nand3_7.VSS
rlabel metal2 8567 20864 8567 20864 1 SARlogic_0.dffrs_10.nand3_6.VDD
rlabel metal1 8977 19738 8977 19738 3 SARlogic_0.dffrs_10.nand3_6.Z
rlabel metal1 7891 19620 7891 19620 7 SARlogic_0.dffrs_10.nand3_6.A
rlabel metal1 7891 19739 7891 19739 7 SARlogic_0.dffrs_10.nand3_6.B
rlabel metal1 7891 19855 7891 19855 7 SARlogic_0.dffrs_10.nand3_6.C
rlabel metal2 8495 18914 8495 18914 5 SARlogic_0.dffrs_10.nand3_6.VSS
rlabel metal2 10053 23069 10053 23069 1 SARlogic_0.dffrs_10.nand3_2.VDD
rlabel metal1 10463 21943 10463 21943 3 SARlogic_0.dffrs_10.nand3_2.Z
rlabel metal1 9377 21825 9377 21825 7 SARlogic_0.dffrs_10.nand3_2.A
rlabel metal1 9377 21944 9377 21944 7 SARlogic_0.dffrs_10.nand3_2.B
rlabel metal1 9377 22060 9377 22060 7 SARlogic_0.dffrs_10.nand3_2.C
rlabel metal2 9981 21119 9981 21119 5 SARlogic_0.dffrs_10.nand3_2.VSS
rlabel metal2 8567 23069 8567 23069 1 SARlogic_0.dffrs_10.nand3_1.VDD
rlabel metal1 8977 21943 8977 21943 3 SARlogic_0.dffrs_10.nand3_1.Z
rlabel metal1 7891 21825 7891 21825 7 SARlogic_0.dffrs_10.nand3_1.A
rlabel metal1 7891 21944 7891 21944 7 SARlogic_0.dffrs_10.nand3_1.B
rlabel metal1 7891 22060 7891 22060 7 SARlogic_0.dffrs_10.nand3_1.C
rlabel metal2 8495 21119 8495 21119 5 SARlogic_0.dffrs_10.nand3_1.VSS
rlabel metal2 8567 25274 8567 25274 1 SARlogic_0.dffrs_10.nand3_0.VDD
rlabel metal1 8977 24148 8977 24148 3 SARlogic_0.dffrs_10.nand3_0.Z
rlabel metal1 7891 24030 7891 24030 7 SARlogic_0.dffrs_10.nand3_0.A
rlabel metal1 7891 24149 7891 24149 7 SARlogic_0.dffrs_10.nand3_0.B
rlabel metal1 7891 24265 7891 24265 7 SARlogic_0.dffrs_10.nand3_0.C
rlabel metal2 8495 23324 8495 23324 5 SARlogic_0.dffrs_10.nand3_0.VSS
rlabel metal1 3361 24265 3361 24265 7 SARlogic_0.dffrs_9.setb
rlabel metal1 3361 21042 3361 21042 7 SARlogic_0.dffrs_9.clk
rlabel metal1 3361 17417 3361 17417 7 SARlogic_0.dffrs_9.d
rlabel metal1 3378 16630 3378 16630 7 SARlogic_0.dffrs_9.resetb
rlabel metal2 6829 21944 6829 21944 3 SARlogic_0.dffrs_9.Q
rlabel metal2 6829 19739 6829 19739 3 SARlogic_0.dffrs_9.Qb
rlabel metal5 5469 25370 5469 25370 1 SARlogic_0.dffrs_9.vdd
rlabel metal4 5577 16591 5577 16591 5 SARlogic_0.dffrs_9.vss
rlabel metal2 4525 18659 4525 18659 1 SARlogic_0.dffrs_9.nand3_8.VDD
rlabel metal1 4935 17533 4935 17533 3 SARlogic_0.dffrs_9.nand3_8.Z
rlabel metal1 3849 17415 3849 17415 7 SARlogic_0.dffrs_9.nand3_8.A
rlabel metal1 3849 17534 3849 17534 7 SARlogic_0.dffrs_9.nand3_8.B
rlabel metal1 3849 17650 3849 17650 7 SARlogic_0.dffrs_9.nand3_8.C
rlabel metal2 4453 16709 4453 16709 5 SARlogic_0.dffrs_9.nand3_8.VSS
rlabel metal2 6011 20865 6011 20865 1 SARlogic_0.dffrs_9.nand3_7.VDD
rlabel metal1 6421 19739 6421 19739 3 SARlogic_0.dffrs_9.nand3_7.Z
rlabel metal1 5335 19621 5335 19621 7 SARlogic_0.dffrs_9.nand3_7.A
rlabel metal1 5335 19740 5335 19740 7 SARlogic_0.dffrs_9.nand3_7.B
rlabel metal1 5335 19856 5335 19856 7 SARlogic_0.dffrs_9.nand3_7.C
rlabel metal2 5939 18915 5939 18915 5 SARlogic_0.dffrs_9.nand3_7.VSS
rlabel metal2 4525 20864 4525 20864 1 SARlogic_0.dffrs_9.nand3_6.VDD
rlabel metal1 4935 19738 4935 19738 3 SARlogic_0.dffrs_9.nand3_6.Z
rlabel metal1 3849 19620 3849 19620 7 SARlogic_0.dffrs_9.nand3_6.A
rlabel metal1 3849 19739 3849 19739 7 SARlogic_0.dffrs_9.nand3_6.B
rlabel metal1 3849 19855 3849 19855 7 SARlogic_0.dffrs_9.nand3_6.C
rlabel metal2 4453 18914 4453 18914 5 SARlogic_0.dffrs_9.nand3_6.VSS
rlabel metal2 6011 23069 6011 23069 1 SARlogic_0.dffrs_9.nand3_2.VDD
rlabel metal1 6421 21943 6421 21943 3 SARlogic_0.dffrs_9.nand3_2.Z
rlabel metal1 5335 21825 5335 21825 7 SARlogic_0.dffrs_9.nand3_2.A
rlabel metal1 5335 21944 5335 21944 7 SARlogic_0.dffrs_9.nand3_2.B
rlabel metal1 5335 22060 5335 22060 7 SARlogic_0.dffrs_9.nand3_2.C
rlabel metal2 5939 21119 5939 21119 5 SARlogic_0.dffrs_9.nand3_2.VSS
rlabel metal2 4525 23069 4525 23069 1 SARlogic_0.dffrs_9.nand3_1.VDD
rlabel metal1 4935 21943 4935 21943 3 SARlogic_0.dffrs_9.nand3_1.Z
rlabel metal1 3849 21825 3849 21825 7 SARlogic_0.dffrs_9.nand3_1.A
rlabel metal1 3849 21944 3849 21944 7 SARlogic_0.dffrs_9.nand3_1.B
rlabel metal1 3849 22060 3849 22060 7 SARlogic_0.dffrs_9.nand3_1.C
rlabel metal2 4453 21119 4453 21119 5 SARlogic_0.dffrs_9.nand3_1.VSS
rlabel metal2 4525 25274 4525 25274 1 SARlogic_0.dffrs_9.nand3_0.VDD
rlabel metal1 4935 24148 4935 24148 3 SARlogic_0.dffrs_9.nand3_0.Z
rlabel metal1 3849 24030 3849 24030 7 SARlogic_0.dffrs_9.nand3_0.A
rlabel metal1 3849 24149 3849 24149 7 SARlogic_0.dffrs_9.nand3_0.B
rlabel metal1 3849 24265 3849 24265 7 SARlogic_0.dffrs_9.nand3_0.C
rlabel metal2 4453 23324 4453 23324 5 SARlogic_0.dffrs_9.nand3_0.VSS
rlabel metal1 15487 24265 15487 24265 7 SARlogic_0.dffrs_12.setb
rlabel metal1 15487 21042 15487 21042 7 SARlogic_0.dffrs_12.clk
rlabel metal1 15487 17417 15487 17417 7 SARlogic_0.dffrs_12.d
rlabel metal1 15504 16630 15504 16630 7 SARlogic_0.dffrs_12.resetb
rlabel metal2 18955 21944 18955 21944 3 SARlogic_0.dffrs_12.Q
rlabel metal2 18955 19739 18955 19739 3 SARlogic_0.dffrs_12.Qb
rlabel metal5 17595 25370 17595 25370 1 SARlogic_0.dffrs_12.vdd
rlabel metal4 17703 16591 17703 16591 5 SARlogic_0.dffrs_12.vss
rlabel metal2 16651 18659 16651 18659 1 SARlogic_0.dffrs_12.nand3_8.VDD
rlabel metal1 17061 17533 17061 17533 3 SARlogic_0.dffrs_12.nand3_8.Z
rlabel metal1 15975 17415 15975 17415 7 SARlogic_0.dffrs_12.nand3_8.A
rlabel metal1 15975 17534 15975 17534 7 SARlogic_0.dffrs_12.nand3_8.B
rlabel metal1 15975 17650 15975 17650 7 SARlogic_0.dffrs_12.nand3_8.C
rlabel metal2 16579 16709 16579 16709 5 SARlogic_0.dffrs_12.nand3_8.VSS
rlabel metal2 18137 20865 18137 20865 1 SARlogic_0.dffrs_12.nand3_7.VDD
rlabel metal1 18547 19739 18547 19739 3 SARlogic_0.dffrs_12.nand3_7.Z
rlabel metal1 17461 19621 17461 19621 7 SARlogic_0.dffrs_12.nand3_7.A
rlabel metal1 17461 19740 17461 19740 7 SARlogic_0.dffrs_12.nand3_7.B
rlabel metal1 17461 19856 17461 19856 7 SARlogic_0.dffrs_12.nand3_7.C
rlabel metal2 18065 18915 18065 18915 5 SARlogic_0.dffrs_12.nand3_7.VSS
rlabel metal2 16651 20864 16651 20864 1 SARlogic_0.dffrs_12.nand3_6.VDD
rlabel metal1 17061 19738 17061 19738 3 SARlogic_0.dffrs_12.nand3_6.Z
rlabel metal1 15975 19620 15975 19620 7 SARlogic_0.dffrs_12.nand3_6.A
rlabel metal1 15975 19739 15975 19739 7 SARlogic_0.dffrs_12.nand3_6.B
rlabel metal1 15975 19855 15975 19855 7 SARlogic_0.dffrs_12.nand3_6.C
rlabel metal2 16579 18914 16579 18914 5 SARlogic_0.dffrs_12.nand3_6.VSS
rlabel metal2 18137 23069 18137 23069 1 SARlogic_0.dffrs_12.nand3_2.VDD
rlabel metal1 18547 21943 18547 21943 3 SARlogic_0.dffrs_12.nand3_2.Z
rlabel metal1 17461 21825 17461 21825 7 SARlogic_0.dffrs_12.nand3_2.A
rlabel metal1 17461 21944 17461 21944 7 SARlogic_0.dffrs_12.nand3_2.B
rlabel metal1 17461 22060 17461 22060 7 SARlogic_0.dffrs_12.nand3_2.C
rlabel metal2 18065 21119 18065 21119 5 SARlogic_0.dffrs_12.nand3_2.VSS
rlabel metal2 16651 23069 16651 23069 1 SARlogic_0.dffrs_12.nand3_1.VDD
rlabel metal1 17061 21943 17061 21943 3 SARlogic_0.dffrs_12.nand3_1.Z
rlabel metal1 15975 21825 15975 21825 7 SARlogic_0.dffrs_12.nand3_1.A
rlabel metal1 15975 21944 15975 21944 7 SARlogic_0.dffrs_12.nand3_1.B
rlabel metal1 15975 22060 15975 22060 7 SARlogic_0.dffrs_12.nand3_1.C
rlabel metal2 16579 21119 16579 21119 5 SARlogic_0.dffrs_12.nand3_1.VSS
rlabel metal2 16651 25274 16651 25274 1 SARlogic_0.dffrs_12.nand3_0.VDD
rlabel metal1 17061 24148 17061 24148 3 SARlogic_0.dffrs_12.nand3_0.Z
rlabel metal1 15975 24030 15975 24030 7 SARlogic_0.dffrs_12.nand3_0.A
rlabel metal1 15975 24149 15975 24149 7 SARlogic_0.dffrs_12.nand3_0.B
rlabel metal1 15975 24265 15975 24265 7 SARlogic_0.dffrs_12.nand3_0.C
rlabel metal2 16579 23324 16579 23324 5 SARlogic_0.dffrs_12.nand3_0.VSS
rlabel metal1 11445 24265 11445 24265 7 SARlogic_0.dffrs_11.setb
rlabel metal1 11445 21042 11445 21042 7 SARlogic_0.dffrs_11.clk
rlabel metal1 11445 17417 11445 17417 7 SARlogic_0.dffrs_11.d
rlabel metal1 11462 16630 11462 16630 7 SARlogic_0.dffrs_11.resetb
rlabel metal2 14913 21944 14913 21944 3 SARlogic_0.dffrs_11.Q
rlabel metal2 14913 19739 14913 19739 3 SARlogic_0.dffrs_11.Qb
rlabel metal5 13553 25370 13553 25370 1 SARlogic_0.dffrs_11.vdd
rlabel metal4 13661 16591 13661 16591 5 SARlogic_0.dffrs_11.vss
rlabel metal2 12609 18659 12609 18659 1 SARlogic_0.dffrs_11.nand3_8.VDD
rlabel metal1 13019 17533 13019 17533 3 SARlogic_0.dffrs_11.nand3_8.Z
rlabel metal1 11933 17415 11933 17415 7 SARlogic_0.dffrs_11.nand3_8.A
rlabel metal1 11933 17534 11933 17534 7 SARlogic_0.dffrs_11.nand3_8.B
rlabel metal1 11933 17650 11933 17650 7 SARlogic_0.dffrs_11.nand3_8.C
rlabel metal2 12537 16709 12537 16709 5 SARlogic_0.dffrs_11.nand3_8.VSS
rlabel metal2 14095 20865 14095 20865 1 SARlogic_0.dffrs_11.nand3_7.VDD
rlabel metal1 14505 19739 14505 19739 3 SARlogic_0.dffrs_11.nand3_7.Z
rlabel metal1 13419 19621 13419 19621 7 SARlogic_0.dffrs_11.nand3_7.A
rlabel metal1 13419 19740 13419 19740 7 SARlogic_0.dffrs_11.nand3_7.B
rlabel metal1 13419 19856 13419 19856 7 SARlogic_0.dffrs_11.nand3_7.C
rlabel metal2 14023 18915 14023 18915 5 SARlogic_0.dffrs_11.nand3_7.VSS
rlabel metal2 12609 20864 12609 20864 1 SARlogic_0.dffrs_11.nand3_6.VDD
rlabel metal1 13019 19738 13019 19738 3 SARlogic_0.dffrs_11.nand3_6.Z
rlabel metal1 11933 19620 11933 19620 7 SARlogic_0.dffrs_11.nand3_6.A
rlabel metal1 11933 19739 11933 19739 7 SARlogic_0.dffrs_11.nand3_6.B
rlabel metal1 11933 19855 11933 19855 7 SARlogic_0.dffrs_11.nand3_6.C
rlabel metal2 12537 18914 12537 18914 5 SARlogic_0.dffrs_11.nand3_6.VSS
rlabel metal2 14095 23069 14095 23069 1 SARlogic_0.dffrs_11.nand3_2.VDD
rlabel metal1 14505 21943 14505 21943 3 SARlogic_0.dffrs_11.nand3_2.Z
rlabel metal1 13419 21825 13419 21825 7 SARlogic_0.dffrs_11.nand3_2.A
rlabel metal1 13419 21944 13419 21944 7 SARlogic_0.dffrs_11.nand3_2.B
rlabel metal1 13419 22060 13419 22060 7 SARlogic_0.dffrs_11.nand3_2.C
rlabel metal2 14023 21119 14023 21119 5 SARlogic_0.dffrs_11.nand3_2.VSS
rlabel metal2 12609 23069 12609 23069 1 SARlogic_0.dffrs_11.nand3_1.VDD
rlabel metal1 13019 21943 13019 21943 3 SARlogic_0.dffrs_11.nand3_1.Z
rlabel metal1 11933 21825 11933 21825 7 SARlogic_0.dffrs_11.nand3_1.A
rlabel metal1 11933 21944 11933 21944 7 SARlogic_0.dffrs_11.nand3_1.B
rlabel metal1 11933 22060 11933 22060 7 SARlogic_0.dffrs_11.nand3_1.C
rlabel metal2 12537 21119 12537 21119 5 SARlogic_0.dffrs_11.nand3_1.VSS
rlabel metal2 12609 25274 12609 25274 1 SARlogic_0.dffrs_11.nand3_0.VDD
rlabel metal1 13019 24148 13019 24148 3 SARlogic_0.dffrs_11.nand3_0.Z
rlabel metal1 11933 24030 11933 24030 7 SARlogic_0.dffrs_11.nand3_0.A
rlabel metal1 11933 24149 11933 24149 7 SARlogic_0.dffrs_11.nand3_0.B
rlabel metal1 11933 24265 11933 24265 7 SARlogic_0.dffrs_11.nand3_0.C
rlabel metal2 12537 23324 12537 23324 5 SARlogic_0.dffrs_11.nand3_0.VSS
rlabel metal2 -12630 27550 -12630 27550 7 inv2_0.in
rlabel metal1 -12335 28819 -12335 28819 1 inv2_0.vdd
rlabel metal2 -12030 27550 -12030 27550 3 inv2_0.out
rlabel metal1 -12325 26679 -12325 26679 5 inv2_0.vss
rlabel metal3 -11840 27546 -11840 27546 7 adc_PISO_0.load
rlabel metal2 -11112 27289 -11112 27289 5 adc_PISO_0.B6
rlabel metal2 -1640 27289 -1640 27289 5 adc_PISO_0.B5
rlabel metal2 7832 27289 7832 27289 5 adc_PISO_0.B4
rlabel metal2 45724 37550 45724 37550 1 adc_PISO_0.serial_out
rlabel metal1 -10921 32152 -10921 32152 7 adc_PISO_0.avdd
rlabel metal2 17304 27290 17304 27290 5 adc_PISO_0.B3
rlabel metal1 -10921 27713 -10921 27713 7 adc_PISO_0.avss
rlabel metal2 26776 27290 26776 27290 5 adc_PISO_0.B2
rlabel metal2 36247 27290 36247 27290 5 adc_PISO_0.B1
rlabel metal3 -8093 33344 -8093 33344 7 adc_PISO_0.clk
rlabel metal2 -11141 30976 -11141 30976 7 adc_PISO_0.2inmux_0.Bit
rlabel metal2 -11141 30820 -11141 30820 7 adc_PISO_0.2inmux_0.Load
rlabel metal1 -10586 32169 -10586 32169 1 adc_PISO_0.2inmux_0.VDD
rlabel metal2 -5767 29723 -5767 29723 3 adc_PISO_0.2inmux_0.OUT
rlabel metal1 -10617 27689 -10617 27689 5 adc_PISO_0.2inmux_0.VSS
rlabel metal2 -11141 28480 -11141 28480 7 adc_PISO_0.2inmux_0.In
rlabel metal2 -1669 30976 -1669 30976 7 adc_PISO_0.2inmux_2.Bit
rlabel metal2 -1669 30820 -1669 30820 7 adc_PISO_0.2inmux_2.Load
rlabel metal1 -1114 32169 -1114 32169 1 adc_PISO_0.2inmux_2.VDD
rlabel metal2 3705 29723 3705 29723 3 adc_PISO_0.2inmux_2.OUT
rlabel metal1 -1145 27689 -1145 27689 5 adc_PISO_0.2inmux_2.VSS
rlabel metal2 -1669 28480 -1669 28480 7 adc_PISO_0.2inmux_2.In
rlabel metal1 -5507 36570 -5507 36570 7 adc_PISO_0.dffrs_0.setb
rlabel metal1 -5507 33347 -5507 33347 7 adc_PISO_0.dffrs_0.clk
rlabel metal1 -5507 29722 -5507 29722 7 adc_PISO_0.dffrs_0.d
rlabel metal1 -5490 28935 -5490 28935 7 adc_PISO_0.dffrs_0.resetb
rlabel metal2 -2039 34249 -2039 34249 3 adc_PISO_0.dffrs_0.Q
rlabel metal2 -2039 32044 -2039 32044 3 adc_PISO_0.dffrs_0.Qb
rlabel metal5 -3399 37675 -3399 37675 1 adc_PISO_0.dffrs_0.vdd
rlabel metal4 -3440 28896 -3440 28896 5 adc_PISO_0.dffrs_0.vss
rlabel metal1 3965 36570 3965 36570 7 adc_PISO_0.dffrs_1.setb
rlabel metal1 3965 33347 3965 33347 7 adc_PISO_0.dffrs_1.clk
rlabel metal1 3965 29722 3965 29722 7 adc_PISO_0.dffrs_1.d
rlabel metal1 3982 28935 3982 28935 7 adc_PISO_0.dffrs_1.resetb
rlabel metal2 7433 34249 7433 34249 3 adc_PISO_0.dffrs_1.Q
rlabel metal2 7433 32044 7433 32044 3 adc_PISO_0.dffrs_1.Qb
rlabel metal5 6073 37675 6073 37675 1 adc_PISO_0.dffrs_1.vdd
rlabel metal4 6032 28896 6032 28896 5 adc_PISO_0.dffrs_1.vss
rlabel metal2 7803 30977 7803 30977 7 adc_PISO_0.2inmux_3.Bit
rlabel metal2 7803 30821 7803 30821 7 adc_PISO_0.2inmux_3.Load
rlabel metal1 8358 32170 8358 32170 1 adc_PISO_0.2inmux_3.VDD
rlabel metal2 13177 29724 13177 29724 3 adc_PISO_0.2inmux_3.OUT
rlabel metal1 8327 27690 8327 27690 5 adc_PISO_0.2inmux_3.VSS
rlabel metal2 7803 28481 7803 28481 7 adc_PISO_0.2inmux_3.In
rlabel metal1 13437 36571 13437 36571 7 adc_PISO_0.dffrs_2.setb
rlabel metal1 13437 33348 13437 33348 7 adc_PISO_0.dffrs_2.clk
rlabel metal1 13437 29723 13437 29723 7 adc_PISO_0.dffrs_2.d
rlabel metal1 13454 28936 13454 28936 7 adc_PISO_0.dffrs_2.resetb
rlabel metal2 16905 34250 16905 34250 3 adc_PISO_0.dffrs_2.Q
rlabel metal2 16905 32045 16905 32045 3 adc_PISO_0.dffrs_2.Qb
rlabel metal5 15545 37676 15545 37676 1 adc_PISO_0.dffrs_2.vdd
rlabel metal4 15504 28897 15504 28897 5 adc_PISO_0.dffrs_2.vss
rlabel metal2 17275 30977 17275 30977 7 adc_PISO_0.2inmux_4.Bit
rlabel metal2 17275 30821 17275 30821 7 adc_PISO_0.2inmux_4.Load
rlabel metal1 17830 32170 17830 32170 1 adc_PISO_0.2inmux_4.VDD
rlabel metal2 22649 29724 22649 29724 3 adc_PISO_0.2inmux_4.OUT
rlabel metal1 17799 27690 17799 27690 5 adc_PISO_0.2inmux_4.VSS
rlabel metal2 17275 28481 17275 28481 7 adc_PISO_0.2inmux_4.In
rlabel metal1 22909 36571 22909 36571 7 adc_PISO_0.dffrs_3.setb
rlabel metal1 22909 33348 22909 33348 7 adc_PISO_0.dffrs_3.clk
rlabel metal1 22909 29723 22909 29723 7 adc_PISO_0.dffrs_3.d
rlabel metal1 22926 28936 22926 28936 7 adc_PISO_0.dffrs_3.resetb
rlabel metal2 26377 34250 26377 34250 3 adc_PISO_0.dffrs_3.Q
rlabel metal2 26377 32045 26377 32045 3 adc_PISO_0.dffrs_3.Qb
rlabel metal5 25017 37676 25017 37676 1 adc_PISO_0.dffrs_3.vdd
rlabel metal4 24976 28897 24976 28897 5 adc_PISO_0.dffrs_3.vss
rlabel metal2 26747 30977 26747 30977 7 adc_PISO_0.2inmux_5.Bit
rlabel metal2 26747 30821 26747 30821 7 adc_PISO_0.2inmux_5.Load
rlabel metal1 27302 32170 27302 32170 1 adc_PISO_0.2inmux_5.VDD
rlabel metal2 32121 29724 32121 29724 3 adc_PISO_0.2inmux_5.OUT
rlabel metal1 27271 27690 27271 27690 5 adc_PISO_0.2inmux_5.VSS
rlabel metal2 26747 28481 26747 28481 7 adc_PISO_0.2inmux_5.In
rlabel metal2 36219 30977 36219 30977 7 adc_PISO_0.2inmux_1.Bit
rlabel metal2 36219 30821 36219 30821 7 adc_PISO_0.2inmux_1.Load
rlabel metal1 36774 32170 36774 32170 1 adc_PISO_0.2inmux_1.VDD
rlabel metal2 41593 29724 41593 29724 3 adc_PISO_0.2inmux_1.OUT
rlabel metal1 36743 27690 36743 27690 5 adc_PISO_0.2inmux_1.VSS
rlabel metal2 36219 28481 36219 28481 7 adc_PISO_0.2inmux_1.In
rlabel metal1 32381 36571 32381 36571 7 adc_PISO_0.dffrs_4.setb
rlabel metal1 32381 33348 32381 33348 7 adc_PISO_0.dffrs_4.clk
rlabel metal1 32381 29723 32381 29723 7 adc_PISO_0.dffrs_4.d
rlabel metal1 32398 28936 32398 28936 7 adc_PISO_0.dffrs_4.resetb
rlabel metal2 35849 34250 35849 34250 3 adc_PISO_0.dffrs_4.Q
rlabel metal2 35849 32045 35849 32045 3 adc_PISO_0.dffrs_4.Qb
rlabel metal5 34489 37676 34489 37676 1 adc_PISO_0.dffrs_4.vdd
rlabel metal4 34448 28897 34448 28897 5 adc_PISO_0.dffrs_4.vss
rlabel metal1 41853 36571 41853 36571 7 adc_PISO_0.dffrs_5.setb
rlabel metal1 41853 33348 41853 33348 7 adc_PISO_0.dffrs_5.clk
rlabel metal1 41853 29723 41853 29723 7 adc_PISO_0.dffrs_5.d
rlabel metal1 41870 28936 41870 28936 7 adc_PISO_0.dffrs_5.resetb
rlabel metal2 45321 34250 45321 34250 3 adc_PISO_0.dffrs_5.Q
rlabel metal2 45321 32045 45321 32045 3 adc_PISO_0.dffrs_5.Qb
rlabel metal5 43961 37676 43961 37676 1 adc_PISO_0.dffrs_5.vdd
rlabel metal4 43920 28897 43920 28897 5 adc_PISO_0.dffrs_5.vss
rlabel metal2 38145 38613 38145 38613 1 Piso_out
port 10 n
rlabel metal2 40721 38313 40721 38313 6 osu_sc_buf_4_flat_0.A
rlabel metal2 40161 38573 40161 38573 6 osu_sc_buf_4_flat_0.Y
rlabel metal1 40851 38993 40851 38993 6 osu_sc_buf_4_flat_0.VDD
rlabel metal1 40851 37913 40851 37913 6 osu_sc_buf_4_flat_0.VSS
<< end >>
