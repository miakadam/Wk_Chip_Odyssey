magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< nwell >>
rect -954 -1710 954 1710
<< pmos >>
rect -704 -1500 -304 1500
rect -200 -1500 200 1500
rect 304 -1500 704 1500
<< pdiff >>
rect -792 1487 -704 1500
rect -792 -1487 -779 1487
rect -733 -1487 -704 1487
rect -792 -1500 -704 -1487
rect -304 1487 -200 1500
rect -304 -1487 -275 1487
rect -229 -1487 -200 1487
rect -304 -1500 -200 -1487
rect 200 1487 304 1500
rect 200 -1487 229 1487
rect 275 -1487 304 1487
rect 200 -1500 304 -1487
rect 704 1487 792 1500
rect 704 -1487 733 1487
rect 779 -1487 792 1487
rect 704 -1500 792 -1487
<< pdiffc >>
rect -779 -1487 -733 1487
rect -275 -1487 -229 1487
rect 229 -1487 275 1487
rect 733 -1487 779 1487
<< nsubdiff >>
rect -930 1614 930 1686
rect -930 1570 -858 1614
rect -930 -1570 -917 1570
rect -871 -1570 -858 1570
rect 858 1570 930 1614
rect -930 -1614 -858 -1570
rect 858 -1570 871 1570
rect 917 -1570 930 1570
rect 858 -1614 930 -1570
rect -930 -1686 930 -1614
<< nsubdiffcont >>
rect -917 -1570 -871 1570
rect 871 -1570 917 1570
<< polysilicon >>
rect -704 1579 -304 1592
rect -704 1533 -691 1579
rect -317 1533 -304 1579
rect -704 1500 -304 1533
rect -200 1579 200 1592
rect -200 1533 -187 1579
rect 187 1533 200 1579
rect -200 1500 200 1533
rect 304 1579 704 1592
rect 304 1533 317 1579
rect 691 1533 704 1579
rect 304 1500 704 1533
rect -704 -1533 -304 -1500
rect -704 -1579 -691 -1533
rect -317 -1579 -304 -1533
rect -704 -1592 -304 -1579
rect -200 -1533 200 -1500
rect -200 -1579 -187 -1533
rect 187 -1579 200 -1533
rect -200 -1592 200 -1579
rect 304 -1533 704 -1500
rect 304 -1579 317 -1533
rect 691 -1579 704 -1533
rect 304 -1592 704 -1579
<< polycontact >>
rect -691 1533 -317 1579
rect -187 1533 187 1579
rect 317 1533 691 1579
rect -691 -1579 -317 -1533
rect -187 -1579 187 -1533
rect 317 -1579 691 -1533
<< metal1 >>
rect -917 1627 917 1673
rect -917 1570 -871 1627
rect -702 1533 -691 1579
rect -317 1533 -306 1579
rect -198 1533 -187 1579
rect 187 1533 198 1579
rect 306 1533 317 1579
rect 691 1533 702 1579
rect 871 1570 917 1627
rect -779 1487 -733 1498
rect -779 -1498 -733 -1487
rect -275 1487 -229 1498
rect -275 -1498 -229 -1487
rect 229 1487 275 1498
rect 229 -1498 275 -1487
rect 733 1487 779 1498
rect 733 -1498 779 -1487
rect -917 -1627 -871 -1570
rect -702 -1579 -691 -1533
rect -317 -1579 -306 -1533
rect -198 -1579 -187 -1533
rect 187 -1579 198 -1533
rect 306 -1579 317 -1533
rect 691 -1579 702 -1533
rect 871 -1627 917 -1570
rect -917 -1673 917 -1627
<< properties >>
string FIXED_BBOX -894 -1650 894 1650
string gencell pfet_03v3
string library gf180mcu
string parameters w 15.0 l 2.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
