magic
tech gf180mcuD
timestamp 1757884890
<< checkpaint >>
rect -154 156 304 190
rect -206 -326 304 156
rect -154 -332 304 -326
<< metal1 >>
rect 0 0 20 20
rect 0 -40 20 -20
rect 0 -80 20 -60
rect 0 -120 20 -100
use nfet_03v3_WAQWUP  XM3
timestamp 0
transform 1 0 23 0 1 -85
box -29 -41 29 41
use pfet_03v3_LSTY94  XM4
timestamp 0
transform 1 0 75 0 1 -71
box -29 -61 29 61
<< labels >>
flabel metal1 0 0 20 20 0 FreeSans 128 0 0 0 avdd
port 0 nsew
flabel metal1 0 -40 20 -20 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 0 -80 20 -60 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 0 -120 20 -100 0 FreeSans 128 0 0 0 avss
port 3 nsew
<< end >>
