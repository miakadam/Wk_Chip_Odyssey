* NGSPICE file created from and2.ext - technology: (null)

.subckt and2 VDD OUT A B VSS
X0 a_n1203_400 B.t0 inv2_0.in.t2 VSS.t3 nfet_03v3
**devattr s=17600,576 d=10400,304
X1 a_n1203_400 A.t0 VSS.t5 VSS.t4 nfet_03v3
**devattr s=17600,576 d=10400,304
X2 inv2_0.in.t3 B.t1 VDD.t1 VDD.t0 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X3 OUT.t1 inv2_0.in.t4 VDD.t3 VDD.t2 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X4 OUT.t0 inv2_0.in.t5 VSS.t7 VSS.t6 nfet_03v3
**devattr s=17600,576 d=17600,576
X5 VSS.t1 A.t1 a_n1203_400 VSS.t0 nfet_03v3
**devattr s=10400,304 d=17600,576
X6 VDD.t5 A.t2 inv2_0.in.t0 VDD.t4 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X7 inv2_0.in.t1 B.t2 a_n1203_400 VSS.t2 nfet_03v3
**devattr s=10400,304 d=17600,576
R0 B.n1 B.t1 34.2529
R1 B.n0 B.t0 19.673
R2 B.n0 B.t2 19.4007
R3 nand2_0.A B.n1 6.43968
R4 B.n1 B.n0 0.106438
R5 nand2_0.A B 0.01175
R6 inv2_0.in.n0 inv2_0.in.t4 34.1797
R7 inv2_0.in.n0 inv2_0.in.t5 19.5798
R8 inv2_0.in.n2 inv2_0.in.t2 18.7717
R9 inv2_0.in.n2 inv2_0.in.t1 9.2885
R10 nand2_0.OUT inv2_0.in.n0 4.67986
R11 inv2_0.in.n1 inv2_0.in.t0 4.23346
R12 inv2_0.in.n1 inv2_0.in.t3 3.85546
R13 inv2_0.in.n3 inv2_0.in.n2 0.4055
R14 inv2_0.in.n3 inv2_0.in.n1 0.352625
R15 inv2_0.in nand2_0.OUT 0.193357
R16 inv2_0.in inv2_0.in.n3 0.0615714
R17 VSS.n13 VSS.n4 491393
R18 VSS.n14 VSS.n13 46157.7
R19 VSS.n13 VSS.n12 12638.9
R20 VSS.t6 VSS.n4 847.827
R21 VSS.n10 VSS.t6 847.827
R22 VSS.t2 VSS.n10 847.827
R23 VSS.n12 VSS.t3 847.827
R24 VSS.n12 VSS.t0 847.827
R25 VSS.n14 VSS.t4 847.827
R26 VSS.t3 VSS.t2 720.653
R27 VSS.t0 VSS.t4 720.653
R28 VSS.n15 VSS.n2 87.3061
R29 VSS.n15 VSS.n3 87.3061
R30 VSS.n6 VSS.n5 67.4727
R31 VSS.n7 VSS.n6 67.4727
R32 VSS.n5 VSS.n2 66.5005
R33 VSS.n7 VSS.n3 66.5005
R34 VSS.n9 VSS.n5 20.8061
R35 VSS.n9 VSS.n7 20.8061
R36 VSS.n11 VSS.n2 20.8061
R37 VSS.n11 VSS.n3 20.8061
R38 VSS.n1 VSS.t1 4.7885
R39 VSS.n8 VSS.t7 4.7885
R40 VSS.n16 VSS.t5 4.7885
R41 VSS.n6 VSS.n0 2.12302
R42 VSS.n9 VSS.n8 1.3005
R43 VSS.n10 VSS.n9 1.3005
R44 VSS.n6 VSS.n4 1.3005
R45 VSS.n11 VSS.n1 1.3005
R46 VSS.n12 VSS.n11 1.3005
R47 VSS.n16 VSS.n15 1.3005
R48 VSS.n15 VSS.n14 1.3005
R49 VSS.n17 VSS.n16 0.771017
R50 VSS.n17 VSS.n1 0.463217
R51 VSS.n8 VSS.n0 0.463217
R52 VSS VSS.n0 0.1787
R53 VSS VSS.n17 0.1301
R54 A.n1 A.t2 34.1066
R55 A.n0 A.t1 19.673
R56 A.n0 A.t0 19.4007
R57 nand2_0.B A.n1 5.09932
R58 A.n1 A.n0 0.252687
R59 nand2_0.B A 0.01175
R60 VDD.t2 VDD.n3 236.083
R61 VDD.n7 VDD.t0 236.083
R62 VDD.n6 VDD.t2 235.294
R63 VDD.t0 VDD.n6 235.294
R64 VDD.n9 VDD.t4 131.589
R65 VDD.n3 VDD.n1 78.2255
R66 VDD.n3 VDD.n2 78.2255
R67 VDD.n7 VDD.n1 78.2255
R68 VDD.n7 VDD.n2 78.2255
R69 VDD.n5 VDD.n1 36.2255
R70 VDD.n5 VDD.n2 36.2255
R71 VDD.n3 VDD.n0 2.00183
R72 VDD.n9 VDD.t5 1.49467
R73 VDD.n8 VDD.t1 1.49467
R74 VDD.n4 VDD.t3 1.47383
R75 VDD.n5 VDD.n4 0.788
R76 VDD.n6 VDD.n5 0.788
R77 VDD.n8 VDD.n7 0.788
R78 VDD.n4 VDD.n0 0.561043
R79 VDD.n11 VDD.n10 0.255287
R80 VDD VDD.n0 0.20525
R81 VDD VDD.n11 0.0509874
R82 VDD.n11 VDD.n8 0.0313054
R83 VDD.n11 VDD.n9 0.0313054
R84 OUT.n0 OUT.t0 9.6935
R85 OUT.n0 OUT.t1 4.35383
R86 inv2_0.out OUT.n0 0.254429
R87 inv2_0.out OUT 0.01175
.ends

