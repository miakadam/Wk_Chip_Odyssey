** sch_path: /foss/designs/comparator/final_magic/nand3/nand3.sch
.subckt nand3 VDD Z A B C VSS
*.PININFO VDD:B VSS:B Z:B A:B B:B C:B
XM1 Z A net1 VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM2 net1 B net2 VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
XM3 Z B VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM4 Z A VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM5 Z C VDD VDD pfet_03v3 L=0.4u W=2.5u nf=1 m=1
XM6 net2 C VSS VSS nfet_03v3 L=0.4u W=1u nf=1 m=1
.ends
