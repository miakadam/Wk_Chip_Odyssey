magic
tech gf180mcuD
magscale 1 5
timestamp 1757862833
<< metal1 >>
rect 840 750 1605 810
rect 910 685 945 750
rect 1360 635 1405 750
rect 1735 685 1855 710
rect 939 576 977 582
rect 939 550 945 576
rect 971 550 977 576
rect 939 544 977 550
rect 1689 571 1727 577
rect 1689 545 1695 571
rect 1721 545 1727 571
rect 1689 539 1727 545
rect 1874 576 1912 582
rect 1874 550 1880 576
rect 1906 550 1912 576
rect 1874 544 1912 550
rect 849 321 887 327
rect 849 295 855 321
rect 881 295 887 321
rect 849 289 887 295
rect 1034 321 1072 327
rect 1034 295 1040 321
rect 1066 295 1072 321
rect 1034 289 1072 295
rect 1779 326 1817 332
rect 1779 300 1785 326
rect 1811 300 1817 326
rect 1779 294 1817 300
rect 900 145 1015 205
rect 930 85 1000 145
rect 1740 140 1855 200
rect 1770 94 1840 140
rect 930 45 1315 85
rect 1435 54 1840 94
rect 930 -20 1000 45
rect 1770 -20 1840 54
rect 905 -80 1020 -20
rect 1750 -80 1865 -20
rect 939 -164 977 -158
rect 939 -190 945 -164
rect 971 -190 977 -164
rect 939 -196 977 -190
rect 1684 -164 1722 -158
rect 1684 -190 1690 -164
rect 1716 -190 1722 -164
rect 1684 -196 1722 -190
rect 1874 -164 1912 -158
rect 1874 -190 1880 -164
rect 1906 -190 1912 -164
rect 1874 -196 1912 -190
rect 849 -419 887 -413
rect 849 -445 855 -419
rect 881 -445 887 -419
rect 849 -451 887 -445
rect 1034 -414 1072 -408
rect 1034 -440 1040 -414
rect 1066 -440 1072 -414
rect 1034 -446 1072 -440
rect 935 -600 975 -565
rect 1365 -600 1400 -305
rect 1779 -419 1817 -413
rect 1779 -445 1785 -419
rect 1811 -445 1817 -419
rect 1779 -451 1817 -445
rect 1750 -595 1875 -560
rect 860 -660 1525 -600
<< via1 >>
rect 945 550 971 576
rect 1695 545 1721 571
rect 1880 550 1906 576
rect 855 295 881 321
rect 1040 295 1066 321
rect 1785 300 1811 326
rect 945 -190 971 -164
rect 1690 -190 1716 -164
rect 1880 -190 1906 -164
rect 855 -445 881 -419
rect 1040 -440 1066 -414
rect 1785 -445 1811 -419
<< metal2 >>
rect 845 576 2020 585
rect 845 550 945 576
rect 971 571 1880 576
rect 971 550 1695 571
rect 845 545 1695 550
rect 1721 550 1880 571
rect 1906 550 2020 576
rect 1721 545 2020 550
rect 845 535 2020 545
rect 840 326 2020 335
rect 840 321 1785 326
rect 840 295 855 321
rect 881 295 1040 321
rect 1066 300 1785 321
rect 1811 300 2020 326
rect 1066 295 2020 300
rect 840 285 2020 295
rect 1360 -150 1405 285
rect 830 -164 2020 -150
rect 830 -190 945 -164
rect 971 -190 1690 -164
rect 1716 -190 1880 -164
rect 1906 -190 2020 -164
rect 830 -200 2020 -190
rect 845 -414 2020 -405
rect 845 -419 1040 -414
rect 845 -445 855 -419
rect 881 -440 1040 -419
rect 1066 -419 2020 -414
rect 1066 -440 1785 -419
rect 881 -445 1785 -440
rect 1811 -445 2020 -419
rect 845 -455 2020 -445
use CDAC_INV_V0  CDAC_INV_V0_0
timestamp 1757701119
transform 1 0 755 0 1 115
box 480 -440 770 546
use nfet_03v3_QETW5R  nfet_03v3_QETW5R_0
timestamp 1757845275
transform 1 0 1801 0 -1 423
box -191 -293 191 293
use pfet_03v3_YXQA8C  pfet_03v3_YXQA8C_0
timestamp 1757845275
transform 1 0 1801 0 -1 -292
box -191 -293 191 293
use nfet_03v3_QETW5R  XM1
timestamp 1757845275
transform 1 0 961 0 1 -292
box -191 -293 191 293
use pfet_03v3_YXQA8C  XM4
timestamp 1757845275
transform 1 0 961 0 1 423
box -191 -293 191 293
<< labels >>
rlabel metal1 900 775 905 795 7 avdd
port 3 w
rlabel metal1 945 50 950 70 7 sw_bit
port 1 w
rlabel metal1 915 -630 920 -610 7 avss
port 2 w
rlabel metal1 1795 -590 1800 -570 7 avdd
rlabel space 1770 695 1775 715 7 avss
rlabel metal2 1165 550 1170 570 7 vreflow
port 5 w
rlabel metal2 1175 -190 1180 -170 7 sw_vout
port 0 w
rlabel metal2 1175 -440 1180 -420 7 sw_Vref
port 4 w
<< end >>
