magic
tech gf180mcuD
magscale 1 10
timestamp 1757649945
<< nwell >>
rect 2613 -735 2681 -734
<< pwell >>
rect 2613 -1472 2681 -860
<< metal1 >>
rect 2102 -71 2178 -38
rect 2286 -71 2362 -38
rect 2470 -71 2546 -38
rect 2008 -190 2088 -188
rect 1933 -310 2020 -190
rect 2076 -310 2088 -190
rect 2008 -312 2088 -310
rect 2376 -190 2456 -188
rect 2376 -310 2388 -190
rect 2444 -310 2456 -190
rect 2376 -312 2456 -310
rect 2698 -190 2778 -188
rect 2698 -311 2710 -190
rect 2766 -311 2778 -190
rect 2698 -313 2778 -311
rect 2192 -490 2272 -488
rect 1933 -610 2057 -490
rect 2192 -610 2204 -490
rect 2260 -610 2272 -490
rect 2192 -612 2272 -610
rect 2560 -490 2640 -488
rect 2560 -610 2572 -490
rect 2628 -610 2640 -490
rect 2560 -612 2640 -610
rect 2100 -742 2112 -686
rect 2168 -742 2180 -686
rect 2100 -756 2180 -742
rect 2284 -742 2296 -686
rect 2352 -742 2364 -686
rect 2284 -756 2364 -742
rect 2468 -742 2480 -686
rect 2536 -742 2548 -686
rect 2468 -756 2548 -742
rect 2100 -836 2180 -834
rect 1712 -892 2112 -836
rect 2168 -892 2180 -836
rect 2100 -894 2180 -892
rect 2284 -952 2364 -950
rect 1712 -1008 2296 -952
rect 2352 -1008 2364 -952
rect 2284 -1010 2364 -1008
rect 2613 -952 2693 -950
rect 2613 -1008 2625 -952
rect 2681 -1008 2798 -952
rect 2613 -1010 2693 -1008
rect 2468 -1068 2548 -1066
rect 1712 -1124 2480 -1068
rect 2536 -1124 2548 -1068
rect 2468 -1126 2548 -1124
rect 2100 -1218 2180 -1204
rect 2100 -1274 2112 -1218
rect 2168 -1274 2180 -1218
rect 2284 -1218 2364 -1204
rect 2284 -1274 2296 -1218
rect 2352 -1274 2364 -1218
rect 2468 -1218 2548 -1204
rect 2468 -1274 2480 -1218
rect 2536 -1274 2548 -1218
rect 1933 -1497 2025 -1323
rect 2560 -1350 2640 -1348
rect 2560 -1470 2572 -1350
rect 2628 -1470 2640 -1350
rect 2560 -1472 2640 -1470
rect 1887 -1725 1933 -1591
rect 2102 -1622 2178 -1589
rect 2286 -1622 2362 -1589
rect 2470 -1622 2546 -1589
rect 2715 -1725 2761 -1591
rect 1875 -1737 1955 -1725
rect 1875 -1793 1887 -1737
rect 1943 -1793 1955 -1737
rect 1875 -1805 1955 -1793
rect 2693 -1737 2771 -1725
rect 2693 -1793 2705 -1737
rect 2761 -1793 2771 -1737
rect 2693 -1805 2771 -1793
<< via1 >>
rect 2020 -310 2076 -190
rect 2388 -310 2444 -190
rect 2710 -311 2766 -190
rect 2204 -610 2260 -490
rect 2572 -610 2628 -490
rect 2112 -742 2168 -686
rect 2296 -742 2352 -686
rect 2480 -742 2536 -686
rect 2112 -892 2168 -836
rect 2296 -1008 2352 -952
rect 2625 -1008 2681 -952
rect 2480 -1124 2536 -1068
rect 2112 -1274 2168 -1218
rect 2296 -1274 2352 -1218
rect 2480 -1274 2536 -1218
rect 2572 -1470 2628 -1350
rect 1887 -1793 1943 -1737
rect 2705 -1793 2761 -1737
<< metal2 >>
rect 2020 65 2766 145
rect 2020 -188 2076 65
rect 2388 -188 2444 65
rect 2710 -188 2766 65
rect 2008 -190 2088 -188
rect 2008 -310 2020 -190
rect 2076 -310 2088 -190
rect 2008 -312 2088 -310
rect 2376 -190 2456 -188
rect 2376 -310 2388 -190
rect 2444 -310 2456 -190
rect 2376 -312 2456 -310
rect 2698 -190 2778 -188
rect 2698 -311 2710 -190
rect 2766 -311 2778 -190
rect 2020 -320 2076 -312
rect 2388 -320 2444 -312
rect 2698 -313 2778 -311
rect 2710 -321 2766 -313
rect 2204 -488 2260 -480
rect 2572 -488 2628 -480
rect 2192 -490 2681 -488
rect 2192 -610 2204 -490
rect 2260 -610 2572 -490
rect 2628 -610 2681 -490
rect 2192 -612 2681 -610
rect 2204 -620 2260 -612
rect 2572 -620 2681 -612
rect 2100 -686 2180 -676
rect 2100 -742 2112 -686
rect 2168 -742 2180 -686
rect 2100 -752 2180 -742
rect 2284 -686 2364 -676
rect 2284 -742 2296 -686
rect 2352 -742 2364 -686
rect 2284 -752 2364 -742
rect 2468 -686 2548 -676
rect 2468 -742 2480 -686
rect 2536 -742 2548 -686
rect 2468 -752 2548 -742
rect 2112 -834 2168 -752
rect 2100 -836 2180 -834
rect 2100 -892 2112 -836
rect 2168 -892 2180 -836
rect 2100 -894 2180 -892
rect 2112 -1208 2168 -894
rect 2296 -950 2352 -752
rect 2284 -952 2364 -950
rect 2284 -1008 2296 -952
rect 2352 -1008 2364 -952
rect 2284 -1010 2364 -1008
rect 2296 -1208 2352 -1010
rect 2480 -1066 2536 -752
rect 2613 -950 2681 -620
rect 2613 -952 2693 -950
rect 2613 -1008 2625 -952
rect 2681 -1008 2693 -952
rect 2613 -1010 2693 -1008
rect 2468 -1068 2548 -1066
rect 2468 -1124 2480 -1068
rect 2536 -1124 2548 -1068
rect 2468 -1126 2548 -1124
rect 2480 -1208 2536 -1126
rect 2100 -1218 2180 -1208
rect 2100 -1274 2112 -1218
rect 2168 -1274 2180 -1218
rect 2100 -1284 2180 -1274
rect 2284 -1218 2364 -1208
rect 2284 -1274 2296 -1218
rect 2352 -1274 2364 -1218
rect 2284 -1284 2364 -1274
rect 2468 -1218 2548 -1208
rect 2468 -1274 2480 -1218
rect 2536 -1274 2548 -1218
rect 2468 -1284 2548 -1274
rect 2613 -1340 2681 -1010
rect 2572 -1348 2681 -1340
rect 2560 -1350 2681 -1348
rect 2560 -1470 2572 -1350
rect 2628 -1470 2681 -1350
rect 2560 -1472 2681 -1470
rect 2572 -1480 2628 -1472
rect 1875 -1737 2771 -1725
rect 1875 -1793 1887 -1737
rect 1943 -1793 2705 -1737
rect 2761 -1793 2771 -1737
rect 1875 -1805 2771 -1793
use nfet_03v3_EPF4UP  M1
timestamp 1757649695
transform 1 0 2324 0 1 -1410
box -474 -310 474 310
use pfet_03v3_54RA84  M3
timestamp 1757649695
transform 1 0 2324 0 1 -400
box -474 -460 474 460
<< labels >>
rlabel metal2 2388 145 2388 145 1 VDD
port 0 n
rlabel metal1 2798 -981 2798 -981 3 Z
port 1 e
rlabel metal1 1712 -1099 1712 -1099 7 A
port 2 w
rlabel metal1 1712 -980 1712 -980 7 B
port 3 w
rlabel metal1 1712 -864 1712 -864 7 C
port 4 w
rlabel metal2 2316 -1805 2316 -1805 5 VSS
port 5 s
<< end >>
