magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -450 -10622 450 10622
<< nmos >>
rect -200 8012 200 10412
rect -200 5380 200 7780
rect -200 2748 200 5148
rect -200 116 200 2516
rect -200 -2516 200 -116
rect -200 -5148 200 -2748
rect -200 -7780 200 -5380
rect -200 -10412 200 -8012
<< ndiff >>
rect -288 10399 -200 10412
rect -288 8025 -275 10399
rect -229 8025 -200 10399
rect -288 8012 -200 8025
rect 200 10399 288 10412
rect 200 8025 229 10399
rect 275 8025 288 10399
rect 200 8012 288 8025
rect -288 7767 -200 7780
rect -288 5393 -275 7767
rect -229 5393 -200 7767
rect -288 5380 -200 5393
rect 200 7767 288 7780
rect 200 5393 229 7767
rect 275 5393 288 7767
rect 200 5380 288 5393
rect -288 5135 -200 5148
rect -288 2761 -275 5135
rect -229 2761 -200 5135
rect -288 2748 -200 2761
rect 200 5135 288 5148
rect 200 2761 229 5135
rect 275 2761 288 5135
rect 200 2748 288 2761
rect -288 2503 -200 2516
rect -288 129 -275 2503
rect -229 129 -200 2503
rect -288 116 -200 129
rect 200 2503 288 2516
rect 200 129 229 2503
rect 275 129 288 2503
rect 200 116 288 129
rect -288 -129 -200 -116
rect -288 -2503 -275 -129
rect -229 -2503 -200 -129
rect -288 -2516 -200 -2503
rect 200 -129 288 -116
rect 200 -2503 229 -129
rect 275 -2503 288 -129
rect 200 -2516 288 -2503
rect -288 -2761 -200 -2748
rect -288 -5135 -275 -2761
rect -229 -5135 -200 -2761
rect -288 -5148 -200 -5135
rect 200 -2761 288 -2748
rect 200 -5135 229 -2761
rect 275 -5135 288 -2761
rect 200 -5148 288 -5135
rect -288 -5393 -200 -5380
rect -288 -7767 -275 -5393
rect -229 -7767 -200 -5393
rect -288 -7780 -200 -7767
rect 200 -5393 288 -5380
rect 200 -7767 229 -5393
rect 275 -7767 288 -5393
rect 200 -7780 288 -7767
rect -288 -8025 -200 -8012
rect -288 -10399 -275 -8025
rect -229 -10399 -200 -8025
rect -288 -10412 -200 -10399
rect 200 -8025 288 -8012
rect 200 -10399 229 -8025
rect 275 -10399 288 -8025
rect 200 -10412 288 -10399
<< ndiffc >>
rect -275 8025 -229 10399
rect 229 8025 275 10399
rect -275 5393 -229 7767
rect 229 5393 275 7767
rect -275 2761 -229 5135
rect 229 2761 275 5135
rect -275 129 -229 2503
rect 229 129 275 2503
rect -275 -2503 -229 -129
rect 229 -2503 275 -129
rect -275 -5135 -229 -2761
rect 229 -5135 275 -2761
rect -275 -7767 -229 -5393
rect 229 -7767 275 -5393
rect -275 -10399 -229 -8025
rect 229 -10399 275 -8025
<< psubdiff >>
rect -426 10526 426 10598
rect -426 10482 -354 10526
rect -426 -10482 -413 10482
rect -367 -10482 -354 10482
rect 354 10482 426 10526
rect -426 -10526 -354 -10482
rect 354 -10482 367 10482
rect 413 -10482 426 10482
rect 354 -10526 426 -10482
rect -426 -10598 426 -10526
<< psubdiffcont >>
rect -413 -10482 -367 10482
rect 367 -10482 413 10482
<< polysilicon >>
rect -200 10491 200 10504
rect -200 10445 -187 10491
rect 187 10445 200 10491
rect -200 10412 200 10445
rect -200 7979 200 8012
rect -200 7933 -187 7979
rect 187 7933 200 7979
rect -200 7920 200 7933
rect -200 7859 200 7872
rect -200 7813 -187 7859
rect 187 7813 200 7859
rect -200 7780 200 7813
rect -200 5347 200 5380
rect -200 5301 -187 5347
rect 187 5301 200 5347
rect -200 5288 200 5301
rect -200 5227 200 5240
rect -200 5181 -187 5227
rect 187 5181 200 5227
rect -200 5148 200 5181
rect -200 2715 200 2748
rect -200 2669 -187 2715
rect 187 2669 200 2715
rect -200 2656 200 2669
rect -200 2595 200 2608
rect -200 2549 -187 2595
rect 187 2549 200 2595
rect -200 2516 200 2549
rect -200 83 200 116
rect -200 37 -187 83
rect 187 37 200 83
rect -200 24 200 37
rect -200 -37 200 -24
rect -200 -83 -187 -37
rect 187 -83 200 -37
rect -200 -116 200 -83
rect -200 -2549 200 -2516
rect -200 -2595 -187 -2549
rect 187 -2595 200 -2549
rect -200 -2608 200 -2595
rect -200 -2669 200 -2656
rect -200 -2715 -187 -2669
rect 187 -2715 200 -2669
rect -200 -2748 200 -2715
rect -200 -5181 200 -5148
rect -200 -5227 -187 -5181
rect 187 -5227 200 -5181
rect -200 -5240 200 -5227
rect -200 -5301 200 -5288
rect -200 -5347 -187 -5301
rect 187 -5347 200 -5301
rect -200 -5380 200 -5347
rect -200 -7813 200 -7780
rect -200 -7859 -187 -7813
rect 187 -7859 200 -7813
rect -200 -7872 200 -7859
rect -200 -7933 200 -7920
rect -200 -7979 -187 -7933
rect 187 -7979 200 -7933
rect -200 -8012 200 -7979
rect -200 -10445 200 -10412
rect -200 -10491 -187 -10445
rect 187 -10491 200 -10445
rect -200 -10504 200 -10491
<< polycontact >>
rect -187 10445 187 10491
rect -187 7933 187 7979
rect -187 7813 187 7859
rect -187 5301 187 5347
rect -187 5181 187 5227
rect -187 2669 187 2715
rect -187 2549 187 2595
rect -187 37 187 83
rect -187 -83 187 -37
rect -187 -2595 187 -2549
rect -187 -2715 187 -2669
rect -187 -5227 187 -5181
rect -187 -5347 187 -5301
rect -187 -7859 187 -7813
rect -187 -7979 187 -7933
rect -187 -10491 187 -10445
<< metal1 >>
rect -413 10539 413 10585
rect -413 10482 -367 10539
rect -198 10445 -187 10491
rect 187 10445 198 10491
rect 367 10482 413 10539
rect -275 10399 -229 10410
rect -275 8014 -229 8025
rect 229 10399 275 10410
rect 229 8014 275 8025
rect -198 7933 -187 7979
rect 187 7933 198 7979
rect -198 7813 -187 7859
rect 187 7813 198 7859
rect -275 7767 -229 7778
rect -275 5382 -229 5393
rect 229 7767 275 7778
rect 229 5382 275 5393
rect -198 5301 -187 5347
rect 187 5301 198 5347
rect -198 5181 -187 5227
rect 187 5181 198 5227
rect -275 5135 -229 5146
rect -275 2750 -229 2761
rect 229 5135 275 5146
rect 229 2750 275 2761
rect -198 2669 -187 2715
rect 187 2669 198 2715
rect -198 2549 -187 2595
rect 187 2549 198 2595
rect -275 2503 -229 2514
rect -275 118 -229 129
rect 229 2503 275 2514
rect 229 118 275 129
rect -198 37 -187 83
rect 187 37 198 83
rect -198 -83 -187 -37
rect 187 -83 198 -37
rect -275 -129 -229 -118
rect -275 -2514 -229 -2503
rect 229 -129 275 -118
rect 229 -2514 275 -2503
rect -198 -2595 -187 -2549
rect 187 -2595 198 -2549
rect -198 -2715 -187 -2669
rect 187 -2715 198 -2669
rect -275 -2761 -229 -2750
rect -275 -5146 -229 -5135
rect 229 -2761 275 -2750
rect 229 -5146 275 -5135
rect -198 -5227 -187 -5181
rect 187 -5227 198 -5181
rect -198 -5347 -187 -5301
rect 187 -5347 198 -5301
rect -275 -5393 -229 -5382
rect -275 -7778 -229 -7767
rect 229 -5393 275 -5382
rect 229 -7778 275 -7767
rect -198 -7859 -187 -7813
rect 187 -7859 198 -7813
rect -198 -7979 -187 -7933
rect 187 -7979 198 -7933
rect -275 -8025 -229 -8014
rect -275 -10410 -229 -10399
rect 229 -8025 275 -8014
rect 229 -10410 275 -10399
rect -413 -10539 -367 -10482
rect -198 -10491 -187 -10445
rect 187 -10491 198 -10445
rect 367 -10539 413 -10482
rect -413 -10585 413 -10539
<< properties >>
string FIXED_BBOX -390 -10562 390 10562
string gencell nfet_03v3
string library gf180mcu
string parameters w 12.0 l 2.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
