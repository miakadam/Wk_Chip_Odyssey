magic
tech gf180mcuD
magscale 1 10
timestamp 1757500055
<< nwell >>
rect -1718 -310 1718 310
<< pmos >>
rect -1468 -100 -1268 100
rect -1164 -100 -964 100
rect -860 -100 -660 100
rect -556 -100 -356 100
rect -252 -100 -52 100
rect 52 -100 252 100
rect 356 -100 556 100
rect 660 -100 860 100
rect 964 -100 1164 100
rect 1268 -100 1468 100
<< pdiff >>
rect -1556 87 -1468 100
rect -1556 -87 -1543 87
rect -1497 -87 -1468 87
rect -1556 -100 -1468 -87
rect -1268 87 -1164 100
rect -1268 -87 -1239 87
rect -1193 -87 -1164 87
rect -1268 -100 -1164 -87
rect -964 87 -860 100
rect -964 -87 -935 87
rect -889 -87 -860 87
rect -964 -100 -860 -87
rect -660 87 -556 100
rect -660 -87 -631 87
rect -585 -87 -556 87
rect -660 -100 -556 -87
rect -356 87 -252 100
rect -356 -87 -327 87
rect -281 -87 -252 87
rect -356 -100 -252 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 252 87 356 100
rect 252 -87 281 87
rect 327 -87 356 87
rect 252 -100 356 -87
rect 556 87 660 100
rect 556 -87 585 87
rect 631 -87 660 87
rect 556 -100 660 -87
rect 860 87 964 100
rect 860 -87 889 87
rect 935 -87 964 87
rect 860 -100 964 -87
rect 1164 87 1268 100
rect 1164 -87 1193 87
rect 1239 -87 1268 87
rect 1164 -100 1268 -87
rect 1468 87 1556 100
rect 1468 -87 1497 87
rect 1543 -87 1556 87
rect 1468 -100 1556 -87
<< pdiffc >>
rect -1543 -87 -1497 87
rect -1239 -87 -1193 87
rect -935 -87 -889 87
rect -631 -87 -585 87
rect -327 -87 -281 87
rect -23 -87 23 87
rect 281 -87 327 87
rect 585 -87 631 87
rect 889 -87 935 87
rect 1193 -87 1239 87
rect 1497 -87 1543 87
<< nsubdiff >>
rect -1694 214 1694 286
rect -1694 170 -1622 214
rect -1694 -170 -1681 170
rect -1635 -170 -1622 170
rect 1622 170 1694 214
rect -1694 -214 -1622 -170
rect 1622 -170 1635 170
rect 1681 -170 1694 170
rect 1622 -214 1694 -170
rect -1694 -286 1694 -214
<< nsubdiffcont >>
rect -1681 -170 -1635 170
rect 1635 -170 1681 170
<< polysilicon >>
rect -1468 179 -1268 192
rect -1468 133 -1455 179
rect -1281 133 -1268 179
rect -1468 100 -1268 133
rect -1164 179 -964 192
rect -1164 133 -1151 179
rect -977 133 -964 179
rect -1164 100 -964 133
rect -860 179 -660 192
rect -860 133 -847 179
rect -673 133 -660 179
rect -860 100 -660 133
rect -556 179 -356 192
rect -556 133 -543 179
rect -369 133 -356 179
rect -556 100 -356 133
rect -252 179 -52 192
rect -252 133 -239 179
rect -65 133 -52 179
rect -252 100 -52 133
rect 52 179 252 192
rect 52 133 65 179
rect 239 133 252 179
rect 52 100 252 133
rect 356 179 556 192
rect 356 133 369 179
rect 543 133 556 179
rect 356 100 556 133
rect 660 179 860 192
rect 660 133 673 179
rect 847 133 860 179
rect 660 100 860 133
rect 964 179 1164 192
rect 964 133 977 179
rect 1151 133 1164 179
rect 964 100 1164 133
rect 1268 179 1468 192
rect 1268 133 1281 179
rect 1455 133 1468 179
rect 1268 100 1468 133
rect -1468 -133 -1268 -100
rect -1468 -179 -1455 -133
rect -1281 -179 -1268 -133
rect -1468 -192 -1268 -179
rect -1164 -133 -964 -100
rect -1164 -179 -1151 -133
rect -977 -179 -964 -133
rect -1164 -192 -964 -179
rect -860 -133 -660 -100
rect -860 -179 -847 -133
rect -673 -179 -660 -133
rect -860 -192 -660 -179
rect -556 -133 -356 -100
rect -556 -179 -543 -133
rect -369 -179 -356 -133
rect -556 -192 -356 -179
rect -252 -133 -52 -100
rect -252 -179 -239 -133
rect -65 -179 -52 -133
rect -252 -192 -52 -179
rect 52 -133 252 -100
rect 52 -179 65 -133
rect 239 -179 252 -133
rect 52 -192 252 -179
rect 356 -133 556 -100
rect 356 -179 369 -133
rect 543 -179 556 -133
rect 356 -192 556 -179
rect 660 -133 860 -100
rect 660 -179 673 -133
rect 847 -179 860 -133
rect 660 -192 860 -179
rect 964 -133 1164 -100
rect 964 -179 977 -133
rect 1151 -179 1164 -133
rect 964 -192 1164 -179
rect 1268 -133 1468 -100
rect 1268 -179 1281 -133
rect 1455 -179 1468 -133
rect 1268 -192 1468 -179
<< polycontact >>
rect -1455 133 -1281 179
rect -1151 133 -977 179
rect -847 133 -673 179
rect -543 133 -369 179
rect -239 133 -65 179
rect 65 133 239 179
rect 369 133 543 179
rect 673 133 847 179
rect 977 133 1151 179
rect 1281 133 1455 179
rect -1455 -179 -1281 -133
rect -1151 -179 -977 -133
rect -847 -179 -673 -133
rect -543 -179 -369 -133
rect -239 -179 -65 -133
rect 65 -179 239 -133
rect 369 -179 543 -133
rect 673 -179 847 -133
rect 977 -179 1151 -133
rect 1281 -179 1455 -133
<< metal1 >>
rect -1681 170 -1635 181
rect -1466 133 -1455 179
rect -1281 133 -1270 179
rect -1162 133 -1151 179
rect -977 133 -966 179
rect -858 133 -847 179
rect -673 133 -662 179
rect -554 133 -543 179
rect -369 133 -358 179
rect -250 133 -239 179
rect -65 133 -54 179
rect 54 133 65 179
rect 239 133 250 179
rect 358 133 369 179
rect 543 133 554 179
rect 662 133 673 179
rect 847 133 858 179
rect 966 133 977 179
rect 1151 133 1162 179
rect 1270 133 1281 179
rect 1455 133 1466 179
rect 1635 170 1681 181
rect -1543 87 -1497 98
rect -1543 -98 -1497 -87
rect -1239 87 -1193 98
rect -1239 -98 -1193 -87
rect -935 87 -889 98
rect -935 -98 -889 -87
rect -631 87 -585 98
rect -631 -98 -585 -87
rect -327 87 -281 98
rect -327 -98 -281 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 281 87 327 98
rect 281 -98 327 -87
rect 585 87 631 98
rect 585 -98 631 -87
rect 889 87 935 98
rect 889 -98 935 -87
rect 1193 87 1239 98
rect 1193 -98 1239 -87
rect 1497 87 1543 98
rect 1497 -98 1543 -87
rect -1681 -181 -1635 -170
rect -1466 -179 -1455 -133
rect -1281 -179 -1270 -133
rect -1162 -179 -1151 -133
rect -977 -179 -966 -133
rect -858 -179 -847 -133
rect -673 -179 -662 -133
rect -554 -179 -543 -133
rect -369 -179 -358 -133
rect -250 -179 -239 -133
rect -65 -179 -54 -133
rect 54 -179 65 -133
rect 239 -179 250 -133
rect 358 -179 369 -133
rect 543 -179 554 -133
rect 662 -179 673 -133
rect 847 -179 858 -133
rect 966 -179 977 -133
rect 1151 -179 1162 -133
rect 1270 -179 1281 -133
rect 1455 -179 1466 -133
rect 1635 -181 1681 -170
<< properties >>
string FIXED_BBOX -1658 -250 1658 250
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
