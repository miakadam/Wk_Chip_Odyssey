magic
tech gf180mcuD
magscale 1 10
timestamp 1755242987
<< pwell >>
rect -350 -1710 350 1710
<< nmos >>
rect -100 -1500 100 1500
<< ndiff >>
rect -188 1487 -100 1500
rect -188 -1487 -175 1487
rect -129 -1487 -100 1487
rect -188 -1500 -100 -1487
rect 100 1487 188 1500
rect 100 -1487 129 1487
rect 175 -1487 188 1487
rect 100 -1500 188 -1487
<< ndiffc >>
rect -175 -1487 -129 1487
rect 129 -1487 175 1487
<< psubdiff >>
rect -326 1614 326 1686
rect -326 1570 -254 1614
rect -326 -1570 -313 1570
rect -267 -1570 -254 1570
rect 254 1570 326 1614
rect -326 -1614 -254 -1570
rect 254 -1570 267 1570
rect 313 -1570 326 1570
rect 254 -1614 326 -1570
rect -326 -1686 326 -1614
<< psubdiffcont >>
rect -313 -1570 -267 1570
rect 267 -1570 313 1570
<< polysilicon >>
rect -100 1579 100 1592
rect -100 1533 -87 1579
rect 87 1533 100 1579
rect -100 1500 100 1533
rect -100 -1533 100 -1500
rect -100 -1579 -87 -1533
rect 87 -1579 100 -1533
rect -100 -1592 100 -1579
<< polycontact >>
rect -87 1533 87 1579
rect -87 -1579 87 -1533
<< metal1 >>
rect -313 1627 313 1673
rect -313 1570 -267 1627
rect -98 1533 -87 1579
rect 87 1533 98 1579
rect 267 1570 313 1627
rect -175 1487 -129 1498
rect -175 -1498 -129 -1487
rect 129 1487 175 1498
rect 129 -1498 175 -1487
rect -313 -1627 -267 -1570
rect -98 -1579 -87 -1533
rect 87 -1579 98 -1533
rect 267 -1627 313 -1570
rect -313 -1673 313 -1627
<< properties >>
string FIXED_BBOX -290 -1650 290 1650
string gencell nfet_03v3
string library gf180mcu
string parameters w 15.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
