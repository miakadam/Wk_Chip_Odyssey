* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dffsr_1.2.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__dffsr_1 D CLK Q QN R VDD VSS S
X0 VSS.t7 a_820_160.t4 a_770_210.t0 VSS.t6 nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X1 a_820_160.t2 a_1370_430.t2 a_1280_210.t0 VSS.t10 nfet_03v3 ad=0.3425p pd=1.7u as=0.225p ps=1.35u w=0.6u l=0.3u
X2 a_1280_720.t1 D.t0 VDD.t19 VDD.t18 pfet_03v3 ad=0.6375p pd=2.45u as=0.85p ps=4.4u w=1.7u l=0.3u
X3 VDD.t7 a_2470_490.t3 QN.t0 VDD.t6 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 VSS.t21 a_250_210.t2 a_2470_490.t1 VSS.t20 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X5 Q.t1 QN.t2 VSS.t29 VSS.t28 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X6 VSS.t19 a_410_720.t3 a_1720_210.t1 VSS.t18 nfet_03v3 ad=0.23375p pd=1.4u as=0.10625p ps=1.1u w=0.85u l=0.3u
X7 a_2340_210.t0 a_1370_430.t3 a_2110_210.t3 VSS.t8 nfet_03v3 ad=0.225p pd=1.35u as=0.3425p ps=1.7u w=0.6u l=0.3u
X8 a_820_160.t1 CLK.t0 a_1280_720.t0 VDD.t0 pfet_03v3 ad=0.7225p pd=2.55u as=0.6375p ps=2.45u w=1.7u l=0.3u
X9 VDD.t21 S.t0 a_570_720.t2 VDD.t20 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 VSS.t12 a_2470_490.t4 a_2340_210.t1 VSS.t11 nfet_03v3 ad=0.215p pd=1.4u as=0.225p ps=1.35u w=0.6u l=0.3u
X11 VDD.t17 a_410_720.t4 a_1720_720.t0 VDD.t16 pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X12 a_2340_720.t1 CLK.t1 a_2110_210.t0 VDD.t5 pfet_03v3 ad=0.6375p pd=2.45u as=0.7225p ps=2.55u w=1.7u l=0.3u
X13 Q.t0 QN.t3 VDD.t27 VDD.t26 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X14 a_2000_210.t0 a_410_720.t5 VSS.t25 VSS.t24 nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
X15 a_250_210.t0 R.t0 VSS.t5 VSS.t4 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X16 a_570_720.t1 a_250_210.t3 a_410_720.t1 VDD.t29 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X17 a_2910_720.t2 S.t1 VDD.t11 VDD.t10 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X18 a_410_720.t2 a_250_210.t4 VSS.t23 VSS.t22 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X19 a_570_720.t0 a_820_160.t5 VDD.t2 VDD.t1 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X20 VDD.t13 a_2470_490.t5 a_2340_720.t0 VDD.t12 pfet_03v3 ad=0.4675p pd=2.25u as=0.6375p ps=2.45u w=1.7u l=0.3u
X21 VDD.t9 a_2110_210.t4 a_2910_720.t1 VDD.t8 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X22 a_1370_430.t1 CLK.t2 VSS.t17 VSS.t16 nfet_03v3 ad=0.425p pd=2.7u as=0.215p ps=1.4u w=0.85u l=0.3u
X23 a_250_210.t1 R.t1 VDD.t23 VDD.t22 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X24 a_2000_720.t0 a_410_720.t6 VDD.t15 VDD.t14 pfet_03v3 ad=0.2125p pd=1.95u as=0.4675p ps=2.25u w=1.7u l=0.3u
X25 a_2110_210.t1 CLK.t3 a_2000_210.t1 VSS.t13 nfet_03v3 ad=0.3425p pd=1.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X26 a_3100_210.t0 a_2110_210.t5 VSS.t1 VSS.t0 nfet_03v3 ad=0.10625p pd=1.1u as=0.425p ps=2.7u w=0.85u l=0.3u
X27 a_2470_490.t2 a_250_210.t5 a_2910_720.t0 VDD.t28 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X28 a_770_210.t1 S.t2 a_410_720.t0 VSS.t9 nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
X29 a_1370_430.t0 CLK.t4 VDD.t4 VDD.t3 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X30 a_2110_210.t2 a_1370_430.t4 a_2000_720.t1 VDD.t25 pfet_03v3 ad=0.7225p pd=2.55u as=0.2125p ps=1.95u w=1.7u l=0.3u
X31 a_1720_210.t0 CLK.t5 a_820_160.t0 VSS.t2 nfet_03v3 ad=0.10625p pd=1.1u as=0.3425p ps=1.7u w=0.85u l=0.3u
X32 a_1720_720.t1 a_1370_430.t5 a_820_160.t3 VDD.t24 pfet_03v3 ad=0.2125p pd=1.95u as=0.7225p ps=2.55u w=1.7u l=0.3u
X33 a_1280_210.t1 D.t1 VSS.t27 VSS.t26 nfet_03v3 ad=0.225p pd=1.35u as=0.3p ps=2.2u w=0.6u l=0.3u
X34 a_2470_490.t0 S.t3 a_3100_210.t1 VSS.t3 nfet_03v3 ad=0.23375p pd=1.4u as=0.10625p ps=1.1u w=0.85u l=0.3u
X35 VSS.t15 a_2470_490.t6 QN.t1 VSS.t14 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
R0 a_820_160.n1 a_820_160.t4 38.0938
R1 a_820_160.n1 a_820_160.t5 25.7243
R2 a_820_160.n2 a_820_160.n1 8.2705
R3 a_820_160.n3 a_820_160.n2 7.33918
R4 a_820_160.n3 a_820_160.t2 3.61374
R5 a_820_160.n2 a_820_160.n0 3.54277
R6 a_820_160.t0 a_820_160.n3 3.1505
R7 a_820_160.n0 a_820_160.t3 1.7505
R8 a_820_160.n0 a_820_160.t1 1.7505
R9 a_770_210.t0 a_770_210.t1 1.85344
R10 VSS.n18 VSS.n17 1238.1
R11 VSS.n35 VSS.n34 1186.51
R12 VSS.t13 VSS.n23 1109.13
R13 VSS.t8 VSS.t11 1083.33
R14 VSS.n13 VSS.t14 1057.54
R15 VSS.n40 VSS.t22 954.365
R16 VSS.t4 VSS.n40 851.191
R17 VSS.n22 VSS.t16 799.604
R18 VSS.n28 VSS.t24 799.604
R19 VSS.n34 VSS.t26 799.604
R20 VSS.t20 VSS.n13 748.016
R21 VSS.n10 VSS.t28 696.429
R22 VSS.n30 VSS.t10 644.841
R23 VSS.n29 VSS.t2 593.255
R24 VSS.t10 VSS.n29 593.255
R25 VSS.n39 VSS.t9 593.255
R26 VSS.t3 VSS.t0 567.461
R27 VSS.t2 VSS.t18 567.461
R28 VSS.t6 VSS.t9 567.461
R29 VSS.t28 VSS.n9 552.189
R30 VSS.n14 VSS.t20 490.079
R31 VSS.n41 VSS.t4 448.892
R32 VSS.n18 VSS.t16 438.493
R33 VSS.n24 VSS.t24 438.493
R34 VSS.n30 VSS.t26 438.493
R35 VSS.n14 VSS.t3 386.906
R36 VSS.n17 VSS.t0 283.731
R37 VSS.t22 VSS.n39 283.731
R38 VSS.n10 VSS.t14 180.556
R39 VSS.n24 VSS.t13 128.969
R40 VSS.t11 VSS.n22 77.3815
R41 VSS.n23 VSS.t8 77.3815
R42 VSS.t18 VSS.n28 77.3815
R43 VSS.n35 VSS.t6 77.3815
R44 VSS.n11 VSS.n10 10.4005
R45 VSS.n13 VSS.n12 10.4005
R46 VSS.n15 VSS.n14 10.4005
R47 VSS.n17 VSS.n16 10.4005
R48 VSS.n19 VSS.n18 10.4005
R49 VSS.n22 VSS.n21 10.4005
R50 VSS.n23 VSS.n4 10.4005
R51 VSS.n25 VSS.n24 10.4005
R52 VSS.n28 VSS.n27 10.4005
R53 VSS.n29 VSS.n2 10.4005
R54 VSS.n31 VSS.n30 10.4005
R55 VSS.n34 VSS.n33 10.4005
R56 VSS.n36 VSS.n35 10.4005
R57 VSS.n39 VSS.n38 10.4005
R58 VSS.n40 VSS.n0 10.4005
R59 VSS.n32 VSS.t27 9.404
R60 VSS.n41 VSS.t5 8.61774
R61 VSS.n6 VSS.t1 8.61774
R62 VSS.n1 VSS.t7 8.55474
R63 VSS.n7 VSS.t21 8.54574
R64 VSS.n37 VSS.t23 8.54574
R65 VSS.n9 VSS.n8 6.5435
R66 VSS.n20 VSS.n5 6.5345
R67 VSS.n26 VSS.n3 6.5075
R68 VSS.n5 VSS.t12 2.888
R69 VSS.n5 VSS.t17 2.27035
R70 VSS.n8 VSS.t29 2.03874
R71 VSS.n8 VSS.t15 2.03874
R72 VSS.n3 VSS.t25 2.03874
R73 VSS.n3 VSS.t19 2.03874
R74 VSS.n41 VSS.n0 0.161214
R75 VSS.n12 VSS.n11 0.154786
R76 VSS.n16 VSS.n15 0.154786
R77 VSS.n21 VSS.n4 0.154786
R78 VSS.n25 VSS.n4 0.154786
R79 VSS.n27 VSS.n2 0.154786
R80 VSS.n31 VSS.n2 0.154786
R81 VSS.n38 VSS.n36 0.154786
R82 VSS.n19 VSS.n6 0.1355
R83 VSS.n15 VSS.n7 0.116214
R84 VSS.n20 VSS.n19 0.109786
R85 VSS.n26 VSS.n25 0.109786
R86 VSS.n32 VSS.n31 0.109786
R87 VSS.n33 VSS.n1 0.103357
R88 VSS.n38 VSS.n37 0.0905
R89 VSS.n37 VSS.n0 0.0647857
R90 VSS.n21 VSS.n20 0.0455
R91 VSS.n27 VSS.n26 0.0455
R92 VSS.n33 VSS.n32 0.0455
R93 VSS.n36 VSS.n1 0.0455
R94 VSS.n12 VSS.n7 0.0390714
R95 VSS.n11 VSS.n9 0.0326429
R96 VSS.n16 VSS.n6 0.0197857
R97 VSS VSS.n41 0.00371429
R98 a_1370_430.n0 a_1370_430.t5 62.9278
R99 a_1370_430.n1 a_1370_430.t4 62.6114
R100 a_1370_430.n0 a_1370_430.t2 22.5088
R101 a_1370_430.n1 a_1370_430.t3 21.9005
R102 a_1370_430.n2 a_1370_430.n0 19.7118
R103 a_1370_430.n3 a_1370_430.t1 8.54574
R104 a_1370_430.n2 a_1370_430.n1 8.0005
R105 a_1370_430.t0 a_1370_430.n3 3.65819
R106 a_1370_430.n3 a_1370_430.n2 0.743643
R107 a_1280_210.t0 a_1280_210.t1 7.8755
R108 D.n0 D.t1 39.8187
R109 D.n0 D.t0 30.0854
R110 D D.n0 12.5005
R111 VDD.n20 VDD.n5 375
R112 VDD.n22 VDD.t25 335.938
R113 VDD.t1 VDD.n34 335.938
R114 VDD.t5 VDD.t12 328.125
R115 VDD.n12 VDD.t6 320.312
R116 VDD.t10 VDD.t8 265.625
R117 VDD.t22 VDD.n40 257.812
R118 VDD.n21 VDD.t3 242.189
R119 VDD.n28 VDD.t14 242.189
R120 VDD.n34 VDD.t18 242.189
R121 VDD.n35 VDD.t20 242.189
R122 VDD.n40 VDD.t29 242.189
R123 VDD.n11 VDD.t26 210.939
R124 VDD.n13 VDD.t28 195.312
R125 VDD.n33 VDD.t0 195.312
R126 VDD.t28 VDD.n12 179.689
R127 VDD.n29 VDD.t24 179.689
R128 VDD.n29 VDD.t0 179.689
R129 VDD.n9 VDD.t26 176.786
R130 VDD.t24 VDD.t16 171.875
R131 VDD.n41 VDD.t22 145.413
R132 VDD.t3 VDD.n20 132.812
R133 VDD.t14 VDD.n27 132.812
R134 VDD.t18 VDD.n33 132.812
R135 VDD.n39 VDD.t20 132.812
R136 VDD.t29 VDD.n39 132.812
R137 VDD.n13 VDD.t10 70.313
R138 VDD.t6 VDD.n11 54.688
R139 VDD.t8 VDD.n5 39.063
R140 VDD.n27 VDD.t25 39.063
R141 VDD.t12 VDD.n21 23.438
R142 VDD.n22 VDD.t5 23.438
R143 VDD.t16 VDD.n28 23.438
R144 VDD.n35 VDD.t1 23.438
R145 VDD.n31 VDD.t19 14.1575
R146 VDD.n11 VDD.n10 12.6005
R147 VDD.n12 VDD.n7 12.6005
R148 VDD.n14 VDD.n13 12.6005
R149 VDD.n16 VDD.n5 12.6005
R150 VDD.n20 VDD.n19 12.6005
R151 VDD.n21 VDD.n4 12.6005
R152 VDD.n23 VDD.n22 12.6005
R153 VDD.n27 VDD.n26 12.6005
R154 VDD.n28 VDD.n3 12.6005
R155 VDD.n30 VDD.n29 12.6005
R156 VDD.n33 VDD.n32 12.6005
R157 VDD.n34 VDD.n2 12.6005
R158 VDD.n36 VDD.n35 12.6005
R159 VDD.n39 VDD.n38 12.6005
R160 VDD.n40 VDD.n0 12.6005
R161 VDD.n18 VDD.n17 5.4075
R162 VDD.n41 VDD.t23 3.29819
R163 VDD.n9 VDD.n8 2.9335
R164 VDD.n25 VDD.n24 2.9245
R165 VDD.n37 VDD.n1 2.8975
R166 VDD.n15 VDD.n6 2.8975
R167 VDD.n1 VDD.t2 1.13285
R168 VDD.n1 VDD.t21 1.13285
R169 VDD.n24 VDD.t15 1.13285
R170 VDD.n24 VDD.t17 1.13285
R171 VDD.n17 VDD.t4 1.13285
R172 VDD.n17 VDD.t13 1.13285
R173 VDD.n6 VDD.t11 1.13285
R174 VDD.n6 VDD.t9 1.13285
R175 VDD.n8 VDD.t27 1.13285
R176 VDD.n8 VDD.t7 1.13285
R177 VDD.n41 VDD.n0 0.161214
R178 VDD.n10 VDD.n7 0.154786
R179 VDD.n14 VDD.n7 0.154786
R180 VDD.n19 VDD.n16 0.154786
R181 VDD.n23 VDD.n4 0.154786
R182 VDD.n26 VDD.n23 0.154786
R183 VDD.n30 VDD.n3 0.154786
R184 VDD.n32 VDD.n30 0.154786
R185 VDD.n38 VDD.n0 0.154786
R186 VDD.n36 VDD.n2 0.148357
R187 VDD.n19 VDD.n18 0.109786
R188 VDD.n26 VDD.n25 0.109786
R189 VDD.n32 VDD.n31 0.109786
R190 VDD.n38 VDD.n37 0.109786
R191 VDD.n15 VDD.n14 0.0840714
R192 VDD.n16 VDD.n15 0.0712143
R193 VDD.n18 VDD.n4 0.0455
R194 VDD.n25 VDD.n3 0.0455
R195 VDD.n31 VDD.n2 0.0455
R196 VDD.n37 VDD.n36 0.0455
R197 VDD.n10 VDD.n9 0.0326429
R198 VDD VDD.n41 0.00371429
R199 a_1280_720.t0 a_1280_720.t1 3.08874
R200 a_2470_490.n2 a_2470_490.t5 40.1505
R201 a_2470_490.n0 a_2470_490.t3 37.3854
R202 a_2470_490.n2 a_2470_490.t4 30.4172
R203 a_2470_490.n0 a_2470_490.t6 29.477
R204 a_2470_490.n3 a_2470_490.n2 19.0987
R205 a_2470_490.n1 a_2470_490.n0 8.263
R206 a_2470_490.n4 a_2470_490.n3 6.4445
R207 a_2470_490.n1 a_2470_490.t2 4.47385
R208 a_2470_490.n4 a_2470_490.t1 2.03874
R209 a_2470_490.t0 a_2470_490.n4 2.03874
R210 a_2470_490.n3 a_2470_490.n1 0.5405
R211 QN.n0 QN.t2 40.0952
R212 QN.n0 QN.t3 27.3202
R213 QN.n1 QN.t1 9.27474
R214 QN.n1 QN.n0 8.0005
R215 QN QN.n2 4.5005
R216 QN.n2 QN.t0 3.39569
R217 QN.n2 QN.n1 0.1325
R218 a_250_210.n0 a_250_210.t5 48.0035
R219 a_250_210.n1 a_250_210.t3 45.6255
R220 a_250_210.n1 a_250_210.t4 20.6838
R221 a_250_210.n0 a_250_210.t2 19.4119
R222 a_250_210.n2 a_250_210.n0 17.2412
R223 a_250_210.n2 a_250_210.n1 12.5005
R224 a_250_210.t0 a_250_210.n3 8.65149
R225 a_250_210.n3 a_250_210.n2 4.87175
R226 a_250_210.n3 a_250_210.t1 3.56294
R227 Q.n0 Q.t1 9.37674
R228 Q Q.n0 4.5005
R229 Q.n0 Q.t0 2.88119
R230 a_410_720.n0 a_410_720.t6 32.5029
R231 a_410_720.n0 a_410_720.t4 31.46
R232 a_410_720.n1 a_410_720.t5 20.4405
R233 a_410_720.n3 a_410_720.n2 18.8364
R234 a_410_720.n1 a_410_720.n0 15.8172
R235 a_410_720.n2 a_410_720.t3 14.9655
R236 a_410_720.n4 a_410_720.n3 6.4085
R237 a_410_720.n3 a_410_720.t1 5.11135
R238 a_410_720.n2 a_410_720.n1 3.6505
R239 a_410_720.t0 a_410_720.n4 2.03874
R240 a_410_720.n4 a_410_720.t2 2.03874
R241 a_1720_210.t0 a_1720_210.t1 1.85344
R242 a_2110_210.n0 a_2110_210.t4 46.2338
R243 a_2110_210.n2 a_2110_210.n0 18.794
R244 a_2110_210.n0 a_2110_210.t5 16.1254
R245 a_2110_210.n2 a_2110_210.n1 10.8864
R246 a_2110_210.n3 a_2110_210.n2 7.82732
R247 a_2110_210.n1 a_2110_210.t3 3.61374
R248 a_2110_210.n1 a_2110_210.t1 3.1505
R249 a_2110_210.t0 a_2110_210.n3 1.7505
R250 a_2110_210.n3 a_2110_210.t2 1.7505
R251 a_2340_210.t0 a_2340_210.t1 7.8755
R252 CLK.n3 CLK.t2 37.1088
R253 CLK.n2 CLK.t1 34.7672
R254 CLK.n0 CLK.t0 34.1124
R255 CLK.n3 CLK.t4 30.4172
R256 CLK.n1 CLK.t3 26.8163
R257 CLK.n0 CLK.t5 24.8905
R258 CLK.n4 CLK.n3 8.0005
R259 CLK CLK.n4 4.5005
R260 CLK.n1 CLK.n0 0.8105
R261 CLK.n4 CLK.n2 0.563
R262 CLK.n2 CLK.n1 0.308
R263 S.n0 S.t2 38.1227
R264 S.n1 S.t3 35.0811
R265 S.n1 S.t1 30.4172
R266 S.n0 S.t0 26.1588
R267 S S.n0 17.4805
R268 S.n2 S.n1 12.5005
R269 S S.n2 0.0275
R270 S.n2 S 0.0275
R271 a_570_720.t0 a_570_720.n0 7.46685
R272 a_570_720.n0 a_570_720.t2 1.13285
R273 a_570_720.n0 a_570_720.t1 1.13285
R274 a_1720_720.t0 a_1720_720.t1 1.02991
R275 a_2340_720.t0 a_2340_720.t1 3.08874
R276 a_2000_210.t0 a_2000_210.t1 1.85344
R277 R.n0 R.t0 36.777
R278 R.n0 R.t1 30.0854
R279 R R.n0 12.5005
R280 a_2910_720.n0 a_2910_720.t1 7.46685
R281 a_2910_720.t0 a_2910_720.n0 1.13285
R282 a_2910_720.n0 a_2910_720.t2 1.13285
R283 a_2000_720.t0 a_2000_720.t1 1.02991
R284 a_3100_210.t0 a_3100_210.t1 1.85344
C0 CLK D 0.07514f
C1 R S 0.00839f
C2 S VDD 0.83909f
C3 R VDD 0.14182f
C4 S QN 0.01523f
C5 QN VDD 0.344f
C6 S D 0.0208f
C7 R D 0.0014f
C8 Q S 0.00694f
C9 D VDD 0.11406f
C10 Q VDD 0.15213f
C11 CLK S 0.01881f
C12 Q QN 0.32436f
C13 CLK VDD 0.5461f
C14 Q VSS 0.31322f
C15 QN VSS 0.61355f
C16 CLK VSS 0.88944f
C17 D VSS 0.31529f
C18 S VSS 0.96909f
C19 R VSS 0.38821f
C20 VDD VSS 8.70612f
.ends

