magic
tech gf180mcuD
magscale 1 10
timestamp 1757543970
<< checkpaint >>
rect -2060 1100 2704 1160
rect -2060 1040 3408 1100
rect -2060 980 4112 1040
rect -2060 -4060 4816 980
rect -1356 -4120 4816 -4060
rect -652 -4180 4816 -4120
rect 52 -4240 4816 -4180
<< error_p >>
rect 8625 2542 8636 2588
rect 8410 2379 8442 2388
rect 8373 2296 8442 2379
rect 8350 2287 8442 2296
rect 8170 2202 8200 2213
rect 8166 2197 8200 2202
rect 8272 2050 8304 2213
rect 8350 2050 8444 2287
rect 8105 1690 8116 1736
rect 8373 1699 8444 2050
rect 8373 1596 8442 1699
rect 8625 1630 8636 1676
rect 8373 1559 8433 1596
<< metal1 >>
rect 1421 1319 2322 1380
rect 2639 1322 3540 1383
rect 1421 992 2322 1053
rect 2639 995 3540 1056
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use CDAC_INV_V0  x1v
timestamp 1757543936
transform 1 0 5376 0 1 2980
box 2537 -1361 3228 577
use nfet_03v3_W5K4UP  XM1
timestamp 0
transform 1 0 322 0 1 -1450
box -382 -610 382 610
use pfet_03v3_LS6D84  XM2
timestamp 0
transform 1 0 2434 0 1 -1630
box -382 -610 382 610
use nfet_03v3_W5K4UP  XM3
timestamp 0
transform 1 0 1026 0 1 -1510
box -382 -610 382 610
use pfet_03v3_LS6D84  XM4
timestamp 0
transform 1 0 1730 0 1 -1570
box -382 -610 382 610
<< labels >>
flabel metal1 0 -2000 200 -1800 0 FreeSans 1280 0 0 0 vreflow
port 5 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 sw_Vref
port 4 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 avdd
port 3 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 avss
port 2 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 sw_bit
port 1 nsew
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 sw_vout
port 0 nsew
<< end >>
