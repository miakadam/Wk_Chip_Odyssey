magic
tech gf180mcuD
magscale 1 10
timestamp 1758003801
<< nwell >>
rect 1250 -450 1850 570
<< pwell >>
rect 1502 -539 1588 -459
rect 1250 -1170 1850 -550
<< nmos >>
rect 1500 -960 1600 -760
<< pmos >>
rect 1500 -240 1600 360
<< ndiff >>
rect 1412 -773 1500 -760
rect 1412 -947 1425 -773
rect 1471 -947 1500 -773
rect 1412 -960 1500 -947
rect 1600 -773 1688 -760
rect 1600 -947 1629 -773
rect 1675 -947 1688 -773
rect 1600 -960 1688 -947
<< pdiff >>
rect 1412 347 1500 360
rect 1412 -227 1425 347
rect 1471 -227 1500 347
rect 1412 -240 1500 -227
rect 1600 347 1688 360
rect 1600 -227 1629 347
rect 1675 -227 1688 347
rect 1600 -240 1688 -227
<< ndiffc >>
rect 1425 -947 1471 -773
rect 1629 -947 1675 -773
<< pdiffc >>
rect 1425 -227 1471 347
rect 1629 -227 1675 347
<< psubdiff >>
rect 1274 -646 1826 -574
rect 1274 -690 1346 -646
rect 1274 -1030 1287 -690
rect 1333 -1030 1346 -690
rect 1754 -690 1826 -646
rect 1274 -1074 1346 -1030
rect 1754 -1030 1767 -690
rect 1813 -1030 1826 -690
rect 1754 -1074 1826 -1030
rect 1274 -1146 1826 -1074
<< nsubdiff >>
rect 1274 474 1826 546
rect 1274 430 1346 474
rect 1274 -310 1287 430
rect 1333 -310 1346 430
rect 1754 430 1826 474
rect 1274 -354 1346 -310
rect 1754 -310 1767 430
rect 1813 -310 1826 430
rect 1754 -354 1826 -310
rect 1274 -426 1826 -354
<< psubdiffcont >>
rect 1287 -1030 1333 -690
rect 1767 -1030 1813 -690
<< nsubdiffcont >>
rect 1287 -310 1333 430
rect 1767 -310 1813 430
<< polysilicon >>
rect 1500 439 1600 452
rect 1500 393 1513 439
rect 1587 393 1600 439
rect 1500 360 1600 393
rect 1500 -273 1600 -240
rect 1500 -319 1513 -273
rect 1587 -319 1600 -273
rect 1500 -332 1600 -319
rect 1500 -681 1600 -668
rect 1500 -727 1513 -681
rect 1587 -727 1600 -681
rect 1500 -760 1600 -727
rect 1500 -993 1600 -960
rect 1500 -1039 1513 -993
rect 1587 -1039 1600 -993
rect 1500 -1052 1600 -1039
<< polycontact >>
rect 1513 393 1587 439
rect 1513 -319 1587 -273
rect 1513 -727 1587 -681
rect 1513 -1039 1587 -993
<< metal1 >>
rect 1250 570 1850 770
rect 1287 430 1333 570
rect 1502 439 1598 470
rect 1502 393 1513 439
rect 1587 393 1598 439
rect 1767 430 1813 570
rect 1333 347 1471 358
rect 1333 -227 1425 347
rect 1629 347 1675 358
rect 1612 63 1629 73
rect 1675 63 1692 73
rect 1612 -177 1624 63
rect 1680 -177 1692 63
rect 1612 -187 1629 -177
rect 1333 -238 1471 -227
rect 1675 -187 1692 -177
rect 1629 -238 1675 -227
rect 1287 -321 1333 -310
rect 1502 -319 1513 -273
rect 1587 -319 1598 -273
rect 1502 -460 1598 -319
rect 1767 -321 1813 -310
rect 1434 -472 1598 -460
rect 1434 -528 1446 -472
rect 1502 -528 1598 -472
rect 1434 -540 1598 -528
rect 1287 -690 1333 -679
rect 1502 -681 1598 -540
rect 1502 -727 1513 -681
rect 1587 -727 1598 -681
rect 1767 -690 1813 -679
rect 1333 -773 1471 -762
rect 1333 -947 1425 -773
rect 1629 -773 1675 -762
rect 1612 -832 1629 -822
rect 1675 -832 1692 -822
rect 1612 -888 1624 -832
rect 1680 -888 1692 -832
rect 1612 -898 1629 -888
rect 1333 -958 1471 -947
rect 1675 -898 1692 -888
rect 1629 -958 1675 -947
rect 1287 -1170 1333 -1030
rect 1502 -1039 1513 -993
rect 1587 -1039 1598 -993
rect 1502 -1070 1598 -1039
rect 1767 -1170 1813 -1030
rect 1250 -1370 1850 -1170
<< via1 >>
rect 1624 -177 1629 63
rect 1629 -177 1675 63
rect 1675 -177 1680 63
rect 1446 -528 1502 -472
rect 1624 -888 1629 -832
rect 1629 -888 1675 -832
rect 1675 -888 1680 -832
<< metal2 >>
rect 1612 63 1692 73
rect 1612 -177 1624 63
rect 1680 -177 1692 63
rect 1434 -472 1504 -460
rect 1250 -528 1446 -472
rect 1502 -528 1504 -472
rect 1434 -540 1504 -528
rect 1612 -472 1692 -177
rect 1612 -528 1850 -472
rect 1612 -832 1692 -528
rect 1612 -888 1624 -832
rect 1680 -888 1692 -832
rect 1612 -898 1692 -888
<< labels >>
rlabel metal2 1250 -499 1250 -499 7 in
port 0 w
rlabel metal1 1545 770 1545 770 1 vdd
port 1 n
rlabel metal2 1850 -499 1850 -499 3 out
port 2 e
rlabel metal1 1555 -1370 1555 -1370 5 vss
port 3 s
<< end >>
