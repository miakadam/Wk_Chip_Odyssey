magic
tech gf180mcuD
magscale 1 10
timestamp 1755250623
<< error_s >>
rect 4324 437 4616 446
rect 4904 437 5196 446
rect 4368 388 4370 400
rect 4380 354 4382 400
rect 4558 398 4560 400
rect 4570 388 4572 400
rect 4948 388 4950 400
rect 4960 366 4966 410
rect 4960 354 4986 366
rect 4370 352 4382 354
rect 4368 340 4382 352
rect 4560 352 4570 354
rect 4950 352 4986 354
rect 4560 342 4572 352
rect 4558 340 4572 342
rect 4948 340 4986 352
rect 5138 354 5140 400
rect 5150 388 5152 400
rect 5138 352 5150 354
rect 5138 340 5152 352
rect 4960 330 4986 340
rect 4858 288 4860 300
rect 4858 180 4860 192
rect 4870 180 4872 192
rect 4928 180 4930 300
rect 4940 288 4942 300
rect 4940 180 4942 192
rect 2754 -63 2936 -54
rect 3454 -63 3636 -54
rect 5864 -63 6036 -44
rect 6674 -63 6846 -54
rect 2798 -112 2800 -100
rect 2810 -146 2812 -100
rect 2878 -134 2880 -100
rect 2890 -112 2892 -100
rect 3498 -112 3500 -100
rect 2800 -157 2825 -146
rect 2864 -157 2890 -134
rect 3510 -144 3512 -100
rect 3578 -124 3580 -100
rect 3590 -112 3592 -100
rect 5908 -102 5922 -90
rect 4578 -122 4580 -110
rect 3544 -134 3580 -124
rect 2800 -158 2837 -157
rect 2798 -170 2837 -158
rect 2859 -158 2890 -157
rect 3500 -157 3525 -144
rect 3534 -157 3590 -134
rect 3500 -158 3590 -157
rect 2859 -170 2892 -158
rect 3498 -170 3592 -158
rect 3544 -180 3580 -170
rect 2745 -268 2791 -192
rect 3588 -202 3590 -190
rect 3600 -257 3602 -190
rect 2905 -268 2928 -257
rect 2910 -290 2928 -268
rect 3468 -268 3491 -257
rect 3590 -258 3628 -257
rect 3468 -280 3490 -268
rect 3588 -270 3628 -258
rect 3658 -270 3660 -190
rect 3670 -202 3672 -190
rect 4590 -254 4592 -110
rect 4660 -122 4662 -110
rect 4848 -122 4850 -110
rect 3670 -270 3672 -258
rect 4590 -264 4616 -254
rect 4860 -264 4862 -110
rect 4928 -254 4930 -110
rect 4940 -122 4942 -110
rect 5910 -124 5922 -102
rect 5978 -124 5980 -90
rect 5990 -102 5992 -90
rect 6718 -112 6732 -100
rect 6720 -124 6732 -112
rect 5910 -148 5956 -124
rect 5908 -160 5956 -148
rect 5964 -148 5990 -124
rect 5964 -157 5992 -148
rect 5959 -160 5992 -157
rect 6720 -157 6746 -124
rect 6788 -146 6790 -100
rect 6800 -112 6802 -100
rect 6781 -157 6800 -146
rect 6720 -158 6747 -157
rect 5920 -170 5956 -160
rect 6718 -170 6747 -158
rect 6769 -158 6800 -157
rect 6769 -170 6802 -158
rect 5818 -202 5820 -190
rect 4904 -264 4930 -254
rect 5898 -257 5900 -190
rect 5910 -202 5912 -190
rect 4580 -268 4626 -264
rect 4578 -280 4626 -268
rect 4660 -280 4662 -268
rect 4860 -278 4940 -264
rect 4324 -288 4341 -280
rect 4580 -290 4626 -280
rect 4848 -290 4850 -278
rect 4860 -290 4942 -278
rect 5179 -288 5196 -277
rect 5818 -280 5820 -268
rect 5868 -270 5910 -257
rect 6005 -268 6028 -257
rect 6010 -270 6028 -268
rect 6664 -268 6701 -244
rect 6815 -268 6861 -192
rect 5868 -280 5912 -270
rect 6664 -280 6700 -268
rect 4590 -300 4626 -290
rect 4860 -300 4930 -290
rect 2814 -349 2825 -303
rect 3514 -349 3525 -303
rect 4368 -332 4370 -320
rect 4368 -371 4370 -368
rect 4380 -371 4382 -320
rect 4558 -371 4560 -320
rect 4570 -332 4572 -320
rect 4570 -371 4572 -368
rect 4368 -380 4572 -371
rect 4600 -380 4626 -300
rect 4894 -320 4920 -300
rect 6708 -302 6710 -290
rect 4948 -332 4976 -320
rect 4950 -368 4976 -332
rect 4948 -371 4976 -368
rect 5138 -371 5140 -320
rect 5150 -332 5152 -320
rect 5914 -349 5925 -303
rect 6708 -351 6710 -348
rect 6720 -351 6722 -290
rect 6788 -351 6790 -290
rect 6800 -302 6802 -290
rect 6800 -351 6802 -348
rect 6708 -360 6802 -351
rect 5150 -371 5152 -368
rect 4948 -380 5152 -371
rect 4314 -743 4626 -734
rect 4680 -770 4686 -604
rect 4884 -734 4910 -724
rect 4884 -743 5206 -734
rect 4620 -780 4626 -770
rect 4884 -780 4910 -743
rect 4358 -792 4360 -780
rect 4370 -826 4372 -780
rect 4568 -814 4570 -780
rect 4580 -792 4582 -780
rect 4938 -792 4966 -780
rect 4940 -814 4966 -792
rect 4544 -826 4570 -814
rect 4804 -824 4986 -814
rect 4360 -828 4383 -826
rect 4358 -837 4383 -828
rect 4544 -828 4580 -826
rect 4358 -840 4387 -837
rect 4544 -840 4582 -828
rect 4804 -840 4996 -824
rect 5148 -826 5150 -780
rect 5160 -792 5162 -780
rect 5137 -828 5160 -826
rect 5137 -837 5162 -828
rect 5133 -840 5162 -837
rect 4544 -850 4570 -840
rect 4620 -850 4626 -840
rect 4950 -850 4986 -840
rect 4600 -1040 4602 -880
rect 4680 -892 4682 -880
rect 4848 -892 4850 -880
rect 4668 -1040 4670 -1038
rect 4680 -1040 4682 -1028
rect 4848 -1040 4850 -1028
rect 4860 -1040 4862 -880
rect 4928 -1040 4930 -880
rect 4940 -892 4942 -880
rect 4940 -1040 4942 -1028
rect 3054 -1351 3236 -1334
rect 6324 -1351 6506 -1334
rect 3098 -1392 3100 -1380
rect 3110 -1434 3112 -1380
rect 3190 -1392 3192 -1380
rect 6368 -1392 6370 -1380
rect 6380 -1434 6382 -1380
rect 6448 -1434 6450 -1380
rect 6460 -1392 6462 -1380
rect 3100 -1438 3125 -1434
rect 3098 -1445 3125 -1438
rect 3171 -1438 3190 -1434
rect 6370 -1438 6395 -1434
rect 3171 -1445 3192 -1438
rect 3098 -1450 3137 -1445
rect 3159 -1450 3192 -1445
rect 6368 -1445 6395 -1438
rect 6441 -1438 6460 -1434
rect 6441 -1445 6462 -1438
rect 6368 -1450 6407 -1445
rect 6429 -1450 6462 -1445
rect 3064 -1556 3091 -1534
rect 3205 -1545 3226 -1534
rect 6344 -1545 6361 -1524
rect 3205 -1556 3228 -1545
rect 3064 -1580 3090 -1556
rect 3110 -1724 3136 -1580
rect 3210 -1637 3228 -1556
rect 6338 -1556 6361 -1545
rect 6475 -1556 6506 -1524
rect 6338 -1591 6360 -1556
rect 6390 -1591 6406 -1570
rect 4278 -1612 4280 -1600
rect 3210 -1665 3226 -1637
rect 3744 -1663 3926 -1654
rect 3090 -1730 3136 -1724
rect 3144 -1711 3180 -1684
rect 3144 -1730 3182 -1711
rect 3210 -1730 3228 -1665
rect 3788 -1710 3790 -1700
rect 3800 -1724 3802 -1700
rect 3880 -1710 3882 -1700
rect 3018 -1870 3020 -1858
rect 3030 -1870 3032 -1730
rect 3098 -1857 3100 -1730
rect 3188 -1742 3228 -1730
rect 3190 -1757 3228 -1742
rect 3190 -1770 3226 -1757
rect 3200 -1857 3202 -1770
rect 3068 -1858 3110 -1857
rect 3190 -1858 3228 -1857
rect 3068 -1870 3112 -1858
rect 3188 -1870 3228 -1858
rect 3268 -1870 3270 -1730
rect 3800 -1738 3836 -1724
rect 3800 -1744 3870 -1738
rect 3790 -1758 3880 -1744
rect 3788 -1770 3882 -1758
rect 3800 -1780 3836 -1770
rect 3890 -1780 3936 -1724
rect 3698 -1802 3700 -1790
rect 3280 -1870 3282 -1858
rect 3698 -1870 3700 -1858
rect 3710 -1870 3712 -1790
rect 3778 -1857 3780 -1790
rect 3790 -1802 3792 -1790
rect 3868 -1802 3870 -1790
rect 3880 -1857 3882 -1790
rect 3748 -1858 3790 -1857
rect 3870 -1858 3908 -1857
rect 3748 -1870 3792 -1858
rect 3868 -1870 3908 -1858
rect 3948 -1870 3950 -1790
rect 3960 -1802 3962 -1790
rect 3960 -1870 3962 -1858
rect 4278 -1870 4280 -1858
rect 4290 -1870 4292 -1600
rect 4348 -1857 4350 -1600
rect 4360 -1612 4362 -1600
rect 5158 -1612 5160 -1600
rect 5170 -1857 5172 -1600
rect 4326 -1858 4360 -1857
rect 5160 -1858 5194 -1857
rect 4326 -1870 4362 -1858
rect 5158 -1870 5194 -1858
rect 5228 -1870 5230 -1600
rect 5240 -1612 5242 -1600
rect 6384 -1637 6406 -1591
rect 5644 -1663 5826 -1654
rect 5688 -1710 5690 -1700
rect 5700 -1714 5746 -1690
rect 5768 -1714 5770 -1700
rect 5780 -1710 5782 -1700
rect 6338 -1711 6360 -1665
rect 6390 -1684 6406 -1637
rect 6390 -1711 6426 -1684
rect 5700 -1744 5770 -1714
rect 5690 -1758 5780 -1744
rect 5688 -1770 5782 -1758
rect 5700 -1780 5746 -1770
rect 5790 -1780 5826 -1770
rect 5608 -1802 5610 -1790
rect 5240 -1870 5242 -1858
rect 5608 -1870 5610 -1858
rect 5620 -1870 5622 -1790
rect 5688 -1857 5690 -1790
rect 5700 -1802 5702 -1790
rect 5778 -1802 5780 -1790
rect 5790 -1857 5792 -1790
rect 5658 -1858 5700 -1857
rect 5780 -1858 5818 -1857
rect 5658 -1870 5702 -1858
rect 5778 -1870 5818 -1858
rect 5858 -1870 5860 -1790
rect 5870 -1802 5872 -1790
rect 5870 -1870 5872 -1858
rect 6288 -1870 6290 -1858
rect 6300 -1870 6302 -1730
rect 6368 -1857 6370 -1730
rect 6380 -1742 6382 -1730
rect 6384 -1757 6426 -1711
rect 6480 -1714 6506 -1556
rect 6460 -1730 6506 -1714
rect 6390 -1760 6426 -1757
rect 6470 -1857 6472 -1730
rect 6338 -1858 6380 -1857
rect 6460 -1858 6498 -1857
rect 6338 -1870 6382 -1858
rect 6458 -1870 6498 -1858
rect 6538 -1870 6540 -1730
rect 6550 -1870 6552 -1858
rect 3114 -1949 3125 -1903
rect 3794 -1949 3805 -1903
rect 5704 -1949 5715 -1903
rect 6384 -1949 6395 -1903
rect 3124 -2384 3135 -2355
rect 3124 -2401 3192 -2384
rect 3804 -2394 3815 -2357
rect 4402 -2377 4436 -2364
rect 5144 -2377 5178 -2364
rect 3861 -2394 3872 -2392
rect 3804 -2403 3872 -2394
rect 5704 -2394 5715 -2357
rect 5761 -2394 5772 -2392
rect 5704 -2403 5772 -2394
rect 4308 -2422 4310 -2410
rect 3028 -2442 3030 -2430
rect 3040 -2570 3042 -2430
rect 3108 -2484 3110 -2430
rect 3120 -2442 3122 -2430
rect 3198 -2442 3200 -2430
rect 3084 -2501 3120 -2484
rect 3078 -2547 3120 -2501
rect 3154 -2530 3200 -2524
rect 3130 -2547 3166 -2530
rect 3108 -2570 3110 -2547
rect 3124 -2570 3166 -2547
rect 3210 -2570 3212 -2430
rect 3278 -2570 3280 -2430
rect 3290 -2442 3292 -2430
rect 3708 -2452 3710 -2440
rect 3788 -2484 3790 -2440
rect 3800 -2452 3802 -2440
rect 3878 -2452 3880 -2440
rect 3764 -2503 3800 -2484
rect 3758 -2549 3800 -2503
rect 3810 -2549 3846 -2530
rect 3124 -2593 3156 -2570
rect 3078 -2667 3110 -2621
rect 3130 -2667 3156 -2593
rect 3124 -2713 3156 -2667
rect 3130 -2720 3156 -2713
rect 3210 -2720 3246 -2570
rect 3720 -2580 3722 -2578
rect 3788 -2580 3790 -2549
rect 3800 -2580 3802 -2568
rect 3804 -2580 3846 -2549
rect 3890 -2580 3892 -2440
rect 3958 -2580 3960 -2440
rect 3970 -2452 3972 -2440
rect 3970 -2580 3972 -2568
rect 3804 -2595 3826 -2580
rect 3758 -2669 3780 -2623
rect 3810 -2669 3826 -2595
rect 3804 -2715 3826 -2669
rect 3810 -2720 3827 -2715
rect 3890 -2720 3926 -2580
rect 4308 -2680 4310 -2668
rect 4320 -2680 4322 -2518
rect 4378 -2680 4380 -2410
rect 4390 -2422 4392 -2410
rect 5188 -2422 5190 -2410
rect 4390 -2680 4392 -2668
rect 5188 -2680 5190 -2668
rect 5200 -2680 5202 -2410
rect 5270 -2422 5272 -2410
rect 5608 -2452 5610 -2440
rect 5258 -2680 5260 -2528
rect 5620 -2580 5622 -2440
rect 5688 -2484 5690 -2440
rect 5700 -2452 5702 -2440
rect 5778 -2452 5780 -2440
rect 5664 -2503 5700 -2484
rect 5658 -2549 5700 -2503
rect 5710 -2549 5746 -2530
rect 5688 -2580 5690 -2549
rect 5700 -2580 5702 -2568
rect 5704 -2580 5746 -2549
rect 5790 -2580 5792 -2440
rect 5858 -2580 5860 -2440
rect 5870 -2452 5872 -2440
rect 5870 -2580 5872 -2568
rect 5704 -2595 5726 -2580
rect 5270 -2680 5272 -2668
rect 5658 -2669 5680 -2623
rect 5710 -2669 5726 -2595
rect 5704 -2715 5726 -2669
rect 5710 -2720 5727 -2715
rect 5790 -2720 5826 -2580
rect 3084 -2813 3110 -2794
rect 3078 -2859 3110 -2813
rect 3130 -2859 3156 -2840
rect 3124 -2905 3156 -2859
rect 3078 -2979 3110 -2933
rect 3130 -2979 3156 -2905
rect 3124 -3025 3156 -2979
rect 3130 -3030 3156 -3025
rect 3210 -3030 3246 -2794
rect 3764 -2815 3781 -2794
rect 3758 -2826 3781 -2815
rect 3758 -2861 3780 -2826
rect 3810 -2861 3826 -2840
rect 3804 -2907 3826 -2861
rect 3758 -2981 3780 -2935
rect 3810 -2981 3826 -2907
rect 3804 -3027 3826 -2981
rect 3810 -3030 3827 -3027
rect 3890 -3030 3926 -2794
rect 5664 -2815 5681 -2804
rect 5658 -2826 5681 -2815
rect 5658 -2861 5680 -2826
rect 5710 -2861 5726 -2850
rect 5704 -2907 5726 -2861
rect 5658 -2981 5680 -2935
rect 5710 -2981 5726 -2907
rect 5704 -3027 5726 -2981
rect 5710 -3040 5727 -3027
rect 5790 -3040 5826 -2804
rect 3084 -3125 3110 -3104
rect 3078 -3171 3110 -3125
rect 3130 -3171 3156 -3150
rect 3124 -3217 3156 -3171
rect 3078 -3291 3110 -3245
rect 3130 -3291 3156 -3217
rect 3124 -3337 3156 -3291
rect 3130 -3340 3156 -3337
rect 3210 -3340 3246 -3104
rect 3754 -3138 3781 -3114
rect 3890 -3127 3916 -3114
rect 5664 -3127 5681 -3114
rect 3754 -3160 3780 -3138
rect 3800 -3339 3826 -3160
rect 3890 -3219 3918 -3127
rect 5658 -3138 5681 -3127
rect 5658 -3173 5680 -3138
rect 5710 -3173 5726 -3160
rect 5704 -3219 5726 -3173
rect 3890 -3247 3916 -3219
rect 3890 -3339 3918 -3247
rect 5658 -3293 5680 -3247
rect 5710 -3293 5726 -3219
rect 5704 -3339 5726 -3293
rect 3800 -3350 3827 -3339
rect 3890 -3350 3916 -3339
rect 5710 -3350 5727 -3339
rect 5790 -3350 5826 -3114
rect 3064 -3450 3110 -3424
rect 3210 -3450 3246 -3424
rect 3754 -3450 3781 -3434
rect 3890 -3439 3895 -3434
rect 5664 -3439 5681 -3424
rect 3108 -3482 3110 -3470
rect 3120 -3472 3122 -3470
rect 3108 -3531 3110 -3528
rect 3188 -3531 3190 -3470
rect 3200 -3482 3202 -3470
rect 3754 -3480 3780 -3450
rect 3200 -3531 3202 -3528
rect 3108 -3540 3202 -3531
rect 3800 -3651 3826 -3480
rect 3890 -3531 3918 -3439
rect 5658 -3450 5681 -3439
rect 5658 -3485 5680 -3450
rect 5710 -3485 5726 -3470
rect 5704 -3531 5726 -3485
rect 3890 -3559 3916 -3531
rect 3890 -3651 3918 -3559
rect 5658 -3605 5680 -3559
rect 5710 -3605 5726 -3531
rect 5704 -3651 5726 -3605
rect 3800 -3670 3827 -3651
rect 3890 -3670 3916 -3651
rect 5710 -3660 5727 -3651
rect 5790 -3660 5826 -3424
rect 6130 -3660 6136 -2224
rect 6374 -2384 6385 -2355
rect 6374 -2401 6442 -2384
rect 6448 -2440 6450 -2430
rect 6290 -2580 6292 -2440
rect 6358 -2580 6360 -2440
rect 6460 -2484 6462 -2430
rect 6450 -2501 6486 -2484
rect 6450 -2570 6488 -2501
rect 6528 -2570 6530 -2430
rect 6540 -2442 6542 -2430
rect 6370 -2720 6406 -2580
rect 6460 -2593 6488 -2570
rect 6460 -2621 6486 -2593
rect 6460 -2713 6488 -2621
rect 6460 -2720 6486 -2713
rect 6324 -2840 6360 -2794
rect 6460 -2813 6486 -2794
rect 6370 -3030 6406 -2840
rect 6460 -2905 6488 -2813
rect 6460 -2933 6486 -2905
rect 6460 -3025 6488 -2933
rect 6460 -3030 6486 -3025
rect 6334 -3125 6360 -3114
rect 6328 -3171 6360 -3125
rect 6380 -3171 6406 -3160
rect 6374 -3217 6406 -3171
rect 6328 -3291 6360 -3245
rect 6380 -3291 6406 -3217
rect 6374 -3337 6406 -3291
rect 6380 -3350 6406 -3337
rect 6460 -3350 6496 -3114
rect 6314 -3450 6360 -3424
rect 6460 -3450 6496 -3424
rect 6358 -3482 6360 -3470
rect 6358 -3531 6360 -3528
rect 6370 -3531 6372 -3470
rect 6438 -3531 6440 -3470
rect 6450 -3482 6452 -3470
rect 6450 -3531 6452 -3528
rect 6358 -3540 6452 -3531
rect 3764 -3751 3781 -3734
rect 3758 -3762 3781 -3751
rect 3758 -3797 3780 -3762
rect 3810 -3797 3826 -3780
rect 3804 -3843 3826 -3797
rect 3758 -3917 3780 -3871
rect 3810 -3917 3826 -3843
rect 3804 -3963 3826 -3917
rect 3810 -3970 3827 -3963
rect 3890 -3970 3926 -3734
rect 5664 -3751 5681 -3734
rect 5658 -3762 5681 -3751
rect 5658 -3797 5680 -3762
rect 5710 -3797 5726 -3780
rect 5704 -3843 5726 -3797
rect 5658 -3917 5680 -3871
rect 5710 -3917 5726 -3843
rect 5704 -3963 5726 -3917
rect 5710 -3970 5727 -3963
rect 5790 -3970 5826 -3734
rect 3764 -4063 3781 -4044
rect 3758 -4074 3781 -4063
rect 3758 -4109 3780 -4074
rect 3810 -4109 3826 -4090
rect 3804 -4155 3826 -4109
rect 3758 -4229 3780 -4183
rect 3810 -4229 3826 -4155
rect 3804 -4275 3826 -4229
rect 3810 -4280 3827 -4275
rect 3890 -4280 3926 -4044
rect 5664 -4063 5681 -4044
rect 5658 -4074 5681 -4063
rect 5658 -4109 5680 -4074
rect 5710 -4109 5726 -4090
rect 5704 -4155 5726 -4109
rect 5658 -4229 5680 -4183
rect 5710 -4229 5726 -4155
rect 5704 -4275 5726 -4229
rect 5710 -4280 5727 -4275
rect 5790 -4280 5826 -4044
rect 3764 -4375 3781 -4364
rect 3758 -4386 3781 -4375
rect 3758 -4421 3780 -4386
rect 3810 -4421 3826 -4410
rect 3804 -4467 3826 -4421
rect 3758 -4541 3780 -4495
rect 3810 -4541 3826 -4467
rect 3804 -4587 3826 -4541
rect 3810 -4600 3827 -4587
rect 3890 -4600 3926 -4364
rect 5664 -4375 5681 -4364
rect 5658 -4386 5681 -4375
rect 5658 -4421 5680 -4386
rect 5710 -4421 5726 -4410
rect 5704 -4467 5726 -4421
rect 5658 -4541 5680 -4495
rect 5710 -4541 5726 -4467
rect 5704 -4587 5726 -4541
rect 5710 -4600 5727 -4587
rect 5790 -4600 5826 -4364
rect 3754 -4698 3781 -4674
rect 3754 -4700 3780 -4698
rect 3890 -4700 3936 -4674
rect 5644 -4698 5681 -4674
rect 5644 -4700 5680 -4698
rect 5790 -4700 5826 -4674
rect 3798 -4732 3800 -4720
rect 3798 -4781 3800 -4778
rect 3810 -4781 3812 -4720
rect 3878 -4722 3880 -4720
rect 3890 -4732 3892 -4720
rect 5688 -4732 5690 -4720
rect 3890 -4781 3892 -4778
rect 3798 -4790 3892 -4781
rect 5688 -4781 5690 -4778
rect 5700 -4781 5702 -4720
rect 5768 -4781 5770 -4720
rect 5780 -4732 5782 -4720
rect 5780 -4781 5782 -4778
rect 5688 -4790 5782 -4781
rect 4608 -5152 4610 -5140
rect 4620 -5364 4622 -5140
rect 4620 -5384 4646 -5364
rect 4344 -5408 4371 -5384
rect 4610 -5398 4646 -5384
rect 4608 -5410 4646 -5398
rect 4678 -5410 4680 -5140
rect 4690 -5152 4692 -5140
rect 4888 -5152 4890 -5140
rect 4900 -5372 4902 -5140
rect 4958 -5364 4960 -5140
rect 4970 -5152 4972 -5140
rect 4934 -5384 4960 -5364
rect 4934 -5398 4970 -5384
rect 4690 -5410 4692 -5398
rect 4888 -5410 4890 -5398
rect 4934 -5410 4972 -5398
rect 5209 -5408 5236 -5384
rect 4620 -5430 4646 -5410
rect 4934 -5420 4960 -5410
rect 4388 -5442 4390 -5430
rect 4388 -5491 4390 -5488
rect 4588 -5491 4590 -5430
rect 4600 -5442 4602 -5430
rect 4978 -5442 4980 -5430
rect 4600 -5491 4602 -5488
rect 4388 -5500 4602 -5491
rect 4978 -5491 4980 -5488
rect 4990 -5491 5016 -5420
rect 5178 -5491 5180 -5430
rect 5190 -5442 5192 -5430
rect 5190 -5491 5192 -5488
rect 4978 -5500 5192 -5491
rect 4620 -5510 4646 -5500
rect 4990 -5510 5016 -5500
rect 4738 -5874 4749 -5841
rect 4738 -5887 4766 -5874
rect 4774 -5887 4806 -5874
rect 4818 -5932 4820 -5920
rect 4830 -5964 4832 -5920
rect 4830 -5984 4866 -5964
rect 4684 -6000 4720 -5984
rect 4820 -5988 4866 -5984
rect 4818 -6000 4866 -5988
rect 4888 -6000 4890 -5928
rect 4900 -5932 4902 -5920
rect 4900 -6000 4902 -5988
rect 4830 -6010 4866 -6000
rect 4728 -6042 4730 -6030
rect 4740 -6032 4742 -6030
rect 4808 -6074 4810 -6030
rect 4820 -6042 4822 -6030
rect 4730 -6088 4820 -6074
rect 4728 -6100 4822 -6088
<< nwell >>
rect 4580 340 4680 390
rect 4860 380 4910 400
rect 4850 190 4910 380
rect 4620 -380 4680 -110
<< pwell >>
rect 4840 -840 4910 -610
rect 4290 -2300 4350 -2030
<< metal1 >>
rect 2610 440 4210 560
rect 2610 290 4190 440
rect 4370 340 4380 400
rect 4560 340 4570 400
rect 4950 340 4960 400
rect 5140 340 5150 400
rect 2610 -50 4330 290
rect 3060 -60 3310 -50
rect 2800 -170 2810 -100
rect 2880 -170 2890 -100
rect 3060 -180 3350 -60
rect 3500 -170 3510 -100
rect 3580 -170 3590 -100
rect 2910 -190 3350 -180
rect 2910 -280 3490 -190
rect 3590 -270 3600 -190
rect 3660 -270 3670 -190
rect 3750 -280 4330 -50
rect 2910 -290 3350 -280
rect 3060 -420 3350 -290
rect 3750 -430 4180 -280
rect 4430 -320 4510 340
rect 4860 180 4870 300
rect 4930 180 4940 300
rect 4580 -280 4590 -110
rect 4650 -280 4660 -110
rect 4850 -290 4860 -110
rect 4930 -290 4940 -110
rect 5010 -320 5090 340
rect 5340 300 5730 520
rect 5190 -180 5730 300
rect 5910 -160 5920 -90
rect 5980 -160 5990 -90
rect 6160 -170 6550 510
rect 6720 -170 6730 -100
rect 6790 -170 6800 -100
rect 5190 -270 5710 -180
rect 5340 -280 5710 -270
rect 5820 -280 5830 -190
rect 5900 -280 5910 -190
rect 6010 -270 6700 -170
rect 6160 -280 6700 -270
rect 6970 -280 7000 -180
rect 4370 -380 4380 -320
rect 4560 -380 4570 -320
rect 4950 -380 4960 -320
rect 5140 -380 5150 -320
rect 5340 -410 5730 -280
rect 6160 -420 6550 -280
rect 6710 -360 6720 -290
rect 6790 -360 6800 -290
rect 4360 -840 4370 -780
rect 4570 -840 4580 -780
rect 4940 -840 4950 -780
rect 5150 -840 5160 -780
rect 3100 -1450 3110 -1380
rect 3180 -1450 3190 -1380
rect 3030 -1730 3090 -1480
rect 3110 -1730 3180 -1580
rect 3210 -1730 3270 -1480
rect 3020 -1870 3030 -1730
rect 3100 -1770 3180 -1730
rect 3100 -1870 3110 -1770
rect 3190 -1870 3200 -1730
rect 3270 -1870 3280 -1730
rect 3790 -1770 3800 -1700
rect 3870 -1770 3880 -1700
rect 3700 -1870 3710 -1790
rect 3780 -1870 3790 -1790
rect 3870 -1870 3880 -1790
rect 3950 -1870 3960 -1790
rect 4280 -1870 4290 -1600
rect 4350 -1870 4360 -1600
rect 4430 -1940 4490 -840
rect 4590 -1040 4600 -880
rect 4670 -1040 4680 -880
rect 4850 -1040 4860 -880
rect 4930 -1040 4940 -880
rect 5020 -1940 5080 -840
rect 6370 -1450 6380 -1380
rect 6450 -1450 6460 -1380
rect 5160 -1870 5170 -1600
rect 5230 -1870 5240 -1600
rect 5690 -1770 5700 -1700
rect 5770 -1770 5780 -1700
rect 6300 -1730 6360 -1480
rect 6390 -1730 6460 -1570
rect 6480 -1730 6540 -1480
rect 5610 -1870 5620 -1790
rect 5690 -1870 5700 -1790
rect 5780 -1870 5790 -1790
rect 5860 -1870 5870 -1790
rect 6290 -1870 6300 -1730
rect 6370 -1870 6380 -1730
rect 6390 -1760 6470 -1730
rect 6460 -1870 6470 -1760
rect 6540 -1870 6550 -1730
rect 3030 -2570 3040 -2430
rect 3110 -2570 3120 -2430
rect 3200 -2530 3210 -2430
rect 3130 -2570 3210 -2530
rect 3280 -2570 3290 -2430
rect 3040 -3450 3110 -2570
rect 3130 -2720 3200 -2570
rect 3130 -3030 3200 -2840
rect 3130 -3340 3200 -3150
rect 3210 -3450 3280 -2570
rect 3710 -2580 3720 -2440
rect 3790 -2580 3800 -2440
rect 3880 -2530 3890 -2440
rect 3810 -2580 3890 -2530
rect 3960 -2580 3970 -2440
rect 3110 -3540 3120 -3470
rect 3190 -3540 3200 -3470
rect 3720 -4700 3780 -2580
rect 3810 -2720 3880 -2580
rect 3810 -3030 3880 -2840
rect 3800 -3350 3870 -3160
rect 3800 -3670 3870 -3480
rect 3810 -3970 3880 -3780
rect 3810 -4280 3880 -4090
rect 3810 -4600 3880 -4410
rect 3890 -4700 3950 -2580
rect 4310 -2680 4320 -2410
rect 4380 -2680 4390 -2410
rect 3800 -4790 3810 -4720
rect 3880 -4790 3890 -4720
rect 4470 -5430 4540 -2350
rect 4610 -5410 4620 -5140
rect 4680 -5410 4690 -5140
rect 4890 -5410 4900 -5140
rect 4960 -5410 4970 -5140
rect 5060 -5430 5130 -2340
rect 5190 -2680 5200 -2410
rect 5260 -2680 5270 -2410
rect 6290 -2440 6360 -2430
rect 5610 -2580 5620 -2440
rect 5690 -2580 5700 -2440
rect 5780 -2530 5790 -2440
rect 5710 -2580 5790 -2530
rect 5860 -2580 5870 -2440
rect 6280 -2580 6290 -2440
rect 6360 -2530 6370 -2440
rect 6360 -2580 6440 -2530
rect 6450 -2570 6460 -2430
rect 6530 -2570 6540 -2430
rect 5620 -4700 5680 -2580
rect 5710 -2720 5780 -2580
rect 5710 -3040 5780 -2850
rect 5710 -3350 5780 -3160
rect 5710 -3660 5780 -3470
rect 5710 -3970 5780 -3780
rect 5710 -4280 5780 -4090
rect 5710 -4600 5780 -4410
rect 5790 -4700 5850 -2580
rect 6290 -3450 6360 -2580
rect 6370 -2720 6440 -2580
rect 6370 -3030 6440 -2840
rect 6380 -3350 6450 -3160
rect 6460 -3450 6530 -2570
rect 6360 -3540 6370 -3470
rect 6440 -3540 6450 -3470
rect 5690 -4790 5700 -4720
rect 5770 -4790 5780 -4720
rect 4390 -5500 4400 -5430
rect 4590 -5500 4600 -5430
rect 4980 -5500 4990 -5430
rect 5180 -5500 5190 -5430
rect 4560 -6000 4720 -5920
rect 4820 -6000 4830 -5920
rect 4890 -6000 4900 -5920
rect 4730 -6100 4740 -6030
rect 4810 -6100 4820 -6030
rect 3100 -6260 4460 -6120
<< via1 >>
rect 4380 340 4560 400
rect 4960 340 5140 400
rect 2810 -170 2880 -100
rect 3510 -170 3580 -100
rect 3600 -270 3660 -190
rect 4870 180 4930 300
rect 4590 -280 4650 -110
rect 4860 -290 4930 -110
rect 5920 -160 5980 -90
rect 6730 -170 6790 -100
rect 5830 -280 5900 -190
rect 4380 -380 4560 -320
rect 4960 -380 5140 -320
rect 6720 -360 6790 -290
rect 4370 -840 4570 -780
rect 4950 -840 5150 -780
rect 3110 -1450 3180 -1380
rect 3030 -1870 3100 -1730
rect 3200 -1870 3270 -1730
rect 3800 -1770 3870 -1700
rect 3710 -1870 3780 -1790
rect 3880 -1870 3950 -1790
rect 4290 -1870 4350 -1600
rect 4600 -1040 4670 -880
rect 4860 -1040 4930 -880
rect 6380 -1450 6450 -1380
rect 5170 -1870 5230 -1600
rect 5700 -1770 5770 -1700
rect 5620 -1870 5690 -1790
rect 5790 -1870 5860 -1790
rect 6300 -1870 6370 -1730
rect 6470 -1870 6540 -1730
rect 3040 -2570 3110 -2430
rect 3210 -2570 3280 -2430
rect 3720 -2580 3790 -2440
rect 3890 -2580 3960 -2440
rect 3120 -3540 3190 -3470
rect 4320 -2680 4380 -2410
rect 3810 -4790 3880 -4720
rect 4620 -5410 4680 -5140
rect 4900 -5410 4960 -5140
rect 5200 -2680 5260 -2410
rect 5620 -2580 5690 -2440
rect 5790 -2580 5860 -2440
rect 6290 -2580 6360 -2440
rect 6460 -2570 6530 -2430
rect 6370 -3540 6440 -3470
rect 5700 -4790 5770 -4720
rect 4400 -5500 4590 -5430
rect 4990 -5500 5180 -5430
rect 4830 -6000 4890 -5920
rect 4740 -6100 4810 -6030
<< metal2 >>
rect 2810 660 2880 720
rect 3510 660 3580 720
rect 2620 580 6790 660
rect 2810 -100 2880 580
rect 2810 -180 2880 -170
rect 3510 -100 3580 580
rect 4380 400 4560 410
rect 4960 400 5140 410
rect 4560 340 4910 400
rect 4380 330 4560 340
rect 4850 310 4910 340
rect 4960 330 5140 340
rect 4850 300 4930 310
rect 4850 190 4870 300
rect 4870 170 4930 180
rect 5920 -90 5980 580
rect 3510 -180 3580 -170
rect 4590 -110 4660 -100
rect 4860 -110 4930 -100
rect 3600 -190 3660 -180
rect 3600 -280 3660 -270
rect 4660 -290 4680 -110
rect 4590 -300 4680 -290
rect 5920 -170 5980 -160
rect 6730 -100 6790 580
rect 6730 -180 6790 -170
rect 5820 -190 5900 -180
rect 5820 -290 5900 -280
rect 6720 -290 6790 -280
rect 4860 -300 4930 -290
rect 4380 -320 4560 -310
rect 4620 -320 4680 -300
rect 4960 -320 5140 -310
rect 4620 -380 4960 -320
rect 4380 -390 4560 -380
rect 4960 -390 5140 -380
rect 6720 -480 6790 -360
rect 4550 -540 4670 -530
rect 4860 -540 4980 -530
rect 4670 -650 4680 -580
rect 4550 -660 4680 -650
rect 6710 -560 6960 -480
rect 4860 -660 4980 -650
rect 4630 -770 4680 -660
rect 4370 -780 4570 -770
rect 2400 -910 3900 -810
rect 4370 -850 4570 -840
rect 4620 -780 5150 -770
rect 4620 -840 4950 -780
rect 4620 -870 4680 -840
rect 4950 -850 5150 -840
rect 3800 -940 3900 -910
rect 4600 -880 4680 -870
rect 2410 -1190 3200 -1080
rect 3110 -1380 3190 -1190
rect 3180 -1450 3190 -1380
rect 3110 -1460 3180 -1450
rect 3800 -1700 3890 -940
rect 4670 -1040 4680 -880
rect 4860 -880 4930 -870
rect 4600 -1050 4670 -1040
rect 4860 -1050 4930 -1040
rect 6380 -1380 6450 -1370
rect 6380 -1460 6450 -1450
rect 3030 -1730 3100 -1720
rect 3030 -1880 3100 -1870
rect 3200 -1730 3270 -1720
rect 3870 -1770 3890 -1700
rect 3800 -1780 3890 -1770
rect 4290 -1600 4350 -1590
rect 3200 -1880 3270 -1870
rect 3040 -2110 3100 -1880
rect 3210 -2110 3270 -1880
rect 3710 -1790 3780 -1780
rect 3710 -1880 3780 -1870
rect 3880 -1790 3950 -1780
rect 3880 -1880 3950 -1870
rect 3710 -2110 3770 -1880
rect 3890 -2110 3950 -1880
rect 4290 -2110 4350 -1870
rect 5170 -1600 5230 -1590
rect 5700 -1700 5770 -1690
rect 5170 -1950 5230 -1870
rect 5620 -1790 5690 -1730
rect 6300 -1730 6370 -1690
rect 5700 -1780 5770 -1770
rect 5170 -2050 5250 -1950
rect 3040 -2200 4350 -2110
rect 3040 -2420 3100 -2200
rect 3210 -2420 3270 -2200
rect 3040 -2430 3110 -2420
rect 3040 -2580 3110 -2570
rect 3210 -2430 3280 -2420
rect 3210 -2580 3280 -2570
rect 3710 -2430 3770 -2200
rect 3890 -2430 3950 -2200
rect 4290 -2250 4350 -2200
rect 5190 -2080 5250 -2050
rect 5190 -2100 5270 -2080
rect 5620 -2100 5690 -1870
rect 5790 -1790 5860 -1770
rect 5790 -2100 5860 -1870
rect 6300 -2100 6370 -1870
rect 6470 -1730 6540 -1710
rect 6470 -2100 6540 -1870
rect 5190 -2180 6540 -2100
rect 5190 -2220 5270 -2180
rect 4290 -2300 4360 -2250
rect 4300 -2400 4360 -2300
rect 5210 -2400 5270 -2220
rect 4300 -2410 4380 -2400
rect 3710 -2440 3790 -2430
rect 3710 -2580 3720 -2440
rect 3720 -2590 3790 -2580
rect 3890 -2440 3960 -2430
rect 4300 -2520 4320 -2410
rect 3890 -2590 3960 -2580
rect 4320 -2690 4380 -2680
rect 5200 -2410 5270 -2400
rect 5260 -2530 5270 -2410
rect 5620 -2440 5690 -2180
rect 5620 -2590 5690 -2580
rect 5790 -2440 5860 -2180
rect 5790 -2590 5860 -2580
rect 6290 -2440 6360 -2180
rect 6460 -2430 6530 -2180
rect 6460 -2580 6530 -2570
rect 6290 -2590 6360 -2580
rect 5200 -2690 5260 -2680
rect 3120 -3470 3190 -3460
rect 3110 -3540 3120 -3470
rect 3110 -3790 3190 -3540
rect 6370 -3470 6440 -3460
rect 6370 -3550 6440 -3540
rect 2590 -3910 3190 -3790
rect 3810 -4720 3880 -4710
rect 5700 -4720 5770 -4710
rect 3880 -4790 3890 -4720
rect 3810 -4960 3890 -4790
rect 5700 -4800 5770 -4790
rect 2540 -5120 3890 -4960
rect 4620 -5140 4680 -5130
rect 4900 -5140 4960 -5130
rect 4390 -5430 4590 -5420
rect 4390 -5510 4590 -5500
rect 4620 -5600 4680 -5410
rect 4890 -5410 4900 -5370
rect 4890 -5600 4960 -5410
rect 4990 -5430 5180 -5420
rect 4990 -5510 5180 -5500
rect 4620 -5650 4960 -5600
rect 4620 -5670 4920 -5650
rect 4830 -5680 4920 -5670
rect 4830 -5920 4900 -5680
rect 4890 -5930 4900 -5920
rect 4830 -6010 4890 -6000
rect 4740 -6030 4810 -6020
rect 4730 -6100 4740 -6030
rect 4730 -6280 4810 -6100
rect 6860 -6280 6960 -560
rect 4730 -6390 7030 -6280
rect 6860 -6400 6960 -6390
<< via2 >>
rect 2810 -170 2880 -100
rect 4380 340 4560 400
rect 4960 340 5140 400
rect 3510 -170 3580 -100
rect 3600 -270 3660 -190
rect 4590 -280 4650 -110
rect 4650 -280 4660 -110
rect 4590 -290 4660 -280
rect 4860 -290 4930 -110
rect 5820 -280 5830 -190
rect 5830 -280 5900 -190
rect 4380 -380 4560 -320
rect 4960 -380 5140 -320
rect 4550 -650 4670 -540
rect 4860 -650 4980 -540
rect 4370 -840 4570 -780
rect 4950 -840 5150 -780
rect 6380 -1450 6450 -1380
rect 5700 -1770 5770 -1700
rect 6370 -3540 6440 -3470
rect 5700 -4790 5770 -4720
rect 4390 -5500 4400 -5430
rect 4400 -5500 4580 -5430
rect 4990 -5500 5180 -5430
<< metal3 >>
rect 2800 -170 2810 -100
rect 2880 -170 2890 -100
rect 3500 -170 3510 -100
rect 3580 -170 3590 -100
rect 3590 -270 3600 -190
rect 3660 -270 3670 -190
rect 3600 -540 3670 -270
rect 3880 -540 4050 830
rect 4370 340 4380 400
rect 4560 340 4570 400
rect 4950 340 4960 400
rect 5140 340 5150 400
rect 4840 -110 4920 -100
rect 4580 -290 4590 -110
rect 4660 -120 4670 -110
rect 4660 -290 4680 -120
rect 4370 -380 4380 -320
rect 4560 -380 4570 -320
rect 4600 -540 4680 -290
rect 3600 -650 4550 -540
rect 4670 -650 4680 -540
rect 4840 -290 4860 -110
rect 4930 -290 4940 -110
rect 4840 -540 4920 -290
rect 4950 -380 4960 -320
rect 5140 -380 5150 -320
rect 5440 -540 5610 820
rect 5800 -280 5820 -190
rect 5900 -280 5910 -190
rect 5800 -540 5900 -280
rect 4840 -650 4860 -540
rect 4980 -650 5900 -540
rect 4840 -770 4910 -650
rect 4560 -780 4910 -770
rect 4360 -840 4370 -780
rect 4570 -840 4910 -780
rect 4940 -840 4950 -780
rect 5150 -840 5160 -780
rect 4840 -880 4910 -840
rect 4840 -930 4860 -880
rect 4850 -1040 4860 -930
rect 4930 -1040 4940 -880
rect 5700 -910 7100 -830
rect 5700 -1700 5780 -910
rect 6380 -1220 7100 -1130
rect 6380 -1380 6480 -1220
rect 6370 -1450 6380 -1380
rect 6450 -1450 6480 -1380
rect 5690 -1770 5700 -1700
rect 5770 -1770 5780 -1700
rect 5700 -1780 5780 -1770
rect 6360 -3540 6370 -3470
rect 6440 -3540 6450 -3470
rect 6380 -3800 6440 -3540
rect 6380 -3890 7130 -3800
rect 5690 -4790 5700 -4720
rect 5770 -4790 5780 -4720
rect 5710 -5030 5780 -4790
rect 5710 -5130 7110 -5030
rect 4380 -5500 4390 -5430
rect 4580 -5500 4590 -5430
rect 4980 -5500 4990 -5430
rect 5180 -5500 5190 -5430
rect 4390 -6490 4490 -5500
rect 5090 -6490 5190 -5500
<< via3 >>
rect 4860 -1040 4930 -880
<< metal4 >>
rect 4860 -880 4930 -870
rect 4860 -1050 4930 -1040
use pfet_03v3_H5R3BY  XM1
timestamp 1755242987
transform 1 0 2848 0 1 -230
box -278 -250 278 250
use pfet_03v3_H5R3BY  XM2
timestamp 1755242987
transform 1 0 3548 0 1 -230
box -278 -250 278 250
use pfet_03v3_669F58  XM3
timestamp 1755242987
transform 1 0 4470 0 1 10
box -350 -510 2560 570
use pfet_03v3_669F58  XM4
timestamp 1755242987
transform 1 0 5050 0 1 10
box -350 -510 2560 570
use pfet_03v3_H5R3BY  XM5
timestamp 1755242987
transform 1 0 5948 0 1 -230
box -278 -250 278 250
use pfet_03v3_H5R3BY  XM6
timestamp 1755242987
transform -1 0 6758 0 1 -230
box -278 -250 278 250
use nfet_03v3_E4SVYL  XM7
timestamp 1755242987
transform 1 0 4470 0 1 -1370
box -350 -710 350 710
use nfet_03v3_E4SVYL  XM8
timestamp 1755242987
transform 1 0 5050 0 1 -1370
box -350 -710 350 710
use nfet_03v3_2KYBZL  XM9
timestamp 1755242987
transform 1 0 4500 0 1 -3910
box -350 -1710 350 1710
use nfet_03v3_2KYBZL  XM10
timestamp 1755242987
transform 1 0 5080 0 1 -3910
box -350 -1710 350 1710
use nfet_03v3_Z8672T  XM11
timestamp 1755250179
transform -1 0 4772 0 1 -5960
box -298 -300 332 250
use pfet_03v3_H5R3BY  XM12
timestamp 1755242987
transform 1 0 5738 0 1 -1830
box -278 -250 278 250
use pfet_03v3_HDLTJN  XM13
timestamp 1755242987
transform 1 0 6418 0 1 -1674
box -278 -406 278 406
use pfet_03v3_GU2533  XM14
timestamp 1755242987
transform 1 0 6408 0 1 -2942
box -278 -718 278 718
use pfet_03v3_HVKTJN  XM15
timestamp 1755242987
transform 1 0 5738 0 1 -3568
box -278 -1342 278 1342
use pfet_03v3_H5R3BY  XM16
timestamp 1755242987
transform 1 0 3828 0 1 -1830
box -278 -250 278 250
use pfet_03v3_HDLTJN  XM17
timestamp 1755242987
transform 1 0 3148 0 1 -1674
box -278 -406 278 406
use pfet_03v3_GU2533  XM18
timestamp 1755242987
transform -1 0 3158 0 1 -2942
box -278 -718 278 718
use pfet_03v3_HVKTJN  XM19
timestamp 1755242987
transform 1 0 3838 0 1 -3568
box -278 -1342 278 1342
<< labels >>
rlabel metal2 2620 620 2620 620 7 Clk
port 0 w
rlabel metal3 4440 -6490 4440 -6490 5 Vin1
port 1 s
rlabel metal3 5140 -6490 5140 -6490 5 Vin2
port 2 s
rlabel metal1 2610 530 2610 530 1 VDD
port 3 n
rlabel metal3 3960 830 3960 830 1 Vout1
port 5 n
rlabel metal3 5530 820 5530 820 1 Vout2
port 6 n
rlabel metal3 7100 -870 7100 -870 1 off5
port 7 n
rlabel metal3 7100 -1180 7100 -1180 3 off6
port 8 e
rlabel metal3 7130 -3850 7130 -3850 3 off7
port 9 e
rlabel metal3 7110 -5080 7110 -5080 3 off8
port 10 e
rlabel metal2 2400 -860 2400 -860 7 off1
port 11 w
rlabel metal2 2410 -1140 2410 -1140 7 off2
port 12 w
rlabel metal2 2590 -3850 2590 -3850 7 off3
port 13 w
rlabel metal2 2540 -5040 2540 -5040 7 off4
port 14 w
rlabel space 5070 -6200 5070 -6200 3 VSS
rlabel space 5050 -6240 5100 -6180 1 remove
rlabel metal1 3100 -6190 3100 -6190 1 VSS
port 4 n
<< end >>
