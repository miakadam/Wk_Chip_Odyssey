magic
tech gf180mcuD
magscale 1 10
timestamp 1757399739
<< pwell >>
rect -1884 -266 1884 266
<< nmos >>
rect -1772 -150 -1572 150
rect -1468 -150 -1268 150
rect -1164 -150 -964 150
rect -860 -150 -660 150
rect -556 -150 -356 150
rect -252 -150 -52 150
rect 52 -150 252 150
rect 356 -150 556 150
rect 660 -150 860 150
rect 964 -150 1164 150
rect 1268 -150 1468 150
rect 1572 -150 1772 150
<< ndiff >>
rect -1860 137 -1772 150
rect -1860 -137 -1847 137
rect -1801 -137 -1772 137
rect -1860 -150 -1772 -137
rect -1572 137 -1468 150
rect -1572 -137 -1543 137
rect -1497 -137 -1468 137
rect -1572 -150 -1468 -137
rect -1268 137 -1164 150
rect -1268 -137 -1239 137
rect -1193 -137 -1164 137
rect -1268 -150 -1164 -137
rect -964 137 -860 150
rect -964 -137 -935 137
rect -889 -137 -860 137
rect -964 -150 -860 -137
rect -660 137 -556 150
rect -660 -137 -631 137
rect -585 -137 -556 137
rect -660 -150 -556 -137
rect -356 137 -252 150
rect -356 -137 -327 137
rect -281 -137 -252 137
rect -356 -150 -252 -137
rect -52 137 52 150
rect -52 -137 -23 137
rect 23 -137 52 137
rect -52 -150 52 -137
rect 252 137 356 150
rect 252 -137 281 137
rect 327 -137 356 137
rect 252 -150 356 -137
rect 556 137 660 150
rect 556 -137 585 137
rect 631 -137 660 137
rect 556 -150 660 -137
rect 860 137 964 150
rect 860 -137 889 137
rect 935 -137 964 137
rect 860 -150 964 -137
rect 1164 137 1268 150
rect 1164 -137 1193 137
rect 1239 -137 1268 137
rect 1164 -150 1268 -137
rect 1468 137 1572 150
rect 1468 -137 1497 137
rect 1543 -137 1572 137
rect 1468 -150 1572 -137
rect 1772 137 1860 150
rect 1772 -137 1801 137
rect 1847 -137 1860 137
rect 1772 -150 1860 -137
<< ndiffc >>
rect -1847 -137 -1801 137
rect -1543 -137 -1497 137
rect -1239 -137 -1193 137
rect -935 -137 -889 137
rect -631 -137 -585 137
rect -327 -137 -281 137
rect -23 -137 23 137
rect 281 -137 327 137
rect 585 -137 631 137
rect 889 -137 935 137
rect 1193 -137 1239 137
rect 1497 -137 1543 137
rect 1801 -137 1847 137
<< polysilicon >>
rect -1772 229 -1572 242
rect -1772 183 -1759 229
rect -1585 183 -1572 229
rect -1772 150 -1572 183
rect -1468 229 -1268 242
rect -1468 183 -1455 229
rect -1281 183 -1268 229
rect -1468 150 -1268 183
rect -1164 229 -964 242
rect -1164 183 -1151 229
rect -977 183 -964 229
rect -1164 150 -964 183
rect -860 229 -660 242
rect -860 183 -847 229
rect -673 183 -660 229
rect -860 150 -660 183
rect -556 229 -356 242
rect -556 183 -543 229
rect -369 183 -356 229
rect -556 150 -356 183
rect -252 229 -52 242
rect -252 183 -239 229
rect -65 183 -52 229
rect -252 150 -52 183
rect 52 229 252 242
rect 52 183 65 229
rect 239 183 252 229
rect 52 150 252 183
rect 356 229 556 242
rect 356 183 369 229
rect 543 183 556 229
rect 356 150 556 183
rect 660 229 860 242
rect 660 183 673 229
rect 847 183 860 229
rect 660 150 860 183
rect 964 229 1164 242
rect 964 183 977 229
rect 1151 183 1164 229
rect 964 150 1164 183
rect 1268 229 1468 242
rect 1268 183 1281 229
rect 1455 183 1468 229
rect 1268 150 1468 183
rect 1572 229 1772 242
rect 1572 183 1585 229
rect 1759 183 1772 229
rect 1572 150 1772 183
rect -1772 -183 -1572 -150
rect -1772 -229 -1759 -183
rect -1585 -229 -1572 -183
rect -1772 -242 -1572 -229
rect -1468 -183 -1268 -150
rect -1468 -229 -1455 -183
rect -1281 -229 -1268 -183
rect -1468 -242 -1268 -229
rect -1164 -183 -964 -150
rect -1164 -229 -1151 -183
rect -977 -229 -964 -183
rect -1164 -242 -964 -229
rect -860 -183 -660 -150
rect -860 -229 -847 -183
rect -673 -229 -660 -183
rect -860 -242 -660 -229
rect -556 -183 -356 -150
rect -556 -229 -543 -183
rect -369 -229 -356 -183
rect -556 -242 -356 -229
rect -252 -183 -52 -150
rect -252 -229 -239 -183
rect -65 -229 -52 -183
rect -252 -242 -52 -229
rect 52 -183 252 -150
rect 52 -229 65 -183
rect 239 -229 252 -183
rect 52 -242 252 -229
rect 356 -183 556 -150
rect 356 -229 369 -183
rect 543 -229 556 -183
rect 356 -242 556 -229
rect 660 -183 860 -150
rect 660 -229 673 -183
rect 847 -229 860 -183
rect 660 -242 860 -229
rect 964 -183 1164 -150
rect 964 -229 977 -183
rect 1151 -229 1164 -183
rect 964 -242 1164 -229
rect 1268 -183 1468 -150
rect 1268 -229 1281 -183
rect 1455 -229 1468 -183
rect 1268 -242 1468 -229
rect 1572 -183 1772 -150
rect 1572 -229 1585 -183
rect 1759 -229 1772 -183
rect 1572 -242 1772 -229
<< polycontact >>
rect -1759 183 -1585 229
rect -1455 183 -1281 229
rect -1151 183 -977 229
rect -847 183 -673 229
rect -543 183 -369 229
rect -239 183 -65 229
rect 65 183 239 229
rect 369 183 543 229
rect 673 183 847 229
rect 977 183 1151 229
rect 1281 183 1455 229
rect 1585 183 1759 229
rect -1759 -229 -1585 -183
rect -1455 -229 -1281 -183
rect -1151 -229 -977 -183
rect -847 -229 -673 -183
rect -543 -229 -369 -183
rect -239 -229 -65 -183
rect 65 -229 239 -183
rect 369 -229 543 -183
rect 673 -229 847 -183
rect 977 -229 1151 -183
rect 1281 -229 1455 -183
rect 1585 -229 1759 -183
<< metal1 >>
rect -1770 183 -1759 229
rect -1585 183 -1574 229
rect -1466 183 -1455 229
rect -1281 183 -1270 229
rect -1162 183 -1151 229
rect -977 183 -966 229
rect -858 183 -847 229
rect -673 183 -662 229
rect -554 183 -543 229
rect -369 183 -358 229
rect -250 183 -239 229
rect -65 183 -54 229
rect 54 183 65 229
rect 239 183 250 229
rect 358 183 369 229
rect 543 183 554 229
rect 662 183 673 229
rect 847 183 858 229
rect 966 183 977 229
rect 1151 183 1162 229
rect 1270 183 1281 229
rect 1455 183 1466 229
rect 1574 183 1585 229
rect 1759 183 1770 229
rect -1847 137 -1801 148
rect -1847 -148 -1801 -137
rect -1543 137 -1497 148
rect -1543 -148 -1497 -137
rect -1239 137 -1193 148
rect -1239 -148 -1193 -137
rect -935 137 -889 148
rect -935 -148 -889 -137
rect -631 137 -585 148
rect -631 -148 -585 -137
rect -327 137 -281 148
rect -327 -148 -281 -137
rect -23 137 23 148
rect -23 -148 23 -137
rect 281 137 327 148
rect 281 -148 327 -137
rect 585 137 631 148
rect 585 -148 631 -137
rect 889 137 935 148
rect 889 -148 935 -137
rect 1193 137 1239 148
rect 1193 -148 1239 -137
rect 1497 137 1543 148
rect 1497 -148 1543 -137
rect 1801 137 1847 148
rect 1801 -148 1847 -137
rect -1770 -229 -1759 -183
rect -1585 -229 -1574 -183
rect -1466 -229 -1455 -183
rect -1281 -229 -1270 -183
rect -1162 -229 -1151 -183
rect -977 -229 -966 -183
rect -858 -229 -847 -183
rect -673 -229 -662 -183
rect -554 -229 -543 -183
rect -369 -229 -358 -183
rect -250 -229 -239 -183
rect -65 -229 -54 -183
rect 54 -229 65 -183
rect 239 -229 250 -183
rect 358 -229 369 -183
rect 543 -229 554 -183
rect 662 -229 673 -183
rect 847 -229 858 -183
rect 966 -229 977 -183
rect 1151 -229 1162 -183
rect 1270 -229 1281 -183
rect 1455 -229 1466 -183
rect 1574 -229 1585 -183
rect 1759 -229 1770 -183
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.5 l 1 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
