magic
tech gf180mcuD
magscale 1 10
timestamp 1757925408
<< pwell >>
rect 1627 -371 1644 -368
rect 1746 -371 1842 -358
rect 1888 -369 1923 -357
rect 2226 -371 2323 -358
<< metal1 >>
rect 1290 880 2778 1080
rect 1542 749 1638 780
rect 1807 668 2261 880
rect 2430 749 2526 780
rect 1448 373 1528 383
rect 1448 133 1460 373
rect 1516 133 1528 373
rect 1448 123 1528 133
rect 1715 72 2353 668
rect 2540 373 2620 383
rect 2540 133 2552 373
rect 2608 133 2620 373
rect 2540 123 2620 133
rect 1542 -84 1638 -9
rect 1542 -140 1562 -84
rect 1618 -140 1638 -84
rect 1542 -358 1638 -140
rect 2430 -228 2526 -9
rect 2362 -240 2526 -228
rect 2362 -296 2374 -240
rect 2430 -296 2526 -240
rect 2362 -308 2526 -296
rect 2430 -358 2526 -308
rect 1542 -371 1842 -358
rect 2226 -371 2526 -358
rect 1638 -404 1746 -371
rect 2322 -404 2452 -371
rect 1363 -648 1505 -452
rect 1652 -522 1732 -512
rect 1652 -578 1664 -522
rect 1720 -578 1732 -522
rect 1652 -588 1732 -578
rect 1873 -648 2015 -452
rect 2132 -522 2212 -512
rect 2132 -578 2144 -522
rect 2200 -578 2212 -522
rect 2132 -588 2212 -578
rect 2336 -522 2416 -512
rect 2336 -578 2348 -522
rect 2404 -578 2416 -522
rect 2336 -588 2416 -578
rect 2540 -522 2620 -512
rect 2540 -578 2552 -522
rect 2608 -578 2620 -522
rect 2540 -588 2620 -578
rect 1327 -860 1373 -731
rect 1542 -760 1638 -729
rect 1746 -760 1842 -729
rect 2011 -860 2057 -731
rect 2226 -760 2322 -729
rect 2430 -760 2526 -729
rect 2695 -860 2741 -720
rect 1290 -1060 2778 -860
<< via1 >>
rect 1460 133 1516 373
rect 2552 133 2608 373
rect 1562 -140 1618 -84
rect 2374 -296 2430 -240
rect 1664 -578 1720 -522
rect 2144 -578 2200 -522
rect 2348 -578 2404 -522
rect 2552 -578 2608 -522
<< metal2 >>
rect 1448 373 2620 383
rect 1448 133 1460 373
rect 1516 133 2552 373
rect 2608 133 2620 373
rect 1448 123 2620 133
rect 1542 -84 1620 -72
rect 1203 -140 1562 -84
rect 1618 -140 1620 -84
rect 1542 -152 1620 -140
rect 2540 -162 2620 123
rect 2540 -218 2778 -162
rect 2362 -240 2432 -228
rect 1203 -296 2374 -240
rect 2430 -296 2432 -240
rect 2362 -308 2432 -296
rect 1652 -522 1732 -512
rect 1652 -578 1664 -522
rect 1720 -578 1732 -522
rect 1652 -764 1732 -578
rect 2132 -522 2212 -512
rect 2132 -578 2144 -522
rect 2200 -578 2212 -522
rect 2132 -588 2212 -578
rect 2336 -522 2416 -512
rect 2336 -578 2348 -522
rect 2404 -578 2416 -522
rect 2336 -764 2416 -578
rect 2540 -522 2620 -218
rect 2540 -578 2552 -522
rect 2608 -578 2620 -522
rect 2540 -588 2620 -578
rect 1652 -836 2416 -764
<< via2 >>
rect 2144 -578 2200 -522
rect 2552 -578 2608 -522
<< metal3 >>
rect 2132 -522 2620 -512
rect 2132 -578 2144 -522
rect 2200 -578 2552 -522
rect 2608 -578 2620 -522
rect 2132 -588 2620 -578
use nfet_03v3_EMCFTP  nfet_03v3_EMCFTP_0
timestamp 1757924681
transform 1 0 2376 0 1 -550
box -402 -310 402 310
use pfet_03v3_LJVJK4  pfet_03v3_LJVJK4_0
timestamp 1757924681
transform 1 0 2478 0 1 370
box -300 -510 300 510
use nfet_03v3_EMCFTP  XM1
timestamp 1757924681
transform 1 0 1692 0 1 -550
box -402 -310 402 310
use pfet_03v3_LJVJK4  XM2
timestamp 1757924681
transform 1 0 1590 0 1 370
box -300 -510 300 510
<< labels >>
rlabel metal1 2026 1080 2026 1080 1 VDD
port 0 n
rlabel metal2 2778 -190 2778 -190 3 OUT
port 1 e
rlabel metal2 1203 -271 1203 -271 7 A
port 2 w
rlabel metal2 1203 -113 1203 -113 7 B
port 3 w
rlabel metal1 2035 -1060 2035 -1060 5 VSS
port 4 s
<< end >>
