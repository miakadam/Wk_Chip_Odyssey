magic
tech gf180mcuD
magscale 1 10
timestamp 1757820791
<< metal1 >>
rect -58 7732 12 7744
rect 4010 7732 4096 7744
rect -58 7676 -46 7732
rect 10 7676 20 7732
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect -58 7664 12 7676
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 3222 5355 4022 5411
rect 7222 5355 8034 5411
rect 11276 5355 12076 5411
rect 15318 5355 16118 5411
rect 19360 5355 20160 5411
rect 23402 5355 24202 5411
rect 3966 5233 4022 5355
rect 7978 5233 8034 5355
rect 12020 5233 12076 5355
rect 16062 5233 16118 5355
rect 20104 5233 20160 5355
rect 24146 5233 24202 5355
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect -330 4509 -260 4521
rect 3682 4509 3752 4521
rect 7694 4509 7764 4521
rect 11736 4509 11806 4521
rect 15778 4509 15848 4521
rect 19820 4509 19890 4521
rect 23862 4509 23932 4521
rect -330 4453 -318 4509
rect -262 4453 418 4509
rect 3682 4453 3694 4509
rect 3750 4453 4032 4509
rect 7694 4453 7706 4509
rect 7762 4453 8080 4509
rect 11736 4453 11748 4509
rect 11804 4453 12107 4509
rect 15778 4453 15790 4509
rect 15846 4453 16149 4509
rect 19820 4453 19832 4509
rect 19888 4453 20191 4509
rect 23862 4453 23874 4509
rect 23930 4453 24236 4509
rect -330 4441 -260 4453
rect 3682 4441 3752 4453
rect 7694 4441 7764 4453
rect 11736 4441 11806 4453
rect 15778 4441 15848 4453
rect 19820 4441 19890 4453
rect 23862 4441 23932 4453
rect -121 885 -41 897
rect 3954 885 4024 897
rect 7966 885 8046 897
rect 12008 885 12088 897
rect 16050 885 16130 897
rect 20092 885 20172 897
rect 24134 885 24214 897
rect -121 829 -109 885
rect -53 829 90 885
rect 3954 829 3966 885
rect 4022 829 4032 885
rect 7966 829 7978 885
rect 8034 829 8081 885
rect 12008 829 12020 885
rect 12076 829 12111 885
rect 16050 829 16062 885
rect 16118 829 16149 885
rect 20092 829 20104 885
rect 20160 829 20191 885
rect 24134 829 24146 885
rect 24202 829 24239 885
rect -121 817 -41 829
rect 3954 817 4024 829
rect 7966 817 8046 829
rect 12008 817 12088 829
rect 16050 817 16130 829
rect 20092 817 20172 829
rect 24134 817 24214 829
rect -121 98 -35 110
rect 3818 98 3888 110
rect 7830 98 7900 110
rect 11872 98 11942 110
rect 15914 98 15984 110
rect 19956 98 20026 110
rect 23998 98 24068 110
rect -121 42 -109 98
rect -53 42 27 98
rect 3818 42 3830 98
rect 3886 42 4039 98
rect 7830 42 7842 98
rect 7898 42 8081 98
rect 11872 42 11884 98
rect 11940 42 12123 98
rect 15914 42 15926 98
rect 15982 42 16165 98
rect 19956 42 19968 98
rect 20024 42 20207 98
rect 23998 42 24010 98
rect 24066 42 24249 98
rect -121 30 -35 42
rect 3818 30 3888 42
rect 7830 30 7900 42
rect 11872 30 11942 42
rect 15914 30 15984 42
rect 19956 30 20026 42
rect 23998 30 24068 42
<< via1 >>
rect -46 7676 10 7732
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect 3966 5167 4022 5223
rect 7978 5167 8034 5223
rect 12020 5167 12076 5223
rect 16062 5167 16118 5223
rect 20104 5167 20160 5223
rect 24146 5167 24202 5223
rect -318 4453 -262 4509
rect 3694 4453 3750 4509
rect 7706 4453 7762 4509
rect 11748 4453 11804 4509
rect 15790 4453 15846 4509
rect 19832 4453 19888 4509
rect 23874 4453 23930 4509
rect -109 829 -53 885
rect 3966 829 4022 885
rect 7978 829 8034 885
rect 12020 829 12076 885
rect 16062 829 16118 885
rect 20104 829 20160 885
rect 24146 829 24202 885
rect -109 42 -53 98
rect 3830 42 3886 98
rect 7842 42 7898 98
rect 11884 42 11940 98
rect 15926 42 15982 98
rect 19968 42 20024 98
rect 24010 42 24066 98
<< metal2 >>
rect -201 9004 10 9014
rect -201 8904 -46 9004
rect -46 7744 10 8904
rect -58 7732 12 7744
rect -58 7676 -46 7732
rect 10 7676 12 7732
rect -58 7664 12 7676
rect -330 4509 -260 4521
rect -330 4453 -318 4509
rect -262 4453 -260 4509
rect -330 4441 -260 4453
rect -318 -245 -262 4441
rect 3558 3207 3614 9863
rect 3830 9007 3886 9017
rect 3682 4509 3752 4521
rect 3682 4453 3694 4509
rect 3750 4453 3752 4509
rect 3682 4441 3752 4453
rect 3478 3151 3614 3207
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
rect 3694 -233 3750 4441
rect 3830 110 3886 8907
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 3954 5223 4034 5233
rect 3954 5167 3966 5223
rect 4022 5167 4034 5223
rect 3954 5165 4034 5167
rect 3966 897 4022 5165
rect 7570 3207 7626 9863
rect 7842 9004 7898 9014
rect 7694 4509 7764 4521
rect 7694 4453 7706 4509
rect 7762 4453 7764 4509
rect 7694 4441 7764 4453
rect 7490 3151 7626 3207
rect 3954 885 4024 897
rect 3954 829 3966 885
rect 4022 829 4024 885
rect 3954 817 4024 829
rect 3818 98 3888 110
rect 3818 42 3830 98
rect 3886 42 3888 98
rect 3818 30 3888 42
rect 7706 -233 7762 4441
rect 7842 110 7898 8904
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 7966 5223 8046 5233
rect 7966 5167 7978 5223
rect 8034 5167 8046 5223
rect 7966 5165 8046 5167
rect 7978 897 8034 5165
rect 11612 3207 11668 9863
rect 11884 9004 11940 9014
rect 11736 4509 11806 4521
rect 11736 4453 11748 4509
rect 11804 4453 11806 4509
rect 11736 4441 11806 4453
rect 11532 3151 11668 3207
rect 7966 885 8046 897
rect 7966 829 7978 885
rect 8034 829 8046 885
rect 7966 817 8046 829
rect 7830 98 7900 110
rect 7830 42 7842 98
rect 7898 42 7900 98
rect 7830 30 7900 42
rect 11748 -233 11804 4441
rect 11884 110 11940 8904
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 12008 5223 12088 5233
rect 12008 5167 12020 5223
rect 12076 5167 12088 5223
rect 12008 5165 12088 5167
rect 12020 897 12076 5165
rect 15654 3207 15710 9863
rect 15926 9004 15982 9014
rect 15778 4509 15848 4521
rect 15778 4453 15790 4509
rect 15846 4453 15848 4509
rect 15778 4441 15848 4453
rect 15574 3151 15710 3207
rect 12008 885 12088 897
rect 12008 829 12020 885
rect 12076 829 12088 885
rect 12008 817 12088 829
rect 11872 98 11942 110
rect 11872 42 11884 98
rect 11940 42 11942 98
rect 11872 30 11942 42
rect 15790 -233 15846 4441
rect 15926 110 15982 8904
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 16050 5223 16130 5233
rect 16050 5167 16062 5223
rect 16118 5167 16130 5223
rect 16050 5165 16130 5167
rect 16062 897 16118 5165
rect 19696 3207 19752 9863
rect 19968 9004 20024 9014
rect 19820 4509 19890 4521
rect 19820 4453 19832 4509
rect 19888 4453 19890 4509
rect 19820 4441 19890 4453
rect 19616 3151 19752 3207
rect 16050 885 16130 897
rect 16050 829 16062 885
rect 16118 829 16130 885
rect 16050 817 16130 829
rect 15914 98 15984 110
rect 15914 42 15926 98
rect 15982 42 15984 98
rect 15914 30 15984 42
rect 19832 -233 19888 4441
rect 19968 110 20024 8904
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 20092 5223 20172 5233
rect 20092 5167 20104 5223
rect 20160 5167 20172 5223
rect 20092 5165 20172 5167
rect 20104 897 20160 5165
rect 23738 3207 23794 9863
rect 24010 9004 24066 9014
rect 23862 4509 23932 4521
rect 23862 4453 23874 4509
rect 23930 4453 23932 4509
rect 23862 4441 23932 4453
rect 23658 3151 23794 3207
rect 20092 885 20172 897
rect 20092 829 20104 885
rect 20160 829 20172 885
rect 20092 817 20172 829
rect 19956 98 20026 110
rect 19956 42 19968 98
rect 20024 42 20026 98
rect 19956 30 20026 42
rect 23874 -233 23930 4441
rect 24010 110 24066 8904
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect 24134 5223 24214 5233
rect 24134 5167 24146 5223
rect 24202 5167 24214 5223
rect 24134 5165 24214 5167
rect 24146 897 24202 5165
rect 24134 885 24214 897
rect 24134 829 24146 885
rect 24202 829 24214 885
rect 24134 817 24214 829
rect 23998 98 24068 110
rect 23998 42 24010 98
rect 24066 42 24068 98
rect 23998 30 24068 42
<< via2 >>
rect -46 8904 10 9004
rect 3830 8907 3886 9007
rect -109 829 -53 885
rect -109 42 -53 98
rect 4022 7676 4078 7732
rect 7842 8904 7898 9004
rect 8064 7676 8120 7732
rect 11884 8904 11940 9004
rect 12106 7676 12162 7732
rect 15926 8904 15982 9004
rect 16148 7676 16204 7732
rect 19968 8904 20024 9004
rect 20190 7676 20246 7732
rect 24010 8904 24066 9004
rect 24232 7676 24288 7732
<< metal3 >>
rect 3820 9004 3830 9007
rect -56 8904 -46 9004
rect 10 8907 3830 9004
rect 3886 9004 3896 9007
rect 3886 8907 7842 9004
rect 10 8904 7842 8907
rect 7898 8904 11884 9004
rect 11940 8904 15926 9004
rect 15982 8904 19968 9004
rect 20024 8904 24010 9004
rect 24066 8904 24076 9004
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect -121 885 -41 897
rect -121 829 -109 885
rect -53 829 -41 885
rect -121 817 -41 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
<< via3 >>
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect -109 829 -53 885
rect -109 42 -53 98
<< metal4 >>
rect 4010 7732 4096 7744
rect 4010 7676 4022 7732
rect 4078 7676 4096 7732
rect 4010 7664 4096 7676
rect 8052 7732 8138 7744
rect 8052 7676 8064 7732
rect 8120 7676 8138 7732
rect 8052 7664 8138 7676
rect 12094 7732 12180 7744
rect 12094 7676 12106 7732
rect 12162 7676 12180 7732
rect 12094 7664 12180 7676
rect 16136 7732 16222 7744
rect 16136 7676 16148 7732
rect 16204 7676 16222 7732
rect 16136 7664 16222 7676
rect 20178 7732 20264 7744
rect 20178 7676 20190 7732
rect 20246 7676 20264 7732
rect 20178 7664 20264 7676
rect 24220 7732 24306 7744
rect 24220 7676 24232 7732
rect 24288 7676 24306 7732
rect 24220 7664 24306 7676
rect -121 885 156 897
rect -121 829 -109 885
rect -53 829 156 885
rect -121 737 156 829
rect -121 98 -35 110
rect -121 42 -109 98
rect -53 42 -35 98
rect -121 30 -35 42
<< via4 >>
rect 4022 7676 4078 7732
rect 8064 7676 8120 7732
rect 12106 7676 12162 7732
rect 16148 7676 16204 7732
rect 20190 7676 20246 7732
rect 24232 7676 24288 7732
rect -109 42 -53 98
<< metal5 >>
rect 4010 7732 4167 7744
rect 4010 7676 4022 7732
rect 4078 7676 4167 7732
rect 4010 7664 4167 7676
rect 8052 7732 8209 7744
rect 8052 7676 8064 7732
rect 8120 7676 8209 7732
rect 8052 7664 8209 7676
rect 12094 7732 12251 7744
rect 12094 7676 12106 7732
rect 12162 7676 12251 7732
rect 12094 7664 12251 7676
rect 16136 7732 16293 7744
rect 16136 7676 16148 7732
rect 16204 7676 16293 7732
rect 16136 7664 16293 7676
rect 20178 7732 20350 7744
rect 20178 7676 20190 7732
rect 20246 7676 20350 7732
rect 20178 7664 20350 7676
rect 24220 7732 24381 7744
rect 24220 7676 24232 7732
rect 24288 7676 24381 7732
rect 24220 7664 24381 7676
rect -121 98 167 190
rect -121 42 -109 98
rect -53 42 167 98
rect -121 30 167 42
use dffrs  dffrs_0 comparator/final_magic/dffrs
timestamp 1757808491
transform 1 0 858 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_1
timestamp 1757808491
transform 1 0 4870 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_2
timestamp 1757808491
transform 1 0 8912 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_3
timestamp 1757808491
transform 1 0 12954 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_4
timestamp 1757808491
transform 1 0 16996 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_5
timestamp 1757808491
transform 1 0 21038 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_6
timestamp 1757808491
transform 1 0 25080 0 1 5928
box -848 -5898 2620 2881
use dffrs  dffrs_7
timestamp 1757808491
transform 1 0 4870 0 1 15507
box -848 -5898 2620 2881
use dffrs  dffrs_8
timestamp 1757808491
transform 1 0 11992 0 1 20024
box -848 -5898 2620 2881
use dffrs  dffrs_9
timestamp 1757808491
transform 1 0 18885 0 1 20203
box -848 -5898 2620 2881
use dffrs  dffrs_10
timestamp 1757808491
transform 1 0 25447 0 1 20254
box -848 -5898 2620 2881
use dffrs  dffrs_11
timestamp 1757808491
transform 1 0 32774 0 1 20203
box -848 -5898 2620 2881
use dffrs  dffrs_12
timestamp 1757808491
transform 1 0 40765 0 1 20178
box -848 -5898 2620 2881
use dffrs  dffrs_13
timestamp 1757808491
transform 1 0 49496 0 1 20178
box -848 -5898 2620 2881
<< end >>
