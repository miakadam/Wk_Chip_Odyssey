** sch_path: /foss/designs/comparator/final_magic/or2/osu_sc_or2_1.sch
.subckt osu_sc_or2_1 B A Y VDD VSS
*.PININFO B:I A:I Y:O VDD:I VSS:I
XM1 net1 B VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM2 net2 A net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM3 net2 B VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM4 net2 A VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
XM5 Y net2 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
XM6 Y net2 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends
.GLOBAL VDD
.GLOBAL VSS
