magic
tech gf180mcuD
magscale 1 10
timestamp 1755276579
<< pwell >>
rect -2236 -1358 2236 1358
<< psubdiff >>
rect -2212 1262 2212 1334
rect -2212 1218 -2140 1262
rect -2212 -1218 -2199 1218
rect -2153 -1218 -2140 1218
rect 2140 1218 2212 1262
rect -2212 -1262 -2140 -1218
rect 2140 -1218 2153 1218
rect 2199 -1218 2212 1218
rect 2140 -1262 2212 -1218
rect -2212 -1334 2212 -1262
<< psubdiffcont >>
rect -2199 -1218 -2153 1218
rect 2153 -1218 2199 1218
<< polysilicon >>
rect -2000 1109 2000 1122
rect -2000 1063 -1987 1109
rect 1987 1063 2000 1109
rect -2000 1000 2000 1063
rect -2000 -1063 2000 -1000
rect -2000 -1109 -1987 -1063
rect 1987 -1109 2000 -1063
rect -2000 -1122 2000 -1109
<< polycontact >>
rect -1987 1063 1987 1109
rect -1987 -1109 1987 -1063
<< nhighres >>
rect -2000 -1000 2000 1000
<< metal1 >>
rect -2199 1275 2199 1321
rect -2199 1218 -2153 1275
rect 2153 1218 2199 1275
rect -1998 1063 -1987 1109
rect 1987 1063 1998 1109
rect -1998 -1109 -1987 -1063
rect 1987 -1109 1998 -1063
rect -2199 -1275 -2153 -1218
rect 2153 -1275 2199 -1218
rect -2199 -1321 2199 -1275
<< properties >>
string FIXED_BBOX -2176 -1298 2176 1298
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 20.0 l 10.0 m 1 nx 1 wmin 1.000 lmin 1.000 class resistor rho 1000 val 500.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
