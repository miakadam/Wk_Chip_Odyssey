magic
tech gf180mcuD
magscale 1 10
timestamp 1757505342
<< error_p >>
rect -314 113 -303 159
rect -130 113 -119 159
rect 54 113 65 159
rect 238 113 249 159
rect -314 -159 -303 -113
rect -130 -159 -119 -113
rect 54 -159 65 -113
rect 238 -159 249 -113
<< nwell >>
rect -566 -290 566 290
<< pmos >>
rect -316 -80 -236 80
rect -132 -80 -52 80
rect 52 -80 132 80
rect 236 -80 316 80
<< pdiff >>
rect -404 67 -316 80
rect -404 -67 -391 67
rect -345 -67 -316 67
rect -404 -80 -316 -67
rect -236 67 -132 80
rect -236 -67 -207 67
rect -161 -67 -132 67
rect -236 -80 -132 -67
rect -52 67 52 80
rect -52 -67 -23 67
rect 23 -67 52 67
rect -52 -80 52 -67
rect 132 67 236 80
rect 132 -67 161 67
rect 207 -67 236 67
rect 132 -80 236 -67
rect 316 67 404 80
rect 316 -67 345 67
rect 391 -67 404 67
rect 316 -80 404 -67
<< pdiffc >>
rect -391 -67 -345 67
rect -207 -67 -161 67
rect -23 -67 23 67
rect 161 -67 207 67
rect 345 -67 391 67
<< nsubdiff >>
rect -542 194 542 266
rect -542 -194 -470 194
rect 470 150 542 194
rect 470 -150 483 150
rect 529 -150 542 150
rect 470 -194 542 -150
rect -542 -266 542 -194
<< nsubdiffcont >>
rect 483 -150 529 150
<< polysilicon >>
rect -316 159 -236 172
rect -316 113 -303 159
rect -249 113 -236 159
rect -316 80 -236 113
rect -132 159 -52 172
rect -132 113 -119 159
rect -65 113 -52 159
rect -132 80 -52 113
rect 52 159 132 172
rect 52 113 65 159
rect 119 113 132 159
rect 52 80 132 113
rect 236 159 316 172
rect 236 113 249 159
rect 303 113 316 159
rect 236 80 316 113
rect -316 -113 -236 -80
rect -316 -159 -303 -113
rect -249 -159 -236 -113
rect -316 -172 -236 -159
rect -132 -113 -52 -80
rect -132 -159 -119 -113
rect -65 -159 -52 -113
rect -132 -172 -52 -159
rect 52 -113 132 -80
rect 52 -159 65 -113
rect 119 -159 132 -113
rect 52 -172 132 -159
rect 236 -113 316 -80
rect 236 -159 249 -113
rect 303 -159 316 -113
rect 236 -172 316 -159
<< polycontact >>
rect -303 113 -249 159
rect -119 113 -65 159
rect 65 113 119 159
rect 249 113 303 159
rect -303 -159 -249 -113
rect -119 -159 -65 -113
rect 65 -159 119 -113
rect 249 -159 303 -113
<< metal1 >>
rect -314 113 -303 159
rect -249 113 -238 159
rect -130 113 -119 159
rect -65 113 -54 159
rect 54 113 65 159
rect 119 113 130 159
rect 238 113 249 159
rect 303 113 314 159
rect 483 150 529 161
rect -391 67 -345 78
rect -391 -78 -345 -67
rect -207 67 -161 78
rect -207 -78 -161 -67
rect -23 67 23 78
rect -23 -78 23 -67
rect 161 67 207 78
rect 161 -78 207 -67
rect 345 67 391 78
rect 345 -78 391 -67
rect -314 -159 -303 -113
rect -249 -159 -238 -113
rect -130 -159 -119 -113
rect -65 -159 -54 -113
rect 54 -159 65 -113
rect 119 -159 130 -113
rect 238 -159 249 -113
rect 303 -159 314 -113
rect 483 -161 529 -150
<< properties >>
string FIXED_BBOX -506 -230 506 230
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.8 l 0.4 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
