magic
tech gf180mcuD
magscale 1 10
timestamp 1758001983
<< error_p >>
rect -48 133 -37 179
rect -48 -179 -37 -133
<< pwell >>
rect -300 -310 300 310
<< nmos >>
rect -50 -100 50 100
<< ndiff >>
rect -138 87 -50 100
rect -138 -87 -125 87
rect -79 -87 -50 87
rect -138 -100 -50 -87
rect 50 87 138 100
rect 50 -87 79 87
rect 125 -87 138 87
rect 50 -100 138 -87
<< ndiffc >>
rect -125 -87 -79 87
rect 79 -87 125 87
<< psubdiff >>
rect -276 214 276 286
rect -276 170 -204 214
rect -276 -170 -263 170
rect -217 -170 -204 170
rect 204 170 276 214
rect -276 -214 -204 -170
rect 204 -170 217 170
rect 263 -170 276 170
rect 204 -214 276 -170
rect -276 -286 276 -214
<< psubdiffcont >>
rect -263 -170 -217 170
rect 217 -170 263 170
<< polysilicon >>
rect -50 179 50 192
rect -50 133 -37 179
rect 37 133 50 179
rect -50 100 50 133
rect -50 -133 50 -100
rect -50 -179 -37 -133
rect 37 -179 50 -133
rect -50 -192 50 -179
<< polycontact >>
rect -37 133 37 179
rect -37 -179 37 -133
<< metal1 >>
rect -263 170 -217 181
rect -48 133 -37 179
rect 37 133 48 179
rect 217 170 263 181
rect -125 87 -79 98
rect -125 -98 -79 -87
rect 79 87 125 98
rect 79 -98 125 -87
rect -263 -181 -217 -170
rect -48 -179 -37 -133
rect 37 -179 48 -133
rect 217 -181 263 -170
<< properties >>
string FIXED_BBOX -240 -250 240 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
