magic
tech gf180mcuD
magscale 1 10
timestamp 1757373041
<< metal1 >>
rect 2547 565 2593 577
rect 2547 519 2642 565
rect 2547 465 2593 519
rect 2570 -56 2711 74
rect 2775 -783 2824 -403
rect 2896 -930 2953 -293
rect 2553 -1090 2719 -958
rect 2537 -1310 2593 -1143
rect 2537 -1360 2677 -1310
rect 2547 -1361 2677 -1360
use nfet_03v3_86US5R  XM3
timestamp 1757365333
transform 1 0 2804 0 1 -1001
box -290 -386 290 386
use pfet_03v3_YPRA8C  XM4
timestamp 1757365333
transform 1 0 2800 0 1 16
box -290 -586 290 586
<< labels >>
rlabel space 2549 10 2549 10 7 avdd
port 0 w
rlabel metal1 2554 -1018 2554 -1018 7 avss
port 1 w
rlabel metal1 2776 -631 2777 -610 1 in
port 2 n
rlabel metal1 2941 -617 2942 -596 1 out
port 3 n
<< end >>
