magic
tech gf180mcuD
magscale 1 10
timestamp 1757649695
<< error_p >>
rect -222 283 -211 329
rect -38 283 -27 329
rect 146 283 157 329
rect -222 -329 -211 -283
rect -38 -329 -27 -283
rect 146 -329 157 -283
<< nwell >>
rect -474 -460 474 460
<< pmos >>
rect -224 -250 -144 250
rect -40 -250 40 250
rect 144 -250 224 250
<< pdiff >>
rect -312 237 -224 250
rect -312 -237 -299 237
rect -253 -237 -224 237
rect -312 -250 -224 -237
rect -144 237 -40 250
rect -144 -237 -115 237
rect -69 -237 -40 237
rect -144 -250 -40 -237
rect 40 237 144 250
rect 40 -237 69 237
rect 115 -237 144 237
rect 40 -250 144 -237
rect 224 237 312 250
rect 224 -237 253 237
rect 299 -237 312 237
rect 224 -250 312 -237
<< pdiffc >>
rect -299 -237 -253 237
rect -115 -237 -69 237
rect 69 -237 115 237
rect 253 -237 299 237
<< nsubdiff >>
rect -450 364 450 436
rect -450 320 -378 364
rect -450 -320 -437 320
rect -391 -320 -378 320
rect 378 320 450 364
rect -450 -364 -378 -320
rect 378 -320 391 320
rect 437 -320 450 320
rect 378 -364 450 -320
rect -450 -436 450 -364
<< nsubdiffcont >>
rect -437 -320 -391 320
rect 391 -320 437 320
<< polysilicon >>
rect -224 329 -144 342
rect -224 283 -211 329
rect -157 283 -144 329
rect -224 250 -144 283
rect -40 329 40 342
rect -40 283 -27 329
rect 27 283 40 329
rect -40 250 40 283
rect 144 329 224 342
rect 144 283 157 329
rect 211 283 224 329
rect 144 250 224 283
rect -224 -283 -144 -250
rect -224 -329 -211 -283
rect -157 -329 -144 -283
rect -224 -342 -144 -329
rect -40 -283 40 -250
rect -40 -329 -27 -283
rect 27 -329 40 -283
rect -40 -342 40 -329
rect 144 -283 224 -250
rect 144 -329 157 -283
rect 211 -329 224 -283
rect 144 -342 224 -329
<< polycontact >>
rect -211 283 -157 329
rect -27 283 27 329
rect 157 283 211 329
rect -211 -329 -157 -283
rect -27 -329 27 -283
rect 157 -329 211 -283
<< metal1 >>
rect -437 320 -391 331
rect -222 283 -211 329
rect -157 283 -146 329
rect -38 283 -27 329
rect 27 283 38 329
rect 146 283 157 329
rect 211 283 222 329
rect 391 320 437 331
rect -299 237 -253 248
rect -299 -248 -253 -237
rect -115 237 -69 248
rect -115 -248 -69 -237
rect 69 237 115 248
rect 69 -248 115 -237
rect 253 237 299 248
rect 253 -248 299 -237
rect -437 -331 -391 -320
rect -222 -329 -211 -283
rect -157 -329 -146 -283
rect -38 -329 -27 -283
rect 27 -329 38 -283
rect 146 -329 157 -283
rect 211 -329 222 -283
rect 391 -331 437 -320
<< properties >>
string FIXED_BBOX -414 -400 414 400
string gencell pfet_03v3
string library gf180mcu
string parameters w 2.5 l 0.4 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
