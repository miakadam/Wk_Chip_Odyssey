magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 73 -23 119
rect 23 73 34 84
rect -105 -38 -59 38
rect 59 -38 105 38
rect -34 -119 -23 -73
<< nwell >>
rect -204 -218 204 218
<< pmos >>
rect -30 -40 30 40
<< pdiff >>
rect -118 27 -30 40
rect -118 -27 -105 27
rect -59 -27 -30 27
rect -118 -40 -30 -27
rect 30 27 118 40
rect 30 -27 59 27
rect 105 -27 118 27
rect 30 -40 118 -27
<< pdiffc >>
rect -105 -27 -59 27
rect 59 -27 105 27
<< polysilicon >>
rect -36 119 36 132
rect -36 73 -23 119
rect 23 73 36 119
rect -36 60 36 73
rect -30 40 30 60
rect -30 -60 30 -40
rect -36 -73 36 -60
rect -36 -119 -23 -73
rect 23 -119 36 -73
rect -36 -132 36 -119
<< polycontact >>
rect -23 73 23 119
rect -23 -119 23 -73
<< metal1 >>
rect -34 73 -23 119
rect 23 73 34 119
rect -105 27 -59 38
rect -105 -38 -59 -27
rect 59 27 105 38
rect 59 -38 105 -27
rect -34 -119 -23 -73
rect 23 -119 34 -73
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.4 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
