* NGSPICE file created from inv2.ext - technology: (null)

.subckt inv2 in vdd out vss
X0 out.t1 in.t0 vdd.t1 vdd.t0 pfet_03v3
**devattr s=52800,1376 d=52800,1376
X1 out.t0 in.t1 vss.t1 vss.t0 nfet_03v3
**devattr s=17600,576 d=17600,576
R0 in.n0 in.t0 34.1797
R1 in.n0 in.t1 19.5798
R2 in in.n0 4.87271
R3 vdd.n0 vdd.t0 118.543
R4 vdd.n0 vdd.t1 1.79661
R5 vdd vdd.n0 0.336853
R6 out.n0 out.t0 9.6935
R7 out.n0 out.t1 4.35383
R8 out out.n0 0.254429
R9 vss.n0 vss.t0 425.248
R10 vss.n0 vss.t1 5.06763
R11 vss vss.n0 0.288334
.ends

