magic
tech gf180mcuD
magscale 1 10
timestamp 1757365333
<< error_p >>
rect -38 233 -27 279
rect -38 -279 -27 -233
<< pwell >>
rect -290 -410 290 410
<< nmos >>
rect -40 -200 40 200
<< ndiff >>
rect -128 187 -40 200
rect -128 -187 -115 187
rect -69 -187 -40 187
rect -128 -200 -40 -187
rect 40 187 128 200
rect 40 -187 69 187
rect 115 -187 128 187
rect 40 -200 128 -187
<< ndiffc >>
rect -115 -187 -69 187
rect 69 -187 115 187
<< psubdiff >>
rect -266 314 266 386
rect -266 270 -194 314
rect -266 -270 -253 270
rect -207 -270 -194 270
rect 194 270 266 314
rect -266 -314 -194 -270
rect 194 -270 207 270
rect 253 -270 266 270
rect 194 -314 266 -270
rect -266 -386 266 -314
<< psubdiffcont >>
rect -253 -270 -207 270
rect 207 -270 253 270
<< polysilicon >>
rect -40 279 40 292
rect -40 233 -27 279
rect 27 233 40 279
rect -40 200 40 233
rect -40 -233 40 -200
rect -40 -279 -27 -233
rect 27 -279 40 -233
rect -40 -292 40 -279
<< polycontact >>
rect -27 233 27 279
rect -27 -279 27 -233
<< metal1 >>
rect -253 327 253 373
rect -253 270 -207 327
rect -38 233 -27 279
rect 27 233 38 279
rect 207 270 253 327
rect -115 187 -69 198
rect -115 -198 -69 -187
rect 69 187 115 198
rect 69 -198 115 -187
rect -253 -327 -207 -270
rect -38 -279 -27 -233
rect 27 -279 38 -233
rect 207 -327 253 -270
rect -253 -373 253 -327
<< properties >>
string FIXED_BBOX -230 -350 230 350
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.0 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
