magic
tech gf180mcuD
magscale 1 10
timestamp 1756957756
<< error_s >>
rect 16432 2139 16520 2152
rect 16432 2085 16507 2139
rect 16432 2072 16520 2085
rect 11666 1962 11706 1984
rect 7382 1821 7393 1867
rect 8039 1841 8050 1887
rect 7439 1821 7450 1832
rect 11394 1807 11405 1853
rect 11451 1807 11462 1818
rect 7313 1710 7359 1786
rect 7473 1710 7519 1786
rect 7963 1730 8009 1806
rect 8137 1730 8183 1806
rect 11325 1696 11371 1772
rect 11485 1696 11531 1772
rect 7382 1629 7393 1675
rect 8039 1649 8050 1695
rect 11394 1615 11405 1661
rect 11786 1484 11826 1962
rect 16370 1873 16381 1919
rect 16427 1873 16438 1884
rect 16494 1859 16530 1883
rect 16532 1872 16543 1918
rect 16602 1859 16638 1883
rect 16494 1840 16538 1859
rect 16482 1839 16538 1840
rect 16594 1839 16638 1859
rect 16494 1838 16640 1839
rect 12030 1785 12041 1831
rect 12087 1785 12098 1796
rect 11961 1674 12007 1750
rect 12121 1674 12167 1750
rect 13618 1749 13629 1795
rect 16301 1762 16347 1838
rect 16461 1762 16640 1838
rect 16494 1760 16640 1762
rect 13675 1749 13686 1760
rect 16492 1759 16640 1760
rect 16492 1758 16582 1759
rect 16494 1739 16538 1758
rect 16539 1757 16540 1758
rect 16594 1739 16638 1759
rect 12030 1593 12041 1639
rect 12832 1607 12843 1653
rect 13549 1638 13595 1714
rect 13709 1638 13755 1714
rect 16370 1681 16381 1727
rect 16494 1714 16530 1739
rect 16532 1680 16543 1726
rect 16602 1715 16638 1739
rect 12889 1607 12900 1618
rect 12763 1496 12809 1572
rect 12923 1496 12969 1572
rect 13618 1557 13629 1603
rect 16370 1561 16381 1607
rect 16427 1561 16438 1572
rect 12832 1415 12843 1461
rect 13618 1437 13629 1483
rect 16301 1450 16347 1526
rect 16461 1450 16507 1526
rect 13675 1437 13686 1448
rect 12832 1295 12843 1341
rect 13549 1326 13595 1402
rect 13709 1326 13755 1402
rect 16370 1369 16381 1415
rect 12889 1295 12900 1306
rect 12763 1184 12809 1260
rect 12923 1184 12969 1260
rect 13618 1245 13629 1291
rect 16370 1249 16381 1295
rect 16427 1249 16438 1260
rect 12832 1103 12843 1149
rect 13618 1125 13629 1171
rect 16301 1138 16347 1214
rect 16461 1138 16507 1214
rect 13675 1125 13686 1136
rect 12832 983 12843 1029
rect 13549 1014 13595 1090
rect 13709 1014 13755 1090
rect 16370 1057 16381 1103
rect 12889 983 12900 994
rect 12763 872 12809 948
rect 12923 872 12969 948
rect 13618 933 13629 979
rect 16370 937 16381 983
rect 16427 937 16438 948
rect 12832 791 12843 837
rect 13618 813 13629 859
rect 16301 826 16347 902
rect 16461 826 16507 902
rect 13675 813 13686 824
rect 12000 671 12011 717
rect 12057 671 12068 682
rect 12832 671 12843 717
rect 13549 702 13595 778
rect 13709 702 13755 778
rect 16370 745 16381 791
rect 12889 671 12900 682
rect 11931 560 11977 636
rect 12091 560 12137 636
rect 12763 560 12809 636
rect 12923 560 12969 636
rect 13618 621 13629 667
rect 16370 625 16381 671
rect 16427 625 16438 636
rect 12000 479 12011 525
rect 12832 479 12843 525
rect 13618 501 13629 547
rect 16301 514 16347 590
rect 16461 514 16507 590
rect 13675 501 13686 512
rect 13549 390 13595 466
rect 13709 390 13755 466
rect 16370 433 16381 479
rect 13618 309 13629 355
rect 16370 313 16381 359
rect 16427 313 16438 324
rect 13618 189 13629 235
rect 13675 189 13686 200
rect 15560 179 15571 225
rect 16301 202 16347 278
rect 16461 202 16507 278
rect 15617 179 15628 190
rect 12004 41 12015 87
rect 13549 78 13595 154
rect 13709 78 13755 154
rect 15491 68 15537 144
rect 15651 68 15697 144
rect 16370 121 16381 167
rect 12061 41 12072 52
rect 11935 -70 11981 6
rect 12095 -70 12141 6
rect 13618 -3 13629 43
rect 15560 -13 15571 33
rect 16370 1 16381 47
rect 16427 1 16438 12
rect 12004 -151 12015 -105
rect 13618 -123 13629 -77
rect 13675 -123 13686 -112
rect 15560 -133 15571 -87
rect 16301 -110 16347 -34
rect 16461 -110 16507 -34
rect 15617 -133 15628 -122
rect 12004 -271 12015 -225
rect 13549 -234 13595 -158
rect 13709 -234 13755 -158
rect 12061 -271 12072 -260
rect 11935 -382 11981 -306
rect 12095 -382 12141 -306
rect 13618 -315 13629 -269
rect 15353 -300 15385 -199
rect 15491 -244 15537 -168
rect 15651 -244 15697 -168
rect 16370 -191 16381 -145
rect 15064 -385 15075 -339
rect 15121 -385 15132 -374
rect 12004 -463 12015 -417
rect 13618 -435 13629 -389
rect 13675 -435 13686 -424
rect 13549 -546 13595 -470
rect 13709 -546 13755 -470
rect 14857 -552 14889 -451
rect 14995 -496 15041 -420
rect 15155 -496 15201 -420
rect 13618 -627 13629 -581
rect 14568 -637 14579 -591
rect 14625 -637 14636 -626
rect 14499 -748 14545 -672
rect 14659 -748 14705 -672
rect 14568 -829 14579 -783
rect 14857 -820 14891 -552
rect 15064 -577 15075 -531
rect 15064 -697 15075 -651
rect 15121 -697 15132 -686
rect 14995 -808 15041 -732
rect 15155 -808 15201 -732
rect 9709 -915 9720 -869
rect 14857 -923 14889 -820
rect 15064 -889 15075 -843
rect 15353 -880 15387 -300
rect 15560 -325 15571 -279
rect 15560 -445 15571 -399
rect 15617 -445 15628 -434
rect 15491 -556 15537 -480
rect 15651 -556 15697 -480
rect 15560 -637 15571 -591
rect 15560 -757 15571 -711
rect 15617 -757 15628 -746
rect 15491 -868 15537 -792
rect 15651 -868 15697 -792
rect 9633 -1026 9679 -950
rect 9807 -1026 9853 -950
rect 15353 -983 15385 -880
rect 15560 -949 15571 -903
rect 9709 -1107 9720 -1061
<< metal1 >>
rect 9734 214 9810 224
rect 9734 -342 9744 214
rect 9800 -342 9810 214
rect 9734 -352 9810 -342
<< via1 >>
rect 9744 -342 9800 214
<< metal2 >>
rect 9734 214 9810 224
rect 9734 -342 9744 214
rect 9800 -342 9810 214
rect 9734 -536 9810 -342
use nfet_03v3_5KTYYT  nfet_03v3_5KTYYT_0
timestamp 1756956737
transform 1 0 10532 0 1 768
box -820 -216 820 216
use nfet_03v3_5KTYYT  nfet_03v3_5KTYYT_1
timestamp 1756956737
transform 1 0 9012 0 1 768
box -820 -216 820 216
use nfet_03v3_58UUYT  nfet_03v3_58UUYT_0
timestamp 1756956737
transform 1 0 10532 0 1 -64
box -820 -416 820 416
use pfet_03v3_KUQE4Y  XM1
timestamp 1756956737
transform 1 0 7416 0 1 1748
box -278 -250 278 250
use pfet_03v3_H5R3BY  XM2
timestamp 1756956737
transform 1 0 12064 0 1 1712
box -278 -250 278 250
use pfet_03v3_V5CHCW  XM3
timestamp 1756956737
transform 1 0 9188 0 1 1794
box -654 -310 654 310
use pfet_03v3_V5CHCW  XM4
timestamp 1756956737
transform 1 0 10376 0 1 1794
box -654 -310 654 310
use pfet_03v3_H5R3BY  XM5
timestamp 1756956737
transform 1 0 11428 0 1 1734
box -278 -250 278 250
use pfet_03v3_KUUUNT  XM6
timestamp 1756956737
transform 1 0 8073 0 1 1768
box -209 -218 209 218
use nfet_03v3_58UUYT  XM9
timestamp 1756956737
transform 1 0 9012 0 1 -64
box -820 -416 820 416
use nfet_03v3_J7ZQZQ  XM11
timestamp 1756956737
transform 1 0 9743 0 1 -988
box -147 -156 147 156
use pfet_03v3_H5R3BY  XM12
timestamp 1756956737
transform 1 0 12034 0 1 598
box -278 -250 278 250
use pfet_03v3_HDLTJN  XM13
timestamp 1756956737
transform 1 0 12038 0 1 -188
box -278 -406 278 406
use pfet_03v3_GU2533  XM14
timestamp 1756956737
transform 1 0 12866 0 1 1066
box -278 -718 278 718
use pfet_03v3_HVKTJN  XM15
timestamp 1756956737
transform 1 0 13652 0 1 584
box -278 -1342 278 1342
use pfet_03v3_H5R3BY  XM16
timestamp 1756956737
transform 1 0 14602 0 1 -710
box -278 -250 278 250
use pfet_03v3_HDLTJN  XM17
timestamp 1756956737
transform 1 0 15098 0 1 -614
box -278 -406 278 406
use pfet_03v3_GU2533  XM18
timestamp 1756956737
transform 1 0 15594 0 1 -362
box -278 -718 278 718
use pfet_03v3_KUCGSX  XM19
timestamp 1756957756
transform 1 0 16404 0 1 1020
box -116 -1224 236 1132
<< end >>
