magic
tech gf180mcuD
magscale 1 10
timestamp 1757566850
<< error_p >>
rect -38 133 -27 179
rect -38 -179 -27 -133
<< pwell >>
rect -290 -310 290 310
<< nmos >>
rect -40 -100 40 100
<< ndiff >>
rect -128 87 -40 100
rect -128 -87 -115 87
rect -69 -87 -40 87
rect -128 -100 -40 -87
rect 40 87 128 100
rect 40 -87 69 87
rect 115 -87 128 87
rect 40 -100 128 -87
<< ndiffc >>
rect -115 -87 -69 87
rect 69 -87 115 87
<< psubdiff >>
rect -266 214 266 286
rect -266 170 -194 214
rect -266 -170 -253 170
rect -207 -170 -194 170
rect 194 170 266 214
rect -266 -214 -194 -170
rect 194 -170 207 170
rect 253 -170 266 170
rect 194 -214 266 -170
rect -266 -286 266 -214
<< psubdiffcont >>
rect -253 -170 -207 170
rect 207 -170 253 170
<< polysilicon >>
rect -40 179 40 192
rect -40 133 -27 179
rect 27 133 40 179
rect -40 100 40 133
rect -40 -133 40 -100
rect -40 -179 -27 -133
rect 27 -179 40 -133
rect -40 -192 40 -179
<< polycontact >>
rect -27 133 27 179
rect -27 -179 27 -133
<< metal1 >>
rect -253 170 -207 181
rect -38 133 -27 179
rect 27 133 38 179
rect 207 170 253 181
rect -115 87 -69 98
rect -115 -98 -69 -87
rect 69 87 115 98
rect 69 -98 115 -87
rect -253 -181 -207 -170
rect -38 -179 -27 -133
rect 27 -179 38 -133
rect 207 -181 253 -170
<< properties >>
string FIXED_BBOX -230 -250 230 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
