** sch_path: /foss/designs/libs/WK_Kadam/CDAC_Switch_V2/c_dac2_switch.sch
.subckt c_dac2_switch sw_vout sw_bit avss avdd sw_Vref vreflow
*.PININFO avdd:B avss:B sw_bit:B sw_vout:B sw_Vref:B vreflow:B
XM1 sw_vout sw_bit sw_Vref avss nfet_03v3 L=0.4u W=4u nf=2 m=1
XM3 sw_vout net1 vreflow avss nfet_03v3 L=0.4u W=4u nf=2 m=1
XM4 vreflow sw_bit sw_vout avdd pfet_03v3 L=0.4u W=4u nf=2 m=1
XM2 sw_Vref net1 sw_vout avdd pfet_03v3 L=0.4u W=4u nf=2 m=1
x1 avdd sw_bit net1 avss CDAC_INV_V0
.ends

* expanding   symbol:  libs/WK_Kadam/MK_INV_v1/CDAC_INV_V0.sym # of pins=4
** sym_path: /foss/designs/libs/WK_Kadam/MK_INV_v1/CDAC_INV_V0.sym
** sch_path: /foss/designs/libs/WK_Kadam/MK_INV_v1/CDAC_INV_V0.sch
.subckt CDAC_INV_V0 avdd in out avss
*.PININFO avdd:B avss:B in:B out:B
XXM3 out in avss avss nfet_03v3 L=0.4u W=2u nf=1 m=1
XXM4 out in avdd avdd pfet_03v3 L=0.4u W=4u nf=1 m=1
.ends

