magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< error_p >>
rect -34 73 -23 119
rect -110 -38 -64 38
rect 64 -38 110 38
rect -34 -119 -23 -73
<< pwell >>
rect -147 -156 147 156
<< nmos >>
rect -35 -40 35 40
<< ndiff >>
rect -123 27 -35 40
rect -123 -27 -110 27
rect -64 -27 -35 27
rect -123 -40 -35 -27
rect 35 27 123 40
rect 35 -27 64 27
rect 110 -27 123 27
rect 35 -40 123 -27
<< ndiffc >>
rect -110 -27 -64 27
rect 64 -27 110 27
<< polysilicon >>
rect -36 119 36 132
rect -36 73 -23 119
rect 23 73 36 119
rect -36 60 36 73
rect -35 40 35 60
rect -35 -60 35 -40
rect -36 -73 36 -60
rect -36 -119 -23 -73
rect 23 -119 36 -73
rect -36 -132 36 -119
<< polycontact >>
rect -23 73 23 119
rect -23 -119 23 -73
<< metal1 >>
rect -34 73 -23 119
rect 23 73 34 119
rect -110 27 -64 38
rect -110 -38 -64 -27
rect 64 27 110 38
rect 64 -38 110 -27
rect -34 -119 -23 -73
rect 23 -119 34 -73
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.4 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
