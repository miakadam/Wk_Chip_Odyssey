magic
tech gf180mcuD
magscale 1 10
timestamp 1758005944
<< nwell >>
rect -1553 910 -953 1930
rect -665 910 415 1930
<< pwell >>
rect 67 821 153 901
rect -1553 190 415 810
<< nmos >>
rect -1303 400 -1203 600
rect -1099 400 -999 600
rect -619 400 -519 600
rect -415 400 -315 600
rect 65 400 165 600
<< pmos >>
rect -1303 1120 -1203 1720
rect -415 1120 -315 1720
rect 65 1120 165 1720
<< ndiff >>
rect -1391 587 -1303 600
rect -1391 413 -1378 587
rect -1332 413 -1303 587
rect -1391 400 -1303 413
rect -1203 587 -1099 600
rect -1203 413 -1174 587
rect -1128 413 -1099 587
rect -1203 400 -1099 413
rect -999 587 -911 600
rect -999 413 -970 587
rect -924 413 -911 587
rect -999 400 -911 413
rect -707 587 -619 600
rect -707 413 -694 587
rect -648 413 -619 587
rect -707 400 -619 413
rect -519 587 -415 600
rect -519 413 -490 587
rect -444 413 -415 587
rect -519 400 -415 413
rect -315 587 -227 600
rect -315 413 -286 587
rect -240 413 -227 587
rect -315 400 -227 413
rect -23 587 65 600
rect -23 413 -10 587
rect 36 413 65 587
rect -23 400 65 413
rect 165 587 253 600
rect 165 413 194 587
rect 240 413 253 587
rect 165 400 253 413
<< pdiff >>
rect -1391 1707 -1303 1720
rect -1391 1133 -1378 1707
rect -1332 1133 -1303 1707
rect -1391 1120 -1303 1133
rect -1203 1707 -1115 1720
rect -1203 1133 -1174 1707
rect -1128 1133 -1115 1707
rect -1203 1120 -1115 1133
rect -503 1707 -415 1720
rect -503 1133 -490 1707
rect -444 1133 -415 1707
rect -503 1120 -415 1133
rect -315 1707 -227 1720
rect -315 1133 -286 1707
rect -240 1133 -227 1707
rect -315 1120 -227 1133
rect -23 1707 65 1720
rect -23 1133 -10 1707
rect 36 1133 65 1707
rect -23 1120 65 1133
rect 165 1707 253 1720
rect 165 1133 194 1707
rect 240 1133 253 1707
rect 165 1120 253 1133
<< ndiffc >>
rect -1378 413 -1332 587
rect -1174 413 -1128 587
rect -970 413 -924 587
rect -694 413 -648 587
rect -490 413 -444 587
rect -286 413 -240 587
rect -10 413 36 587
rect 194 413 240 587
<< pdiffc >>
rect -1378 1133 -1332 1707
rect -1174 1133 -1128 1707
rect -490 1133 -444 1707
rect -286 1133 -240 1707
rect -10 1133 36 1707
rect 194 1133 240 1707
<< psubdiff >>
rect -1529 714 391 786
rect -1529 670 -1457 714
rect -1529 330 -1516 670
rect -1470 330 -1457 670
rect -845 670 -773 714
rect -1529 286 -1457 330
rect -845 330 -832 670
rect -786 330 -773 670
rect -161 670 -89 714
rect -845 286 -773 330
rect -161 330 -148 670
rect -102 330 -89 670
rect 319 670 391 714
rect -161 286 -89 330
rect 319 330 332 670
rect 378 330 391 670
rect 319 286 391 330
rect -1529 214 391 286
<< nsubdiff >>
rect -1529 1834 -977 1906
rect -1529 1790 -1457 1834
rect -1529 1050 -1516 1790
rect -1470 1050 -1457 1790
rect -1049 1790 -977 1834
rect -1529 1006 -1457 1050
rect -1049 1050 -1036 1790
rect -990 1050 -977 1790
rect -1049 1006 -977 1050
rect -1529 934 -977 1006
rect -641 1834 391 1906
rect -641 1790 -569 1834
rect -641 1050 -628 1790
rect -582 1050 -569 1790
rect -161 1790 -89 1834
rect -641 1006 -569 1050
rect -161 1050 -148 1790
rect -102 1050 -89 1790
rect 319 1790 391 1834
rect -161 1006 -89 1050
rect 319 1050 332 1790
rect 378 1050 391 1790
rect 319 1006 391 1050
rect -641 934 391 1006
<< psubdiffcont >>
rect -1516 330 -1470 670
rect -832 330 -786 670
rect -148 330 -102 670
rect 332 330 378 670
<< nsubdiffcont >>
rect -1516 1050 -1470 1790
rect -1036 1050 -990 1790
rect -628 1050 -582 1790
rect -148 1050 -102 1790
rect 332 1050 378 1790
<< polysilicon >>
rect -1303 1799 -1203 1812
rect -1303 1753 -1290 1799
rect -1216 1753 -1203 1799
rect -1303 1720 -1203 1753
rect -1303 1087 -1203 1120
rect -1303 1041 -1290 1087
rect -1216 1041 -1203 1087
rect -1303 1028 -1203 1041
rect -415 1799 -315 1812
rect -415 1753 -402 1799
rect -328 1753 -315 1799
rect -415 1720 -315 1753
rect -415 1087 -315 1120
rect -415 1041 -402 1087
rect -328 1041 -315 1087
rect -415 1028 -315 1041
rect 65 1799 165 1812
rect 65 1753 78 1799
rect 152 1753 165 1799
rect 65 1720 165 1753
rect 65 1087 165 1120
rect 65 1041 78 1087
rect 152 1041 165 1087
rect 65 1028 165 1041
rect -1303 679 -1203 692
rect -1303 633 -1290 679
rect -1216 633 -1203 679
rect -1303 600 -1203 633
rect -1099 679 -999 692
rect -1099 633 -1086 679
rect -1012 633 -999 679
rect -1099 600 -999 633
rect -1303 367 -1203 400
rect -1303 321 -1290 367
rect -1216 321 -1203 367
rect -1303 308 -1203 321
rect -1099 367 -999 400
rect -1099 321 -1086 367
rect -1012 321 -999 367
rect -1099 308 -999 321
rect -619 679 -519 692
rect -619 633 -606 679
rect -532 633 -519 679
rect -619 600 -519 633
rect -415 679 -315 692
rect -415 633 -402 679
rect -328 633 -315 679
rect -415 600 -315 633
rect -619 367 -519 400
rect -619 321 -606 367
rect -532 321 -519 367
rect -619 308 -519 321
rect -415 367 -315 400
rect -415 321 -402 367
rect -328 321 -315 367
rect -415 308 -315 321
rect 65 679 165 692
rect 65 633 78 679
rect 152 633 165 679
rect 65 600 165 633
rect 65 367 165 400
rect 65 321 78 367
rect 152 321 165 367
rect 65 308 165 321
<< polycontact >>
rect -1290 1753 -1216 1799
rect -1290 1041 -1216 1087
rect -402 1753 -328 1799
rect -402 1041 -328 1087
rect 78 1753 152 1799
rect 78 1041 152 1087
rect -1290 633 -1216 679
rect -1086 633 -1012 679
rect -1290 321 -1216 367
rect -1086 321 -1012 367
rect -606 633 -532 679
rect -402 633 -328 679
rect -606 321 -532 367
rect -402 321 -328 367
rect 78 633 152 679
rect 78 321 152 367
<< metal1 >>
rect -1553 1930 415 2130
rect -1516 1790 -1470 1801
rect -1301 1799 -1205 1830
rect -1301 1753 -1290 1799
rect -1216 1753 -1205 1799
rect -1036 1790 -582 1930
rect -1378 1707 -1332 1718
rect -1395 1423 -1378 1433
rect -1174 1707 -1036 1718
rect -1332 1423 -1315 1433
rect -1395 1183 -1383 1423
rect -1327 1183 -1315 1423
rect -1395 1173 -1378 1183
rect -1332 1173 -1315 1183
rect -1378 1122 -1332 1133
rect -1128 1133 -1036 1707
rect -1174 1122 -1036 1133
rect -1516 1039 -1470 1050
rect -1301 1041 -1290 1087
rect -1216 1041 -1205 1087
rect -1301 966 -1205 1041
rect -990 1122 -628 1790
rect -1036 1039 -990 1050
rect -413 1799 -317 1830
rect -413 1753 -402 1799
rect -328 1753 -317 1799
rect -148 1790 -102 1930
rect -582 1707 -444 1718
rect -582 1133 -490 1707
rect -286 1707 -240 1718
rect -303 1423 -286 1433
rect -240 1423 -223 1433
rect -303 1183 -291 1423
rect -235 1183 -223 1423
rect -303 1173 -286 1183
rect -582 1122 -444 1133
rect -240 1173 -223 1183
rect -286 1122 -240 1133
rect -628 1039 -582 1050
rect -413 1041 -402 1087
rect -328 1041 -317 1087
rect -1301 910 -1281 966
rect -1225 910 -1205 966
rect -1301 692 -1205 910
rect -413 822 -317 1041
rect 67 1799 163 1830
rect 67 1753 78 1799
rect 152 1753 163 1799
rect 332 1790 378 1930
rect -102 1707 36 1718
rect -102 1133 -10 1707
rect 194 1707 240 1718
rect 177 1423 194 1433
rect 240 1423 257 1433
rect 177 1183 189 1423
rect 245 1183 257 1423
rect 177 1173 194 1183
rect -102 1122 36 1133
rect 240 1173 257 1183
rect 194 1122 240 1133
rect -148 1039 -102 1050
rect 67 1041 78 1087
rect 152 1041 163 1087
rect 67 900 163 1041
rect 332 1039 378 1050
rect -481 810 -317 822
rect -1 888 163 900
rect -1 832 11 888
rect 67 832 163 888
rect -1 820 163 832
rect -481 754 -469 810
rect -413 754 -317 810
rect -481 742 -317 754
rect -413 692 -317 742
rect -1516 670 -1470 681
rect -1301 679 -1001 692
rect -1301 633 -1290 679
rect -1216 646 -1086 679
rect -1216 633 -1205 646
rect -1097 633 -1086 646
rect -1012 633 -1001 679
rect -832 670 -786 681
rect -1470 587 -1332 598
rect -1470 413 -1378 587
rect -1174 587 -1128 598
rect -1191 528 -1174 538
rect -970 587 -832 598
rect -1128 528 -1111 538
rect -1191 472 -1179 528
rect -1123 472 -1111 528
rect -1191 462 -1174 472
rect -1470 402 -1332 413
rect -1128 462 -1111 472
rect -1174 402 -1128 413
rect -924 413 -832 587
rect -970 402 -832 413
rect -1516 190 -1470 330
rect -1301 321 -1290 367
rect -1216 321 -1205 367
rect -1301 290 -1205 321
rect -1097 321 -1086 367
rect -1012 321 -1001 367
rect -1097 290 -1001 321
rect -617 679 -317 692
rect -617 633 -606 679
rect -532 646 -402 679
rect -532 633 -521 646
rect -413 633 -402 646
rect -328 633 -317 679
rect -148 670 -102 681
rect -694 587 -648 598
rect -711 528 -694 538
rect -490 587 -444 598
rect -648 528 -631 538
rect -711 472 -699 528
rect -643 472 -631 528
rect -711 462 -694 472
rect -648 462 -631 472
rect -507 528 -490 538
rect -286 587 -240 598
rect -444 528 -427 538
rect -507 472 -495 528
rect -439 472 -427 528
rect -507 462 -490 472
rect -694 402 -648 413
rect -444 462 -427 472
rect -303 528 -286 538
rect -240 528 -223 538
rect -303 472 -291 528
rect -235 472 -223 528
rect -303 462 -286 472
rect -490 402 -444 413
rect -240 462 -223 472
rect -286 402 -240 413
rect -832 190 -786 330
rect -617 321 -606 367
rect -532 321 -521 367
rect -617 290 -521 321
rect -413 321 -402 367
rect -328 321 -317 367
rect -413 290 -317 321
rect 67 679 163 820
rect 67 633 78 679
rect 152 633 163 679
rect 332 670 378 681
rect -102 587 36 598
rect -102 413 -10 587
rect 194 587 240 598
rect 177 528 194 538
rect 240 528 257 538
rect 177 472 189 528
rect 245 472 257 528
rect 177 462 194 472
rect -102 402 36 413
rect 240 462 257 472
rect 194 402 240 413
rect -148 190 -102 330
rect 67 321 78 367
rect 152 321 163 367
rect 67 290 163 321
rect 332 190 378 330
rect -1553 -10 415 190
<< via1 >>
rect -1383 1183 -1378 1423
rect -1378 1183 -1332 1423
rect -1332 1183 -1327 1423
rect -291 1183 -286 1423
rect -286 1183 -240 1423
rect -240 1183 -235 1423
rect -1281 910 -1225 966
rect 189 1183 194 1423
rect 194 1183 240 1423
rect 240 1183 245 1423
rect 11 832 67 888
rect -469 754 -413 810
rect -1179 472 -1174 528
rect -1174 472 -1128 528
rect -1128 472 -1123 528
rect -699 472 -694 528
rect -694 472 -648 528
rect -648 472 -643 528
rect -495 472 -490 528
rect -490 472 -444 528
rect -444 472 -439 528
rect -291 472 -286 528
rect -286 472 -240 528
rect -240 472 -235 528
rect 189 472 194 528
rect 194 472 240 528
rect 240 472 245 528
<< metal2 >>
rect -1395 1423 -223 1433
rect -1395 1183 -1383 1423
rect -1327 1183 -291 1423
rect -235 1183 -223 1423
rect -1395 1173 -223 1183
rect -1301 966 -1223 978
rect -1647 910 -1281 966
rect -1225 910 -1223 966
rect -1301 898 -1223 910
rect -303 888 -223 1173
rect 177 1423 257 1433
rect 177 1183 189 1423
rect 245 1183 257 1423
rect -1 888 69 900
rect -303 832 11 888
rect 67 832 69 888
rect -481 810 -411 822
rect -1647 754 -469 810
rect -413 754 -411 810
rect -481 742 -411 754
rect -1191 528 -1111 538
rect -1191 472 -1179 528
rect -1123 472 -1111 528
rect -1191 286 -1111 472
rect -711 528 -631 538
rect -711 472 -699 528
rect -643 472 -631 528
rect -711 462 -631 472
rect -507 528 -427 538
rect -507 472 -495 528
rect -439 472 -427 528
rect -507 286 -427 472
rect -303 528 -223 832
rect -1 820 69 832
rect 177 888 257 1183
rect 177 832 422 888
rect -303 472 -291 528
rect -235 472 -223 528
rect -303 462 -223 472
rect 177 528 257 832
rect 177 472 189 528
rect 245 472 257 528
rect 177 462 257 472
rect -1191 214 -427 286
<< via2 >>
rect -699 472 -643 528
rect -291 472 -235 528
<< metal3 >>
rect -711 528 -223 538
rect -711 472 -699 528
rect -643 472 -291 528
rect -235 472 -223 528
rect -711 462 -223 472
<< labels >>
rlabel metal1 -580 2130 -580 2130 1 VDD
port 0 n
rlabel metal2 422 858 422 858 3 OUT
port 1 e
rlabel metal2 -1647 937 -1647 937 7 A
port 2 w
rlabel metal2 -1647 782 -1647 782 7 B
port 3 w
rlabel metal1 -521 -10 -521 -10 5 VSS
port 4 s
<< end >>
