magic
tech gf180mcuD
magscale 1 10
timestamp 1755269198
<< error_s >>
rect 1164 257 1346 266
rect 544 176 555 209
rect 1208 208 1210 220
rect 1220 218 1222 220
rect 1288 196 1290 220
rect 1300 208 1302 220
rect 1254 176 1290 196
rect 544 163 576 176
rect 584 163 612 176
rect 1210 163 1235 176
rect 1210 162 1247 163
rect 1208 150 1247 162
rect 1254 162 1300 176
rect 1254 150 1302 162
rect 1254 140 1290 150
rect 448 118 450 130
rect 448 -30 450 -18
rect 460 -30 462 130
rect 518 16 520 130
rect 530 118 532 130
rect 1298 118 1300 130
rect 484 -4 520 16
rect 484 -18 530 -4
rect 484 -30 532 -18
rect 630 -30 666 -4
rect 1310 -17 1312 130
rect 1178 -28 1201 -17
rect 1300 -18 1338 -17
rect 1178 -30 1200 -28
rect 1298 -30 1338 -18
rect 1368 -30 1370 130
rect 1380 118 1382 130
rect 1380 -30 1382 -18
rect 484 -40 520 -30
rect 528 -62 530 -50
rect 528 -111 530 -108
rect 540 -111 576 -40
rect 608 -52 610 -50
rect 620 -62 622 -50
rect 620 -111 622 -108
rect 1224 -109 1235 -63
rect 528 -120 622 -111
rect 540 -130 576 -120
rect 594 -504 605 -471
rect 594 -517 626 -504
rect 651 -517 662 -504
rect 1174 -517 1185 -471
rect 1204 -517 1242 -504
rect 498 -562 500 -550
rect 498 -710 500 -698
rect 510 -710 512 -550
rect 568 -664 570 -550
rect 580 -562 582 -550
rect 1248 -562 1250 -550
rect 534 -674 570 -664
rect 524 -684 570 -674
rect 1260 -664 1262 -550
rect 1260 -674 1306 -664
rect 1260 -684 1316 -674
rect 524 -698 580 -684
rect 524 -710 582 -698
rect 685 -708 726 -684
rect 690 -710 726 -708
rect 1114 -708 1151 -684
rect 1250 -698 1316 -684
rect 1114 -710 1150 -708
rect 1248 -710 1316 -698
rect 1318 -710 1320 -550
rect 1330 -562 1332 -550
rect 1330 -710 1332 -698
rect 524 -720 570 -710
rect 1260 -720 1316 -710
rect 578 -742 580 -730
rect 590 -732 592 -730
rect 668 -732 670 -730
rect 680 -742 682 -730
rect 1158 -742 1160 -730
rect 1170 -732 1172 -730
rect 1248 -732 1250 -730
rect 1260 -742 1262 -730
rect 580 -798 680 -791
rect 1160 -798 1260 -791
rect 578 -810 682 -798
rect 1158 -810 1262 -798
<< metal1 >>
rect 300 270 1540 510
rect 780 130 1060 270
rect 1210 150 1220 220
rect 1290 150 1300 220
rect 450 -30 460 130
rect 520 -30 530 130
rect 630 -30 1200 130
rect 1300 -30 1310 130
rect 1370 -30 1380 130
rect 530 -120 540 -50
rect 610 -120 620 -50
rect 780 -200 1060 -30
rect 830 -550 1000 -380
rect 500 -710 510 -550
rect 570 -710 580 -550
rect 690 -710 1150 -550
rect 1250 -710 1260 -550
rect 1320 -710 1330 -550
rect 580 -810 590 -730
rect 670 -810 680 -730
rect 830 -850 1000 -710
rect 1160 -810 1170 -730
rect 1250 -810 1260 -730
rect 340 -1080 1490 -850
<< via1 >>
rect 1220 150 1290 220
rect 460 -30 520 130
rect 1310 -30 1370 130
rect 540 -120 610 -50
rect 510 -710 570 -550
rect 1260 -710 1320 -550
rect 590 -810 670 -730
rect 1170 -810 1250 -730
<< metal2 >>
rect 1220 220 1290 230
rect 460 150 1220 220
rect 460 130 520 150
rect 1220 140 1290 150
rect 460 -260 520 -30
rect 1310 130 1370 140
rect 540 -50 610 -40
rect 1310 -50 1370 -30
rect 610 -120 1370 -50
rect 540 -130 610 -120
rect 20 -270 520 -260
rect 1310 -260 1370 -120
rect 1310 -270 1810 -260
rect 20 -330 570 -270
rect 510 -550 570 -330
rect 510 -720 570 -710
rect 1260 -330 1810 -270
rect 1260 -550 1320 -330
rect 1260 -720 1320 -710
rect 590 -730 670 -720
rect 1170 -730 1250 -720
rect 580 -810 590 -730
rect 670 -810 680 -730
rect 580 -1240 680 -810
rect 1160 -810 1170 -730
rect 1250 -810 1260 -730
rect 1160 -1240 1260 -810
use nfet_03v3_5QDTWG  XM1
timestamp 1755268346
transform 1 0 628 0 1 -630
box -278 -290 278 290
use nfet_03v3_5QDTWG  XM2
timestamp 1755268346
transform 1 0 1208 0 1 -630
box -278 -290 278 290
use pfet_03v3_YBHBCY  XM3
timestamp 1755268346
transform 1 0 578 0 1 50
box -278 -290 278 290
use pfet_03v3_YBHBCY  XM4
timestamp 1755268346
transform 1 0 1258 0 1 50
box -278 -290 278 290
<< labels >>
rlabel metal1 300 480 300 480 1 VDD
port 0 n
rlabel metal1 340 -1020 340 -1020 1 VSS
port 1 n
rlabel metal2 630 -1240 630 -1240 5 Vin1
port 2 s
rlabel metal2 1210 -1240 1210 -1240 5 Vin2
port 3 s
rlabel metal2 20 -300 20 -300 7 Vout1
port 4 w
rlabel metal2 1810 -300 1810 -300 3 Vout2
port 5 e
<< end >>
