magic
tech gf180mcuD
magscale 1 10
timestamp 1757406152
<< pwell >>
rect -1262 -310 1262 310
<< nmos >>
rect -1012 -100 -812 100
rect -708 -100 -508 100
rect -404 -100 -204 100
rect -100 -100 100 100
rect 204 -100 404 100
rect 508 -100 708 100
rect 812 -100 1012 100
<< ndiff >>
rect -1100 87 -1012 100
rect -1100 -87 -1087 87
rect -1041 -87 -1012 87
rect -1100 -100 -1012 -87
rect -812 87 -708 100
rect -812 -87 -783 87
rect -737 -87 -708 87
rect -812 -100 -708 -87
rect -508 87 -404 100
rect -508 -87 -479 87
rect -433 -87 -404 87
rect -508 -100 -404 -87
rect -204 87 -100 100
rect -204 -87 -175 87
rect -129 -87 -100 87
rect -204 -100 -100 -87
rect 100 87 204 100
rect 100 -87 129 87
rect 175 -87 204 87
rect 100 -100 204 -87
rect 404 87 508 100
rect 404 -87 433 87
rect 479 -87 508 87
rect 404 -100 508 -87
rect 708 87 812 100
rect 708 -87 737 87
rect 783 -87 812 87
rect 708 -100 812 -87
rect 1012 87 1100 100
rect 1012 -87 1041 87
rect 1087 -87 1100 87
rect 1012 -100 1100 -87
<< ndiffc >>
rect -1087 -87 -1041 87
rect -783 -87 -737 87
rect -479 -87 -433 87
rect -175 -87 -129 87
rect 129 -87 175 87
rect 433 -87 479 87
rect 737 -87 783 87
rect 1041 -87 1087 87
<< psubdiff >>
rect -1238 214 1238 286
rect -1238 170 -1166 214
rect -1238 -170 -1225 170
rect -1179 -170 -1166 170
rect 1166 170 1238 214
rect -1238 -214 -1166 -170
rect 1166 -170 1179 170
rect 1225 -170 1238 170
rect 1166 -214 1238 -170
rect -1238 -286 1238 -214
<< psubdiffcont >>
rect -1225 -170 -1179 170
rect 1179 -170 1225 170
<< polysilicon >>
rect -1012 179 -812 192
rect -1012 133 -999 179
rect -825 133 -812 179
rect -1012 100 -812 133
rect -708 179 -508 192
rect -708 133 -695 179
rect -521 133 -508 179
rect -708 100 -508 133
rect -404 179 -204 192
rect -404 133 -391 179
rect -217 133 -204 179
rect -404 100 -204 133
rect -100 179 100 192
rect -100 133 -87 179
rect 87 133 100 179
rect -100 100 100 133
rect 204 179 404 192
rect 204 133 217 179
rect 391 133 404 179
rect 204 100 404 133
rect 508 179 708 192
rect 508 133 521 179
rect 695 133 708 179
rect 508 100 708 133
rect 812 179 1012 192
rect 812 133 825 179
rect 999 133 1012 179
rect 812 100 1012 133
rect -1012 -133 -812 -100
rect -1012 -179 -999 -133
rect -825 -179 -812 -133
rect -1012 -192 -812 -179
rect -708 -133 -508 -100
rect -708 -179 -695 -133
rect -521 -179 -508 -133
rect -708 -192 -508 -179
rect -404 -133 -204 -100
rect -404 -179 -391 -133
rect -217 -179 -204 -133
rect -404 -192 -204 -179
rect -100 -133 100 -100
rect -100 -179 -87 -133
rect 87 -179 100 -133
rect -100 -192 100 -179
rect 204 -133 404 -100
rect 204 -179 217 -133
rect 391 -179 404 -133
rect 204 -192 404 -179
rect 508 -133 708 -100
rect 508 -179 521 -133
rect 695 -179 708 -133
rect 508 -192 708 -179
rect 812 -133 1012 -100
rect 812 -179 825 -133
rect 999 -179 1012 -133
rect 812 -192 1012 -179
<< polycontact >>
rect -999 133 -825 179
rect -695 133 -521 179
rect -391 133 -217 179
rect -87 133 87 179
rect 217 133 391 179
rect 521 133 695 179
rect 825 133 999 179
rect -999 -179 -825 -133
rect -695 -179 -521 -133
rect -391 -179 -217 -133
rect -87 -179 87 -133
rect 217 -179 391 -133
rect 521 -179 695 -133
rect 825 -179 999 -133
<< metal1 >>
rect -1225 170 -1179 181
rect -1010 133 -999 179
rect -825 133 -814 179
rect -706 133 -695 179
rect -521 133 -510 179
rect -402 133 -391 179
rect -217 133 -206 179
rect -98 133 -87 179
rect 87 133 98 179
rect 206 133 217 179
rect 391 133 402 179
rect 510 133 521 179
rect 695 133 706 179
rect 814 133 825 179
rect 999 133 1010 179
rect 1179 170 1225 181
rect -1087 87 -1041 98
rect -1087 -98 -1041 -87
rect -783 87 -737 98
rect -783 -98 -737 -87
rect -479 87 -433 98
rect -479 -98 -433 -87
rect -175 87 -129 98
rect -175 -98 -129 -87
rect 129 87 175 98
rect 129 -98 175 -87
rect 433 87 479 98
rect 433 -98 479 -87
rect 737 87 783 98
rect 737 -98 783 -87
rect 1041 87 1087 98
rect 1041 -98 1087 -87
rect -1225 -181 -1179 -170
rect -1010 -179 -999 -133
rect -825 -179 -814 -133
rect -706 -179 -695 -133
rect -521 -179 -510 -133
rect -402 -179 -391 -133
rect -217 -179 -206 -133
rect -98 -179 -87 -133
rect 87 -179 98 -133
rect 206 -179 217 -133
rect 391 -179 402 -133
rect 510 -179 521 -133
rect 695 -179 706 -133
rect 814 -179 825 -133
rect 999 -179 1010 -133
rect 1179 -181 1225 -170
<< properties >>
string FIXED_BBOX -1202 -250 1202 250
string gencell nfet_03v3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
