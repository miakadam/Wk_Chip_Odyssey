magic
tech gf180mcuD
magscale 1 10
timestamp 1756956737
<< pwell >>
rect -820 -416 820 416
<< nmos >>
rect -708 -300 -508 300
rect -404 -300 -204 300
rect -100 -300 100 300
rect 204 -300 404 300
rect 508 -300 708 300
<< ndiff >>
rect -796 287 -708 300
rect -796 -287 -783 287
rect -737 -287 -708 287
rect -796 -300 -708 -287
rect -508 287 -404 300
rect -508 -287 -479 287
rect -433 -287 -404 287
rect -508 -300 -404 -287
rect -204 287 -100 300
rect -204 -287 -175 287
rect -129 -287 -100 287
rect -204 -300 -100 -287
rect 100 287 204 300
rect 100 -287 129 287
rect 175 -287 204 287
rect 100 -300 204 -287
rect 404 287 508 300
rect 404 -287 433 287
rect 479 -287 508 287
rect 404 -300 508 -287
rect 708 287 796 300
rect 708 -287 737 287
rect 783 -287 796 287
rect 708 -300 796 -287
<< ndiffc >>
rect -783 -287 -737 287
rect -479 -287 -433 287
rect -175 -287 -129 287
rect 129 -287 175 287
rect 433 -287 479 287
rect 737 -287 783 287
<< polysilicon >>
rect -708 379 -508 392
rect -708 333 -695 379
rect -521 333 -508 379
rect -708 300 -508 333
rect -404 379 -204 392
rect -404 333 -391 379
rect -217 333 -204 379
rect -404 300 -204 333
rect -100 379 100 392
rect -100 333 -87 379
rect 87 333 100 379
rect -100 300 100 333
rect 204 379 404 392
rect 204 333 217 379
rect 391 333 404 379
rect 204 300 404 333
rect 508 379 708 392
rect 508 333 521 379
rect 695 333 708 379
rect 508 300 708 333
rect -708 -333 -508 -300
rect -708 -379 -695 -333
rect -521 -379 -508 -333
rect -708 -392 -508 -379
rect -404 -333 -204 -300
rect -404 -379 -391 -333
rect -217 -379 -204 -333
rect -404 -392 -204 -379
rect -100 -333 100 -300
rect -100 -379 -87 -333
rect 87 -379 100 -333
rect -100 -392 100 -379
rect 204 -333 404 -300
rect 204 -379 217 -333
rect 391 -379 404 -333
rect 204 -392 404 -379
rect 508 -333 708 -300
rect 508 -379 521 -333
rect 695 -379 708 -333
rect 508 -392 708 -379
<< polycontact >>
rect -695 333 -521 379
rect -391 333 -217 379
rect -87 333 87 379
rect 217 333 391 379
rect 521 333 695 379
rect -695 -379 -521 -333
rect -391 -379 -217 -333
rect -87 -379 87 -333
rect 217 -379 391 -333
rect 521 -379 695 -333
<< metal1 >>
rect -706 333 -695 379
rect -521 333 -510 379
rect -402 333 -391 379
rect -217 333 -206 379
rect -98 333 -87 379
rect 87 333 98 379
rect 206 333 217 379
rect 391 333 402 379
rect 510 333 521 379
rect 695 333 706 379
rect -783 287 -737 298
rect -783 -298 -737 -287
rect -479 287 -433 298
rect -479 -298 -433 -287
rect -175 287 -129 298
rect -175 -298 -129 -287
rect 129 287 175 298
rect 129 -298 175 -287
rect 433 287 479 298
rect 433 -298 479 -287
rect 737 287 783 298
rect 737 -298 783 -287
rect -706 -379 -695 -333
rect -521 -379 -510 -333
rect -402 -379 -391 -333
rect -217 -379 -206 -333
rect -98 -379 -87 -333
rect 87 -379 98 -333
rect 206 -379 217 -333
rect 391 -379 402 -333
rect 510 -379 521 -333
rect 695 -379 706 -333
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 3.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
