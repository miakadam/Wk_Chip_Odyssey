magic
tech gf180mcuD
magscale 1 10
timestamp 1758254207
<< nwell >>
rect -11031 3790 -9891 4430
rect -9651 2352 -9071 3524
rect -8681 3457 -7641 4077
rect -7251 2352 -6671 3524
rect -9879 887 -6443 907
rect -11199 307 -10619 887
rect -10339 307 -5983 887
rect -5703 307 -5123 887
rect -9879 287 -6443 307
<< pwell >>
rect -8681 2637 -7641 3257
rect -7101 2324 -7061 2350
rect -6953 2324 -6913 2344
rect -9651 1552 -9071 2324
rect -7251 1552 -6671 2324
rect -10017 -869 -6305 -49
rect -6681 -1207 -6601 -1085
rect -10379 -4003 -5943 -1207
<< nmos >>
rect -10831 3370 -10771 3540
rect -10661 3370 -10601 3540
rect -10491 3370 -10431 3540
rect -10321 3370 -10261 3540
rect -10151 3370 -10091 3540
rect -8431 2847 -8351 3047
rect -7971 2847 -7891 3047
rect -9401 1714 -9321 2114
rect -7001 1714 -6921 2114
rect -9767 -659 -9567 -259
rect -9463 -659 -9263 -259
rect -9159 -659 -8959 -259
rect -8855 -659 -8655 -259
rect -8551 -659 -8351 -259
rect -7971 -659 -7771 -259
rect -7667 -659 -7467 -259
rect -7363 -659 -7163 -259
rect -7059 -659 -6859 -259
rect -6755 -659 -6555 -259
rect -9933 -2044 -9733 -1744
rect -9629 -2044 -9429 -1744
rect -9325 -2044 -9125 -1744
rect -9021 -2044 -8821 -1744
rect -8717 -2044 -8517 -1744
rect -8413 -2044 -8213 -1744
rect -8109 -2044 -7909 -1744
rect -7805 -2044 -7605 -1744
rect -7501 -2044 -7301 -1744
rect -7197 -2044 -6997 -1744
rect -6893 -2044 -6693 -1744
rect -6589 -2044 -6389 -1744
rect -9933 -3007 -9733 -2707
rect -9629 -3007 -9429 -2707
rect -9325 -3007 -9125 -2707
rect -9021 -3007 -8821 -2707
rect -8717 -3007 -8517 -2707
rect -8413 -3007 -8213 -2707
rect -8109 -3007 -7909 -2707
rect -7805 -3007 -7605 -2707
rect -7501 -3007 -7301 -2707
rect -7197 -3007 -6997 -2707
rect -6893 -3007 -6693 -2707
rect -6589 -3007 -6389 -2707
rect -8385 -3793 -8305 -3633
rect -8201 -3793 -8121 -3633
rect -8017 -3793 -7937 -3633
<< pmos >>
rect -10831 3880 -10771 4220
rect -10661 3880 -10601 4220
rect -10491 3880 -10431 4220
rect -10321 3880 -10261 4220
rect -10151 3880 -10091 4220
rect -8431 3667 -8351 3867
rect -7971 3667 -7891 3867
rect -9401 2562 -9321 3362
rect -7001 2562 -6921 3362
rect -10949 517 -10869 677
rect -10089 517 -10009 677
rect -9629 497 -9429 697
rect -9325 497 -9125 697
rect -9021 497 -8821 697
rect -8717 497 -8517 697
rect -8413 497 -8213 697
rect -8109 497 -7909 697
rect -7805 497 -7605 697
rect -7501 497 -7301 697
rect -7197 497 -6997 697
rect -6893 497 -6693 697
rect -6313 517 -6233 677
rect -5453 517 -5373 677
<< ndiff >>
rect -10931 3478 -10831 3540
rect -10931 3432 -10909 3478
rect -10863 3432 -10831 3478
rect -10931 3370 -10831 3432
rect -10771 3478 -10661 3540
rect -10771 3432 -10739 3478
rect -10693 3432 -10661 3478
rect -10771 3370 -10661 3432
rect -10601 3478 -10491 3540
rect -10601 3432 -10569 3478
rect -10523 3432 -10491 3478
rect -10601 3370 -10491 3432
rect -10431 3478 -10321 3540
rect -10431 3432 -10399 3478
rect -10353 3432 -10321 3478
rect -10431 3370 -10321 3432
rect -10261 3478 -10151 3540
rect -10261 3432 -10229 3478
rect -10183 3432 -10151 3478
rect -10261 3370 -10151 3432
rect -10091 3478 -9991 3540
rect -10091 3432 -10059 3478
rect -10013 3432 -9991 3478
rect -10091 3370 -9991 3432
rect -8519 3034 -8431 3047
rect -8519 2860 -8506 3034
rect -8460 2860 -8431 3034
rect -8519 2847 -8431 2860
rect -8351 3034 -8263 3047
rect -8351 2860 -8322 3034
rect -8276 2860 -8263 3034
rect -8351 2847 -8263 2860
rect -8059 3034 -7971 3047
rect -8059 2860 -8046 3034
rect -8000 2860 -7971 3034
rect -8059 2847 -7971 2860
rect -7891 3034 -7803 3047
rect -7891 2860 -7862 3034
rect -7816 2860 -7803 3034
rect -7891 2847 -7803 2860
rect -9489 2101 -9401 2114
rect -9489 1727 -9476 2101
rect -9430 1727 -9401 2101
rect -9489 1714 -9401 1727
rect -9321 2101 -9233 2114
rect -9321 1727 -9292 2101
rect -9246 1727 -9233 2101
rect -9321 1714 -9233 1727
rect -7089 2101 -7001 2114
rect -7089 1727 -7076 2101
rect -7030 1727 -7001 2101
rect -7089 1714 -7001 1727
rect -6921 2101 -6833 2114
rect -6921 1727 -6892 2101
rect -6846 1727 -6833 2101
rect -6921 1714 -6833 1727
rect -9855 -272 -9767 -259
rect -9855 -646 -9842 -272
rect -9796 -646 -9767 -272
rect -9855 -659 -9767 -646
rect -9567 -272 -9463 -259
rect -9567 -646 -9538 -272
rect -9492 -646 -9463 -272
rect -9567 -659 -9463 -646
rect -9263 -272 -9159 -259
rect -9263 -646 -9234 -272
rect -9188 -646 -9159 -272
rect -9263 -659 -9159 -646
rect -8959 -272 -8855 -259
rect -8959 -646 -8930 -272
rect -8884 -646 -8855 -272
rect -8959 -659 -8855 -646
rect -8655 -272 -8551 -259
rect -8655 -646 -8626 -272
rect -8580 -646 -8551 -272
rect -8655 -659 -8551 -646
rect -8351 -272 -8263 -259
rect -8351 -646 -8322 -272
rect -8276 -646 -8263 -272
rect -8351 -659 -8263 -646
rect -8059 -272 -7971 -259
rect -8059 -646 -8046 -272
rect -8000 -646 -7971 -272
rect -8059 -659 -7971 -646
rect -7771 -272 -7667 -259
rect -7771 -646 -7742 -272
rect -7696 -646 -7667 -272
rect -7771 -659 -7667 -646
rect -7467 -272 -7363 -259
rect -7467 -646 -7438 -272
rect -7392 -646 -7363 -272
rect -7467 -659 -7363 -646
rect -7163 -272 -7059 -259
rect -7163 -646 -7134 -272
rect -7088 -646 -7059 -272
rect -7163 -659 -7059 -646
rect -6859 -272 -6755 -259
rect -6859 -646 -6830 -272
rect -6784 -646 -6755 -272
rect -6859 -659 -6755 -646
rect -6555 -272 -6467 -259
rect -6555 -646 -6526 -272
rect -6480 -646 -6467 -272
rect -6555 -659 -6467 -646
rect -10021 -1757 -9933 -1744
rect -10021 -2031 -10008 -1757
rect -9962 -2031 -9933 -1757
rect -10021 -2044 -9933 -2031
rect -9733 -1757 -9629 -1744
rect -9733 -2031 -9704 -1757
rect -9658 -2031 -9629 -1757
rect -9733 -2044 -9629 -2031
rect -9429 -1757 -9325 -1744
rect -9429 -2031 -9400 -1757
rect -9354 -2031 -9325 -1757
rect -9429 -2044 -9325 -2031
rect -9125 -1757 -9021 -1744
rect -9125 -2031 -9096 -1757
rect -9050 -2031 -9021 -1757
rect -9125 -2044 -9021 -2031
rect -8821 -1757 -8717 -1744
rect -8821 -2031 -8792 -1757
rect -8746 -2031 -8717 -1757
rect -8821 -2044 -8717 -2031
rect -8517 -1757 -8413 -1744
rect -8517 -2031 -8488 -1757
rect -8442 -2031 -8413 -1757
rect -8517 -2044 -8413 -2031
rect -8213 -1757 -8109 -1744
rect -8213 -2031 -8184 -1757
rect -8138 -2031 -8109 -1757
rect -8213 -2044 -8109 -2031
rect -7909 -1757 -7805 -1744
rect -7909 -2031 -7880 -1757
rect -7834 -2031 -7805 -1757
rect -7909 -2044 -7805 -2031
rect -7605 -1757 -7501 -1744
rect -7605 -2031 -7576 -1757
rect -7530 -2031 -7501 -1757
rect -7605 -2044 -7501 -2031
rect -7301 -1757 -7197 -1744
rect -7301 -2031 -7272 -1757
rect -7226 -2031 -7197 -1757
rect -7301 -2044 -7197 -2031
rect -6997 -1757 -6893 -1744
rect -6997 -2031 -6968 -1757
rect -6922 -2031 -6893 -1757
rect -6997 -2044 -6893 -2031
rect -6693 -1757 -6589 -1744
rect -6693 -2031 -6664 -1757
rect -6618 -2031 -6589 -1757
rect -6693 -2044 -6589 -2031
rect -6389 -1757 -6301 -1744
rect -6389 -2031 -6360 -1757
rect -6314 -2031 -6301 -1757
rect -6389 -2044 -6301 -2031
rect -10021 -2720 -9933 -2707
rect -10021 -2994 -10008 -2720
rect -9962 -2994 -9933 -2720
rect -10021 -3007 -9933 -2994
rect -9733 -2720 -9629 -2707
rect -9733 -2994 -9704 -2720
rect -9658 -2994 -9629 -2720
rect -9733 -3007 -9629 -2994
rect -9429 -2720 -9325 -2707
rect -9429 -2994 -9400 -2720
rect -9354 -2994 -9325 -2720
rect -9429 -3007 -9325 -2994
rect -9125 -2720 -9021 -2707
rect -9125 -2994 -9096 -2720
rect -9050 -2994 -9021 -2720
rect -9125 -3007 -9021 -2994
rect -8821 -2720 -8717 -2707
rect -8821 -2994 -8792 -2720
rect -8746 -2994 -8717 -2720
rect -8821 -3007 -8717 -2994
rect -8517 -2720 -8413 -2707
rect -8517 -2994 -8488 -2720
rect -8442 -2994 -8413 -2720
rect -8517 -3007 -8413 -2994
rect -8213 -2720 -8109 -2707
rect -8213 -2994 -8184 -2720
rect -8138 -2994 -8109 -2720
rect -8213 -3007 -8109 -2994
rect -7909 -2720 -7805 -2707
rect -7909 -2994 -7880 -2720
rect -7834 -2994 -7805 -2720
rect -7909 -3007 -7805 -2994
rect -7605 -2720 -7501 -2707
rect -7605 -2994 -7576 -2720
rect -7530 -2994 -7501 -2720
rect -7605 -3007 -7501 -2994
rect -7301 -2720 -7197 -2707
rect -7301 -2994 -7272 -2720
rect -7226 -2994 -7197 -2720
rect -7301 -3007 -7197 -2994
rect -6997 -2720 -6893 -2707
rect -6997 -2994 -6968 -2720
rect -6922 -2994 -6893 -2720
rect -6997 -3007 -6893 -2994
rect -6693 -2720 -6589 -2707
rect -6693 -2994 -6664 -2720
rect -6618 -2994 -6589 -2720
rect -6693 -3007 -6589 -2994
rect -6389 -2720 -6301 -2707
rect -6389 -2994 -6360 -2720
rect -6314 -2994 -6301 -2720
rect -6389 -3007 -6301 -2994
rect -8473 -3646 -8385 -3633
rect -8473 -3780 -8460 -3646
rect -8414 -3780 -8385 -3646
rect -8473 -3793 -8385 -3780
rect -8305 -3646 -8201 -3633
rect -8305 -3780 -8276 -3646
rect -8230 -3780 -8201 -3646
rect -8305 -3793 -8201 -3780
rect -8121 -3646 -8017 -3633
rect -8121 -3780 -8092 -3646
rect -8046 -3780 -8017 -3646
rect -8121 -3793 -8017 -3780
rect -7937 -3646 -7849 -3633
rect -7937 -3780 -7908 -3646
rect -7862 -3780 -7849 -3646
rect -7937 -3793 -7849 -3780
<< pdiff >>
rect -10931 4167 -10831 4220
rect -10931 3933 -10909 4167
rect -10863 3933 -10831 4167
rect -10931 3880 -10831 3933
rect -10771 4192 -10661 4220
rect -10771 3958 -10739 4192
rect -10693 3958 -10661 4192
rect -10771 3880 -10661 3958
rect -10601 4167 -10491 4220
rect -10601 3933 -10569 4167
rect -10523 3933 -10491 4167
rect -10601 3880 -10491 3933
rect -10431 4192 -10321 4220
rect -10431 3958 -10399 4192
rect -10353 3958 -10321 4192
rect -10431 3880 -10321 3958
rect -10261 4167 -10151 4220
rect -10261 3933 -10229 4167
rect -10183 3933 -10151 4167
rect -10261 3880 -10151 3933
rect -10091 4167 -9991 4220
rect -10091 3933 -10059 4167
rect -10013 3933 -9991 4167
rect -10091 3880 -9991 3933
rect -8519 3854 -8431 3867
rect -8519 3680 -8506 3854
rect -8460 3680 -8431 3854
rect -8519 3667 -8431 3680
rect -8351 3854 -8263 3867
rect -8351 3680 -8322 3854
rect -8276 3680 -8263 3854
rect -8351 3667 -8263 3680
rect -8059 3854 -7971 3867
rect -8059 3680 -8046 3854
rect -8000 3680 -7971 3854
rect -8059 3667 -7971 3680
rect -7891 3854 -7803 3867
rect -7891 3680 -7862 3854
rect -7816 3680 -7803 3854
rect -7891 3667 -7803 3680
rect -9489 3349 -9401 3362
rect -9489 2575 -9476 3349
rect -9430 2575 -9401 3349
rect -9489 2562 -9401 2575
rect -9321 3349 -9233 3362
rect -9321 2575 -9292 3349
rect -9246 2575 -9233 3349
rect -9321 2562 -9233 2575
rect -7089 3349 -7001 3362
rect -7089 2575 -7076 3349
rect -7030 2575 -7001 3349
rect -7089 2562 -7001 2575
rect -6921 3349 -6833 3362
rect -6921 2575 -6892 3349
rect -6846 2575 -6833 3349
rect -6921 2562 -6833 2575
rect -11037 664 -10949 677
rect -11037 530 -11024 664
rect -10978 530 -10949 664
rect -11037 517 -10949 530
rect -10869 664 -10781 677
rect -10869 530 -10840 664
rect -10794 530 -10781 664
rect -10869 517 -10781 530
rect -10177 664 -10089 677
rect -10177 530 -10164 664
rect -10118 530 -10089 664
rect -10177 517 -10089 530
rect -10009 664 -9921 677
rect -10009 530 -9980 664
rect -9934 530 -9921 664
rect -10009 517 -9921 530
rect -9717 684 -9629 697
rect -9717 510 -9704 684
rect -9658 510 -9629 684
rect -9717 497 -9629 510
rect -9429 684 -9325 697
rect -9429 510 -9400 684
rect -9354 510 -9325 684
rect -9429 497 -9325 510
rect -9125 684 -9021 697
rect -9125 510 -9096 684
rect -9050 510 -9021 684
rect -9125 497 -9021 510
rect -8821 684 -8717 697
rect -8821 510 -8792 684
rect -8746 510 -8717 684
rect -8821 497 -8717 510
rect -8517 684 -8413 697
rect -8517 510 -8488 684
rect -8442 510 -8413 684
rect -8517 497 -8413 510
rect -8213 684 -8109 697
rect -8213 510 -8184 684
rect -8138 510 -8109 684
rect -8213 497 -8109 510
rect -7909 684 -7805 697
rect -7909 510 -7880 684
rect -7834 510 -7805 684
rect -7909 497 -7805 510
rect -7605 684 -7501 697
rect -7605 510 -7576 684
rect -7530 510 -7501 684
rect -7605 497 -7501 510
rect -7301 684 -7197 697
rect -7301 510 -7272 684
rect -7226 510 -7197 684
rect -7301 497 -7197 510
rect -6997 684 -6893 697
rect -6997 510 -6968 684
rect -6922 510 -6893 684
rect -6997 497 -6893 510
rect -6693 684 -6605 697
rect -6693 510 -6664 684
rect -6618 510 -6605 684
rect -6693 497 -6605 510
rect -6401 664 -6313 677
rect -6401 530 -6388 664
rect -6342 530 -6313 664
rect -6401 517 -6313 530
rect -6233 664 -6145 677
rect -6233 530 -6204 664
rect -6158 530 -6145 664
rect -6233 517 -6145 530
rect -5541 664 -5453 677
rect -5541 530 -5528 664
rect -5482 530 -5453 664
rect -5541 517 -5453 530
rect -5373 664 -5285 677
rect -5373 530 -5344 664
rect -5298 530 -5285 664
rect -5373 517 -5285 530
<< ndiffc >>
rect -10909 3432 -10863 3478
rect -10739 3432 -10693 3478
rect -10569 3432 -10523 3478
rect -10399 3432 -10353 3478
rect -10229 3432 -10183 3478
rect -10059 3432 -10013 3478
rect -8506 2860 -8460 3034
rect -8322 2860 -8276 3034
rect -8046 2860 -8000 3034
rect -7862 2860 -7816 3034
rect -9476 1727 -9430 2101
rect -9292 1727 -9246 2101
rect -7076 1727 -7030 2101
rect -6892 1727 -6846 2101
rect -9842 -646 -9796 -272
rect -9538 -646 -9492 -272
rect -9234 -646 -9188 -272
rect -8930 -646 -8884 -272
rect -8626 -646 -8580 -272
rect -8322 -646 -8276 -272
rect -8046 -646 -8000 -272
rect -7742 -646 -7696 -272
rect -7438 -646 -7392 -272
rect -7134 -646 -7088 -272
rect -6830 -646 -6784 -272
rect -6526 -646 -6480 -272
rect -10008 -2031 -9962 -1757
rect -9704 -2031 -9658 -1757
rect -9400 -2031 -9354 -1757
rect -9096 -2031 -9050 -1757
rect -8792 -2031 -8746 -1757
rect -8488 -2031 -8442 -1757
rect -8184 -2031 -8138 -1757
rect -7880 -2031 -7834 -1757
rect -7576 -2031 -7530 -1757
rect -7272 -2031 -7226 -1757
rect -6968 -2031 -6922 -1757
rect -6664 -2031 -6618 -1757
rect -6360 -2031 -6314 -1757
rect -10008 -2994 -9962 -2720
rect -9704 -2994 -9658 -2720
rect -9400 -2994 -9354 -2720
rect -9096 -2994 -9050 -2720
rect -8792 -2994 -8746 -2720
rect -8488 -2994 -8442 -2720
rect -8184 -2994 -8138 -2720
rect -7880 -2994 -7834 -2720
rect -7576 -2994 -7530 -2720
rect -7272 -2994 -7226 -2720
rect -6968 -2994 -6922 -2720
rect -6664 -2994 -6618 -2720
rect -6360 -2994 -6314 -2720
rect -8460 -3780 -8414 -3646
rect -8276 -3780 -8230 -3646
rect -8092 -3780 -8046 -3646
rect -7908 -3780 -7862 -3646
<< pdiffc >>
rect -10909 3933 -10863 4167
rect -10739 3958 -10693 4192
rect -10569 3933 -10523 4167
rect -10399 3958 -10353 4192
rect -10229 3933 -10183 4167
rect -10059 3933 -10013 4167
rect -8506 3680 -8460 3854
rect -8322 3680 -8276 3854
rect -8046 3680 -8000 3854
rect -7862 3680 -7816 3854
rect -9476 2575 -9430 3349
rect -9292 2575 -9246 3349
rect -7076 2575 -7030 3349
rect -6892 2575 -6846 3349
rect -11024 530 -10978 664
rect -10840 530 -10794 664
rect -10164 530 -10118 664
rect -9980 530 -9934 664
rect -9704 510 -9658 684
rect -9400 510 -9354 684
rect -9096 510 -9050 684
rect -8792 510 -8746 684
rect -8488 510 -8442 684
rect -8184 510 -8138 684
rect -7880 510 -7834 684
rect -7576 510 -7530 684
rect -7272 510 -7226 684
rect -6968 510 -6922 684
rect -6664 510 -6618 684
rect -6388 530 -6342 664
rect -6204 530 -6158 664
rect -5528 530 -5482 664
rect -5344 530 -5298 664
<< psubdiff >>
rect -10831 3278 -10681 3300
rect -10831 3232 -10779 3278
rect -10733 3232 -10681 3278
rect -10831 3210 -10681 3232
rect -10591 3278 -10441 3300
rect -10591 3232 -10539 3278
rect -10493 3232 -10441 3278
rect -10591 3210 -10441 3232
rect -10351 3278 -10201 3300
rect -10351 3232 -10299 3278
rect -10253 3232 -10201 3278
rect -10351 3210 -10201 3232
rect -10111 3278 -9961 3300
rect -10111 3232 -10059 3278
rect -10013 3232 -9961 3278
rect -10111 3210 -9961 3232
rect -8657 3161 -7665 3233
rect -8657 3117 -8585 3161
rect -8657 2777 -8644 3117
rect -8598 2777 -8585 3117
rect -8197 3117 -8125 3161
rect -8657 2733 -8585 2777
rect -8197 2777 -8184 3117
rect -8138 2777 -8125 3117
rect -7737 3117 -7665 3161
rect -8197 2733 -8125 2777
rect -7737 2777 -7724 3117
rect -7678 2777 -7665 3117
rect -7737 2733 -7665 2777
rect -8657 2661 -7665 2733
rect -9627 2228 -9095 2300
rect -9627 1648 -9555 2228
rect -9167 1648 -9095 2228
rect -9627 1635 -9095 1648
rect -9627 1589 -9511 1635
rect -9211 1589 -9095 1635
rect -9627 1576 -9095 1589
rect -7227 2228 -6695 2300
rect -7227 1648 -7155 2228
rect -6767 1648 -6695 2228
rect -7227 1635 -6695 1648
rect -7227 1589 -7111 1635
rect -6811 1589 -6695 1635
rect -7227 1576 -6695 1589
rect -9993 -145 -6329 -73
rect -9993 -189 -9921 -145
rect -9993 -729 -9980 -189
rect -9934 -729 -9921 -189
rect -8197 -189 -8125 -145
rect -9993 -773 -9921 -729
rect -8197 -729 -8184 -189
rect -8138 -729 -8125 -189
rect -6401 -189 -6329 -145
rect -8197 -773 -8125 -729
rect -6401 -729 -6388 -189
rect -6342 -729 -6329 -189
rect -6401 -773 -6329 -729
rect -9993 -845 -6329 -773
rect -10354 -1304 -5968 -1232
rect -10354 -1403 -10154 -1304
rect -10354 -1903 -10304 -1403
rect -10204 -1903 -10154 -1403
rect -6168 -1403 -5968 -1304
rect -10354 -2848 -10154 -1903
rect -6168 -1903 -6118 -1403
rect -6018 -1903 -5968 -1403
rect -10354 -3348 -10304 -2848
rect -10204 -3348 -10154 -2848
rect -6168 -2848 -5968 -1903
rect -10354 -3447 -10154 -3348
rect -6168 -3348 -6118 -2848
rect -6018 -3348 -5968 -2848
rect -6168 -3447 -5968 -3348
rect -10354 -3519 -5968 -3447
rect -8611 -3563 -8539 -3519
rect -8611 -3863 -8598 -3563
rect -8552 -3863 -8539 -3563
rect -7783 -3563 -7711 -3519
rect -8611 -3907 -8539 -3863
rect -7783 -3863 -7770 -3563
rect -7724 -3863 -7711 -3563
rect -7783 -3907 -7711 -3863
rect -8611 -3979 -7711 -3907
<< nsubdiff >>
rect -10831 4358 -10681 4380
rect -10831 4312 -10779 4358
rect -10733 4312 -10681 4358
rect -10831 4290 -10681 4312
rect -10591 4358 -10441 4380
rect -10591 4312 -10539 4358
rect -10493 4312 -10441 4358
rect -10591 4290 -10441 4312
rect -10351 4358 -10201 4380
rect -10351 4312 -10299 4358
rect -10253 4312 -10201 4358
rect -10351 4290 -10201 4312
rect -10111 4358 -9961 4380
rect -10111 4312 -10059 4358
rect -10013 4312 -9961 4358
rect -10111 4290 -9961 4312
rect -8657 3981 -7665 4053
rect -8657 3937 -8585 3981
rect -8657 3597 -8644 3937
rect -8598 3597 -8585 3937
rect -8197 3937 -8125 3981
rect -8657 3553 -8585 3597
rect -8197 3597 -8184 3937
rect -8138 3597 -8125 3937
rect -7737 3937 -7665 3981
rect -8197 3553 -8125 3597
rect -7737 3597 -7724 3937
rect -7678 3597 -7665 3937
rect -7737 3553 -7665 3597
rect -9627 3487 -9095 3500
rect -9627 3441 -9511 3487
rect -9211 3441 -9095 3487
rect -8657 3481 -7665 3553
rect -7227 3487 -6695 3500
rect -9627 3428 -9095 3441
rect -9627 2448 -9555 3428
rect -9167 2448 -9095 3428
rect -7227 3441 -7111 3487
rect -6811 3441 -6695 3487
rect -7227 3428 -6695 3441
rect -9627 2376 -9095 2448
rect -7227 2448 -7155 3428
rect -6767 2448 -6695 3428
rect -7227 2376 -6695 2448
rect -9855 863 -6467 883
rect -11175 791 -10643 863
rect -11175 747 -11103 791
rect -11175 447 -11162 747
rect -11116 447 -11103 747
rect -10715 747 -10643 791
rect -11175 403 -11103 447
rect -10715 447 -10702 747
rect -10656 447 -10643 747
rect -10715 403 -10643 447
rect -11175 331 -10643 403
rect -10315 811 -6007 863
rect -10315 791 -9783 811
rect -10315 747 -10243 791
rect -10315 447 -10302 747
rect -10256 447 -10243 747
rect -9855 767 -9783 791
rect -6539 791 -6007 811
rect -10315 403 -10243 447
rect -9855 427 -9842 767
rect -9796 427 -9783 767
rect -6539 767 -6467 791
rect -9855 403 -9783 427
rect -6539 427 -6526 767
rect -6480 427 -6467 767
rect -6079 747 -6007 791
rect -10315 383 -9783 403
rect -6539 403 -6467 427
rect -6079 447 -6066 747
rect -6020 447 -6007 747
rect -6079 403 -6007 447
rect -6539 383 -6007 403
rect -10315 331 -6007 383
rect -5679 791 -5147 863
rect -5679 747 -5607 791
rect -5679 447 -5666 747
rect -5620 447 -5607 747
rect -5219 747 -5147 791
rect -5679 403 -5607 447
rect -5219 447 -5206 747
rect -5160 447 -5147 747
rect -5219 403 -5147 447
rect -5679 331 -5147 403
rect -9855 311 -6467 331
<< psubdiffcont >>
rect -10779 3232 -10733 3278
rect -10539 3232 -10493 3278
rect -10299 3232 -10253 3278
rect -10059 3232 -10013 3278
rect -8644 2777 -8598 3117
rect -8184 2777 -8138 3117
rect -7724 2777 -7678 3117
rect -9511 1589 -9211 1635
rect -7111 1589 -6811 1635
rect -9980 -729 -9934 -189
rect -8184 -729 -8138 -189
rect -6388 -729 -6342 -189
rect -10304 -1903 -10204 -1403
rect -6118 -1903 -6018 -1403
rect -10304 -3348 -10204 -2848
rect -6118 -3348 -6018 -2848
rect -8598 -3863 -8552 -3563
rect -7770 -3863 -7724 -3563
<< nsubdiffcont >>
rect -10779 4312 -10733 4358
rect -10539 4312 -10493 4358
rect -10299 4312 -10253 4358
rect -10059 4312 -10013 4358
rect -8644 3597 -8598 3937
rect -8184 3597 -8138 3937
rect -7724 3597 -7678 3937
rect -9511 3441 -9211 3487
rect -7111 3441 -6811 3487
rect -11162 447 -11116 747
rect -10702 447 -10656 747
rect -10302 447 -10256 747
rect -9842 427 -9796 767
rect -6526 427 -6480 767
rect -6066 447 -6020 747
rect -5666 447 -5620 747
rect -5206 447 -5160 747
<< polysilicon >>
rect -10831 4220 -10771 4270
rect -10661 4220 -10601 4270
rect -10491 4220 -10431 4270
rect -10321 4220 -10261 4270
rect -10151 4220 -10091 4270
rect -10831 3860 -10771 3880
rect -10661 3860 -10601 3880
rect -10491 3860 -10431 3880
rect -10321 3860 -10261 3880
rect -10831 3850 -10261 3860
rect -10831 3823 -10201 3850
rect -10831 3800 -10274 3823
rect -10661 3620 -10601 3800
rect -10321 3777 -10274 3800
rect -10228 3777 -10201 3823
rect -10321 3750 -10201 3777
rect -10321 3620 -10261 3750
rect -10151 3700 -10091 3880
rect -10831 3560 -10261 3620
rect -10211 3673 -10091 3700
rect -10211 3627 -10184 3673
rect -10138 3627 -10091 3673
rect -10211 3600 -10091 3627
rect -10831 3540 -10771 3560
rect -10661 3540 -10601 3560
rect -10491 3540 -10431 3560
rect -10321 3540 -10261 3560
rect -10151 3540 -10091 3600
rect -8431 3946 -8351 3959
rect -8431 3900 -8418 3946
rect -8364 3900 -8351 3946
rect -8431 3867 -8351 3900
rect -8431 3634 -8351 3667
rect -8431 3588 -8418 3634
rect -8364 3588 -8351 3634
rect -8431 3575 -8351 3588
rect -7971 3946 -7891 3959
rect -7971 3900 -7958 3946
rect -7904 3900 -7891 3946
rect -7971 3867 -7891 3900
rect -7971 3634 -7891 3667
rect -7971 3588 -7958 3634
rect -7904 3588 -7891 3634
rect -7971 3575 -7891 3588
rect -10831 3320 -10771 3370
rect -10661 3320 -10601 3370
rect -10491 3320 -10431 3370
rect -10321 3320 -10261 3370
rect -10151 3320 -10091 3370
rect -9401 3362 -9321 3406
rect -9401 2529 -9321 2562
rect -9401 2483 -9388 2529
rect -9334 2483 -9321 2529
rect -9401 2470 -9321 2483
rect -8431 3126 -8351 3139
rect -8431 3080 -8418 3126
rect -8364 3080 -8351 3126
rect -8431 3047 -8351 3080
rect -8431 2814 -8351 2847
rect -8431 2768 -8418 2814
rect -8364 2768 -8351 2814
rect -8431 2755 -8351 2768
rect -7971 3126 -7891 3139
rect -7971 3080 -7958 3126
rect -7904 3080 -7891 3126
rect -7971 3047 -7891 3080
rect -7971 2814 -7891 2847
rect -7971 2768 -7958 2814
rect -7904 2768 -7891 2814
rect -7971 2755 -7891 2768
rect -7001 3362 -6921 3406
rect -7001 2529 -6921 2562
rect -7001 2483 -6988 2529
rect -6934 2483 -6921 2529
rect -7001 2470 -6921 2483
rect -9401 2193 -9321 2206
rect -9401 2147 -9388 2193
rect -9334 2147 -9321 2193
rect -9401 2114 -9321 2147
rect -9401 1670 -9321 1714
rect -7001 2193 -6921 2206
rect -7001 2147 -6988 2193
rect -6934 2147 -6921 2193
rect -7001 2114 -6921 2147
rect -7001 1670 -6921 1714
rect -10949 756 -10869 769
rect -10949 710 -10936 756
rect -10882 710 -10869 756
rect -10949 677 -10869 710
rect -10949 484 -10869 517
rect -10949 438 -10936 484
rect -10882 438 -10869 484
rect -10949 425 -10869 438
rect -10089 756 -10009 769
rect -10089 710 -10076 756
rect -10022 710 -10009 756
rect -10089 677 -10009 710
rect -10089 484 -10009 517
rect -10089 438 -10076 484
rect -10022 438 -10009 484
rect -10089 425 -10009 438
rect -9629 776 -9429 789
rect -9629 730 -9616 776
rect -9442 730 -9429 776
rect -9629 697 -9429 730
rect -9325 776 -9125 789
rect -9325 730 -9312 776
rect -9138 730 -9125 776
rect -9325 697 -9125 730
rect -9021 776 -8821 789
rect -9021 730 -9008 776
rect -8834 730 -8821 776
rect -9021 697 -8821 730
rect -8717 776 -8517 789
rect -8717 730 -8704 776
rect -8530 730 -8517 776
rect -8717 697 -8517 730
rect -8413 776 -8213 789
rect -8413 730 -8400 776
rect -8226 730 -8213 776
rect -8413 697 -8213 730
rect -8109 776 -7909 789
rect -8109 730 -8096 776
rect -7922 730 -7909 776
rect -8109 697 -7909 730
rect -7805 776 -7605 789
rect -7805 730 -7792 776
rect -7618 730 -7605 776
rect -7805 697 -7605 730
rect -7501 776 -7301 789
rect -7501 730 -7488 776
rect -7314 730 -7301 776
rect -7501 697 -7301 730
rect -7197 776 -6997 789
rect -7197 730 -7184 776
rect -7010 730 -6997 776
rect -7197 697 -6997 730
rect -6893 776 -6693 789
rect -6893 730 -6880 776
rect -6706 730 -6693 776
rect -6893 697 -6693 730
rect -9629 464 -9429 497
rect -9629 418 -9616 464
rect -9442 418 -9429 464
rect -9629 405 -9429 418
rect -9325 464 -9125 497
rect -9325 418 -9312 464
rect -9138 418 -9125 464
rect -9325 405 -9125 418
rect -9021 464 -8821 497
rect -9021 418 -9008 464
rect -8834 418 -8821 464
rect -9021 405 -8821 418
rect -8717 464 -8517 497
rect -8717 418 -8704 464
rect -8530 418 -8517 464
rect -8717 405 -8517 418
rect -8413 464 -8213 497
rect -8413 418 -8400 464
rect -8226 418 -8213 464
rect -8413 405 -8213 418
rect -8109 464 -7909 497
rect -8109 418 -8096 464
rect -7922 418 -7909 464
rect -8109 405 -7909 418
rect -7805 464 -7605 497
rect -7805 418 -7792 464
rect -7618 418 -7605 464
rect -7805 405 -7605 418
rect -7501 464 -7301 497
rect -7501 418 -7488 464
rect -7314 418 -7301 464
rect -7501 405 -7301 418
rect -7197 464 -6997 497
rect -7197 418 -7184 464
rect -7010 418 -6997 464
rect -7197 405 -6997 418
rect -6893 464 -6693 497
rect -6893 418 -6880 464
rect -6706 418 -6693 464
rect -6893 405 -6693 418
rect -6313 756 -6233 769
rect -6313 710 -6300 756
rect -6246 710 -6233 756
rect -6313 677 -6233 710
rect -6313 484 -6233 517
rect -6313 438 -6300 484
rect -6246 438 -6233 484
rect -6313 425 -6233 438
rect -5453 756 -5373 769
rect -5453 710 -5440 756
rect -5386 710 -5373 756
rect -5453 677 -5373 710
rect -5453 484 -5373 517
rect -5453 438 -5440 484
rect -5386 438 -5373 484
rect -5453 425 -5373 438
rect -9767 -180 -9567 -167
rect -9767 -226 -9754 -180
rect -9580 -226 -9567 -180
rect -9767 -259 -9567 -226
rect -9463 -180 -9263 -167
rect -9463 -226 -9450 -180
rect -9276 -226 -9263 -180
rect -9463 -259 -9263 -226
rect -9159 -180 -8959 -167
rect -9159 -226 -9146 -180
rect -8972 -226 -8959 -180
rect -9159 -259 -8959 -226
rect -8855 -180 -8655 -167
rect -8855 -226 -8842 -180
rect -8668 -226 -8655 -180
rect -8855 -259 -8655 -226
rect -8551 -180 -8351 -167
rect -8551 -226 -8538 -180
rect -8364 -226 -8351 -180
rect -8551 -259 -8351 -226
rect -9767 -692 -9567 -659
rect -9767 -738 -9754 -692
rect -9580 -738 -9567 -692
rect -9767 -751 -9567 -738
rect -9463 -692 -9263 -659
rect -9463 -738 -9450 -692
rect -9276 -738 -9263 -692
rect -9463 -751 -9263 -738
rect -9159 -692 -8959 -659
rect -9159 -738 -9146 -692
rect -8972 -738 -8959 -692
rect -9159 -751 -8959 -738
rect -8855 -692 -8655 -659
rect -8855 -738 -8842 -692
rect -8668 -738 -8655 -692
rect -8855 -751 -8655 -738
rect -8551 -692 -8351 -659
rect -8551 -738 -8538 -692
rect -8364 -738 -8351 -692
rect -8551 -751 -8351 -738
rect -7971 -180 -7771 -167
rect -7971 -226 -7958 -180
rect -7784 -226 -7771 -180
rect -7971 -259 -7771 -226
rect -7667 -180 -7467 -167
rect -7667 -226 -7654 -180
rect -7480 -226 -7467 -180
rect -7667 -259 -7467 -226
rect -7363 -180 -7163 -167
rect -7363 -226 -7350 -180
rect -7176 -226 -7163 -180
rect -7363 -259 -7163 -226
rect -7059 -180 -6859 -167
rect -7059 -226 -7046 -180
rect -6872 -226 -6859 -180
rect -7059 -259 -6859 -226
rect -6755 -180 -6555 -167
rect -6755 -226 -6742 -180
rect -6568 -226 -6555 -180
rect -6755 -259 -6555 -226
rect -7971 -692 -7771 -659
rect -7971 -738 -7958 -692
rect -7784 -738 -7771 -692
rect -7971 -751 -7771 -738
rect -7667 -692 -7467 -659
rect -7667 -738 -7654 -692
rect -7480 -738 -7467 -692
rect -7667 -751 -7467 -738
rect -7363 -692 -7163 -659
rect -7363 -738 -7350 -692
rect -7176 -738 -7163 -692
rect -7363 -751 -7163 -738
rect -7059 -692 -6859 -659
rect -7059 -738 -7046 -692
rect -6872 -738 -6859 -692
rect -7059 -751 -6859 -738
rect -6755 -692 -6555 -659
rect -6755 -738 -6742 -692
rect -6568 -738 -6555 -692
rect -6755 -751 -6555 -738
rect -9933 -1665 -9733 -1652
rect -9933 -1711 -9920 -1665
rect -9746 -1711 -9733 -1665
rect -9933 -1744 -9733 -1711
rect -9629 -1665 -9429 -1652
rect -9629 -1711 -9616 -1665
rect -9442 -1711 -9429 -1665
rect -9629 -1744 -9429 -1711
rect -9325 -1665 -9125 -1652
rect -9325 -1711 -9312 -1665
rect -9138 -1711 -9125 -1665
rect -9325 -1744 -9125 -1711
rect -9021 -1665 -8821 -1652
rect -9021 -1711 -9008 -1665
rect -8834 -1711 -8821 -1665
rect -9021 -1744 -8821 -1711
rect -8717 -1665 -8517 -1652
rect -8717 -1711 -8704 -1665
rect -8530 -1711 -8517 -1665
rect -8717 -1744 -8517 -1711
rect -8413 -1665 -8213 -1652
rect -8413 -1711 -8400 -1665
rect -8226 -1711 -8213 -1665
rect -8413 -1744 -8213 -1711
rect -8109 -1665 -7909 -1652
rect -8109 -1711 -8096 -1665
rect -7922 -1711 -7909 -1665
rect -8109 -1744 -7909 -1711
rect -7805 -1665 -7605 -1652
rect -7805 -1711 -7792 -1665
rect -7618 -1711 -7605 -1665
rect -7805 -1744 -7605 -1711
rect -7501 -1665 -7301 -1652
rect -7501 -1711 -7488 -1665
rect -7314 -1711 -7301 -1665
rect -7501 -1744 -7301 -1711
rect -7197 -1665 -6997 -1652
rect -7197 -1711 -7184 -1665
rect -7010 -1711 -6997 -1665
rect -7197 -1744 -6997 -1711
rect -6893 -1665 -6693 -1652
rect -6893 -1711 -6880 -1665
rect -6706 -1711 -6693 -1665
rect -6893 -1744 -6693 -1711
rect -6589 -1665 -6389 -1652
rect -6589 -1711 -6576 -1665
rect -6402 -1711 -6389 -1665
rect -6589 -1744 -6389 -1711
rect -9933 -2077 -9733 -2044
rect -9933 -2123 -9920 -2077
rect -9746 -2123 -9733 -2077
rect -9933 -2136 -9733 -2123
rect -9629 -2077 -9429 -2044
rect -9629 -2123 -9616 -2077
rect -9442 -2123 -9429 -2077
rect -9629 -2136 -9429 -2123
rect -9325 -2077 -9125 -2044
rect -9325 -2123 -9312 -2077
rect -9138 -2123 -9125 -2077
rect -9325 -2136 -9125 -2123
rect -9021 -2077 -8821 -2044
rect -9021 -2123 -9008 -2077
rect -8834 -2123 -8821 -2077
rect -9021 -2136 -8821 -2123
rect -8717 -2077 -8517 -2044
rect -8717 -2123 -8704 -2077
rect -8530 -2123 -8517 -2077
rect -8717 -2136 -8517 -2123
rect -8413 -2077 -8213 -2044
rect -8413 -2123 -8400 -2077
rect -8226 -2123 -8213 -2077
rect -8413 -2136 -8213 -2123
rect -8109 -2077 -7909 -2044
rect -8109 -2123 -8096 -2077
rect -7922 -2123 -7909 -2077
rect -8109 -2136 -7909 -2123
rect -7805 -2077 -7605 -2044
rect -7805 -2123 -7792 -2077
rect -7618 -2123 -7605 -2077
rect -7805 -2136 -7605 -2123
rect -7501 -2077 -7301 -2044
rect -7501 -2123 -7488 -2077
rect -7314 -2123 -7301 -2077
rect -7501 -2136 -7301 -2123
rect -7197 -2077 -6997 -2044
rect -7197 -2123 -7184 -2077
rect -7010 -2123 -6997 -2077
rect -7197 -2136 -6997 -2123
rect -6893 -2077 -6693 -2044
rect -6893 -2123 -6880 -2077
rect -6706 -2123 -6693 -2077
rect -6893 -2136 -6693 -2123
rect -6589 -2077 -6389 -2044
rect -6589 -2123 -6576 -2077
rect -6402 -2123 -6389 -2077
rect -6589 -2136 -6389 -2123
rect -9271 -2138 -9181 -2136
rect -9933 -2628 -9733 -2615
rect -9933 -2674 -9920 -2628
rect -9746 -2674 -9733 -2628
rect -9933 -2707 -9733 -2674
rect -9629 -2628 -9429 -2615
rect -9629 -2674 -9616 -2628
rect -9442 -2674 -9429 -2628
rect -9629 -2707 -9429 -2674
rect -9325 -2628 -9125 -2615
rect -9325 -2674 -9312 -2628
rect -9138 -2674 -9125 -2628
rect -9325 -2707 -9125 -2674
rect -9021 -2628 -8821 -2615
rect -9021 -2674 -9008 -2628
rect -8834 -2674 -8821 -2628
rect -9021 -2707 -8821 -2674
rect -8717 -2628 -8517 -2615
rect -8717 -2674 -8704 -2628
rect -8530 -2674 -8517 -2628
rect -8717 -2707 -8517 -2674
rect -8413 -2628 -8213 -2615
rect -8413 -2674 -8400 -2628
rect -8226 -2674 -8213 -2628
rect -8413 -2707 -8213 -2674
rect -8109 -2628 -7909 -2615
rect -8109 -2674 -8096 -2628
rect -7922 -2674 -7909 -2628
rect -8109 -2707 -7909 -2674
rect -7805 -2628 -7605 -2615
rect -7805 -2674 -7792 -2628
rect -7618 -2674 -7605 -2628
rect -7805 -2707 -7605 -2674
rect -7501 -2628 -7301 -2615
rect -7501 -2674 -7488 -2628
rect -7314 -2674 -7301 -2628
rect -7501 -2707 -7301 -2674
rect -7197 -2628 -6997 -2615
rect -7197 -2674 -7184 -2628
rect -7010 -2674 -6997 -2628
rect -7197 -2707 -6997 -2674
rect -6893 -2628 -6693 -2615
rect -6893 -2674 -6880 -2628
rect -6706 -2674 -6693 -2628
rect -6893 -2707 -6693 -2674
rect -6589 -2628 -6389 -2615
rect -6589 -2674 -6576 -2628
rect -6402 -2674 -6389 -2628
rect -6589 -2707 -6389 -2674
rect -9933 -3040 -9733 -3007
rect -9933 -3086 -9920 -3040
rect -9746 -3086 -9733 -3040
rect -9933 -3099 -9733 -3086
rect -9629 -3040 -9429 -3007
rect -9629 -3086 -9616 -3040
rect -9442 -3086 -9429 -3040
rect -9629 -3099 -9429 -3086
rect -9325 -3040 -9125 -3007
rect -9325 -3086 -9312 -3040
rect -9138 -3086 -9125 -3040
rect -9325 -3099 -9125 -3086
rect -9021 -3040 -8821 -3007
rect -9021 -3086 -9008 -3040
rect -8834 -3086 -8821 -3040
rect -9021 -3099 -8821 -3086
rect -8717 -3040 -8517 -3007
rect -8717 -3086 -8704 -3040
rect -8530 -3086 -8517 -3040
rect -8717 -3099 -8517 -3086
rect -8413 -3040 -8213 -3007
rect -8413 -3086 -8400 -3040
rect -8226 -3086 -8213 -3040
rect -8413 -3099 -8213 -3086
rect -8109 -3040 -7909 -3007
rect -8109 -3086 -8096 -3040
rect -7922 -3086 -7909 -3040
rect -8109 -3099 -7909 -3086
rect -7805 -3040 -7605 -3007
rect -7805 -3086 -7792 -3040
rect -7618 -3086 -7605 -3040
rect -7805 -3099 -7605 -3086
rect -7501 -3040 -7301 -3007
rect -7501 -3086 -7488 -3040
rect -7314 -3086 -7301 -3040
rect -7501 -3099 -7301 -3086
rect -7197 -3040 -6997 -3007
rect -7197 -3086 -7184 -3040
rect -7010 -3086 -6997 -3040
rect -7197 -3099 -6997 -3086
rect -6893 -3040 -6693 -3007
rect -6893 -3086 -6880 -3040
rect -6706 -3086 -6693 -3040
rect -6893 -3099 -6693 -3086
rect -6589 -3040 -6389 -3007
rect -6589 -3086 -6576 -3040
rect -6402 -3086 -6389 -3040
rect -6589 -3099 -6389 -3086
rect -8385 -3554 -8305 -3541
rect -8385 -3600 -8372 -3554
rect -8318 -3600 -8305 -3554
rect -8385 -3633 -8305 -3600
rect -8201 -3554 -8121 -3541
rect -8201 -3600 -8188 -3554
rect -8134 -3600 -8121 -3554
rect -8201 -3633 -8121 -3600
rect -8017 -3554 -7937 -3541
rect -8017 -3600 -8004 -3554
rect -7950 -3600 -7937 -3554
rect -8017 -3633 -7937 -3600
rect -8385 -3826 -8305 -3793
rect -8385 -3872 -8372 -3826
rect -8318 -3872 -8305 -3826
rect -8385 -3885 -8305 -3872
rect -8201 -3826 -8121 -3793
rect -8201 -3872 -8188 -3826
rect -8134 -3872 -8121 -3826
rect -8201 -3885 -8121 -3872
rect -8017 -3826 -7937 -3793
rect -8017 -3872 -8004 -3826
rect -7950 -3872 -7937 -3826
rect -8017 -3885 -7937 -3872
<< polycontact >>
rect -10274 3777 -10228 3823
rect -10184 3627 -10138 3673
rect -8418 3900 -8364 3946
rect -8418 3588 -8364 3634
rect -7958 3900 -7904 3946
rect -7958 3588 -7904 3634
rect -9388 2483 -9334 2529
rect -8418 3080 -8364 3126
rect -8418 2768 -8364 2814
rect -7958 3080 -7904 3126
rect -7958 2768 -7904 2814
rect -6988 2483 -6934 2529
rect -9388 2147 -9334 2193
rect -6988 2147 -6934 2193
rect -10936 710 -10882 756
rect -10936 438 -10882 484
rect -10076 710 -10022 756
rect -10076 438 -10022 484
rect -9616 730 -9442 776
rect -9312 730 -9138 776
rect -9008 730 -8834 776
rect -8704 730 -8530 776
rect -8400 730 -8226 776
rect -8096 730 -7922 776
rect -7792 730 -7618 776
rect -7488 730 -7314 776
rect -7184 730 -7010 776
rect -6880 730 -6706 776
rect -9616 418 -9442 464
rect -9312 418 -9138 464
rect -9008 418 -8834 464
rect -8704 418 -8530 464
rect -8400 418 -8226 464
rect -8096 418 -7922 464
rect -7792 418 -7618 464
rect -7488 418 -7314 464
rect -7184 418 -7010 464
rect -6880 418 -6706 464
rect -6300 710 -6246 756
rect -6300 438 -6246 484
rect -5440 710 -5386 756
rect -5440 438 -5386 484
rect -9754 -226 -9580 -180
rect -9450 -226 -9276 -180
rect -9146 -226 -8972 -180
rect -8842 -226 -8668 -180
rect -8538 -226 -8364 -180
rect -9754 -738 -9580 -692
rect -9450 -738 -9276 -692
rect -9146 -738 -8972 -692
rect -8842 -738 -8668 -692
rect -8538 -738 -8364 -692
rect -7958 -226 -7784 -180
rect -7654 -226 -7480 -180
rect -7350 -226 -7176 -180
rect -7046 -226 -6872 -180
rect -6742 -226 -6568 -180
rect -7958 -738 -7784 -692
rect -7654 -738 -7480 -692
rect -7350 -738 -7176 -692
rect -7046 -738 -6872 -692
rect -6742 -738 -6568 -692
rect -9920 -1711 -9746 -1665
rect -9616 -1711 -9442 -1665
rect -9312 -1711 -9138 -1665
rect -9008 -1711 -8834 -1665
rect -8704 -1711 -8530 -1665
rect -8400 -1711 -8226 -1665
rect -8096 -1711 -7922 -1665
rect -7792 -1711 -7618 -1665
rect -7488 -1711 -7314 -1665
rect -7184 -1711 -7010 -1665
rect -6880 -1711 -6706 -1665
rect -6576 -1711 -6402 -1665
rect -9920 -2123 -9746 -2077
rect -9616 -2123 -9442 -2077
rect -9312 -2123 -9138 -2077
rect -9008 -2123 -8834 -2077
rect -8704 -2123 -8530 -2077
rect -8400 -2123 -8226 -2077
rect -8096 -2123 -7922 -2077
rect -7792 -2123 -7618 -2077
rect -7488 -2123 -7314 -2077
rect -7184 -2123 -7010 -2077
rect -6880 -2123 -6706 -2077
rect -6576 -2123 -6402 -2077
rect -9920 -2674 -9746 -2628
rect -9616 -2674 -9442 -2628
rect -9312 -2674 -9138 -2628
rect -9008 -2674 -8834 -2628
rect -8704 -2674 -8530 -2628
rect -8400 -2674 -8226 -2628
rect -8096 -2674 -7922 -2628
rect -7792 -2674 -7618 -2628
rect -7488 -2674 -7314 -2628
rect -7184 -2674 -7010 -2628
rect -6880 -2674 -6706 -2628
rect -6576 -2674 -6402 -2628
rect -9920 -3086 -9746 -3040
rect -9616 -3086 -9442 -3040
rect -9312 -3086 -9138 -3040
rect -9008 -3086 -8834 -3040
rect -8704 -3086 -8530 -3040
rect -8400 -3086 -8226 -3040
rect -8096 -3086 -7922 -3040
rect -7792 -3086 -7618 -3040
rect -7488 -3086 -7314 -3040
rect -7184 -3086 -7010 -3040
rect -6880 -3086 -6706 -3040
rect -6576 -3086 -6402 -3040
rect -8372 -3600 -8318 -3554
rect -8188 -3600 -8134 -3554
rect -8004 -3600 -7950 -3554
rect -8372 -3872 -8318 -3826
rect -8188 -3872 -8134 -3826
rect -8004 -3872 -7950 -3826
<< metal1 >>
rect -13117 11494 -13047 11506
rect -13117 11438 -13105 11494
rect -13049 11438 -12960 11494
rect -13117 11426 -13047 11438
rect -12442 5434 -2430 5477
rect -12442 5134 -4454 5434
rect -2454 5134 -2430 5434
rect -12442 5097 -2430 5134
rect -13680 3940 -13603 3954
rect -12380 3940 -12294 3954
rect -13680 3939 -12366 3940
rect -13680 3881 -13665 3939
rect -13607 3881 -12366 3939
rect -13680 3880 -12366 3881
rect -12306 3880 -12294 3940
rect -13680 3867 -13603 3880
rect -12380 3866 -12294 3880
rect -12085 2179 -12007 5097
rect -10476 4430 -10396 5097
rect -11031 4358 -9891 4430
rect -11031 4312 -10779 4358
rect -10733 4312 -10539 4358
rect -10493 4312 -10299 4358
rect -10253 4312 -10059 4358
rect -10013 4312 -9891 4358
rect -11031 4290 -9891 4312
rect -10911 4167 -10861 4290
rect -10911 3933 -10909 4167
rect -10863 3933 -10861 4167
rect -10741 4192 -10691 4220
rect -10741 3958 -10739 4192
rect -10693 3958 -10691 4192
rect -10741 3940 -10691 3958
rect -10571 4167 -10521 4290
rect -10911 3880 -10861 3933
rect -10771 3936 -10671 3940
rect -10771 3884 -10747 3936
rect -10695 3884 -10671 3936
rect -10771 3880 -10671 3884
rect -10571 3933 -10569 4167
rect -10523 3933 -10521 4167
rect -10571 3880 -10521 3933
rect -10401 4192 -10351 4220
rect -10401 3958 -10399 4192
rect -10353 3958 -10351 4192
rect -10741 3830 -10691 3880
rect -10401 3830 -10351 3958
rect -10231 4167 -10181 4290
rect -10231 3933 -10229 4167
rect -10183 3933 -10181 4167
rect -10231 3880 -10181 3933
rect -10061 4167 -10011 4220
rect -10061 3933 -10059 4167
rect -10013 3933 -10011 4167
rect -10061 3830 -10011 3933
rect -10741 3770 -10351 3830
rect -10301 3823 -10011 3830
rect -10301 3777 -10274 3823
rect -10228 3777 -10011 3823
rect -10301 3770 -10011 3777
rect -10741 3650 -10691 3770
rect -10401 3650 -10351 3770
rect -10741 3590 -10351 3650
rect -10211 3676 -10111 3680
rect -10211 3624 -10187 3676
rect -10135 3624 -10111 3676
rect -10211 3620 -10111 3624
rect -10911 3478 -10861 3540
rect -10911 3432 -10909 3478
rect -10863 3432 -10861 3478
rect -10911 3300 -10861 3432
rect -10741 3478 -10691 3590
rect -10741 3432 -10739 3478
rect -10693 3432 -10691 3478
rect -10741 3370 -10691 3432
rect -10571 3478 -10521 3540
rect -10571 3432 -10569 3478
rect -10523 3432 -10521 3478
rect -10571 3300 -10521 3432
rect -10401 3478 -10351 3590
rect -10401 3432 -10399 3478
rect -10353 3432 -10351 3478
rect -10401 3370 -10351 3432
rect -10231 3478 -10181 3540
rect -10231 3432 -10229 3478
rect -10183 3432 -10181 3478
rect -10231 3300 -10181 3432
rect -10061 3478 -10011 3770
rect -9396 3487 -9316 5097
rect -8216 4157 -8136 5097
rect -8644 4077 -7678 4157
rect -8644 3937 -8598 4077
rect -8429 3946 -8353 3979
rect -8429 3900 -8418 3946
rect -8364 3900 -8353 3946
rect -8184 3937 -8138 3948
rect -8506 3854 -8460 3865
rect -8598 3680 -8506 3854
rect -8322 3854 -8276 3865
rect -8339 3795 -8322 3805
rect -8276 3795 -8259 3805
rect -8339 3739 -8327 3795
rect -8271 3739 -8259 3795
rect -8339 3729 -8322 3739
rect -8506 3669 -8460 3680
rect -8276 3729 -8259 3739
rect -8322 3669 -8276 3680
rect -8644 3586 -8598 3597
rect -8429 3588 -8418 3634
rect -8364 3588 -8353 3634
rect -7969 3946 -7893 3979
rect -7969 3900 -7958 3946
rect -7904 3900 -7893 3946
rect -7724 3937 -7678 4077
rect -8046 3854 -8000 3865
rect -8063 3795 -8046 3805
rect -7862 3854 -7816 3865
rect -8000 3795 -7983 3805
rect -8063 3739 -8051 3795
rect -7995 3739 -7983 3795
rect -8063 3729 -8046 3739
rect -8000 3729 -7983 3739
rect -8046 3669 -8000 3680
rect -7816 3680 -7724 3854
rect -7862 3669 -7816 3680
rect -9522 3486 -9511 3487
rect -10061 3432 -10059 3478
rect -10013 3432 -10011 3478
rect -9593 3441 -9511 3486
rect -9211 3486 -9200 3487
rect -9211 3441 -9143 3486
rect -9593 3434 -9143 3441
rect -10061 3370 -10011 3432
rect -9585 3426 -9143 3434
rect -9485 3349 -9425 3426
rect -8419 3401 -8363 3588
rect -8184 3586 -8138 3597
rect -7969 3588 -7958 3634
rect -7904 3588 -7893 3634
rect -8201 3537 -8131 3539
rect -7959 3537 -7903 3588
rect -7724 3586 -7678 3597
rect -8201 3481 -8189 3537
rect -8133 3481 -7903 3537
rect -6996 3487 -6916 5097
rect -7122 3486 -7111 3487
rect -8201 3479 -8131 3481
rect -7179 3441 -7111 3486
rect -6811 3486 -6800 3487
rect -6811 3441 -6729 3486
rect -7179 3434 -6729 3441
rect -7179 3426 -6737 3434
rect -8419 3399 -8121 3401
rect -11031 3278 -9891 3300
rect -11031 3232 -10779 3278
rect -10733 3232 -10539 3278
rect -10493 3232 -10299 3278
rect -10253 3232 -10059 3278
rect -10013 3232 -9891 3278
rect -11031 3160 -9891 3232
rect -9485 3202 -9476 3349
rect -9430 3202 -9425 3349
rect -9292 3358 -9246 3360
rect -9292 3349 -9209 3358
rect -9476 2564 -9430 2575
rect -9246 2575 -9209 3349
rect -8419 3343 -8189 3399
rect -8133 3343 -8121 3399
rect -7076 3358 -7030 3360
rect -8419 3341 -8121 3343
rect -7113 3349 -7030 3358
rect -9292 2564 -9209 2575
rect -9399 2502 -9388 2529
rect -9401 2483 -9388 2502
rect -9334 2502 -9323 2529
rect -9334 2483 -9321 2502
rect -10531 2376 -10437 2388
rect -9401 2376 -9321 2483
rect -10531 2300 -10519 2376
rect -10439 2300 -9321 2376
rect -10531 2298 -10437 2300
rect -9401 2193 -9321 2300
rect -9401 2182 -9388 2193
rect -12086 1978 -12006 2179
rect -9399 2147 -9388 2182
rect -9334 2182 -9321 2193
rect -9273 2446 -9209 2564
rect -8644 3117 -8598 3128
rect -8429 3126 -8353 3159
rect -8429 3080 -8418 3126
rect -8364 3080 -8353 3126
rect -8184 3117 -8138 3128
rect -8506 3034 -8460 3045
rect -8598 2860 -8506 3034
rect -8322 3034 -8276 3045
rect -8339 2975 -8322 2985
rect -8276 2975 -8259 2985
rect -8339 2919 -8327 2975
rect -8271 2919 -8259 2975
rect -8339 2909 -8322 2919
rect -8506 2849 -8460 2860
rect -8276 2909 -8259 2919
rect -8322 2849 -8276 2860
rect -8429 2809 -8418 2814
rect -8644 2637 -8598 2777
rect -8431 2799 -8418 2809
rect -8364 2809 -8353 2814
rect -8364 2799 -8351 2809
rect -8431 2743 -8419 2799
rect -8363 2743 -8351 2799
rect -7969 3126 -7893 3159
rect -7969 3080 -7958 3126
rect -7904 3080 -7893 3126
rect -7724 3117 -7678 3128
rect -8046 3034 -8000 3045
rect -8063 2975 -8046 2985
rect -7862 3034 -7816 3045
rect -8000 2975 -7983 2985
rect -8063 2919 -8051 2975
rect -7995 2919 -7983 2975
rect -8063 2909 -8046 2919
rect -8000 2909 -7983 2919
rect -8046 2849 -8000 2860
rect -7816 2860 -7724 3034
rect -7862 2849 -7816 2860
rect -7969 2809 -7958 2814
rect -8184 2766 -8138 2777
rect -7971 2799 -7958 2809
rect -7904 2809 -7893 2814
rect -7904 2799 -7891 2809
rect -8431 2733 -8351 2743
rect -7971 2743 -7959 2799
rect -7903 2743 -7891 2799
rect -7971 2733 -7891 2743
rect -7724 2637 -7678 2777
rect -8644 2557 -7678 2637
rect -7113 2575 -7076 3349
rect -6897 3349 -6837 3426
rect -6897 3202 -6892 3349
rect -7113 2564 -7030 2575
rect -6846 3202 -6837 3349
rect -6892 2564 -6846 2575
rect -9273 2376 -9205 2446
rect -8421 2376 -8349 2378
rect -9273 2300 -8419 2376
rect -8363 2300 -8349 2376
rect -9334 2147 -9323 2182
rect -9273 2112 -9205 2300
rect -8421 2288 -8349 2300
rect -9476 2101 -9430 2112
rect -12103 1961 -11990 1978
rect -12103 1883 -12086 1961
rect -12006 1883 -11990 1961
rect -12103 1872 -11990 1883
rect -9477 1727 -9476 1810
rect -9292 2101 -9205 2112
rect -9430 1727 -9429 1810
rect -9477 1643 -9429 1727
rect -9246 1730 -9205 2101
rect -9292 1716 -9246 1727
rect -11227 1640 -8625 1643
rect -8205 1640 -8139 2557
rect -7113 2446 -7049 2564
rect -6999 2502 -6988 2529
rect -7973 2376 -7901 2378
rect -7117 2376 -7049 2446
rect -7973 2300 -7959 2376
rect -7903 2300 -7049 2376
rect -7973 2288 -7901 2300
rect -7117 2112 -7049 2300
rect -7001 2483 -6988 2502
rect -6934 2502 -6923 2529
rect -6934 2483 -6921 2502
rect -7001 2376 -6921 2483
rect -5895 2376 -5791 2388
rect -7001 2300 -5883 2376
rect -5803 2300 -5791 2376
rect -7001 2193 -6921 2300
rect -5895 2298 -5791 2300
rect -5675 2197 -5597 5097
rect -7001 2182 -6988 2193
rect -6999 2147 -6988 2182
rect -6934 2182 -6921 2193
rect -6934 2147 -6923 2182
rect -7117 2101 -7030 2112
rect -7117 1730 -7076 2101
rect -6892 2101 -6846 2112
rect -7076 1716 -7030 1727
rect -6893 1727 -6892 1810
rect -5676 2027 -5596 2197
rect -5696 1847 -5576 2027
rect -6846 1727 -6845 1810
rect -5696 1787 -5676 1847
rect -5596 1787 -5576 1847
rect -6893 1643 -6845 1727
rect -4791 1649 -4633 1664
rect -4791 1643 -4764 1649
rect -6914 1642 -4764 1643
rect -7131 1640 -4764 1642
rect -11700 1635 -4764 1640
rect -11700 1589 -9511 1635
rect -9211 1589 -7111 1635
rect -6811 1589 -4764 1635
rect -11700 1580 -4764 1589
rect -11700 1551 -11497 1580
rect -11227 1578 -4764 1580
rect -11700 1462 -11642 1551
rect -11551 1462 -11497 1551
rect -4791 1542 -4764 1578
rect -4655 1542 -4633 1649
rect -4791 1531 -4633 1542
rect -11700 1433 -11497 1462
rect -11391 1432 -11287 1446
rect -5035 1432 -4931 1444
rect -11391 1356 -11379 1432
rect -11299 1356 -5023 1432
rect -4943 1356 -4931 1432
rect -11391 1346 -11287 1356
rect -11162 747 -11116 758
rect -10947 756 -10871 1356
rect -10947 710 -10936 756
rect -10882 710 -10871 756
rect -10702 747 -10656 758
rect -11024 666 -10978 675
rect -10840 666 -10794 675
rect -11116 664 -10961 666
rect -11116 530 -11029 664
rect -10973 530 -10961 664
rect -11116 528 -10961 530
rect -10857 664 -10777 666
rect -10857 530 -10845 664
rect -10789 530 -10777 664
rect -10857 528 -10777 530
rect -10719 664 -10702 666
rect -10302 747 -10256 758
rect -10656 664 -10639 666
rect -10719 530 -10707 664
rect -10651 530 -10639 664
rect -10719 528 -10702 530
rect -11024 519 -10978 528
rect -10840 519 -10794 528
rect -11162 436 -11116 447
rect -10947 438 -10936 484
rect -10882 438 -10871 484
rect -10947 408 -10871 438
rect -10656 528 -10639 530
rect -10702 436 -10656 447
rect -10087 756 -10011 1356
rect -10087 710 -10076 756
rect -10022 710 -10011 756
rect -9842 767 -9796 778
rect -9323 776 -8823 832
rect -10164 666 -10118 675
rect -9980 666 -9934 675
rect -10256 664 -10101 666
rect -10256 530 -10169 664
rect -10113 530 -10101 664
rect -10256 528 -10101 530
rect -9997 664 -9917 666
rect -9997 530 -9985 664
rect -9929 530 -9917 664
rect -9997 528 -9917 530
rect -9859 664 -9842 666
rect -9627 730 -9616 776
rect -9442 730 -9431 776
rect -9323 730 -9312 776
rect -9138 730 -9127 776
rect -9019 730 -9008 776
rect -8834 730 -8823 776
rect -8715 776 -8215 832
rect -8715 730 -8704 776
rect -8530 730 -8519 776
rect -8411 730 -8400 776
rect -8226 730 -8215 776
rect -8107 776 -7607 832
rect -8107 730 -8096 776
rect -7922 730 -7911 776
rect -7803 730 -7792 776
rect -7618 730 -7607 776
rect -7499 776 -6999 832
rect -7499 730 -7488 776
rect -7314 730 -7303 776
rect -7195 730 -7184 776
rect -7010 730 -6999 776
rect -6891 730 -6880 776
rect -6706 730 -6695 776
rect -6526 767 -6480 778
rect -9704 684 -9658 695
rect -9796 664 -9779 666
rect -9859 530 -9847 664
rect -9791 530 -9779 664
rect -9859 528 -9842 530
rect -10164 519 -10118 528
rect -9980 519 -9934 528
rect -10302 436 -10256 447
rect -10087 438 -10076 484
rect -10022 438 -10011 484
rect -10087 408 -10011 438
rect -9796 528 -9779 530
rect -9400 684 -9354 695
rect -9417 677 -9400 679
rect -9096 684 -9050 695
rect -9354 677 -9337 679
rect -9417 533 -9405 677
rect -9349 533 -9337 677
rect -9417 531 -9400 533
rect -9704 499 -9658 510
rect -9354 531 -9337 533
rect -9113 576 -9096 586
rect -8792 684 -8746 695
rect -8809 677 -8792 679
rect -8488 684 -8442 695
rect -8746 677 -8729 679
rect -9050 576 -9033 586
rect -9113 520 -9101 576
rect -9045 520 -9033 576
rect -8809 533 -8797 677
rect -8741 533 -8729 677
rect -8809 531 -8792 533
rect -9113 510 -9096 520
rect -9050 510 -9033 520
rect -8746 531 -8729 533
rect -8505 576 -8488 586
rect -8184 684 -8138 695
rect -8201 677 -8184 679
rect -7880 684 -7834 695
rect -8138 677 -8121 679
rect -8442 576 -8425 586
rect -8505 520 -8493 576
rect -8437 520 -8425 576
rect -8201 533 -8189 677
rect -8133 533 -8121 677
rect -8201 531 -8184 533
rect -8505 510 -8488 520
rect -8442 510 -8425 520
rect -8138 531 -8121 533
rect -7897 576 -7880 586
rect -7576 684 -7530 695
rect -7593 677 -7576 679
rect -7272 684 -7226 695
rect -7530 677 -7513 679
rect -7834 576 -7817 586
rect -7897 520 -7885 576
rect -7829 520 -7817 576
rect -7593 533 -7581 677
rect -7525 533 -7513 677
rect -7593 531 -7576 533
rect -7897 510 -7880 520
rect -7834 510 -7817 520
rect -7530 531 -7513 533
rect -7289 576 -7272 586
rect -6968 684 -6922 695
rect -6985 677 -6968 679
rect -6664 684 -6618 695
rect -6922 677 -6905 679
rect -7226 576 -7209 586
rect -7289 520 -7277 576
rect -7221 520 -7209 576
rect -6985 533 -6973 677
rect -6917 533 -6905 677
rect -6985 531 -6968 533
rect -7289 510 -7272 520
rect -7226 510 -7209 520
rect -6922 531 -6905 533
rect -9400 499 -9354 510
rect -9096 499 -9050 510
rect -8792 499 -8746 510
rect -8488 499 -8442 510
rect -8184 499 -8138 510
rect -7880 499 -7834 510
rect -7576 499 -7530 510
rect -7272 499 -7226 510
rect -6968 499 -6922 510
rect -6543 664 -6526 666
rect -6311 756 -6235 1356
rect -6311 710 -6300 756
rect -6246 710 -6235 756
rect -6066 747 -6020 758
rect -6388 666 -6342 675
rect -6204 666 -6158 675
rect -6480 664 -6463 666
rect -6543 530 -6531 664
rect -6475 530 -6463 664
rect -6543 528 -6526 530
rect -6664 499 -6618 510
rect -8310 469 -8230 479
rect -8310 464 -8298 469
rect -8242 464 -8230 469
rect -8092 469 -8012 479
rect -8092 464 -8080 469
rect -8024 464 -8012 469
rect -9842 416 -9796 427
rect -9627 418 -9616 464
rect -9442 418 -9431 464
rect -9323 418 -9312 464
rect -9138 453 -9127 464
rect -9019 453 -9008 464
rect -9138 418 -9008 453
rect -8834 418 -8823 464
rect -8715 418 -8704 464
rect -8530 418 -8519 464
rect -8411 418 -8400 464
rect -8226 418 -8215 464
rect -8107 418 -8096 464
rect -7922 418 -7911 464
rect -7803 418 -7792 464
rect -7618 418 -7607 464
rect -7499 418 -7488 464
rect -7314 453 -7303 464
rect -7195 453 -7184 464
rect -7314 418 -7184 453
rect -7010 418 -6999 464
rect -6891 418 -6880 464
rect -6706 418 -6695 464
rect -6480 528 -6463 530
rect -6405 664 -6325 666
rect -6405 530 -6393 664
rect -6337 530 -6325 664
rect -6405 528 -6325 530
rect -6221 664 -6066 666
rect -6221 530 -6209 664
rect -6153 530 -6066 664
rect -6221 528 -6066 530
rect -6388 519 -6342 528
rect -6204 519 -6158 528
rect -9263 407 -8823 418
rect -8310 413 -8298 418
rect -8242 413 -8230 418
rect -10531 161 -10427 173
rect -10009 161 -9905 171
rect -9263 161 -9159 407
rect -8310 403 -8230 413
rect -8092 413 -8080 418
rect -8024 413 -8012 418
rect -8092 403 -8012 413
rect -7499 407 -7059 418
rect -6526 416 -6480 427
rect -6311 438 -6300 484
rect -6246 438 -6235 484
rect -6311 408 -6235 438
rect -5666 747 -5620 758
rect -5683 664 -5666 666
rect -5451 756 -5375 1356
rect -5035 1344 -4931 1356
rect -5451 710 -5440 756
rect -5386 710 -5375 756
rect -5206 747 -5160 758
rect -5528 666 -5482 675
rect -5344 666 -5298 675
rect -5620 664 -5603 666
rect -5683 530 -5671 664
rect -5615 530 -5603 664
rect -5683 528 -5666 530
rect -6066 436 -6020 447
rect -5620 528 -5603 530
rect -5545 664 -5465 666
rect -5545 530 -5533 664
rect -5477 530 -5465 664
rect -5545 528 -5465 530
rect -5361 664 -5206 666
rect -5361 530 -5349 664
rect -5293 530 -5206 664
rect -5361 528 -5206 530
rect -5528 519 -5482 528
rect -5344 519 -5298 528
rect -5666 436 -5620 447
rect -5451 438 -5440 484
rect -5386 438 -5375 484
rect -5451 408 -5375 438
rect -5206 436 -5160 447
rect -8655 161 -8415 169
rect -10531 77 -10519 161
rect -10439 77 -9997 161
rect -9917 159 -8415 161
rect -9917 79 -9251 159
rect -9171 79 -8643 159
rect -8563 79 -8505 159
rect -8425 79 -8415 159
rect -9917 77 -8415 79
rect -10531 67 -10427 77
rect -10009 67 -9905 77
rect -9263 65 -9159 77
rect -8655 65 -8415 77
rect -7909 161 -7667 169
rect -7163 161 -7059 407
rect -6417 161 -6313 171
rect -5895 161 -5791 171
rect -7909 159 -6405 161
rect -7909 79 -7897 159
rect -7817 79 -7759 159
rect -7679 79 -7151 159
rect -7071 79 -6405 159
rect -7909 77 -6405 79
rect -6325 77 -5883 161
rect -5803 77 -5791 161
rect -7909 65 -7667 77
rect -7163 66 -7059 77
rect -6417 67 -6313 77
rect -5895 67 -5791 77
rect -9461 -135 -8657 -120
rect -9980 -189 -9934 -178
rect -9461 -180 -8842 -135
rect -8762 -180 -8657 -135
rect -7665 -135 -6861 -120
rect -9997 -585 -9980 -575
rect -9765 -226 -9754 -180
rect -9580 -226 -9569 -180
rect -9461 -226 -9450 -180
rect -9276 -226 -9265 -180
rect -9157 -226 -9146 -180
rect -8972 -226 -8961 -180
rect -8853 -226 -8842 -180
rect -8668 -226 -8657 -180
rect -8549 -226 -8538 -180
rect -8364 -226 -8353 -180
rect -8184 -189 -8138 -178
rect -7665 -180 -7560 -135
rect -7480 -180 -6861 -135
rect -9842 -272 -9796 -261
rect -9934 -585 -9917 -575
rect -9997 -729 -9985 -585
rect -9929 -729 -9917 -585
rect -9538 -272 -9492 -261
rect -9555 -495 -9538 -493
rect -9234 -272 -9188 -261
rect -9251 -279 -9234 -277
rect -8930 -272 -8884 -261
rect -9188 -279 -9171 -277
rect -9251 -423 -9239 -279
rect -9183 -423 -9171 -279
rect -9251 -425 -9234 -423
rect -9492 -495 -9475 -493
rect -9555 -639 -9543 -495
rect -9487 -639 -9475 -495
rect -9555 -641 -9538 -639
rect -9842 -657 -9796 -646
rect -9492 -641 -9475 -639
rect -9538 -657 -9492 -646
rect -9188 -425 -9171 -423
rect -8947 -495 -8930 -493
rect -8626 -272 -8580 -261
rect -8643 -279 -8626 -277
rect -8322 -272 -8276 -261
rect -8580 -279 -8563 -277
rect -8643 -423 -8631 -279
rect -8575 -423 -8563 -279
rect -8643 -425 -8626 -423
rect -8884 -495 -8867 -493
rect -8947 -639 -8935 -495
rect -8879 -639 -8867 -495
rect -8947 -641 -8930 -639
rect -9234 -657 -9188 -646
rect -8884 -641 -8867 -639
rect -8930 -657 -8884 -646
rect -8580 -425 -8563 -423
rect -8626 -657 -8580 -646
rect -8322 -657 -8276 -646
rect -9997 -740 -9917 -729
rect -9765 -738 -9754 -692
rect -9580 -738 -9569 -692
rect -9461 -738 -9450 -692
rect -9276 -738 -9265 -692
rect -9157 -738 -9146 -692
rect -8972 -738 -8961 -692
rect -8853 -738 -8842 -692
rect -8668 -738 -8657 -692
rect -8549 -738 -8538 -692
rect -8364 -738 -8353 -692
rect -7969 -226 -7958 -180
rect -7784 -226 -7773 -180
rect -7665 -226 -7654 -180
rect -7480 -226 -7469 -180
rect -7361 -226 -7350 -180
rect -7176 -226 -7165 -180
rect -7057 -226 -7046 -180
rect -6872 -226 -6861 -180
rect -6753 -226 -6742 -180
rect -6568 -226 -6557 -180
rect -6388 -189 -6342 -178
rect -8046 -272 -8000 -261
rect -7742 -272 -7696 -261
rect -7759 -279 -7742 -277
rect -7438 -272 -7392 -261
rect -7696 -279 -7679 -277
rect -7759 -423 -7747 -279
rect -7691 -423 -7679 -279
rect -7759 -425 -7742 -423
rect -8046 -657 -8000 -646
rect -7696 -425 -7679 -423
rect -7455 -495 -7438 -493
rect -7134 -272 -7088 -261
rect -7151 -279 -7134 -277
rect -6830 -272 -6784 -261
rect -7088 -279 -7071 -277
rect -7151 -423 -7139 -279
rect -7083 -423 -7071 -279
rect -7151 -425 -7134 -423
rect -7392 -495 -7375 -493
rect -7455 -639 -7443 -495
rect -7387 -639 -7375 -495
rect -7455 -641 -7438 -639
rect -7742 -657 -7696 -646
rect -7392 -641 -7375 -639
rect -7438 -657 -7392 -646
rect -7088 -425 -7071 -423
rect -6847 -495 -6830 -493
rect -6526 -272 -6480 -261
rect -6784 -495 -6767 -493
rect -6847 -639 -6835 -495
rect -6779 -639 -6767 -495
rect -6847 -641 -6830 -639
rect -7134 -657 -7088 -646
rect -6784 -641 -6767 -639
rect -6830 -657 -6784 -646
rect -6526 -657 -6480 -646
rect -6405 -585 -6388 -575
rect -6342 -585 -6325 -575
rect -8184 -740 -8138 -729
rect -7969 -738 -7958 -692
rect -7784 -738 -7773 -692
rect -7665 -738 -7654 -692
rect -7480 -738 -7469 -692
rect -7361 -738 -7350 -692
rect -7176 -738 -7165 -692
rect -7057 -738 -7046 -692
rect -6872 -738 -6861 -692
rect -6753 -738 -6742 -692
rect -6568 -738 -6557 -692
rect -6405 -729 -6393 -585
rect -6337 -729 -6325 -585
rect -6405 -740 -6325 -729
rect -10869 -1005 -10765 -995
rect -9733 -1005 -9629 -993
rect -9567 -1005 -9463 -993
rect -8959 -1005 -8855 -993
rect -10869 -1085 -10857 -1005
rect -10777 -1085 -9721 -1005
rect -9641 -1085 -9555 -1005
rect -9475 -1085 -8947 -1005
rect -8867 -1085 -8855 -1005
rect -10869 -1095 -10765 -1085
rect -9733 -1097 -9629 -1085
rect -9567 -1097 -9463 -1085
rect -8959 -1097 -8855 -1085
rect -7467 -1005 -7363 -993
rect -6859 -1005 -6755 -993
rect -6693 -1005 -6589 -993
rect -5557 -1005 -5453 -995
rect -7467 -1085 -7455 -1005
rect -7375 -1085 -6847 -1005
rect -6767 -1085 -6681 -1005
rect -6601 -1085 -5545 -1005
rect -5465 -1085 -5453 -1005
rect -7467 -1097 -7363 -1085
rect -6859 -1097 -6755 -1085
rect -6693 -1097 -6589 -1085
rect -5557 -1095 -5453 -1085
rect -10315 -1403 -10193 -1392
rect -10315 -1903 -10304 -1403
rect -10204 -1903 -10193 -1403
rect -6129 -1403 -6007 -1392
rect -9931 -1711 -9920 -1665
rect -9746 -1711 -9735 -1665
rect -9627 -1711 -9616 -1665
rect -9442 -1711 -9431 -1665
rect -9323 -1711 -9312 -1665
rect -9138 -1711 -9127 -1665
rect -9019 -1711 -9008 -1665
rect -8834 -1711 -8823 -1665
rect -8715 -1711 -8704 -1665
rect -8530 -1711 -8519 -1665
rect -8411 -1711 -8400 -1665
rect -8226 -1711 -8215 -1665
rect -8107 -1711 -8096 -1665
rect -7922 -1711 -7911 -1665
rect -7803 -1711 -7792 -1665
rect -7618 -1711 -7607 -1665
rect -7499 -1711 -7488 -1665
rect -7314 -1711 -7303 -1665
rect -7195 -1711 -7184 -1665
rect -7010 -1711 -6999 -1665
rect -6891 -1711 -6880 -1665
rect -6706 -1711 -6695 -1665
rect -6587 -1711 -6576 -1665
rect -6402 -1711 -6391 -1665
rect -10315 -1914 -10193 -1903
rect -10008 -1757 -9962 -1746
rect -9704 -1757 -9658 -1746
rect -9721 -1813 -9704 -1803
rect -9400 -1757 -9354 -1746
rect -9658 -1813 -9641 -1803
rect -9721 -1974 -9709 -1813
rect -9653 -1974 -9641 -1813
rect -9721 -1984 -9704 -1974
rect -10008 -2042 -9962 -2031
rect -9658 -1984 -9641 -1974
rect -9417 -1861 -9400 -1851
rect -9096 -1757 -9050 -1746
rect -9113 -1777 -9096 -1767
rect -8792 -1757 -8746 -1746
rect -9050 -1777 -9033 -1767
rect -9354 -1861 -9337 -1851
rect -9704 -2042 -9658 -2031
rect -9417 -2022 -9405 -1861
rect -9349 -2022 -9337 -1861
rect -9113 -1994 -9101 -1777
rect -9045 -1994 -9033 -1777
rect -9113 -2002 -9096 -1994
rect -9417 -2031 -9400 -2022
rect -9354 -2031 -9337 -2022
rect -9417 -2032 -9337 -2031
rect -9050 -2002 -9033 -1994
rect -8809 -1861 -8792 -1851
rect -8488 -1757 -8442 -1746
rect -8505 -1777 -8488 -1767
rect -8184 -1757 -8138 -1746
rect -8442 -1777 -8425 -1767
rect -8505 -1833 -8493 -1777
rect -8437 -1833 -8425 -1777
rect -8505 -1843 -8488 -1833
rect -8746 -1861 -8729 -1851
rect -9400 -2042 -9354 -2032
rect -9096 -2042 -9050 -2031
rect -8809 -2022 -8797 -1861
rect -8741 -2022 -8729 -1861
rect -8809 -2031 -8792 -2022
rect -8746 -2031 -8729 -2022
rect -8809 -2032 -8729 -2031
rect -8442 -1843 -8425 -1833
rect -8792 -2042 -8746 -2032
rect -8488 -2042 -8442 -2031
rect -8201 -1861 -8184 -1851
rect -7880 -1757 -7834 -1746
rect -7897 -1777 -7880 -1767
rect -7576 -1757 -7530 -1746
rect -7834 -1777 -7817 -1767
rect -7897 -1833 -7885 -1777
rect -7829 -1833 -7817 -1777
rect -7897 -1843 -7880 -1833
rect -8138 -1861 -8121 -1851
rect -8201 -2022 -8189 -1861
rect -8133 -2022 -8121 -1861
rect -8201 -2031 -8184 -2022
rect -8138 -2031 -8121 -2022
rect -8201 -2032 -8121 -2031
rect -7834 -1843 -7817 -1833
rect -8184 -2042 -8138 -2032
rect -7880 -2042 -7834 -2031
rect -7593 -1861 -7576 -1851
rect -7272 -1757 -7226 -1746
rect -7289 -1777 -7272 -1767
rect -6968 -1757 -6922 -1746
rect -7226 -1777 -7209 -1767
rect -7530 -1861 -7513 -1851
rect -7593 -2022 -7581 -1861
rect -7525 -2022 -7513 -1861
rect -7593 -2031 -7576 -2022
rect -7530 -2031 -7513 -2022
rect -7593 -2032 -7513 -2031
rect -7289 -2022 -7277 -1777
rect -7221 -2022 -7209 -1777
rect -7289 -2031 -7272 -2022
rect -7226 -2031 -7209 -2022
rect -7289 -2032 -7209 -2031
rect -6985 -1861 -6968 -1851
rect -6664 -1757 -6618 -1746
rect -6681 -1813 -6664 -1803
rect -6360 -1757 -6314 -1746
rect -6618 -1813 -6601 -1803
rect -6922 -1861 -6905 -1851
rect -6985 -2022 -6973 -1861
rect -6917 -2022 -6905 -1861
rect -6681 -1974 -6669 -1813
rect -6613 -1974 -6601 -1813
rect -6681 -1984 -6664 -1974
rect -6985 -2031 -6968 -2022
rect -6922 -2031 -6905 -2022
rect -6985 -2032 -6905 -2031
rect -6618 -1984 -6601 -1974
rect -7576 -2042 -7530 -2032
rect -7272 -2042 -7226 -2032
rect -6968 -2042 -6922 -2032
rect -6664 -2042 -6618 -2031
rect -6129 -1903 -6118 -1403
rect -6018 -1903 -6007 -1403
rect -6129 -1914 -6007 -1903
rect -6360 -2042 -6314 -2031
rect -9276 -2077 -9261 -2068
rect -9191 -2077 -9176 -2068
rect -8971 -2077 -8956 -2068
rect -8886 -2077 -8871 -2068
rect -8061 -2077 -8046 -2068
rect -7976 -2077 -7961 -2068
rect -7756 -2077 -7741 -2068
rect -7671 -2077 -7656 -2068
rect -6841 -2077 -6826 -2068
rect -6756 -2077 -6741 -2068
rect -9931 -2123 -9920 -2077
rect -9746 -2123 -9735 -2077
rect -9627 -2123 -9616 -2077
rect -9442 -2123 -9431 -2077
rect -9323 -2123 -9312 -2077
rect -9138 -2123 -9127 -2077
rect -9019 -2123 -9008 -2077
rect -8834 -2123 -8823 -2077
rect -8715 -2123 -8704 -2077
rect -8530 -2123 -8519 -2077
rect -8411 -2123 -8400 -2077
rect -8226 -2123 -8215 -2077
rect -8107 -2123 -8096 -2077
rect -7922 -2123 -7911 -2077
rect -7803 -2123 -7792 -2077
rect -7618 -2123 -7607 -2077
rect -7499 -2123 -7488 -2077
rect -7314 -2123 -7303 -2077
rect -7195 -2123 -7184 -2077
rect -7010 -2123 -6999 -2077
rect -6891 -2123 -6880 -2077
rect -6706 -2123 -6695 -2077
rect -6587 -2123 -6576 -2077
rect -6402 -2123 -6391 -2077
rect -13722 -2178 -13632 -2166
rect -9626 -2178 -9431 -2123
rect -9321 -2128 -9261 -2123
rect -9191 -2128 -9136 -2123
rect -8971 -2128 -8956 -2123
rect -8886 -2128 -8871 -2123
rect -8716 -2178 -8521 -2123
rect -8411 -2178 -8216 -2123
rect -8061 -2128 -8046 -2123
rect -7976 -2128 -7961 -2123
rect -7756 -2128 -7741 -2123
rect -7671 -2128 -7656 -2123
rect -7496 -2178 -7301 -2123
rect -7196 -2178 -7001 -2123
rect -6841 -2128 -6826 -2123
rect -6756 -2128 -6741 -2123
rect -13722 -2179 -6031 -2178
rect -13722 -2252 -13707 -2179
rect -13634 -2193 -6031 -2179
rect -13634 -2226 -6511 -2193
rect -13634 -2252 -9254 -2226
rect -13722 -2253 -9254 -2252
rect -13722 -2266 -13632 -2253
rect -9266 -2282 -9254 -2253
rect -9198 -2253 -8039 -2226
rect -9198 -2282 -9186 -2253
rect -9266 -2292 -9186 -2282
rect -8051 -2282 -8039 -2253
rect -7983 -2253 -6511 -2226
rect -6451 -2253 -6031 -2193
rect -7983 -2282 -7971 -2253
rect -8051 -2292 -7971 -2282
rect -8961 -2474 -8881 -2464
rect -13717 -2503 -13627 -2491
rect -8961 -2503 -8949 -2474
rect -13717 -2504 -8949 -2503
rect -13717 -2577 -13704 -2504
rect -13631 -2530 -8949 -2504
rect -8893 -2503 -8881 -2474
rect -7746 -2474 -7666 -2464
rect -7746 -2503 -7734 -2474
rect -8893 -2530 -7734 -2503
rect -7678 -2503 -7666 -2474
rect -7678 -2530 -6251 -2503
rect -13631 -2563 -6251 -2530
rect -6191 -2563 -6031 -2503
rect -13631 -2577 -6031 -2563
rect -13717 -2578 -6031 -2577
rect -13717 -2591 -13627 -2578
rect -9626 -2628 -9431 -2578
rect -8716 -2628 -8521 -2578
rect -8411 -2628 -8216 -2578
rect -7501 -2628 -7306 -2578
rect -7196 -2628 -7001 -2578
rect -9931 -2674 -9920 -2628
rect -9746 -2674 -9735 -2628
rect -9627 -2674 -9616 -2628
rect -9442 -2674 -9431 -2628
rect -9323 -2674 -9312 -2628
rect -9138 -2674 -9127 -2628
rect -9019 -2674 -9008 -2628
rect -8834 -2674 -8823 -2628
rect -8715 -2674 -8704 -2628
rect -8530 -2674 -8519 -2628
rect -8411 -2674 -8400 -2628
rect -8226 -2674 -8215 -2628
rect -8107 -2674 -8096 -2628
rect -7922 -2674 -7911 -2628
rect -7803 -2674 -7792 -2628
rect -7618 -2674 -7607 -2628
rect -7499 -2674 -7488 -2628
rect -7314 -2674 -7303 -2628
rect -7195 -2674 -7184 -2628
rect -7010 -2674 -6999 -2628
rect -6891 -2674 -6880 -2628
rect -6706 -2674 -6695 -2628
rect -6587 -2674 -6576 -2628
rect -6402 -2674 -6391 -2628
rect -9276 -2688 -9261 -2674
rect -9191 -2688 -9176 -2674
rect -8971 -2688 -8956 -2674
rect -8886 -2688 -8871 -2674
rect -8061 -2688 -8046 -2674
rect -7976 -2688 -7961 -2674
rect -7756 -2688 -7741 -2674
rect -7671 -2688 -7656 -2674
rect -6841 -2688 -6826 -2674
rect -6756 -2688 -6741 -2674
rect -10008 -2720 -9962 -2709
rect -10315 -2848 -10193 -2837
rect -10315 -3348 -10304 -2848
rect -10204 -3348 -10193 -2848
rect -9704 -2720 -9658 -2709
rect -9721 -2921 -9704 -2911
rect -9400 -2720 -9354 -2709
rect -9417 -2732 -9400 -2722
rect -9096 -2720 -9050 -2709
rect -9354 -2732 -9337 -2722
rect -9417 -2893 -9405 -2732
rect -9349 -2893 -9337 -2732
rect -9417 -2903 -9400 -2893
rect -9658 -2921 -9641 -2911
rect -9721 -2977 -9709 -2921
rect -9653 -2977 -9641 -2921
rect -9721 -2987 -9704 -2977
rect -10008 -3005 -9962 -2994
rect -9658 -2987 -9641 -2977
rect -9704 -3005 -9658 -2994
rect -9354 -2903 -9337 -2893
rect -9113 -2766 -9096 -2756
rect -8792 -2720 -8746 -2709
rect -8809 -2732 -8792 -2722
rect -8488 -2720 -8442 -2709
rect -8746 -2732 -8729 -2722
rect -9050 -2766 -9033 -2756
rect -9113 -2977 -9101 -2766
rect -9045 -2977 -9033 -2766
rect -8809 -2893 -8797 -2732
rect -8741 -2893 -8729 -2732
rect -8809 -2903 -8792 -2893
rect -9113 -2987 -9096 -2977
rect -9400 -3005 -9354 -2994
rect -9050 -2987 -9033 -2977
rect -9096 -3005 -9050 -2994
rect -8746 -2903 -8729 -2893
rect -8505 -2732 -8488 -2722
rect -8184 -2720 -8138 -2709
rect -8442 -2732 -8425 -2722
rect -8505 -2977 -8493 -2732
rect -8437 -2977 -8425 -2732
rect -8201 -2732 -8184 -2722
rect -7880 -2720 -7834 -2709
rect -8138 -2732 -8121 -2722
rect -8201 -2893 -8189 -2732
rect -8133 -2893 -8121 -2732
rect -8201 -2903 -8184 -2893
rect -8505 -2987 -8488 -2977
rect -8792 -3005 -8746 -2994
rect -8442 -2987 -8425 -2977
rect -8488 -3005 -8442 -2994
rect -8138 -2903 -8121 -2893
rect -7897 -2766 -7880 -2756
rect -7576 -2720 -7530 -2709
rect -7593 -2732 -7576 -2722
rect -7272 -2720 -7226 -2709
rect -7530 -2732 -7513 -2722
rect -7834 -2766 -7817 -2756
rect -7897 -2977 -7885 -2766
rect -7829 -2977 -7817 -2766
rect -7593 -2893 -7581 -2732
rect -7525 -2893 -7513 -2732
rect -7593 -2903 -7576 -2893
rect -7897 -2987 -7880 -2977
rect -8184 -3005 -8138 -2994
rect -7834 -2987 -7817 -2977
rect -7880 -3005 -7834 -2994
rect -7530 -2903 -7513 -2893
rect -7289 -2732 -7272 -2722
rect -6968 -2720 -6922 -2709
rect -7226 -2732 -7209 -2722
rect -7289 -2977 -7277 -2732
rect -7221 -2977 -7209 -2732
rect -7289 -2987 -7272 -2977
rect -7576 -3005 -7530 -2994
rect -7226 -2987 -7209 -2977
rect -6985 -2732 -6968 -2722
rect -6664 -2720 -6618 -2709
rect -6922 -2732 -6905 -2722
rect -6985 -2977 -6973 -2732
rect -6917 -2977 -6905 -2732
rect -6985 -2987 -6968 -2977
rect -7272 -3005 -7226 -2994
rect -6922 -2987 -6905 -2977
rect -6681 -2920 -6664 -2910
rect -6360 -2720 -6314 -2709
rect -6618 -2920 -6601 -2910
rect -6681 -2977 -6669 -2920
rect -6613 -2977 -6601 -2920
rect -6681 -2987 -6664 -2977
rect -6968 -3005 -6922 -2994
rect -6618 -2987 -6601 -2977
rect -6664 -3005 -6618 -2994
rect -6360 -3005 -6314 -2994
rect -6129 -2848 -6007 -2837
rect -9931 -3086 -9920 -3040
rect -9746 -3086 -9735 -3040
rect -9627 -3086 -9616 -3040
rect -9442 -3086 -9431 -3040
rect -9323 -3086 -9312 -3040
rect -9138 -3086 -9127 -3040
rect -9019 -3086 -9008 -3040
rect -8834 -3086 -8823 -3040
rect -8715 -3086 -8704 -3040
rect -8530 -3086 -8519 -3040
rect -8411 -3086 -8400 -3040
rect -8226 -3086 -8215 -3040
rect -8107 -3086 -8096 -3040
rect -7922 -3086 -7911 -3040
rect -7803 -3086 -7792 -3040
rect -7618 -3086 -7607 -3040
rect -7499 -3086 -7488 -3040
rect -7314 -3086 -7303 -3040
rect -7195 -3086 -7184 -3040
rect -7010 -3086 -6999 -3040
rect -6891 -3086 -6880 -3040
rect -6706 -3086 -6695 -3040
rect -6587 -3086 -6576 -3040
rect -6402 -3086 -6391 -3040
rect -6129 -3144 -6118 -2848
rect -6143 -3160 -6118 -3144
rect -6018 -3144 -6007 -2848
rect -6143 -3297 -6129 -3160
rect -10315 -3359 -10193 -3348
rect -6144 -3370 -6129 -3297
rect -6018 -3308 -6002 -3144
rect -6018 -3348 -6007 -3308
rect -6024 -3370 -6007 -3348
rect -6144 -3388 -6007 -3370
rect -8598 -3563 -8552 -3552
rect -8615 -3652 -8598 -3650
rect -8383 -3554 -8307 -3524
rect -8383 -3600 -8372 -3554
rect -8318 -3600 -8307 -3554
rect -8199 -3554 -8123 -3524
rect -8199 -3600 -8188 -3554
rect -8134 -3600 -8123 -3554
rect -8015 -3554 -7939 -3524
rect -8015 -3600 -8004 -3554
rect -7950 -3600 -7939 -3554
rect -7770 -3563 -7724 -3552
rect -8460 -3646 -8414 -3635
rect -8552 -3652 -8535 -3650
rect -8615 -3774 -8603 -3652
rect -8547 -3774 -8535 -3652
rect -8615 -3776 -8598 -3774
rect -8552 -3776 -8535 -3774
rect -8276 -3646 -8230 -3635
rect -8293 -3652 -8276 -3650
rect -8092 -3646 -8046 -3635
rect -8230 -3652 -8213 -3650
rect -8293 -3774 -8281 -3652
rect -8225 -3774 -8213 -3652
rect -8293 -3776 -8276 -3774
rect -8460 -3791 -8414 -3780
rect -8230 -3776 -8213 -3774
rect -8109 -3652 -8092 -3650
rect -7908 -3646 -7862 -3635
rect -8046 -3652 -8029 -3650
rect -8109 -3774 -8097 -3652
rect -8041 -3774 -8029 -3652
rect -8109 -3776 -8092 -3774
rect -8276 -3791 -8230 -3780
rect -8046 -3776 -8029 -3774
rect -8092 -3791 -8046 -3780
rect -7908 -3791 -7862 -3780
rect -8598 -3874 -8552 -3863
rect -8383 -3872 -8372 -3826
rect -8318 -3872 -8307 -3826
rect -8383 -3902 -8307 -3872
rect -8199 -3872 -8188 -3826
rect -8134 -3872 -8123 -3826
rect -13382 -4003 -13286 -3992
rect -11391 -4003 -11287 -3993
rect -8199 -4003 -8123 -3872
rect -8015 -3872 -8004 -3826
rect -7950 -3872 -7939 -3826
rect -8015 -3902 -7939 -3872
rect -7770 -3874 -7724 -3863
rect -5035 -4003 -4931 -3993
rect -13382 -4004 -11379 -4003
rect -13382 -4082 -13368 -4004
rect -13290 -4082 -11379 -4004
rect -13382 -4083 -11379 -4082
rect -11299 -4083 -5023 -4003
rect -4943 -4083 -4931 -4003
rect -13382 -4096 -13286 -4083
rect -11391 -4093 -11287 -4083
rect -5035 -4093 -4931 -4083
rect -12534 -4363 -2407 -4321
rect -12534 -4375 -4454 -4363
rect -12534 -4376 -6132 -4375
rect -12534 -4443 -10639 -4376
rect -12534 -4530 -11640 -4443
rect -11555 -4463 -10639 -4443
rect -10550 -4381 -6132 -4376
rect -10550 -4463 -10083 -4381
rect -11555 -4530 -10083 -4463
rect -12534 -4592 -10083 -4530
rect -9728 -4578 -6132 -4381
rect -6018 -4429 -4454 -4375
rect -6018 -4531 -5654 -4429
rect -5550 -4451 -4454 -4429
rect -5550 -4531 -4764 -4451
rect -6018 -4558 -4764 -4531
rect -4655 -4558 -4454 -4451
rect -6018 -4578 -4454 -4558
rect -9728 -4592 -4454 -4578
rect -12534 -4663 -4454 -4592
rect -2454 -4663 -2407 -4363
rect -12534 -4701 -2407 -4663
<< via1 >>
rect -13105 11438 -13049 11494
rect -4454 5134 -2454 5434
rect -13665 3881 -13607 3939
rect -12366 3880 -12306 3940
rect -10747 3884 -10695 3936
rect -10187 3673 -10135 3676
rect -10187 3627 -10184 3673
rect -10184 3627 -10138 3673
rect -10138 3627 -10135 3673
rect -10187 3624 -10135 3627
rect -8327 3739 -8322 3795
rect -8322 3739 -8276 3795
rect -8276 3739 -8271 3795
rect -8051 3739 -8046 3795
rect -8046 3739 -8000 3795
rect -8000 3739 -7995 3795
rect -8189 3481 -8133 3537
rect -8189 3343 -8133 3399
rect -10519 2300 -10439 2376
rect -8327 2919 -8322 2975
rect -8322 2919 -8276 2975
rect -8276 2919 -8271 2975
rect -8419 2768 -8418 2799
rect -8418 2768 -8364 2799
rect -8364 2768 -8363 2799
rect -8419 2743 -8363 2768
rect -8051 2919 -8046 2975
rect -8046 2919 -8000 2975
rect -8000 2919 -7995 2975
rect -7959 2768 -7958 2799
rect -7958 2768 -7904 2799
rect -7904 2768 -7903 2799
rect -7959 2743 -7903 2768
rect -8419 2300 -8363 2376
rect -12086 1883 -12006 1961
rect -7959 2300 -7903 2376
rect -5883 2300 -5803 2376
rect -5676 1787 -5596 1847
rect -11642 1462 -11551 1551
rect -4764 1542 -4655 1649
rect -11379 1356 -11299 1432
rect -5023 1356 -4943 1432
rect -11029 530 -11024 664
rect -11024 530 -10978 664
rect -10978 530 -10973 664
rect -10845 530 -10840 664
rect -10840 530 -10794 664
rect -10794 530 -10789 664
rect -10707 530 -10702 664
rect -10702 530 -10656 664
rect -10656 530 -10651 664
rect -10169 530 -10164 664
rect -10164 530 -10118 664
rect -10118 530 -10113 664
rect -9985 530 -9980 664
rect -9980 530 -9934 664
rect -9934 530 -9929 664
rect -9847 530 -9842 664
rect -9842 530 -9796 664
rect -9796 530 -9791 664
rect -9405 533 -9400 677
rect -9400 533 -9354 677
rect -9354 533 -9349 677
rect -9101 520 -9096 576
rect -9096 520 -9050 576
rect -9050 520 -9045 576
rect -8797 533 -8792 677
rect -8792 533 -8746 677
rect -8746 533 -8741 677
rect -8493 520 -8488 576
rect -8488 520 -8442 576
rect -8442 520 -8437 576
rect -8189 533 -8184 677
rect -8184 533 -8138 677
rect -8138 533 -8133 677
rect -7885 520 -7880 576
rect -7880 520 -7834 576
rect -7834 520 -7829 576
rect -7581 533 -7576 677
rect -7576 533 -7530 677
rect -7530 533 -7525 677
rect -7277 520 -7272 576
rect -7272 520 -7226 576
rect -7226 520 -7221 576
rect -6973 533 -6968 677
rect -6968 533 -6922 677
rect -6922 533 -6917 677
rect -6531 530 -6526 664
rect -6526 530 -6480 664
rect -6480 530 -6475 664
rect -8298 464 -8242 469
rect -8080 464 -8024 469
rect -8298 418 -8242 464
rect -8080 418 -8024 464
rect -6393 530 -6388 664
rect -6388 530 -6342 664
rect -6342 530 -6337 664
rect -6209 530 -6204 664
rect -6204 530 -6158 664
rect -6158 530 -6153 664
rect -8298 413 -8242 418
rect -8080 413 -8024 418
rect -5671 530 -5666 664
rect -5666 530 -5620 664
rect -5620 530 -5615 664
rect -5533 530 -5528 664
rect -5528 530 -5482 664
rect -5482 530 -5477 664
rect -5349 530 -5344 664
rect -5344 530 -5298 664
rect -5298 530 -5293 664
rect -10519 77 -10439 161
rect -9997 77 -9917 161
rect -9251 79 -9171 159
rect -8643 79 -8563 159
rect -8505 79 -8425 159
rect -7897 79 -7817 159
rect -7759 79 -7679 159
rect -7151 79 -7071 159
rect -6405 77 -6325 161
rect -5883 77 -5803 161
rect -8842 -180 -8762 -135
rect -8842 -215 -8762 -180
rect -7560 -180 -7480 -135
rect -9985 -729 -9980 -585
rect -9980 -729 -9934 -585
rect -9934 -729 -9929 -585
rect -9239 -423 -9234 -279
rect -9234 -423 -9188 -279
rect -9188 -423 -9183 -279
rect -9543 -639 -9538 -495
rect -9538 -639 -9492 -495
rect -9492 -639 -9487 -495
rect -8631 -423 -8626 -279
rect -8626 -423 -8580 -279
rect -8580 -423 -8575 -279
rect -8935 -639 -8930 -495
rect -8930 -639 -8884 -495
rect -8884 -639 -8879 -495
rect -7560 -215 -7480 -180
rect -7747 -423 -7742 -279
rect -7742 -423 -7696 -279
rect -7696 -423 -7691 -279
rect -7139 -423 -7134 -279
rect -7134 -423 -7088 -279
rect -7088 -423 -7083 -279
rect -7443 -639 -7438 -495
rect -7438 -639 -7392 -495
rect -7392 -639 -7387 -495
rect -6835 -639 -6830 -495
rect -6830 -639 -6784 -495
rect -6784 -639 -6779 -495
rect -6393 -729 -6388 -585
rect -6388 -729 -6342 -585
rect -6342 -729 -6337 -585
rect -10857 -1085 -10777 -1005
rect -9721 -1085 -9641 -1005
rect -9555 -1085 -9475 -1005
rect -8947 -1085 -8867 -1005
rect -7455 -1085 -7375 -1005
rect -6847 -1085 -6767 -1005
rect -6681 -1085 -6601 -1005
rect -5545 -1085 -5465 -1005
rect -10304 -1564 -10204 -1403
rect -9709 -1974 -9704 -1813
rect -9704 -1974 -9658 -1813
rect -9658 -1974 -9653 -1813
rect -9405 -2022 -9400 -1861
rect -9400 -2022 -9354 -1861
rect -9354 -2022 -9349 -1861
rect -9101 -1994 -9096 -1777
rect -9096 -1994 -9050 -1777
rect -9050 -1994 -9045 -1777
rect -8493 -1833 -8488 -1777
rect -8488 -1833 -8442 -1777
rect -8442 -1833 -8437 -1777
rect -8797 -2022 -8792 -1861
rect -8792 -2022 -8746 -1861
rect -8746 -2022 -8741 -1861
rect -7885 -1833 -7880 -1777
rect -7880 -1833 -7834 -1777
rect -7834 -1833 -7829 -1777
rect -8189 -2022 -8184 -1861
rect -8184 -2022 -8138 -1861
rect -8138 -2022 -8133 -1861
rect -7581 -2022 -7576 -1861
rect -7576 -2022 -7530 -1861
rect -7530 -2022 -7525 -1861
rect -7277 -2022 -7272 -1777
rect -7272 -2022 -7226 -1777
rect -7226 -2022 -7221 -1777
rect -6973 -2022 -6968 -1861
rect -6968 -2022 -6922 -1861
rect -6922 -2022 -6917 -1861
rect -6669 -1974 -6664 -1813
rect -6664 -1974 -6618 -1813
rect -6618 -1974 -6613 -1813
rect -6118 -1564 -6018 -1403
rect -9261 -2077 -9191 -2068
rect -8956 -2077 -8886 -2068
rect -8046 -2077 -7976 -2068
rect -7741 -2077 -7671 -2068
rect -6826 -2077 -6756 -2068
rect -9261 -2123 -9191 -2077
rect -8956 -2123 -8886 -2077
rect -8046 -2123 -7976 -2077
rect -7741 -2123 -7671 -2077
rect -6826 -2123 -6756 -2077
rect -9261 -2128 -9191 -2123
rect -8956 -2128 -8886 -2123
rect -8046 -2128 -7976 -2123
rect -7741 -2128 -7671 -2123
rect -6826 -2128 -6756 -2123
rect -13707 -2252 -13634 -2179
rect -9254 -2282 -9198 -2226
rect -8039 -2282 -7983 -2226
rect -6511 -2253 -6451 -2193
rect -13704 -2577 -13631 -2504
rect -8949 -2530 -8893 -2474
rect -7734 -2530 -7678 -2474
rect -6251 -2563 -6191 -2503
rect -9261 -2674 -9191 -2628
rect -8956 -2674 -8886 -2628
rect -8046 -2674 -7976 -2628
rect -7741 -2674 -7671 -2628
rect -6826 -2674 -6756 -2628
rect -9261 -2688 -9191 -2674
rect -8956 -2688 -8886 -2674
rect -8046 -2688 -7976 -2674
rect -7741 -2688 -7671 -2674
rect -6826 -2688 -6756 -2674
rect -10304 -3348 -10204 -3187
rect -9405 -2893 -9400 -2732
rect -9400 -2893 -9354 -2732
rect -9354 -2893 -9349 -2732
rect -9709 -2977 -9704 -2921
rect -9704 -2977 -9658 -2921
rect -9658 -2977 -9653 -2921
rect -9101 -2977 -9096 -2766
rect -9096 -2977 -9050 -2766
rect -9050 -2977 -9045 -2766
rect -8797 -2893 -8792 -2732
rect -8792 -2893 -8746 -2732
rect -8746 -2893 -8741 -2732
rect -8493 -2977 -8488 -2732
rect -8488 -2977 -8442 -2732
rect -8442 -2977 -8437 -2732
rect -8189 -2893 -8184 -2732
rect -8184 -2893 -8138 -2732
rect -8138 -2893 -8133 -2732
rect -7885 -2977 -7880 -2766
rect -7880 -2977 -7834 -2766
rect -7834 -2977 -7829 -2766
rect -7581 -2893 -7576 -2732
rect -7576 -2893 -7530 -2732
rect -7530 -2893 -7525 -2732
rect -7277 -2977 -7272 -2732
rect -7272 -2977 -7226 -2732
rect -7226 -2977 -7221 -2732
rect -6973 -2977 -6968 -2732
rect -6968 -2977 -6922 -2732
rect -6922 -2977 -6917 -2732
rect -6669 -2977 -6664 -2920
rect -6664 -2977 -6618 -2920
rect -6618 -2977 -6613 -2920
rect -6129 -3348 -6118 -3160
rect -6118 -3348 -6024 -3160
rect -6129 -3370 -6024 -3348
rect -8603 -3774 -8598 -3652
rect -8598 -3774 -8552 -3652
rect -8552 -3774 -8547 -3652
rect -8281 -3774 -8276 -3652
rect -8276 -3774 -8230 -3652
rect -8230 -3774 -8225 -3652
rect -8097 -3774 -8092 -3652
rect -8092 -3774 -8046 -3652
rect -8046 -3774 -8041 -3652
rect -13368 -4082 -13290 -4004
rect -11379 -4083 -11299 -4003
rect -5023 -4083 -4943 -4003
rect -11640 -4530 -11555 -4443
rect -10639 -4463 -10550 -4376
rect -10083 -4592 -9728 -4381
rect -6132 -4578 -6018 -4375
rect -5654 -4531 -5550 -4429
rect -4764 -4558 -4655 -4451
rect -4454 -4663 -2454 -4363
<< metal2 >>
rect -8093 38010 -8037 38726
rect 4049 38341 4105 38603
rect 4045 38285 18990 38341
rect -13170 27521 -12770 27577
rect -13224 16389 -12960 16509
rect -13233 15879 -12960 15999
rect -13117 11494 -13047 11506
rect -13117 11438 -13105 11494
rect -13049 11438 -13047 11494
rect -13117 11426 -13047 11438
rect -13105 6930 -13049 11426
rect -13369 6920 -13049 6930
rect -13369 6820 -13105 6920
rect -13369 6810 -13049 6820
rect -13369 6770 -13289 6810
rect -4464 5434 -2430 5477
rect -4464 5134 -4454 5434
rect -2454 5134 -2430 5434
rect -4464 5097 -2430 5134
rect -13680 3940 -13603 3954
rect -13894 3939 -13603 3940
rect -13894 3881 -13665 3939
rect -13607 3881 -13603 3939
rect -13894 3880 -13603 3881
rect -13680 3867 -13603 3880
rect -12380 3940 -12294 3954
rect -10771 3940 -10671 3950
rect -12380 3880 -12366 3940
rect -12306 3936 -10671 3940
rect -12306 3884 -10747 3936
rect -10695 3884 -10671 3936
rect -12306 3880 -10671 3884
rect -12380 3866 -12294 3880
rect -10771 3870 -10671 3880
rect -8339 3795 -8259 3805
rect -8339 3739 -8327 3795
rect -8271 3739 -8259 3795
rect -8339 3729 -8259 3739
rect -8063 3795 -7983 3805
rect -8063 3739 -8051 3795
rect -7995 3739 -7983 3795
rect -8063 3729 -7983 3739
rect -10201 3680 -10121 3690
rect -10211 3676 -10111 3680
rect -10211 3624 -10187 3676
rect -10135 3624 -8820 3676
rect -10211 3620 -8820 3624
rect -10201 3610 -10121 3620
rect -8876 3289 -8820 3620
rect -8327 3537 -8271 3729
rect -8202 3537 -8122 3549
rect -8327 3481 -8189 3537
rect -8133 3481 -8122 3537
rect -8327 3289 -8271 3481
rect -8202 3469 -8122 3481
rect -8201 3399 -8121 3409
rect -8051 3399 -7995 3729
rect -8201 3343 -8189 3399
rect -8133 3343 -7995 3399
rect -8201 3333 -8121 3343
rect -8876 3233 -8271 3289
rect -8327 2985 -8271 3233
rect -8051 3289 -7995 3343
rect -8051 3233 -7451 3289
rect -8051 2985 -7995 3233
rect -8339 2975 -8259 2985
rect -8339 2919 -8327 2975
rect -8271 2919 -8259 2975
rect -8339 2909 -8259 2919
rect -8063 2975 -7983 2985
rect -8063 2919 -8051 2975
rect -7995 2919 -7983 2975
rect -8063 2909 -7983 2919
rect -8431 2799 -8351 2809
rect -8431 2743 -8419 2799
rect -8363 2743 -8351 2799
rect -8431 2733 -8351 2743
rect -7971 2799 -7891 2809
rect -7971 2743 -7959 2799
rect -7903 2743 -7891 2799
rect -7971 2733 -7891 2743
rect -10531 2376 -10437 2388
rect -8419 2378 -8363 2733
rect -7959 2378 -7903 2733
rect -10531 2300 -10519 2376
rect -10439 2300 -10437 2376
rect -10531 2298 -10437 2300
rect -8421 2376 -8349 2378
rect -8421 2300 -8419 2376
rect -8363 2300 -8349 2376
rect -12103 1961 -11990 1978
rect -12103 1883 -12086 1961
rect -12006 1883 -11990 1961
rect -12103 1872 -11990 1883
rect -12086 1417 -12006 1872
rect -11650 1551 -11541 1564
rect -11650 1462 -11642 1551
rect -11551 1462 -11541 1551
rect -11650 1455 -11541 1462
rect -12096 1397 -11996 1417
rect -12096 1317 -12086 1397
rect -12006 1317 -11996 1397
rect -12096 1307 -11996 1317
rect -11642 79 -11551 1455
rect -11391 1432 -11287 1446
rect -11391 1356 -11379 1432
rect -11299 1356 -11287 1432
rect -11391 1346 -11287 1356
rect -13722 -2177 -13632 -2166
rect -13880 -2179 -13632 -2177
rect -13880 -2252 -13707 -2179
rect -13634 -2252 -13632 -2179
rect -13722 -2266 -13632 -2252
rect -13717 -2502 -13627 -2491
rect -13878 -2504 -13627 -2502
rect -13878 -2577 -13704 -2504
rect -13631 -2577 -13627 -2504
rect -13717 -2591 -13627 -2577
rect -13382 -4004 -13286 -3992
rect -13784 -4082 -13368 -4004
rect -13290 -4082 -13286 -4004
rect -13382 -4096 -13286 -4082
rect -11640 -4421 -11553 79
rect -11379 -3993 -11299 1346
rect -11051 1123 -10951 1133
rect -11051 1043 -11041 1123
rect -10961 1043 -10951 1123
rect -11051 1033 -10951 1043
rect -10729 1123 -10629 1133
rect -10729 1043 -10719 1123
rect -10639 1043 -10629 1123
rect -10729 1033 -10629 1043
rect -11041 664 -10961 1033
rect -10845 666 -10789 674
rect -11041 530 -11029 664
rect -10973 530 -10961 664
rect -11041 528 -10961 530
rect -10857 664 -10777 666
rect -10857 530 -10845 664
rect -10789 530 -10777 664
rect -11029 520 -10973 528
rect -10857 -995 -10777 530
rect -10719 664 -10639 1033
rect -10719 530 -10707 664
rect -10651 530 -10639 664
rect -10719 528 -10639 530
rect -10707 520 -10651 528
rect -10519 173 -10439 2298
rect -8421 2288 -8349 2300
rect -7973 2376 -7901 2378
rect -7973 2300 -7959 2376
rect -7903 2300 -7901 2376
rect -7973 2288 -7901 2300
rect -5895 2376 -5791 2388
rect -5895 2300 -5883 2376
rect -5803 2300 -5791 2376
rect -5895 2298 -5791 2300
rect -10191 1123 -10091 1133
rect -10191 1043 -10181 1123
rect -10101 1043 -10091 1123
rect -10191 1033 -10091 1043
rect -9869 1123 -9769 1133
rect -9869 1043 -9859 1123
rect -9779 1043 -9769 1123
rect -9869 1033 -9769 1043
rect -9427 1123 -9327 1133
rect -9427 1043 -9417 1123
rect -9337 1043 -9327 1123
rect -9427 1033 -9327 1043
rect -8819 1123 -8719 1133
rect -8819 1043 -8809 1123
rect -8729 1043 -8719 1123
rect -8819 1033 -8719 1043
rect -8211 1123 -8111 1133
rect -8211 1043 -8201 1123
rect -8121 1043 -8111 1123
rect -8211 1033 -8111 1043
rect -7603 1123 -7503 1133
rect -7603 1043 -7593 1123
rect -7513 1043 -7503 1123
rect -7603 1033 -7503 1043
rect -6995 1123 -6895 1133
rect -6995 1043 -6985 1123
rect -6905 1043 -6895 1123
rect -6995 1033 -6895 1043
rect -6553 1123 -6453 1133
rect -6553 1043 -6543 1123
rect -6463 1043 -6453 1123
rect -6553 1033 -6453 1043
rect -6231 1123 -6131 1133
rect -6231 1043 -6221 1123
rect -6141 1043 -6131 1123
rect -6231 1033 -6131 1043
rect -10181 664 -10101 1033
rect -9985 666 -9929 674
rect -10181 530 -10169 664
rect -10113 530 -10101 664
rect -10181 528 -10101 530
rect -9997 664 -9917 666
rect -9997 530 -9985 664
rect -9929 530 -9917 664
rect -10169 520 -10113 528
rect -10531 161 -10427 173
rect -9997 171 -9917 530
rect -9859 664 -9779 1033
rect -9859 530 -9847 664
rect -9791 530 -9779 664
rect -9417 677 -9337 1033
rect -9417 533 -9405 677
rect -9349 533 -9337 677
rect -8809 677 -8729 1033
rect -9417 531 -9337 533
rect -9113 576 -9033 586
rect -9859 528 -9779 530
rect -9847 520 -9791 528
rect -9405 523 -9349 531
rect -9113 520 -9101 576
rect -9045 520 -9033 576
rect -8809 533 -8797 677
rect -8741 533 -8729 677
rect -8201 677 -8121 1033
rect -8809 531 -8729 533
rect -8505 576 -8425 586
rect -8797 523 -8741 531
rect -9113 510 -9033 520
rect -8505 520 -8493 576
rect -8437 520 -8425 576
rect -8201 533 -8189 677
rect -8133 533 -8121 677
rect -7593 677 -7513 1033
rect -8201 531 -8121 533
rect -7897 576 -7817 586
rect -8189 523 -8133 531
rect -10531 77 -10519 161
rect -10439 77 -10427 161
rect -10531 67 -10427 77
rect -10009 161 -9905 171
rect -8505 169 -8425 520
rect -7897 520 -7885 576
rect -7829 520 -7817 576
rect -7593 533 -7581 677
rect -7525 533 -7513 677
rect -6985 677 -6905 1033
rect -7593 531 -7513 533
rect -7289 576 -7209 586
rect -7581 523 -7525 531
rect -8310 469 -8230 479
rect -8310 413 -8298 469
rect -8242 413 -8230 469
rect -8310 339 -8230 413
rect -8092 469 -8012 479
rect -8092 413 -8080 469
rect -8024 413 -8012 469
rect -8320 329 -8220 339
rect -8320 249 -8310 329
rect -8230 249 -8220 329
rect -8320 239 -8220 249
rect -8092 169 -8012 413
rect -7897 339 -7817 520
rect -7289 520 -7277 576
rect -7221 520 -7209 576
rect -6985 533 -6973 677
rect -6917 533 -6905 677
rect -6985 531 -6905 533
rect -6543 664 -6463 1033
rect -6393 666 -6337 674
rect -6973 523 -6917 531
rect -6543 530 -6531 664
rect -6475 530 -6463 664
rect -6543 528 -6463 530
rect -6405 664 -6325 666
rect -6405 530 -6393 664
rect -6337 530 -6325 664
rect -6531 520 -6475 528
rect -7289 510 -7209 520
rect -7907 329 -7807 339
rect -7907 249 -7897 329
rect -7817 249 -7807 329
rect -7907 239 -7807 249
rect -7897 169 -7817 239
rect -6405 171 -6325 530
rect -6221 664 -6141 1033
rect -6221 530 -6209 664
rect -6153 530 -6141 664
rect -6221 528 -6141 530
rect -6209 520 -6153 528
rect -5883 171 -5803 2298
rect -5696 1887 -5576 1907
rect -5696 1787 -5676 1887
rect -5596 1787 -5576 1887
rect -5696 1767 -5576 1787
rect -4791 1649 -4633 1664
rect -4791 1542 -4764 1649
rect -4655 1542 -4633 1649
rect -4791 1531 -4633 1542
rect -5035 1432 -4931 1444
rect -5035 1356 -5023 1432
rect -4943 1356 -4931 1432
rect -5035 1344 -4931 1356
rect -5693 1123 -5593 1133
rect -5693 1043 -5683 1123
rect -5603 1043 -5593 1123
rect -5693 1033 -5593 1043
rect -5371 1123 -5271 1133
rect -5371 1043 -5361 1123
rect -5281 1043 -5271 1123
rect -5371 1033 -5271 1043
rect -5683 664 -5603 1033
rect -5533 666 -5477 674
rect -5683 530 -5671 664
rect -5615 530 -5603 664
rect -5683 528 -5603 530
rect -5545 664 -5465 666
rect -5545 530 -5533 664
rect -5477 530 -5465 664
rect -5671 520 -5615 528
rect -10009 77 -9997 161
rect -9917 77 -9905 161
rect -10009 67 -9905 77
rect -9263 159 -9159 169
rect -9263 79 -9251 159
rect -9171 79 -9159 159
rect -9263 65 -9159 79
rect -8655 159 -8415 169
rect -8102 159 -8002 169
rect -8655 79 -8643 159
rect -8563 79 -8505 159
rect -8425 79 -8092 159
rect -8012 79 -8002 159
rect -8655 65 -8415 79
rect -8102 69 -8002 79
rect -7909 159 -7667 169
rect -7909 79 -7897 159
rect -7817 79 -7759 159
rect -7679 79 -7667 159
rect -7909 65 -7667 79
rect -7163 159 -7059 170
rect -7163 79 -7151 159
rect -7071 79 -7059 159
rect -7163 66 -7059 79
rect -6417 161 -6313 171
rect -6417 77 -6405 161
rect -6325 77 -6313 161
rect -6417 67 -6313 77
rect -5895 161 -5791 171
rect -5895 77 -5883 161
rect -5803 77 -5791 161
rect -5895 67 -5791 77
rect -9251 -279 -9171 65
rect -8852 -135 -8752 -125
rect -8852 -215 -8842 -135
rect -8762 -215 -8752 -135
rect -8852 -225 -8752 -215
rect -9251 -423 -9239 -279
rect -9183 -423 -9171 -279
rect -9251 -425 -9171 -423
rect -8643 -279 -8563 65
rect -8643 -423 -8631 -279
rect -8575 -423 -8563 -279
rect -8643 -425 -8563 -423
rect -7759 -279 -7679 65
rect -7570 -135 -7470 -125
rect -7570 -215 -7560 -135
rect -7480 -215 -7470 -135
rect -7570 -225 -7470 -215
rect -7759 -423 -7747 -279
rect -7691 -423 -7679 -279
rect -7759 -425 -7679 -423
rect -7151 -279 -7071 66
rect -7151 -423 -7139 -279
rect -7083 -423 -7071 -279
rect -7151 -425 -7071 -423
rect -9239 -433 -9183 -425
rect -8631 -433 -8575 -425
rect -7747 -433 -7691 -425
rect -7139 -433 -7083 -425
rect -9543 -493 -9487 -485
rect -8935 -493 -8879 -485
rect -7443 -493 -7387 -485
rect -6835 -493 -6779 -485
rect -9555 -495 -9475 -493
rect -9997 -585 -9917 -575
rect -10306 -729 -9985 -585
rect -9929 -729 -9917 -585
rect -10869 -1005 -10765 -995
rect -10869 -1085 -10857 -1005
rect -10777 -1085 -10765 -1005
rect -10869 -1095 -10765 -1085
rect -10306 -1265 -10202 -729
rect -9997 -740 -9917 -729
rect -9555 -639 -9543 -495
rect -9487 -639 -9475 -495
rect -9555 -993 -9475 -639
rect -8947 -495 -8867 -493
rect -8947 -639 -8935 -495
rect -8879 -639 -8867 -495
rect -8947 -993 -8867 -639
rect -7455 -495 -7375 -493
rect -7455 -639 -7443 -495
rect -7387 -639 -7375 -495
rect -7455 -993 -7375 -639
rect -6847 -495 -6767 -493
rect -6847 -639 -6835 -495
rect -6779 -639 -6767 -495
rect -6847 -993 -6767 -639
rect -6405 -585 -6325 -575
rect -6405 -729 -6393 -585
rect -6337 -729 -6016 -585
rect -6405 -740 -6325 -729
rect -9733 -1005 -9629 -993
rect -9733 -1085 -9721 -1005
rect -9641 -1085 -9629 -1005
rect -9733 -1097 -9629 -1085
rect -9567 -1005 -9463 -993
rect -9567 -1085 -9555 -1005
rect -9475 -1085 -9463 -1005
rect -9567 -1097 -9463 -1085
rect -8959 -1005 -8855 -993
rect -8959 -1085 -8947 -1005
rect -8867 -1085 -8855 -1005
rect -8959 -1097 -8855 -1085
rect -7467 -1005 -7363 -993
rect -7467 -1085 -7455 -1005
rect -7375 -1085 -7363 -1005
rect -7467 -1097 -7363 -1085
rect -6859 -1005 -6755 -993
rect -6859 -1085 -6847 -1005
rect -6767 -1085 -6755 -1005
rect -6859 -1097 -6755 -1085
rect -6693 -1005 -6589 -993
rect -6693 -1085 -6681 -1005
rect -6601 -1085 -6589 -1005
rect -6693 -1097 -6589 -1085
rect -10647 -1369 -10202 -1265
rect -11391 -4003 -11287 -3993
rect -11391 -4083 -11379 -4003
rect -11299 -4083 -11287 -4003
rect -11391 -4093 -11287 -4083
rect -10639 -4123 -10550 -1369
rect -10306 -1403 -10202 -1369
rect -10306 -1564 -10304 -1403
rect -10204 -1564 -10202 -1403
rect -10306 -1576 -10202 -1564
rect -9721 -1813 -9641 -1097
rect -6681 -1575 -6601 -1097
rect -9721 -1974 -9709 -1813
rect -9653 -1974 -9641 -1813
rect -9113 -1631 -6601 -1575
rect -6120 -1256 -6016 -729
rect -5545 -995 -5465 530
rect -5361 664 -5281 1033
rect -5361 530 -5349 664
rect -5293 530 -5281 664
rect -5361 528 -5281 530
rect -5349 520 -5293 528
rect -5557 -1005 -5453 -995
rect -5557 -1085 -5545 -1005
rect -5465 -1085 -5453 -1005
rect -5557 -1095 -5453 -1085
rect -6120 -1360 -5550 -1256
rect -6120 -1403 -6016 -1360
rect -6120 -1564 -6118 -1403
rect -6018 -1564 -6016 -1403
rect -6120 -1576 -6016 -1564
rect -9113 -1777 -9033 -1631
rect -9721 -1984 -9641 -1974
rect -9417 -1861 -9337 -1851
rect -9417 -2022 -9405 -1861
rect -9349 -2022 -9337 -1861
rect -9113 -1994 -9101 -1777
rect -9045 -1994 -9033 -1777
rect -8505 -1777 -8425 -1767
rect -8505 -1833 -8493 -1777
rect -8437 -1833 -8425 -1777
rect -8505 -1843 -8425 -1833
rect -7897 -1777 -7817 -1631
rect -7897 -1833 -7885 -1777
rect -7829 -1833 -7817 -1777
rect -7897 -1843 -7817 -1833
rect -7289 -1777 -7209 -1767
rect -9113 -2002 -9033 -1994
rect -8809 -1861 -8729 -1851
rect -9417 -2352 -9337 -2022
rect -8809 -2022 -8797 -1861
rect -8741 -2022 -8729 -1861
rect -9276 -2068 -8871 -2058
rect -9276 -2128 -9261 -2068
rect -9191 -2128 -8956 -2068
rect -8886 -2128 -8871 -2068
rect -9276 -2138 -8871 -2128
rect -9266 -2226 -9186 -2216
rect -9266 -2282 -9254 -2226
rect -9198 -2282 -9186 -2226
rect -9266 -2292 -9186 -2282
rect -8809 -2352 -8729 -2022
rect -8201 -1861 -8121 -1851
rect -8201 -2022 -8189 -1861
rect -8133 -2022 -8121 -1861
rect -8201 -2352 -8121 -2022
rect -7593 -1861 -7513 -1851
rect -7593 -2022 -7581 -1861
rect -7525 -2022 -7513 -1861
rect -8061 -2068 -7656 -2058
rect -8061 -2128 -8046 -2068
rect -7976 -2128 -7741 -2068
rect -7671 -2128 -7656 -2068
rect -8061 -2138 -7656 -2128
rect -8051 -2226 -7971 -2216
rect -8051 -2282 -8039 -2226
rect -7983 -2282 -7971 -2226
rect -8051 -2292 -7971 -2282
rect -7593 -2352 -7513 -2022
rect -7289 -2022 -7277 -1777
rect -7221 -2022 -7209 -1777
rect -6681 -1813 -6601 -1631
rect -7289 -2032 -7209 -2022
rect -6985 -1861 -6905 -1851
rect -6985 -2022 -6973 -1861
rect -6917 -2022 -6905 -1861
rect -6681 -1974 -6669 -1813
rect -6613 -1974 -6601 -1813
rect -6681 -1984 -6601 -1974
rect -6985 -2352 -6905 -2022
rect -6841 -2068 -6741 -2058
rect -6547 -2068 -6321 -2067
rect -6841 -2128 -6826 -2068
rect -6756 -2127 -6321 -2068
rect -6756 -2128 -6582 -2127
rect -6841 -2138 -6741 -2128
rect -6526 -2193 -6441 -2183
rect -6526 -2253 -6511 -2193
rect -6451 -2253 -6441 -2193
rect -6526 -2268 -6441 -2253
rect -9417 -2408 -6905 -2352
rect -9417 -2732 -9337 -2408
rect -8961 -2474 -8881 -2464
rect -8961 -2530 -8949 -2474
rect -8893 -2530 -8881 -2474
rect -8961 -2540 -8881 -2530
rect -9276 -2628 -8871 -2618
rect -9276 -2688 -9261 -2628
rect -9191 -2688 -8956 -2628
rect -8886 -2688 -8871 -2628
rect -9276 -2698 -8871 -2688
rect -9417 -2893 -9405 -2732
rect -9349 -2893 -9337 -2732
rect -8809 -2732 -8729 -2408
rect -9721 -2921 -9641 -2911
rect -9721 -2977 -9709 -2921
rect -9653 -2977 -9641 -2921
rect -9721 -2987 -9641 -2977
rect -10306 -3187 -10202 -3175
rect -10306 -3348 -10304 -3187
rect -10204 -3348 -10202 -3187
rect -9417 -3239 -9337 -2893
rect -9113 -2766 -9033 -2756
rect -9113 -2977 -9101 -2766
rect -9045 -2977 -9033 -2766
rect -8809 -2893 -8797 -2732
rect -8741 -2893 -8729 -2732
rect -8809 -2903 -8729 -2893
rect -8505 -2732 -8425 -2722
rect -9113 -3123 -9033 -2977
rect -8505 -2977 -8493 -2732
rect -8437 -2977 -8425 -2732
rect -8201 -2732 -8121 -2408
rect -7746 -2474 -7666 -2464
rect -7746 -2530 -7734 -2474
rect -7678 -2530 -7666 -2474
rect -7746 -2540 -7666 -2530
rect -8061 -2628 -7656 -2618
rect -8061 -2688 -8046 -2628
rect -7976 -2688 -7741 -2628
rect -7671 -2688 -7656 -2628
rect -8061 -2698 -7656 -2688
rect -8201 -2893 -8189 -2732
rect -8133 -2893 -8121 -2732
rect -7593 -2732 -7513 -2408
rect -8201 -2903 -8121 -2893
rect -7897 -2766 -7817 -2756
rect -8505 -2987 -8425 -2977
rect -7897 -2977 -7885 -2766
rect -7829 -2977 -7817 -2766
rect -7593 -2893 -7581 -2732
rect -7525 -2893 -7513 -2732
rect -7593 -2903 -7513 -2893
rect -7289 -2732 -7209 -2722
rect -7897 -3123 -7817 -2977
rect -7289 -2977 -7277 -2732
rect -7221 -2977 -7209 -2732
rect -7289 -2987 -7209 -2977
rect -6985 -2732 -6905 -2408
rect -6511 -2408 -6451 -2268
rect -6381 -2288 -6321 -2127
rect -6381 -2348 -6191 -2288
rect -6511 -2468 -6321 -2408
rect -6841 -2628 -6741 -2618
rect -6381 -2628 -6321 -2468
rect -6251 -2493 -6191 -2348
rect -6261 -2503 -6181 -2493
rect -6261 -2563 -6251 -2503
rect -6191 -2563 -6181 -2503
rect -6261 -2573 -6181 -2563
rect -6841 -2688 -6826 -2628
rect -6756 -2688 -6321 -2628
rect -6841 -2698 -6741 -2688
rect -6985 -2977 -6973 -2732
rect -6917 -2977 -6905 -2732
rect -6985 -2987 -6905 -2977
rect -6681 -2920 -6601 -2910
rect -6681 -2977 -6669 -2920
rect -6613 -2977 -6601 -2920
rect -6681 -3123 -6601 -2977
rect -9113 -3179 -6601 -3123
rect -6143 -3160 -6002 -3144
rect -9417 -3250 -6895 -3239
rect -9417 -3306 -6985 -3250
rect -6905 -3306 -6895 -3250
rect -6143 -3297 -6129 -3160
rect -9417 -3316 -6895 -3306
rect -10306 -3650 -10202 -3348
rect -10306 -3652 -8213 -3650
rect -10306 -3774 -8603 -3652
rect -8547 -3774 -8281 -3652
rect -8225 -3774 -8213 -3652
rect -10306 -3776 -8213 -3774
rect -8109 -3652 -8029 -3316
rect -6144 -3370 -6129 -3297
rect -6024 -3308 -6002 -3160
rect -6024 -3370 -6007 -3308
rect -6144 -3388 -6007 -3370
rect -8109 -3774 -8097 -3652
rect -8041 -3774 -8029 -3652
rect -8109 -3776 -8029 -3774
rect -10665 -4376 -10513 -4123
rect -10078 -4372 -9728 -3776
rect -6126 -4311 -6027 -3388
rect -6126 -4356 -6009 -4311
rect -6136 -4367 -6009 -4356
rect -11664 -4443 -11529 -4421
rect -11664 -4530 -11640 -4443
rect -11555 -4530 -11529 -4443
rect -10665 -4463 -10639 -4376
rect -10550 -4463 -10513 -4376
rect -10665 -4496 -10513 -4463
rect -10097 -4381 -9707 -4372
rect -11664 -4545 -11529 -4530
rect -10097 -4592 -10083 -4381
rect -9728 -4592 -9707 -4381
rect -10097 -4613 -9707 -4592
rect -6136 -4375 -6010 -4367
rect -6136 -4578 -6132 -4375
rect -6018 -4578 -6010 -4375
rect -5654 -4419 -5550 -1360
rect -5023 -3993 -4943 1344
rect -5035 -4003 -4931 -3993
rect -5035 -4083 -5023 -4003
rect -4943 -4083 -4931 -4003
rect -5035 -4093 -4931 -4083
rect -5665 -4429 -5537 -4419
rect -5665 -4531 -5654 -4429
rect -5550 -4531 -5537 -4429
rect -4764 -4439 -4655 1531
rect -4464 -4363 -2407 -4321
rect -5665 -4565 -5537 -4531
rect -4774 -4451 -4646 -4439
rect -4774 -4558 -4764 -4451
rect -4655 -4558 -4646 -4451
rect -6136 -4597 -6010 -4578
rect -4774 -4580 -4646 -4558
rect -4464 -4663 -4454 -4363
rect -2454 -4663 -2407 -4363
rect -4464 -4701 -2407 -4663
<< via2 >>
rect -13105 6820 -13049 6920
rect -4454 5134 -2454 5434
rect -12086 1317 -12006 1397
rect -11041 1043 -10961 1123
rect -10719 1043 -10639 1123
rect -10181 1043 -10101 1123
rect -9859 1043 -9779 1123
rect -9417 1043 -9337 1123
rect -8809 1043 -8729 1123
rect -8201 1043 -8121 1123
rect -7593 1043 -7513 1123
rect -6985 1043 -6905 1123
rect -6543 1043 -6463 1123
rect -6221 1043 -6141 1123
rect -9101 520 -9045 576
rect -8493 520 -8437 576
rect -8310 249 -8230 329
rect -7277 520 -7221 576
rect -7897 249 -7817 329
rect -5676 1847 -5596 1887
rect -5676 1807 -5596 1847
rect -5683 1043 -5603 1123
rect -5361 1043 -5281 1123
rect -8092 79 -8012 159
rect -8842 -215 -8762 -135
rect -7560 -215 -7480 -135
rect -9709 -1974 -9653 -1813
rect -9101 -1994 -9045 -1938
rect -8493 -1833 -8437 -1777
rect -8949 -2126 -8893 -2070
rect -9254 -2282 -9198 -2226
rect -7734 -2126 -7678 -2070
rect -8039 -2282 -7983 -2226
rect -7277 -2022 -7221 -1777
rect -6669 -1974 -6613 -1813
rect -8949 -2530 -8893 -2474
rect -9254 -2686 -9198 -2630
rect -9709 -2977 -9653 -2921
rect -9101 -2822 -9045 -2766
rect -8493 -2977 -8437 -2732
rect -7734 -2530 -7678 -2474
rect -8039 -2686 -7983 -2630
rect -7885 -2822 -7829 -2766
rect -7277 -2977 -7221 -2732
rect -6973 -2977 -6917 -2732
rect -6985 -3306 -6905 -3250
rect -4454 -4663 -2454 -4363
<< metal3 >>
rect -13115 6820 -13105 6920
rect -13049 6820 -12960 6920
rect -4464 5434 -2430 5477
rect -4464 5134 -4454 5434
rect -2454 5134 -2430 5434
rect -4464 5097 -2430 5134
rect -5696 1887 -5576 1907
rect -5696 1807 -5676 1887
rect -5596 1807 -5576 1887
rect -5696 1787 -5576 1807
rect -12096 1397 -11996 1417
rect -12096 1317 -12086 1397
rect -12006 1317 -11996 1397
rect -12096 1307 -11996 1317
rect -12086 1123 -12006 1307
rect -11051 1123 -10951 1133
rect -10729 1123 -10629 1133
rect -10191 1123 -10091 1133
rect -9869 1123 -9769 1133
rect -9427 1123 -9327 1133
rect -8211 1123 -8111 1243
rect -5676 1133 -5596 1787
rect -7603 1123 -7503 1133
rect -6995 1123 -6895 1133
rect -6553 1123 -6453 1133
rect -6231 1123 -6131 1133
rect -5693 1123 -5593 1133
rect -5371 1123 -5271 1133
rect -12086 1043 -11041 1123
rect -10961 1043 -10719 1123
rect -10639 1043 -10181 1123
rect -10101 1043 -9859 1123
rect -9779 1043 -9417 1123
rect -9337 1043 -8809 1123
rect -8729 1043 -8201 1123
rect -8121 1043 -7593 1123
rect -7513 1043 -6985 1123
rect -6905 1043 -6543 1123
rect -6463 1043 -6221 1123
rect -6141 1043 -5683 1123
rect -5603 1043 -5361 1123
rect -5281 1043 -5271 1123
rect -11051 1033 -10951 1043
rect -10729 1033 -10629 1043
rect -10191 1033 -10091 1043
rect -9869 1033 -9769 1043
rect -9427 1033 -9327 1043
rect -8819 1033 -8719 1043
rect -8211 1033 -8111 1043
rect -7603 1033 -7503 1043
rect -6995 1033 -6895 1043
rect -6553 1033 -6453 1043
rect -6231 1033 -6131 1043
rect -5693 1033 -5593 1043
rect -5371 1033 -5271 1043
rect -9113 576 -9033 586
rect -9113 520 -9101 576
rect -9045 520 -9033 576
rect -9113 510 -9033 520
rect -8505 576 -8425 586
rect -7289 576 -7209 586
rect -8505 520 -8493 576
rect -8437 520 -7277 576
rect -7221 520 -7209 576
rect -8505 510 -8425 520
rect -7289 510 -7209 520
rect -9101 329 -9045 510
rect -8320 329 -8220 339
rect -7907 329 -7807 339
rect -9101 249 -8310 329
rect -8230 249 -7897 329
rect -7817 249 -7807 329
rect -8852 -135 -8752 249
rect -8320 239 -8220 249
rect -7907 239 -7807 249
rect -8102 159 -8002 169
rect -8102 79 -8092 159
rect -8012 79 -8002 159
rect -8102 31 -8002 79
rect -8102 -49 -7480 31
rect -7560 -125 -7480 -49
rect -8852 -215 -8842 -135
rect -8762 -215 -8752 -135
rect -8852 -225 -8752 -215
rect -7570 -135 -7470 -125
rect -7570 -215 -7560 -135
rect -7480 -215 -7470 -135
rect -7570 -225 -7470 -215
rect -9721 -1777 -7209 -1767
rect -9721 -1813 -8493 -1777
rect -9721 -1974 -9709 -1813
rect -9653 -1833 -8493 -1813
rect -8437 -1833 -7277 -1777
rect -9653 -1843 -7277 -1833
rect -9653 -1974 -9641 -1843
rect -9721 -1984 -9641 -1974
rect -9113 -1938 -9033 -1928
rect -9714 -2408 -9649 -1984
rect -9113 -1994 -9101 -1938
rect -9045 -1994 -9033 -1938
rect -9266 -2226 -9186 -2216
rect -9266 -2282 -9254 -2226
rect -9198 -2282 -9186 -2226
rect -9266 -2292 -9186 -2282
rect -9113 -2292 -9033 -1994
rect -7289 -2022 -7277 -1843
rect -7221 -2022 -7209 -1777
rect -6681 -1813 -6601 -1803
rect -6681 -1974 -6669 -1813
rect -6613 -1974 -6601 -1813
rect -6681 -1984 -6601 -1974
rect -8971 -2070 -8871 -2058
rect -8971 -2126 -8949 -2070
rect -8893 -2126 -8871 -2070
rect -8971 -2138 -8871 -2126
rect -7756 -2070 -7656 -2058
rect -7756 -2126 -7734 -2070
rect -7678 -2126 -7656 -2070
rect -7756 -2138 -7656 -2126
rect -8051 -2226 -7971 -2216
rect -8051 -2282 -8039 -2226
rect -7983 -2282 -7971 -2226
rect -8051 -2292 -7971 -2282
rect -7289 -2292 -7209 -2022
rect -9113 -2352 -8425 -2292
rect -9714 -2468 -9033 -2408
rect -9276 -2630 -9176 -2618
rect -9276 -2686 -9254 -2630
rect -9198 -2686 -9176 -2630
rect -9276 -2698 -9176 -2686
rect -9113 -2766 -9033 -2468
rect -8961 -2474 -8881 -2464
rect -8961 -2530 -8949 -2474
rect -8893 -2530 -8881 -2474
rect -8961 -2540 -8881 -2530
rect -9113 -2822 -9101 -2766
rect -9045 -2822 -9033 -2766
rect -9113 -2832 -9033 -2822
rect -8505 -2732 -8425 -2352
rect -7897 -2352 -7209 -2292
rect -8061 -2630 -7961 -2618
rect -8061 -2686 -8039 -2630
rect -7983 -2686 -7961 -2630
rect -8061 -2698 -7961 -2686
rect -8505 -2911 -8493 -2732
rect -9721 -2921 -8493 -2911
rect -9721 -2977 -9709 -2921
rect -9653 -2977 -8493 -2921
rect -8437 -2911 -8425 -2732
rect -7897 -2766 -7817 -2352
rect -6674 -2408 -6609 -1984
rect -7746 -2474 -7666 -2464
rect -7746 -2530 -7734 -2474
rect -7678 -2530 -7666 -2474
rect -7746 -2540 -7666 -2530
rect -7289 -2468 -6609 -2408
rect -7897 -2822 -7885 -2766
rect -7829 -2822 -7817 -2766
rect -7897 -2832 -7817 -2822
rect -7289 -2732 -7209 -2468
rect -7289 -2911 -7277 -2732
rect -8437 -2977 -7277 -2911
rect -7221 -2977 -7209 -2732
rect -9721 -2987 -7209 -2977
rect -6985 -2732 -6905 -2722
rect -6985 -2977 -6973 -2732
rect -6917 -2977 -6905 -2732
rect -6985 -3239 -6905 -2977
rect -6995 -3250 -6895 -3239
rect -6995 -3306 -6985 -3250
rect -6905 -3306 -6895 -3250
rect -6995 -3316 -6895 -3306
rect -4464 -4363 -2407 -4321
rect -4464 -4663 -4454 -4363
rect -2454 -4663 -2407 -4363
rect -4464 -4701 -2407 -4663
<< via3 >>
rect -4454 5134 -2454 5434
rect -9254 -2282 -9198 -2226
rect -8949 -2126 -8893 -2070
rect -7734 -2126 -7678 -2070
rect -8039 -2282 -7983 -2226
rect -9254 -2686 -9198 -2630
rect -8949 -2530 -8893 -2474
rect -8039 -2686 -7983 -2630
rect -7734 -2530 -7678 -2474
rect -4454 -4663 -2454 -4363
<< metal4 >>
rect -4464 5434 -2430 5477
rect -4464 5134 -4454 5434
rect -2454 5134 -2430 5434
rect -4464 5097 -2430 5134
rect -8971 -2070 -8871 -2058
rect -8971 -2126 -8949 -2070
rect -8893 -2126 -8871 -2070
rect -8971 -2138 -8871 -2126
rect -7756 -2070 -7656 -2058
rect -7756 -2126 -7734 -2070
rect -7678 -2126 -7656 -2070
rect -7756 -2138 -7656 -2126
rect -9266 -2226 -9186 -2216
rect -9266 -2282 -9254 -2226
rect -9198 -2282 -9186 -2226
rect -9266 -2292 -9186 -2282
rect -9254 -2618 -9198 -2292
rect -8949 -2464 -8893 -2138
rect -8051 -2226 -7971 -2216
rect -8051 -2282 -8039 -2226
rect -7983 -2282 -7971 -2226
rect -8051 -2292 -7971 -2282
rect -8961 -2474 -8881 -2464
rect -8961 -2530 -8949 -2474
rect -8893 -2530 -8881 -2474
rect -8961 -2540 -8881 -2530
rect -8039 -2618 -7983 -2292
rect -7734 -2464 -7678 -2138
rect -7746 -2474 -7666 -2464
rect -7746 -2530 -7734 -2474
rect -7678 -2530 -7666 -2474
rect -7746 -2540 -7666 -2530
rect -9276 -2630 -9176 -2618
rect -9276 -2686 -9254 -2630
rect -9198 -2686 -9176 -2630
rect -9276 -2698 -9176 -2686
rect -8061 -2630 -7961 -2618
rect -8061 -2686 -8039 -2630
rect -7983 -2686 -7961 -2630
rect -8061 -2698 -7961 -2686
rect -4464 -4322 30646 -4321
rect 32519 -4322 34291 5770
rect -4464 -4363 34291 -4322
rect -4464 -4663 -4454 -4363
rect -2454 -4663 34291 -4363
rect -4464 -4701 34291 -4663
rect 30646 -4702 34291 -4701
<< via4 >>
rect -4454 5134 -2454 5434
<< metal5 >>
rect 22821 5477 24776 5770
rect -4464 5434 24776 5477
rect -4464 5134 -4454 5434
rect -2454 5134 24776 5434
rect -4464 5097 24776 5134
rect 22821 -4206 24776 5097
<< labels >>
rlabel metal2 -13233 15938 -13233 15938 7 Reset
port 6 w
rlabel metal2 -13224 16448 -13224 16448 7 SAR_in
port 7 w
rlabel metal2 -13170 27549 -13170 27549 7 Load
port 8 w
rlabel metal2 4077 38603 4077 38603 1 Piso_out
port 10 n
rlabel metal2 -8063 38726 -8063 38726 1 Clk_piso
port 9 n
rlabel metal2 -13260 6872 -13260 6872 7 SARlogic_0.clk
rlabel metal2 -12988 15939 -12988 15939 7 SARlogic_0.reset
rlabel metal2 -12988 16447 -12988 16447 7 SARlogic_0.comp_in
rlabel metal2 -13784 -4047 -13784 -4047 7 Clk
port 2 w
rlabel metal5 24711 -4206 24711 -4206 5 Vdd
port 0 s
rlabel metal4 34239 -4702 34239 -4702 5 Vss
port 1 s
rlabel metal2 -13880 -2213 -13880 -2213 7 Vin1
port 3 w
rlabel metal2 -13878 -2540 -13878 -2540 7 Vin2
port 4 w
rlabel metal2 -13894 3909 -13894 3909 7 Comp_out
port 5 w
<< end >>
