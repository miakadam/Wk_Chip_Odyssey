magic
tech gf180mcuD
magscale 1 10
timestamp 1757046296
<< pwell >>
rect 9945 3495 10040 3814
rect 13040 3485 13135 3804
rect 13055 3235 13120 3250
rect 10430 3135 10520 3205
rect 10430 3125 10520 3130
rect 10588 2140 10668 2235
<< polysilicon >>
rect 10430 3135 10520 3205
rect 10430 3125 10520 3130
<< metal1 >>
rect 10588 3486 10668 3496
rect 9900 3260 9960 3485
rect 10025 3260 10035 3485
rect 9900 3255 10035 3260
rect 10284 3402 10364 3412
rect 10284 3241 10296 3402
rect 10352 3241 10364 3402
rect 10588 3269 10600 3486
rect 10656 3269 10668 3486
rect 11196 3486 11276 3496
rect 11196 3430 11208 3486
rect 11264 3430 11276 3486
rect 11196 3420 11276 3430
rect 11804 3486 11884 3496
rect 11804 3430 11816 3486
rect 11872 3430 11884 3486
rect 11804 3420 11884 3430
rect 12412 3486 12492 3496
rect 10588 3261 10668 3269
rect 10892 3402 10972 3412
rect 10284 3231 10364 3241
rect 10892 3241 10904 3402
rect 10960 3241 10972 3402
rect 10892 3231 10972 3241
rect 11500 3402 11580 3412
rect 11500 3241 11512 3402
rect 11568 3241 11580 3402
rect 11500 3231 11580 3241
rect 12108 3402 12188 3412
rect 12108 3241 12120 3402
rect 12176 3241 12188 3402
rect 12108 3231 12188 3241
rect 12412 3241 12424 3486
rect 12480 3241 12492 3486
rect 12412 3231 12492 3241
rect 12716 3402 12796 3412
rect 12716 3241 12728 3402
rect 12784 3241 12796 3402
rect 13045 3260 13055 3485
rect 13120 3260 13180 3485
rect 13045 3255 13180 3260
rect 12716 3231 12796 3241
rect 10425 3140 10440 3195
rect 10075 3085 10270 3140
rect 10380 3135 10440 3140
rect 10510 3140 10525 3195
rect 10510 3135 10565 3140
rect 10730 3135 10745 3195
rect 10815 3135 10830 3195
rect 10985 3085 11180 3140
rect 11290 3085 11485 3140
rect 11640 3135 11655 3195
rect 11725 3135 11740 3195
rect 11945 3135 11960 3195
rect 12030 3135 12045 3195
rect 12205 3085 12400 3140
rect 12505 3085 12700 3140
rect 12860 3135 12875 3195
rect 12945 3135 12960 3195
rect 10075 3070 13670 3085
rect 10075 3010 13190 3070
rect 13250 3010 13670 3070
rect 10075 2700 13450 2760
rect 13510 2700 13670 2760
rect 10075 2685 13670 2700
rect 10075 2635 10270 2685
rect 10985 2635 11180 2685
rect 11290 2635 11485 2685
rect 12200 2635 12395 2685
rect 12505 2635 12700 2685
rect 10430 2590 10440 2635
rect 10425 2575 10440 2590
rect 10510 2590 10520 2635
rect 10735 2590 10745 2635
rect 10510 2575 10525 2590
rect 10730 2575 10745 2590
rect 10815 2590 10825 2635
rect 11645 2590 11655 2635
rect 10815 2575 10830 2590
rect 11640 2575 11655 2590
rect 11725 2590 11735 2635
rect 11950 2590 11960 2635
rect 11725 2575 11740 2590
rect 11945 2575 11960 2590
rect 12030 2590 12040 2635
rect 12865 2590 12875 2635
rect 12030 2575 12045 2590
rect 12860 2575 12875 2590
rect 12945 2590 12955 2635
rect 12945 2575 12960 2590
rect 10284 2531 10364 2541
rect 10284 2370 10296 2531
rect 10352 2370 10364 2531
rect 10892 2531 10972 2541
rect 10284 2360 10364 2370
rect 10588 2497 10668 2507
rect 9980 2342 10060 2352
rect 9980 2286 9992 2342
rect 10048 2286 10060 2342
rect 9980 2276 10060 2286
rect 10588 2286 10600 2497
rect 10656 2286 10668 2497
rect 10892 2370 10904 2531
rect 10960 2370 10972 2531
rect 10892 2360 10972 2370
rect 11196 2531 11276 2541
rect 10588 2276 10668 2286
rect 11196 2286 11208 2531
rect 11264 2286 11276 2531
rect 11500 2531 11580 2541
rect 11500 2370 11512 2531
rect 11568 2370 11580 2531
rect 12108 2531 12188 2541
rect 11500 2360 11580 2370
rect 11804 2497 11884 2507
rect 11196 2276 11276 2286
rect 11804 2286 11816 2497
rect 11872 2286 11884 2497
rect 12108 2370 12120 2531
rect 12176 2370 12188 2531
rect 12108 2360 12188 2370
rect 12412 2531 12492 2541
rect 11804 2276 11884 2286
rect 12412 2286 12424 2531
rect 12480 2286 12492 2531
rect 12412 2276 12492 2286
rect 12716 2531 12796 2541
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2276 12796 2286
rect 13020 2343 13100 2353
rect 13020 2286 13032 2343
rect 13088 2286 13100 2343
rect 13020 2276 13100 2286
<< via1 >>
rect 9960 3260 10025 3485
rect 10296 3241 10352 3402
rect 10600 3269 10656 3486
rect 11208 3430 11264 3486
rect 11816 3430 11872 3486
rect 10904 3241 10960 3402
rect 11512 3241 11568 3402
rect 12120 3241 12176 3402
rect 12424 3241 12480 3486
rect 12728 3241 12784 3402
rect 13055 3260 13120 3485
rect 10440 3135 10510 3195
rect 10745 3135 10815 3195
rect 11655 3135 11725 3195
rect 11960 3135 12030 3195
rect 12875 3135 12945 3195
rect 13190 3010 13250 3070
rect 13450 2700 13510 2760
rect 10440 2575 10510 2635
rect 10745 2575 10815 2635
rect 11655 2575 11725 2635
rect 11960 2575 12030 2635
rect 12875 2575 12945 2635
rect 10296 2370 10352 2531
rect 9992 2286 10048 2342
rect 10600 2286 10656 2497
rect 10904 2370 10960 2531
rect 11208 2286 11264 2531
rect 11512 2370 11568 2531
rect 11816 2286 11872 2497
rect 12120 2370 12176 2531
rect 12424 2286 12480 2531
rect 12728 2286 12784 2531
rect 13032 2286 13088 2343
<< metal2 >>
rect 9945 3485 10040 3814
rect 13040 3688 13135 3804
rect 9945 3260 9960 3485
rect 10025 3260 10040 3485
rect 10588 3632 13135 3688
rect 10588 3486 10668 3632
rect 9945 3255 10040 3260
rect 10284 3402 10364 3412
rect 10284 3241 10296 3402
rect 10352 3241 10364 3402
rect 10588 3269 10600 3486
rect 10656 3269 10668 3486
rect 11196 3486 11276 3496
rect 11196 3430 11208 3486
rect 11264 3430 11276 3486
rect 11196 3420 11276 3430
rect 11804 3486 11884 3632
rect 11804 3430 11816 3486
rect 11872 3430 11884 3486
rect 11804 3420 11884 3430
rect 12412 3486 12492 3496
rect 10588 3261 10668 3269
rect 10892 3402 10972 3412
rect 10284 2911 10364 3241
rect 10892 3241 10904 3402
rect 10960 3241 10972 3402
rect 10425 3195 10830 3205
rect 10425 3135 10440 3195
rect 10510 3135 10745 3195
rect 10815 3135 10830 3195
rect 10425 3125 10830 3135
rect 10892 2911 10972 3241
rect 11500 3402 11580 3412
rect 11500 3241 11512 3402
rect 11568 3241 11580 3402
rect 11500 2911 11580 3241
rect 12108 3402 12188 3412
rect 12108 3241 12120 3402
rect 12176 3241 12188 3402
rect 11640 3195 12045 3205
rect 11640 3135 11655 3195
rect 11725 3135 11960 3195
rect 12030 3135 12045 3195
rect 11640 3125 12045 3135
rect 12108 2911 12188 3241
rect 12412 3241 12424 3486
rect 12480 3241 12492 3486
rect 13040 3485 13135 3632
rect 12412 3231 12492 3241
rect 12716 3402 12796 3412
rect 12716 3241 12728 3402
rect 12784 3241 12796 3402
rect 13040 3260 13055 3485
rect 13120 3260 13135 3485
rect 13040 3255 13135 3260
rect 12716 2911 12796 3241
rect 12860 3195 12960 3205
rect 13154 3195 13380 3196
rect 12860 3135 12875 3195
rect 12945 3136 13380 3195
rect 12945 3135 13119 3136
rect 12860 3125 12960 3135
rect 13175 3070 13260 3080
rect 13175 3010 13190 3070
rect 13250 3010 13260 3070
rect 13175 2995 13260 3010
rect 10284 2855 12796 2911
rect 10284 2531 10364 2855
rect 10425 2635 10830 2645
rect 10425 2575 10440 2635
rect 10510 2575 10745 2635
rect 10815 2575 10830 2635
rect 10425 2565 10830 2575
rect 10284 2370 10296 2531
rect 10352 2370 10364 2531
rect 10892 2531 10972 2855
rect 9980 2342 10060 2352
rect 9980 2286 9992 2342
rect 10048 2286 10060 2342
rect 9980 2276 10060 2286
rect 10284 2024 10364 2370
rect 10588 2497 10668 2507
rect 10588 2286 10600 2497
rect 10656 2286 10668 2497
rect 10892 2370 10904 2531
rect 10960 2370 10972 2531
rect 10892 2360 10972 2370
rect 11196 2531 11276 2541
rect 10588 2140 10668 2286
rect 11196 2286 11208 2531
rect 11264 2286 11276 2531
rect 11500 2531 11580 2855
rect 11640 2635 12045 2645
rect 11640 2575 11655 2635
rect 11725 2575 11960 2635
rect 12030 2575 12045 2635
rect 11640 2565 12045 2575
rect 11500 2370 11512 2531
rect 11568 2370 11580 2531
rect 12108 2531 12188 2855
rect 11500 2360 11580 2370
rect 11804 2497 11884 2507
rect 11196 2276 11276 2286
rect 11804 2286 11816 2497
rect 11872 2286 11884 2497
rect 12108 2370 12120 2531
rect 12176 2370 12188 2531
rect 12108 2360 12188 2370
rect 12412 2531 12492 2541
rect 11804 2140 11884 2286
rect 12412 2286 12424 2531
rect 12480 2286 12492 2531
rect 12412 2276 12492 2286
rect 12716 2531 12796 2855
rect 13190 2855 13250 2995
rect 13320 2975 13380 3136
rect 13320 2915 13510 2975
rect 13190 2795 13380 2855
rect 12860 2635 12960 2645
rect 13320 2635 13380 2795
rect 13450 2770 13510 2915
rect 13440 2760 13520 2770
rect 13440 2700 13450 2760
rect 13510 2700 13520 2760
rect 13440 2690 13520 2700
rect 12860 2575 12875 2635
rect 12945 2575 13380 2635
rect 12860 2565 12960 2575
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2276 12796 2286
rect 13020 2343 13100 2353
rect 13020 2286 13032 2343
rect 13088 2286 13100 2343
rect 13020 2140 13100 2286
rect 10588 2084 13100 2140
rect 10284 2013 12806 2024
rect 10284 1957 12716 2013
rect 12796 1957 12806 2013
rect 10284 1947 12806 1957
<< via2 >>
rect 9960 3260 10025 3485
rect 10600 3269 10656 3325
rect 11208 3430 11264 3486
rect 12424 3241 12480 3486
rect 13055 3260 13120 3485
rect 9992 2286 10048 2342
rect 10600 2441 10656 2497
rect 11208 2286 11264 2531
rect 11816 2441 11872 2497
rect 12424 2286 12480 2531
rect 12728 2286 12784 2531
rect 12716 1957 12796 2013
<< metal3 >>
rect 10035 3486 12492 3496
rect 10035 3485 11208 3486
rect 9950 3260 9960 3485
rect 10025 3430 11208 3485
rect 11264 3430 12424 3486
rect 10025 3420 12424 3430
rect 10025 3260 10035 3420
rect 10588 3325 10668 3335
rect 10588 3269 10600 3325
rect 10656 3269 10668 3325
rect 9960 2855 10025 3260
rect 10588 2971 10668 3269
rect 12412 3241 12424 3420
rect 12480 3241 12492 3486
rect 13045 3260 13055 3485
rect 13120 3260 13130 3485
rect 13045 3255 13130 3260
rect 12412 2971 12492 3241
rect 10588 2911 11276 2971
rect 9960 2795 10668 2855
rect 10588 2497 10668 2795
rect 10588 2441 10600 2497
rect 10656 2441 10668 2497
rect 10588 2431 10668 2441
rect 11196 2531 11276 2911
rect 11196 2352 11208 2531
rect 9980 2342 11208 2352
rect 9980 2286 9992 2342
rect 10048 2286 11208 2342
rect 11264 2352 11276 2531
rect 11804 2911 12492 2971
rect 11804 2497 11884 2911
rect 13055 2855 13120 3255
rect 11804 2441 11816 2497
rect 11872 2441 11884 2497
rect 11804 2431 11884 2441
rect 12412 2795 13120 2855
rect 12412 2531 12492 2795
rect 12412 2352 12424 2531
rect 11264 2286 12424 2352
rect 12480 2286 12492 2531
rect 9980 2276 12492 2286
rect 12716 2531 12796 2541
rect 12716 2286 12728 2531
rect 12784 2286 12796 2531
rect 12716 2024 12796 2286
rect 12706 2013 12806 2024
rect 12706 1957 12716 2013
rect 12796 1957 12806 2013
rect 12706 1947 12806 1957
use nfet_03v3_RPTYYZ  nfet_03v3_RPTYYZ_0
timestamp 1756981609
transform 1 0 12300 0 1 3366
box -820 -266 820 266
use nfet_03v3_RPTYYZ  XM9
timestamp 1756981609
transform 1 0 10780 0 1 2406
box -820 -266 820 266
use nfet_03v3_RPTYYZ  XM10
timestamp 1756981609
transform 1 0 12300 0 1 2406
box -820 -266 820 266
use nfet_03v3_RPTYYZ  XM20
timestamp 1756981609
transform 1 0 10780 0 1 3366
box -820 -266 820 266
<< labels >>
rlabel metal2 11592 1947 11592 1947 5 VSS
port 2 s
rlabel metal1 13668 2721 13668 2721 3 Vin1
port 1 e
rlabel metal2 13092 3804 13092 3804 1 Vd1
port 3 n
rlabel metal2 9996 3813 9996 3813 1 Vd2
port 4 n
rlabel metal1 13668 3048 13668 3048 3 Vin2
port 5 e
<< end >>
