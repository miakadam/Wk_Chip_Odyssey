magic
tech gf180mcuD
magscale 1 10
timestamp 1758001989
<< nwell >>
rect 2812 -216 3016 -163
rect 2050 -265 2053 -262
<< pwell >>
rect 3030 -692 3110 -510
rect 2906 -768 3110 -692
<< nsubdiff >>
rect 2050 -265 2053 -262
<< metal1 >>
rect 1780 700 3268 900
rect 1817 571 1863 700
rect 2032 569 2128 600
rect 2236 569 2332 600
rect 2501 571 2547 700
rect 2716 569 2812 600
rect 2920 569 3016 600
rect 3185 571 3231 700
rect 1862 -108 1957 488
rect 2142 237 2154 477
rect 2210 237 2222 477
rect 2408 -108 2503 488
rect 2826 237 2838 477
rect 2894 237 2906 477
rect 2622 -97 2634 143
rect 2690 -97 2702 143
rect 3030 -97 3042 143
rect 3098 -97 3110 143
rect 2128 -189 2332 -163
rect 2812 -189 3016 -163
rect 2032 -216 2332 -189
rect 2716 -216 3016 -189
rect 2032 -264 2128 -216
rect 2032 -320 2052 -264
rect 2108 -320 2128 -264
rect 2032 -551 2128 -320
rect 2716 -420 2812 -216
rect 2716 -476 2736 -420
rect 2792 -476 2812 -420
rect 1938 -702 2018 -692
rect 1938 -758 1950 -702
rect 2006 -758 2018 -702
rect 1938 -768 2018 -758
rect 2204 -828 2301 -632
rect 1817 -1040 1863 -911
rect 2032 -940 2128 -909
rect 2343 -1040 2501 -549
rect 2716 -551 2812 -476
rect 2546 -828 2643 -632
rect 2826 -702 2906 -692
rect 2826 -758 2838 -702
rect 2894 -758 2906 -702
rect 2826 -768 2906 -758
rect 2716 -940 2812 -909
rect 2981 -1040 3027 -911
rect 1780 -1240 3064 -1040
<< via1 >>
rect 2154 237 2210 477
rect 2838 237 2894 477
rect 2634 -97 2690 143
rect 3042 -97 3098 143
rect 2052 -320 2108 -264
rect 2736 -476 2792 -420
rect 1950 -758 2006 -702
rect 2838 -758 2894 -702
<< metal2 >>
rect 2142 477 2906 487
rect 2142 237 2154 477
rect 2210 237 2838 477
rect 2894 237 2906 477
rect 2142 227 2906 237
rect 2622 143 3110 153
rect 2622 -97 2634 143
rect 2690 -97 3042 143
rect 3098 -97 3110 143
rect 2622 -107 3110 -97
rect 2032 -264 2128 -252
rect 1724 -320 2052 -264
rect 2108 -320 2128 -264
rect 2032 -332 2128 -320
rect 3030 -342 3110 -107
rect 3030 -398 3268 -342
rect 2716 -420 2812 -410
rect 1724 -476 2736 -420
rect 2792 -476 2812 -420
rect 2716 -486 2812 -476
rect 3030 -692 3110 -398
rect 1938 -702 3110 -692
rect 1938 -758 1950 -702
rect 2006 -758 2838 -702
rect 2894 -758 3110 -702
rect 1938 -768 3110 -758
use nfet_03v3_EKBWUP  nfet_03v3_EKBWUP_0
timestamp 1758001983
transform 1 0 2764 0 1 -730
box -300 -310 300 310
use pfet_03v3_LJLJK4  pfet_03v3_LJLJK4_0
timestamp 1758001983
transform 1 0 2866 0 1 190
box -402 -510 402 510
use nfet_03v3_EKBWUP  XM1
timestamp 1758001983
transform 1 0 2080 0 1 -730
box -300 -310 300 310
use pfet_03v3_LJLJK4  XM3
timestamp 1758001983
transform 1 0 2182 0 1 190
box -402 -510 402 510
<< labels >>
rlabel metal1 2525 900 2525 900 1 VDD
port 0 n
rlabel metal1 2418 -1240 2418 -1240 5 VSS
port 1 s
rlabel metal2 3268 -371 3268 -371 3 OUT
port 2 e
rlabel metal2 1724 -291 1724 -291 7 A
port 3 w
rlabel metal2 1724 -448 1724 -448 7 B
port 4 w
<< end >>
