magic
tech gf180mcuD
magscale 1 10
timestamp 1757405367
<< error_p >>
rect -222 113 -211 159
rect -38 113 -27 159
rect 146 113 157 159
rect -222 -159 -211 -113
rect -38 -159 -27 -113
rect 146 -159 157 -113
<< pwell >>
rect -474 -290 474 290
<< nmos >>
rect -224 -80 -144 80
rect -40 -80 40 80
rect 144 -80 224 80
<< ndiff >>
rect -312 67 -224 80
rect -312 -67 -299 67
rect -253 -67 -224 67
rect -312 -80 -224 -67
rect -144 67 -40 80
rect -144 -67 -115 67
rect -69 -67 -40 67
rect -144 -80 -40 -67
rect 40 67 144 80
rect 40 -67 69 67
rect 115 -67 144 67
rect 40 -80 144 -67
rect 224 67 312 80
rect 224 -67 253 67
rect 299 -67 312 67
rect 224 -80 312 -67
<< ndiffc >>
rect -299 -67 -253 67
rect -115 -67 -69 67
rect 69 -67 115 67
rect 253 -67 299 67
<< psubdiff >>
rect -450 194 450 266
rect -450 150 -378 194
rect -450 -150 -437 150
rect -391 -150 -378 150
rect 378 150 450 194
rect -450 -194 -378 -150
rect 378 -150 391 150
rect 437 -150 450 150
rect 378 -194 450 -150
rect -450 -266 450 -194
<< psubdiffcont >>
rect -437 -150 -391 150
rect 391 -150 437 150
<< polysilicon >>
rect -224 159 -144 172
rect -224 113 -211 159
rect -157 113 -144 159
rect -224 80 -144 113
rect -40 159 40 172
rect -40 113 -27 159
rect 27 113 40 159
rect -40 80 40 113
rect 144 159 224 172
rect 144 113 157 159
rect 211 113 224 159
rect 144 80 224 113
rect -224 -113 -144 -80
rect -224 -159 -211 -113
rect -157 -159 -144 -113
rect -224 -172 -144 -159
rect -40 -113 40 -80
rect -40 -159 -27 -113
rect 27 -159 40 -113
rect -40 -172 40 -159
rect 144 -113 224 -80
rect 144 -159 157 -113
rect 211 -159 224 -113
rect 144 -172 224 -159
<< polycontact >>
rect -211 113 -157 159
rect -27 113 27 159
rect 157 113 211 159
rect -211 -159 -157 -113
rect -27 -159 27 -113
rect 157 -159 211 -113
<< metal1 >>
rect -437 207 437 253
rect -437 150 -391 207
rect -222 113 -211 159
rect -157 113 -146 159
rect -38 113 -27 159
rect 27 113 38 159
rect 146 113 157 159
rect 211 113 222 159
rect 391 150 437 207
rect -299 67 -253 78
rect -299 -78 -253 -67
rect -115 67 -69 78
rect -115 -78 -69 -67
rect 69 67 115 78
rect 69 -78 115 -67
rect 253 67 299 78
rect 253 -78 299 -67
rect -437 -207 -391 -150
rect -222 -159 -211 -113
rect -157 -159 -146 -113
rect -38 -159 -27 -113
rect 27 -159 38 -113
rect 146 -159 157 -113
rect 211 -159 222 -113
rect 391 -207 437 -150
rect -437 -253 437 -207
<< properties >>
string FIXED_BBOX -414 -230 414 230
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.8 l 0.4 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
