* SPICE3 file created from 2inmux.ext - technology: (null)

.option scale=5n

X0 a_256_1130.t1 Load.t0 VDD.t21 VDD.t20 pfet_03v3
X1 VSS.t19 or2_0.A a_2484_n766 VSS.t18 nfet_03v3
X2 a_2672_n46 or2_0.B a_2484_n766 VDD.t11 pfet_03v3
X3 a_444_n1930 In.t0 a_256_n1210.t3 VSS.t9 nfet_03v3
X4 a_444_410 Bit.t0 VSS.t15 VSS.t14 nfet_03v3
X5 a_2484_n766 or2_0.B a_2672_n46 VDD.t10 pfet_03v3
X6 OUT.t0 a_2484_n766 VDD.t5 VDD.t4 pfet_03v3
X7 VSS.t17 Bit.t1 a_444_410 VSS.t16 nfet_03v3
X8 a_2672_n46 or2_0.A VDD.t17 VDD.t16 pfet_03v3
X9 a_256_n1210.t1 In.t1 VDD.t13 VDD.t12 pfet_03v3
X10 a_2484_n766 or2_0.B VSS.t11 VSS.t10 nfet_03v3
X11 VSS.t7 inv2_0.out a_444_n1930 VSS.t6 nfet_03v3
X12 or2_0.B a_256_n1210.t4 VDD.t3 VDD.t2 pfet_03v3
X13 VDD.t15 or2_0.A a_2672_n46 VDD.t14 pfet_03v3
X14 a_444_410 Load.t1 a_256_1130.t3 VSS.t23 nfet_03v3
X15 inv2_0.out Load.t2 VSS.t22 VSS.t21 nfet_03v3
X16 OUT.t1 a_2484_n766 VSS.t1 VSS.t0 nfet_03v3
X17 VDD.t1 Bit.t2 a_256_1130.t0 VDD.t0 pfet_03v3
X18 or2_0.A a_256_1130.t4 VDD.t9 VDD.t8 pfet_03v3
X19 a_256_1130.t2 Load.t3 a_444_410 VSS.t20 nfet_03v3
X20 or2_0.A a_256_1130.t5 VSS.t13 VSS.t12 nfet_03v3
X21 VDD.t7 inv2_0.out a_256_n1210.t0 VDD.t6 pfet_03v3
X22 a_256_n1210.t2 In.t2 a_444_n1930 VSS.t8 nfet_03v3
X23 or2_0.B a_256_n1210.t5 VSS.t3 VSS.t2 nfet_03v3
X24 a_444_n1930 inv2_0.out VSS.t5 VSS.t4 nfet_03v3
X25 inv2_0.out Load.t4 VDD.t19 VDD.t18 pfet_03v3
R0 Load.n1 Load.t0 34.2529
R1 Load.n2 Load.t4 34.1797
R2 Load.n0 Load.t1 19.673
R3 Load.n2 Load.t2 19.5798
R4 Load.n0 Load.t3 19.4007
R5 and2_0.B Load.n1 6.45093
R6 inv2_0.in Load.n2 4.87271
R7 Load.n3 inv2_0.in 2.20229
R8 and2_0.B Load.n3 1.42121
R9 Load.n3 Load 0.2255
R10 Load.n1 Load.n0 0.106438
R11 VDD.n37 VDD.t8 236.083
R12 VDD.t20 VDD.n34 236.083
R13 VDD.t2 VDD.n17 236.083
R14 VDD.n23 VDD.t12 236.083
R15 VDD.n15 VDD.t4 236.083
R16 VDD.n9 VDD.t16 236.083
R17 VDD.t8 VDD.n36 235.294
R18 VDD.n36 VDD.t20 235.294
R19 VDD.n22 VDD.t2 235.294
R20 VDD.t12 VDD.n22 235.294
R21 VDD.t4 VDD.n14 235.294
R22 VDD.n14 VDD.t10 235.294
R23 VDD.t11 VDD.n12 235.294
R24 VDD.n12 VDD.t14 235.294
R25 VDD.t10 VDD.t11 200
R26 VDD.t16 VDD.t14 200
R27 VDD.n1 VDD.t0 131.589
R28 VDD.n25 VDD.t6 131.589
R29 VDD.n42 VDD.t18 118.543
R30 VDD.n9 VDD.n8 96.0755
R31 VDD.n10 VDD.n9 96.0755
R32 VDD.n19 VDD.n17 78.2255
R33 VDD.n23 VDD.n19 78.2255
R34 VDD.n23 VDD.n20 78.2255
R35 VDD.n20 VDD.n17 78.2255
R36 VDD.n15 VDD.n6 78.2255
R37 VDD.n15 VDD.n7 78.2255
R38 VDD.n37 VDD.n32 78.2255
R39 VDD.n37 VDD.n33 78.2255
R40 VDD.n34 VDD.n32 78.2255
R41 VDD.n34 VDD.n33 78.2255
R42 VDD.n8 VDD.n6 59.8505
R43 VDD.n10 VDD.n7 59.8505
R44 VDD.n21 VDD.n19 36.2255
R45 VDD.n21 VDD.n20 36.2255
R46 VDD.n11 VDD.n8 36.2255
R47 VDD.n11 VDD.n10 36.2255
R48 VDD.n13 VDD.n6 36.2255
R49 VDD.n13 VDD.n7 36.2255
R50 VDD.n35 VDD.n32 36.2255
R51 VDD.n35 VDD.n33 36.2255
R52 VDD.n29 VDD.n28 2.49936
R53 VDD.n28 VDD.n17 1.93883
R54 VDD.n16 VDD.n15 1.81722
R55 VDD.n38 VDD.n37 1.78583
R56 VDD.n42 VDD.t19 1.74654
R57 VDD.n1 VDD.t1 1.49467
R58 VDD.n25 VDD.t7 1.49467
R59 VDD.n24 VDD.t13 1.49467
R60 VDD.n0 VDD.t21 1.49467
R61 VDD.n18 VDD.t3 1.47383
R62 VDD.n3 VDD.t17 1.47383
R63 VDD.n4 VDD.t15 1.47383
R64 VDD.n5 VDD.t5 1.47383
R65 VDD.n2 VDD.t9 1.47383
R66 VDD.n21 VDD.n18 0.788
R67 VDD.n22 VDD.n21 0.788
R68 VDD.n24 VDD.n23 0.788
R69 VDD.n11 VDD.n4 0.788
R70 VDD.n12 VDD.n11 0.788
R71 VDD.n13 VDD.n5 0.788
R72 VDD.n14 VDD.n13 0.788
R73 VDD.n9 VDD.n3 0.788
R74 VDD.n35 VDD.n2 0.788
R75 VDD.n36 VDD.n35 0.788
R76 VDD.n34 VDD.n0 0.788
R77 VDD.n27 VDD.n18 0.561043
R78 VDD.n31 VDD.n3 0.561043
R79 VDD.n30 VDD.n4 0.561043
R80 VDD.n16 VDD.n5 0.561043
R81 VDD.n39 VDD.n2 0.561043
R82 VDD.n41 VDD.n40 0.415037
R83 inv2_0.vdd VDD.n42 0.313534
R84 VDD.n27 VDD.n26 0.255737
R85 VDD.n40 VDD.n39 0.255737
R86 VDD.n39 VDD.n38 0.2165
R87 inv2_0.vdd VDD.n41 0.1985
R88 VDD.n38 VDD.n31 0.148424
R89 VDD.n28 VDD.n27 0.0635
R90 VDD.n31 VDD.n30 0.0452384
R91 VDD.n26 VDD.n24 0.0313054
R92 VDD.n26 VDD.n25 0.0313054
R93 VDD.n40 VDD.n0 0.0313054
R94 VDD.n40 VDD.n1 0.0313054
R95 VDD.n29 VDD.n16 0.0295407
R96 VDD.n30 or2_0.VDD 0.0157398
R97 VDD.n41 VDD 0.0155
R98 or2_0.VDD VDD.n29 0.000957849
R99 a_256_1130.n0 a_256_1130.t4 34.1797
R100 a_256_1130.n0 a_256_1130.t5 19.5798
R101 a_256_1130.n1 a_256_1130.t3 18.7717
R102 a_256_1130.n1 a_256_1130.t2 9.2885
R103 a_256_1130.n2 a_256_1130.n0 4.93379
R104 a_256_1130.t0 a_256_1130.n3 4.23346
R105 a_256_1130.n3 a_256_1130.t1 3.85546
R106 a_256_1130.n2 a_256_1130.n1 0.4055
R107 a_256_1130.n3 a_256_1130.n2 0.352625
R108 VSS.n19 VSS.n17 60109.5
R109 VSS.n17 VSS.n16 24900
R110 VSS.n36 VSS.n35 19475
R111 VSS.n16 VSS.n12 17479.3
R112 VSS.n52 VSS.n12 16004
R113 VSS.n36 VSS.n17 14900
R114 VSS.n43 VSS.n16 12638.9
R115 VSS.n44 VSS.n43 11510.4
R116 VSS.n35 VSS.n34 7486.96
R117 VSS.n57 VSS.n56 1105.44
R118 VSS.n34 VSS.t2 847.827
R119 VSS.n45 VSS.t2 847.827
R120 VSS.n45 VSS.t8 847.827
R121 VSS.t9 VSS.n44 847.827
R122 VSS.n44 VSS.t6 847.827
R123 VSS.n50 VSS.t4 847.827
R124 VSS.t8 VSS.t9 720.653
R125 VSS.t6 VSS.t4 720.653
R126 VSS.t12 VSS.n37 590.909
R127 VSS.n41 VSS.t12 590.909
R128 VSS.t20 VSS.n41 590.909
R129 VSS.n43 VSS.t23 590.909
R130 VSS.n43 VSS.t16 590.909
R131 VSS.n58 VSS.t14 590.909
R132 VSS.n58 VSS.n57 509.659
R133 VSS.t23 VSS.t20 502.274
R134 VSS.t16 VSS.t14 502.274
R135 VSS.n56 VSS.n50 471.603
R136 VSS.n55 VSS.t21 423.913
R137 VSS.n52 VSS.t21 423.913
R138 VSS.n19 VSS.t0 374.281
R139 VSS.n24 VSS.t0 374.281
R140 VSS.n25 VSS.t10 374.281
R141 VSS.n29 VSS.t10 374.281
R142 VSS.t18 VSS.n32 374.281
R143 VSS.n33 VSS.t18 374.281
R144 VSS.n56 VSS.n55 365.625
R145 VSS.n25 VSS.n24 318.139
R146 VSS.n32 VSS.n29 318.139
R147 VSS.n57 VSS.n12 236.952
R148 VSS.n37 VSS.n36 147.727
R149 VSS.n35 VSS.n33 93.5706
R150 VSS.n59 VSS.n10 87.3061
R151 VSS.n59 VSS.n11 87.3061
R152 VSS.n49 VSS.n13 87.3061
R153 VSS.n49 VSS.n48 87.3061
R154 VSS.n38 VSS.n7 67.4727
R155 VSS.n39 VSS.n7 67.4727
R156 VSS.n15 VSS.n4 67.4727
R157 VSS.n47 VSS.n4 67.4727
R158 VSS.n38 VSS.n10 66.5005
R159 VSS.n39 VSS.n11 66.5005
R160 VSS.n15 VSS.n13 66.5005
R161 VSS.n48 VSS.n47 66.5005
R162 VSS.n54 VSS.n53 44.1404
R163 VSS.n31 VSS.n5 44.1394
R164 VSS.n28 VSS.n26 44.1394
R165 VSS.n23 VSS.n20 44.1394
R166 VSS.n42 VSS.n10 20.8061
R167 VSS.n42 VSS.n11 20.8061
R168 VSS.n40 VSS.n38 20.8061
R169 VSS.n40 VSS.n39 20.8061
R170 VSS.n46 VSS.n15 20.8061
R171 VSS.n47 VSS.n46 20.8061
R172 VSS.n14 VSS.n13 20.8061
R173 VSS.n48 VSS.n14 20.8061
R174 VSS.n30 VSS.t19 4.84702
R175 VSS.n27 VSS.t11 4.84702
R176 VSS.n8 VSS.t13 4.7885
R177 VSS.n9 VSS.t17 4.7885
R178 VSS.n60 VSS.t15 4.7885
R179 VSS.n2 VSS.t7 4.7885
R180 VSS.n3 VSS.t3 4.7885
R181 VSS.n1 VSS.t5 4.7885
R182 VSS.n22 VSS.t1 4.7885
R183 VSS.n51 VSS.t22 4.7885
R184 VSS.n64 VSS.n63 3.51467
R185 VSS.n63 VSS.n7 2.06002
R186 VSS.n21 VSS.n20 1.93869
R187 VSS.n67 VSS.n4 1.90702
R188 VSS.n26 VSS.n18 1.90702
R189 VSS.n66 VSS.n5 1.90702
R190 VSS.n54 VSS.n0 1.90702
R191 VSS.n46 VSS.n3 1.3005
R192 VSS.n46 VSS.n45 1.3005
R193 VSS.n34 VSS.n4 1.3005
R194 VSS.n14 VSS.n2 1.3005
R195 VSS.n44 VSS.n14 1.3005
R196 VSS.n49 VSS.n1 1.3005
R197 VSS.n50 VSS.n49 1.3005
R198 VSS.n20 VSS.n19 1.3005
R199 VSS.n23 VSS.n22 1.3005
R200 VSS.n24 VSS.n23 1.3005
R201 VSS.n26 VSS.n25 1.3005
R202 VSS.n28 VSS.n27 1.3005
R203 VSS.n29 VSS.n28 1.3005
R204 VSS.n31 VSS.n30 1.3005
R205 VSS.n32 VSS.n31 1.3005
R206 VSS.n33 VSS.n5 1.3005
R207 VSS.n37 VSS.n7 1.3005
R208 VSS.n40 VSS.n8 1.3005
R209 VSS.n41 VSS.n40 1.3005
R210 VSS.n42 VSS.n9 1.3005
R211 VSS.n43 VSS.n42 1.3005
R212 VSS.n60 VSS.n59 1.3005
R213 VSS.n59 VSS.n58 1.3005
R214 VSS.n53 VSS.n51 1.3005
R215 VSS.n53 VSS.n52 1.3005
R216 VSS.n55 VSS.n54 1.3005
R217 VSS.n61 VSS.n60 0.771017
R218 VSS.n62 VSS.n8 0.463217
R219 VSS.n61 VSS.n9 0.463217
R220 VSS.n69 VSS.n2 0.463217
R221 VSS.n68 VSS.n3 0.463217
R222 VSS.n70 VSS.n1 0.463217
R223 VSS.n22 VSS.n21 0.463217
R224 VSS.n51 VSS.n0 0.463217
R225 VSS.n62 VSS.n61 0.3083
R226 VSS.n69 VSS.n68 0.3083
R227 VSS.n70 VSS.n69 0.3083
R228 VSS.n68 VSS.n67 0.2165
R229 VSS.n71 VSS.n70 0.1598
R230 VSS.n67 VSS.n66 0.148459
R231 inv2_0.vss VSS.n71 0.1235
R232 VSS.n65 VSS.n6 0.073981
R233 VSS.n63 VSS.n62 0.0635
R234 VSS.n66 VSS.n65 0.0389018
R235 inv2_0.vss VSS.n0 0.0305
R236 VSS.n27 VSS.n6 0.0258591
R237 VSS.n30 VSS.n6 0.0258591
R238 VSS.n65 VSS.n64 0.023066
R239 VSS.n18 or2_0.VSS 0.0158079
R240 VSS.n71 VSS 0.0155
R241 VSS.n21 VSS.n18 0.0139604
R242 VSS.n64 or2_0.VSS 0.00102786
R243 In.n1 In.t1 34.2529
R244 In.n0 In.t0 19.673
R245 In.n0 In.t2 19.4007
R246 and2_1.B In.n1 6.45093
R247 and2_1.B In 1.64621
R248 In.n1 In.n0 0.106438
R249 a_256_n1210.n0 a_256_n1210.t4 34.1797
R250 a_256_n1210.n0 a_256_n1210.t5 19.5798
R251 a_256_n1210.n1 a_256_n1210.t3 18.7717
R252 a_256_n1210.n1 a_256_n1210.t2 9.2885
R253 a_256_n1210.n2 a_256_n1210.n0 4.93379
R254 a_256_n1210.t0 a_256_n1210.n3 4.23346
R255 a_256_n1210.n3 a_256_n1210.t1 3.85546
R256 a_256_n1210.n2 a_256_n1210.n1 0.4055
R257 a_256_n1210.n3 a_256_n1210.n2 0.352625
R258 Bit.n1 Bit.t2 34.1066
R259 Bit.n0 Bit.t1 19.673
R260 Bit.n0 Bit.t0 19.4007
R261 and2_0.A Bit.n1 5.11057
R262 and2_0.A Bit 1.64621
R263 Bit.n1 Bit.n0 0.252687
R264 OUT.n0 OUT.t1 9.6935
R265 OUT.n0 OUT.t0 4.35383
R266 or2_0.OUT OUT.n0 0.260857
R267 or2_0.OUT OUT 0.0905
C0 a_256_n1210.t4 0 0.15843f **FLOATING
C1 a_256_n1210.t5 0 0.07081f **FLOATING
C2 a_256_n1210.n0 0 0.20989f **FLOATING
C3 a_256_n1210.t3 0 0.08492f **FLOATING
C4 a_256_n1210.t2 0 0.04534f **FLOATING
C5 a_256_n1210.n1 0 0.14994f **FLOATING
C6 a_256_n1210.n2 0 0.12745f **FLOATING
C7 a_256_n1210.t1 0 0.144f **FLOATING
C8 a_256_n1210.n3 0 0.92376f **FLOATING
C9 a_256_n1210.t0 0 0.18548f **FLOATING
C10 a_256_1130.t4 0 0.15843f **FLOATING
C11 a_256_1130.t5 0 0.07081f **FLOATING
C12 a_256_1130.n0 0 0.20989f **FLOATING
C13 a_256_1130.t3 0 0.08492f **FLOATING
C14 a_256_1130.t2 0 0.04534f **FLOATING
C15 a_256_1130.n1 0 0.14994f **FLOATING
C16 a_256_1130.n2 0 0.12745f **FLOATING
C17 a_256_1130.t1 0 0.144f **FLOATING
C18 a_256_1130.n3 0 0.92376f **FLOATING
C19 a_256_1130.t0 0 0.18548f **FLOATING
C20 VDD.t21 0 0.00922f **FLOATING
C21 VDD.n0 0 0.04011f **FLOATING
C22 VDD.t1 0 0.00922f **FLOATING
C23 VDD.t0 0 0.07126f **FLOATING
C24 VDD.n1 0 0.15486f **FLOATING
C25 VDD.t9 0 0.00899f **FLOATING
C26 VDD.n2 0 0.02821f **FLOATING
C27 VDD.t17 0 0.00899f **FLOATING
C28 VDD.n3 0 0.02821f **FLOATING
C29 VDD.t15 0 0.00899f **FLOATING
C30 VDD.n4 0 0.02821f **FLOATING
C31 VDD.t5 0 0.00899f **FLOATING
C32 VDD.n5 0 0.02821f **FLOATING
C33 VDD.n6 0 0.01748f **FLOATING
C34 VDD.n7 0 0.01748f **FLOATING
C35 VDD.t14 0 0.0543f **FLOATING
C36 VDD.n8 0 0.01919f **FLOATING
C37 VDD.t16 0 0.05445f **FLOATING
C38 VDD.n9 0 0.06361f **FLOATING
C39 VDD.n10 0 0.01919f **FLOATING
C40 VDD.n11 0 0.00715f **FLOATING
C41 VDD.n12 0 0.0587f **FLOATING
C42 VDD.t11 0 0.0543f **FLOATING
C43 VDD.t10 0 0.0543f **FLOATING
C44 VDD.n13 0 0.00715f **FLOATING
C45 VDD.n14 0 0.0587f **FLOATING
C46 VDD.t4 0 0.05885f **FLOATING
C47 VDD.n15 0 0.06572f **FLOATING
C48 VDD.n16 0 0.25872f **FLOATING
C49 VDD.n17 0 0.06524f **FLOATING
C50 VDD.t3 0 0.00899f **FLOATING
C51 VDD.n18 0 0.02821f **FLOATING
C52 VDD.t13 0 0.00922f **FLOATING
C53 VDD.n19 0 0.01959f **FLOATING
C54 VDD.n20 0 0.01959f **FLOATING
C55 VDD.t2 0 0.05885f **FLOATING
C56 VDD.n21 0 0.00715f **FLOATING
C57 VDD.n22 0 0.0587f **FLOATING
C58 VDD.t12 0 0.05885f **FLOATING
C59 VDD.n23 0 0.05998f **FLOATING
C60 VDD.n24 0 0.04011f **FLOATING
C61 VDD.t7 0 0.00922f **FLOATING
C62 VDD.t6 0 0.07126f **FLOATING
C63 VDD.n25 0 0.15486f **FLOATING
C64 VDD.n26 0 0.05587f **FLOATING
C65 VDD.n27 0 0.02181f **FLOATING
C66 VDD.n28 0 0.1946f **FLOATING
C67 VDD.n29 0 0.6186f **FLOATING
C68 or2_0.VDD 0 0.0396f **FLOATING
C69 VDD.n30 0 0.15447f **FLOATING
C70 VDD.n31 0 0.14304f **FLOATING
C71 VDD.n32 0 0.01959f **FLOATING
C72 VDD.n33 0 0.01959f **FLOATING
C73 VDD.n34 0 0.05998f **FLOATING
C74 VDD.t20 0 0.05885f **FLOATING
C75 VDD.n35 0 0.00715f **FLOATING
C76 VDD.n36 0 0.0587f **FLOATING
C77 VDD.t8 0 0.05885f **FLOATING
C78 VDD.n37 0 0.06391f **FLOATING
C79 VDD.n38 0 0.02556f **FLOATING
C80 VDD.n39 0 0.02996f **FLOATING
C81 VDD.n40 0 0.09644f **FLOATING
C82 VDD 0 0.00719f **FLOATING
C83 VDD.n41 0 0.12527f **FLOATING
C84 VDD.t18 0 0.05975f **FLOATING
C85 VDD.t19 0 0.02365f **FLOATING
C86 VDD.n42 0 0.09385f **FLOATING
C87 inv2_0.vdd 0 0.19111f **FLOATING
